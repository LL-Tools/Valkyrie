

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4368, n4369, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496;

  INV_X4 U4873 ( .A(n8945), .ZN(n8924) );
  AND2_X1 U4874 ( .A1(n9844), .A2(n9833), .ZN(n9814) );
  INV_X1 U4875 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n8489) );
  INV_X1 U4876 ( .A(n5643), .ZN(n5683) );
  INV_X1 U4877 ( .A(n9157), .ZN(n8295) );
  BUF_X1 U4878 ( .A(n6371), .Z(n4388) );
  INV_X1 U4879 ( .A(n7780), .ZN(n9647) );
  BUF_X2 U4881 ( .A(n5177), .Z(n5819) );
  CLKBUF_X2 U4882 ( .A(n5127), .Z(n4393) );
  INV_X1 U4883 ( .A(n10391), .ZN(n7352) );
  INV_X1 U4884 ( .A(n4397), .ZN(n6727) );
  INV_X1 U4885 ( .A(n8489), .ZN(n4368) );
  INV_X1 U4886 ( .A(n4368), .ZN(n4369) );
  INV_X1 U4887 ( .A(n4368), .ZN(P2_U3152) );
  NAND2_X1 U4888 ( .A1(n7335), .A2(n6810), .ZN(n5831) );
  NAND2_X1 U4889 ( .A1(n7024), .A2(n9159), .ZN(n7299) );
  OR2_X1 U4890 ( .A1(n6172), .A2(n6872), .ZN(n6183) );
  NAND2_X1 U4891 ( .A1(n8175), .A2(n8179), .ZN(n8916) );
  INV_X2 U4892 ( .A(n7299), .ZN(n7733) );
  NAND2_X1 U4893 ( .A1(n6393), .A2(n9550), .ZN(n7018) );
  INV_X1 U4895 ( .A(n5826), .ZN(n5525) );
  AND2_X1 U4896 ( .A1(n5160), .A2(n4829), .ZN(n7570) );
  INV_X1 U4897 ( .A(n6829), .ZN(n6401) );
  CLKBUF_X3 U4898 ( .A(n6077), .Z(n6829) );
  NAND2_X1 U4899 ( .A1(n9982), .A2(n9965), .ZN(n9964) );
  OAI211_X1 U4900 ( .C1(n9409), .C2(n6731), .A(n6089), .B(n6088), .ZN(n7972)
         );
  NAND2_X1 U4901 ( .A1(n5582), .A2(n5581), .ZN(n8987) );
  NAND2_X2 U4902 ( .A1(n5306), .A2(n5305), .ZN(n9052) );
  INV_X1 U4903 ( .A(n10400), .ZN(n10424) );
  NAND2_X1 U4904 ( .A1(n9516), .A2(n9514), .ZN(n9899) );
  NAND2_X1 U4905 ( .A1(n9556), .A2(n9555), .ZN(n9583) );
  AOI21_X1 U4907 ( .B1(n9771), .B2(n9981), .A(n9770), .ZN(n10065) );
  XNOR2_X1 U4908 ( .A(n6031), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6032) );
  INV_X1 U4909 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10198) );
  NAND4_X1 U4910 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n8604)
         );
  INV_X2 U4911 ( .A(n10036), .ZN(n10021) );
  OR2_X1 U4912 ( .A1(n8250), .A2(n9277), .ZN(n4371) );
  AND2_X2 U4913 ( .A1(n6189), .A2(n6000), .ZN(n4372) );
  AND2_X1 U4914 ( .A1(n9235), .A2(n8236), .ZN(n4373) );
  AND2_X2 U4915 ( .A1(n9400), .A2(n9399), .ZN(n9577) );
  OR2_X2 U4916 ( .A1(n9210), .A2(n9211), .ZN(n4743) );
  BUF_X1 U4917 ( .A(n5289), .Z(n4390) );
  AOI21_X2 U4918 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4813) );
  NAND2_X2 U4919 ( .A1(n5300), .A2(n4656), .ZN(n4659) );
  OAI211_X2 U4920 ( .C1(n7778), .C2(n4880), .A(n4877), .B(n9440), .ZN(n8022)
         );
  NAND2_X1 U4921 ( .A1(n6809), .A2(n6810), .ZN(n7045) );
  NAND2_X2 U4922 ( .A1(n4776), .A2(n4781), .ZN(n5655) );
  XNOR2_X2 U4923 ( .A(n5375), .B(n5009), .ZN(n6779) );
  BUF_X2 U4925 ( .A(n8969), .Z(n4375) );
  NAND2_X1 U4926 ( .A1(n5642), .A2(n5641), .ZN(n8969) );
  OR2_X1 U4927 ( .A1(n9052), .A2(n8455), .ZN(n5895) );
  AOI22_X2 U4928 ( .A1(n8003), .A2(n8002), .B1(n9052), .B2(n8601), .ZN(n8004)
         );
  NAND2_X1 U4929 ( .A1(n5043), .A2(n4818), .ZN(n4376) );
  OAI21_X1 U4930 ( .B1(n4812), .B2(n4810), .A(n4809), .ZN(n4808) );
  AND2_X2 U4931 ( .A1(n7507), .A2(n8874), .ZN(n5989) );
  OAI21_X1 U4932 ( .B1(n5865), .B2(n5872), .A(n5864), .ZN(n5866) );
  INV_X2 U4933 ( .A(n7571), .ZN(n8607) );
  NAND2_X2 U4934 ( .A1(n6223), .A2(n6222), .ZN(n10136) );
  NAND2_X2 U4935 ( .A1(n4755), .A2(n4754), .ZN(n5434) );
  NAND2_X2 U4936 ( .A1(n5691), .A2(n5690), .ZN(n8959) );
  AOI211_X2 U4937 ( .C1(n4400), .C2(n5939), .A(n8730), .B(n8706), .ZN(n5947)
         );
  NAND2_X2 U4938 ( .A1(n5340), .A2(n5339), .ZN(n9046) );
  XNOR2_X2 U4939 ( .A(n5448), .B(n5011), .ZN(n6802) );
  AOI22_X2 U4940 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .B1(n10199), .B2(n10198), .ZN(n10492) );
  OR2_X2 U4941 ( .A1(n10067), .A2(n9800), .ZN(n9531) );
  NAND2_X2 U4942 ( .A1(n6373), .A2(n6372), .ZN(n9757) );
  OAI22_X2 U4943 ( .A1(n8149), .A2(n4995), .B1(n4996), .B2(n4997), .ZN(n8334)
         );
  NAND2_X2 U4944 ( .A1(n8005), .A2(n8004), .ZN(n8149) );
  NAND2_X2 U4945 ( .A1(n5032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5028) );
  XNOR2_X2 U4946 ( .A(n5051), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5851) );
  XNOR2_X2 U4947 ( .A(n5618), .B(n5614), .ZN(n7950) );
  INV_X2 U4948 ( .A(n7733), .ZN(n8297) );
  INV_X1 U4949 ( .A(n7972), .ZN(n10267) );
  OAI21_X2 U4950 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10449), .ZN(n10478) );
  NAND2_X1 U4951 ( .A1(n8729), .A2(n8352), .ZN(n8707) );
  NAND2_X1 U4952 ( .A1(n4380), .A2(n8349), .ZN(n8784) );
  NAND2_X1 U4953 ( .A1(n9535), .A2(n9764), .ZN(n9605) );
  NAND2_X1 U4954 ( .A1(n4532), .A2(n4531), .ZN(n5948) );
  AND2_X2 U4955 ( .A1(n9531), .A2(n9532), .ZN(n9780) );
  OR2_X1 U4956 ( .A1(n10072), .A2(n9215), .ZN(n9527) );
  INV_X1 U4957 ( .A(n9876), .ZN(n4377) );
  NAND2_X1 U4958 ( .A1(n8234), .A2(n8233), .ZN(n9238) );
  OR2_X1 U4959 ( .A1(n6376), .A2(n6375), .ZN(n6398) );
  NAND2_X1 U4960 ( .A1(n6286), .A2(n6285), .ZN(n10108) );
  NAND2_X1 U4961 ( .A1(n4480), .A2(n4479), .ZN(n5002) );
  NAND2_X1 U4962 ( .A1(n10128), .A2(n9997), .ZN(n9433) );
  MUX2_X1 U4963 ( .A(n5860), .B(n5869), .S(n5976), .Z(n5872) );
  NAND2_X1 U4964 ( .A1(n10298), .A2(n7876), .ZN(n9454) );
  AND2_X1 U4965 ( .A1(n9558), .A2(n9371), .ZN(n9581) );
  INV_X1 U4966 ( .A(n8217), .ZN(n4378) );
  AND2_X1 U4967 ( .A1(n10265), .A2(n8015), .ZN(n8013) );
  INV_X2 U4968 ( .A(n7615), .ZN(n7075) );
  AND4_X1 U4969 ( .A1(n6109), .A2(n6108), .A3(n6106), .A4(n6107), .ZN(n6139)
         );
  NAND4_X1 U4970 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n7614)
         );
  INV_X1 U4971 ( .A(n8938), .ZN(n7270) );
  NAND2_X1 U4972 ( .A1(n10380), .A2(n10381), .ZN(n7335) );
  INV_X1 U4973 ( .A(n5137), .ZN(n4379) );
  NOR2_X1 U4974 ( .A1(n10475), .A2(n10207), .ZN(n10208) );
  CLKBUF_X2 U4975 ( .A(n4620), .Z(n6350) );
  OR2_X1 U4976 ( .A1(n6065), .A2(n6770), .ZN(n6055) );
  INV_X1 U4977 ( .A(n9409), .ZN(n6371) );
  XNOR2_X1 U4978 ( .A(n6014), .B(n6013), .ZN(n6397) );
  NAND2_X2 U4979 ( .A1(n6727), .A2(P1_U3084), .ZN(n10182) );
  AND2_X1 U4980 ( .A1(n6427), .A2(n6231), .ZN(n6241) );
  NOR2_X1 U4981 ( .A1(n4568), .A2(n6009), .ZN(n4566) );
  CLKBUF_X2 U4982 ( .A(n5249), .Z(n4396) );
  CLKBUF_X3 U4983 ( .A(n5249), .Z(n4391) );
  CLKBUF_X3 U4984 ( .A(n5249), .Z(n4392) );
  NAND3_X1 U4985 ( .A1(n8644), .A2(n4789), .A3(n4788), .ZN(n4787) );
  NOR2_X1 U4986 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6007) );
  AND2_X1 U4987 ( .A1(n5982), .A2(n7507), .ZN(n5984) );
  OAI21_X1 U4988 ( .B1(n8962), .B2(n8924), .A(n4894), .ZN(n4893) );
  OR2_X1 U4989 ( .A1(n8975), .A2(n8974), .ZN(n9070) );
  AND2_X1 U4990 ( .A1(n4542), .A2(n9625), .ZN(n4541) );
  AOI21_X1 U4991 ( .B1(n4743), .B2(n4739), .A(n9340), .ZN(n4602) );
  OR2_X1 U4992 ( .A1(n9624), .A2(n9623), .ZN(n4542) );
  NAND2_X1 U4993 ( .A1(n9546), .A2(n9545), .ZN(n4546) );
  NOR2_X1 U4994 ( .A1(n8701), .A2(n8700), .ZN(n8967) );
  OR2_X1 U4995 ( .A1(n4681), .A2(n4687), .ZN(n4680) );
  AOI21_X1 U4996 ( .B1(n4682), .B2(n4688), .A(n4471), .ZN(n4681) );
  OR3_X1 U4997 ( .A1(n9610), .A2(n10061), .A3(n9609), .ZN(n9612) );
  AOI21_X1 U4998 ( .B1(n9784), .B2(n9981), .A(n9783), .ZN(n10070) );
  NAND2_X1 U4999 ( .A1(n8292), .A2(n8291), .ZN(n9289) );
  NOR2_X1 U5000 ( .A1(n5962), .A2(n5955), .ZN(n4690) );
  NAND2_X1 U5001 ( .A1(n8725), .A2(n8726), .ZN(n8724) );
  NOR2_X1 U5002 ( .A1(n4689), .A2(n8652), .ZN(n4688) );
  NAND2_X1 U5003 ( .A1(n5968), .A2(n5969), .ZN(n8657) );
  OR2_X1 U5004 ( .A1(n10043), .A2(n9749), .ZN(n9606) );
  NAND2_X1 U5005 ( .A1(n9411), .A2(n9410), .ZN(n10043) );
  AND2_X1 U5006 ( .A1(n5782), .A2(n5963), .ZN(n8677) );
  NOR2_X1 U5007 ( .A1(n9760), .A2(n10050), .ZN(n9759) );
  NAND2_X1 U5008 ( .A1(n5798), .A2(n5797), .ZN(n8652) );
  NAND2_X1 U5009 ( .A1(n5821), .A2(n5820), .ZN(n8952) );
  OR2_X1 U5010 ( .A1(n8662), .A2(n7511), .ZN(n5968) );
  NAND2_X1 U5011 ( .A1(n8784), .A2(n4986), .ZN(n4985) );
  NAND2_X1 U5012 ( .A1(n5791), .A2(n5790), .ZN(n8662) );
  AND2_X1 U5013 ( .A1(n9780), .A2(n4861), .ZN(n4860) );
  NAND2_X1 U5014 ( .A1(n9345), .A2(n9344), .ZN(n10050) );
  XNOR2_X1 U5015 ( .A(n5796), .B(n5795), .ZN(n9401) );
  NOR2_X1 U5016 ( .A1(n8959), .A2(n8699), .ZN(n5955) );
  NAND2_X1 U5017 ( .A1(n8756), .A2(n4826), .ZN(n8755) );
  OR2_X1 U5018 ( .A1(n9757), .A2(n9769), .ZN(n9535) );
  INV_X1 U5019 ( .A(n9797), .ZN(n9603) );
  NAND2_X1 U5020 ( .A1(n4974), .A2(n4975), .ZN(n4380) );
  NAND2_X1 U5021 ( .A1(n5948), .A2(n8695), .ZN(n8706) );
  AND2_X1 U5022 ( .A1(n4885), .A2(n9347), .ZN(n4884) );
  NOR2_X1 U5023 ( .A1(n9807), .A2(n9808), .ZN(n6415) );
  NAND2_X1 U5024 ( .A1(n8964), .A2(n8354), .ZN(n5956) );
  XNOR2_X1 U5025 ( .A(n5815), .B(n5789), .ZN(n9342) );
  NAND2_X1 U5026 ( .A1(n8711), .A2(n5829), .ZN(n8730) );
  NAND2_X1 U5027 ( .A1(n9527), .A2(n9528), .ZN(n9797) );
  INV_X1 U5028 ( .A(n5944), .ZN(n5775) );
  OR2_X1 U5029 ( .A1(n8976), .A2(n8502), .ZN(n8711) );
  NAND2_X1 U5030 ( .A1(n5788), .A2(n5787), .ZN(n5815) );
  AND2_X1 U5031 ( .A1(n8692), .A2(n8595), .ZN(n8676) );
  NAND2_X1 U5032 ( .A1(n8805), .A2(n5919), .ZN(n8789) );
  NAND2_X1 U5033 ( .A1(n4375), .A2(n8698), .ZN(n8695) );
  NAND2_X1 U5034 ( .A1(n6364), .A2(n6363), .ZN(n10067) );
  NAND2_X1 U5035 ( .A1(n4473), .A2(n6351), .ZN(n10072) );
  AND2_X1 U5036 ( .A1(n8748), .A2(n8757), .ZN(n5944) );
  INV_X1 U5037 ( .A(n4624), .ZN(n4623) );
  OAI21_X1 U5038 ( .B1(n8422), .B2(n5478), .A(n5505), .ZN(n8437) );
  AND2_X1 U5039 ( .A1(n8982), .A2(n8499), .ZN(n5939) );
  NAND2_X1 U5040 ( .A1(n9098), .A2(n5819), .ZN(n5642) );
  NOR3_X1 U5041 ( .A1(n9907), .A2(n4399), .A3(n4417), .ZN(n4622) );
  OR2_X1 U5042 ( .A1(n9836), .A2(n9852), .ZN(n9572) );
  NAND2_X1 U5043 ( .A1(n5588), .A2(n5587), .ZN(n8982) );
  XNOR2_X1 U5044 ( .A(n5686), .B(n5685), .ZN(n9095) );
  NAND2_X1 U5045 ( .A1(n4775), .A2(n4773), .ZN(n5686) );
  NAND2_X1 U5046 ( .A1(n4845), .A2(n4842), .ZN(n10111) );
  NAND2_X1 U5047 ( .A1(n6321), .A2(n6320), .ZN(n10089) );
  OR2_X1 U5048 ( .A1(n10092), .A2(n9886), .ZN(n9864) );
  NAND2_X1 U5049 ( .A1(n5557), .A2(n5556), .ZN(n8992) );
  AND2_X1 U5050 ( .A1(n4844), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U5051 ( .A1(n6310), .A2(n6309), .ZN(n10092) );
  AND2_X1 U5052 ( .A1(n6018), .A2(n6017), .ZN(n9876) );
  AND2_X1 U5053 ( .A1(n5765), .A2(n8825), .ZN(n8859) );
  NAND2_X1 U5054 ( .A1(n5537), .A2(n5536), .ZN(n9000) );
  AND2_X1 U5055 ( .A1(n6360), .A2(n6359), .ZN(n9215) );
  OR2_X1 U5056 ( .A1(n10103), .A2(n9917), .ZN(n9516) );
  AOI21_X1 U5057 ( .B1(n4867), .B2(n4870), .A(n4864), .ZN(n4863) );
  INV_X1 U5058 ( .A(n5771), .ZN(n9004) );
  NOR2_X1 U5059 ( .A1(n4847), .A2(n9943), .ZN(n4846) );
  NAND2_X1 U5060 ( .A1(n6298), .A2(n6297), .ZN(n10103) );
  AND2_X1 U5061 ( .A1(n9435), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U5062 ( .A1(n5458), .A2(n5457), .ZN(n9014) );
  NAND2_X1 U5063 ( .A1(n6352), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U5064 ( .A1(n5489), .A2(n5488), .ZN(n8837) );
  AOI21_X2 U5065 ( .B1(n7835), .B2(n7836), .A(n5237), .ZN(n7863) );
  NAND2_X1 U5066 ( .A1(n6271), .A2(n6270), .ZN(n10113) );
  AOI21_X1 U5067 ( .B1(n4586), .B2(n4584), .A(n4444), .ZN(n4583) );
  AOI21_X1 U5068 ( .B1(n4734), .B2(n4736), .A(n4732), .ZN(n4731) );
  NOR2_X1 U5069 ( .A1(n8201), .A2(n4587), .ZN(n4586) );
  OR2_X1 U5070 ( .A1(n9024), .A2(n8487), .ZN(n5830) );
  NAND2_X1 U5071 ( .A1(n5470), .A2(n5469), .ZN(n9020) );
  NAND2_X1 U5072 ( .A1(n6234), .A2(n6233), .ZN(n10125) );
  OAI21_X1 U5073 ( .B1(n7752), .B2(n4736), .A(n8064), .ZN(n4735) );
  INV_X1 U5074 ( .A(n5904), .ZN(n5760) );
  NAND2_X1 U5075 ( .A1(n5417), .A2(n5416), .ZN(n9024) );
  NAND2_X1 U5076 ( .A1(n6258), .A2(n6257), .ZN(n10119) );
  AND2_X1 U5077 ( .A1(n5899), .A2(n5900), .ZN(n8148) );
  NAND2_X1 U5078 ( .A1(n6245), .A2(n6244), .ZN(n10128) );
  AND2_X1 U5079 ( .A1(n8180), .A2(n8458), .ZN(n5904) );
  NAND2_X1 U5080 ( .A1(n5440), .A2(n5439), .ZN(n9030) );
  NAND2_X1 U5081 ( .A1(n5380), .A2(n5379), .ZN(n9035) );
  OR2_X1 U5082 ( .A1(n9046), .A2(n8153), .ZN(n5899) );
  NAND2_X1 U5083 ( .A1(n6210), .A2(n6209), .ZN(n10141) );
  NAND2_X1 U5084 ( .A1(n5364), .A2(n5363), .ZN(n8180) );
  AND2_X1 U5085 ( .A1(n5881), .A2(n7677), .ZN(n4890) );
  AND2_X1 U5086 ( .A1(n5890), .A2(n8125), .ZN(n7921) );
  CLKBUF_X1 U5087 ( .A(n10422), .Z(n4523) );
  NAND2_X1 U5088 ( .A1(n6181), .A2(n6180), .ZN(n10031) );
  NAND2_X1 U5089 ( .A1(n5226), .A2(n5225), .ZN(n10422) );
  NAND2_X1 U5090 ( .A1(n7382), .A2(n7381), .ZN(n7691) );
  AND2_X1 U5091 ( .A1(n5288), .A2(n5287), .ZN(n8142) );
  XNOR2_X1 U5092 ( .A(n5328), .B(n5323), .ZN(n6746) );
  NAND2_X1 U5093 ( .A1(n5257), .A2(n5256), .ZN(n9061) );
  AND2_X1 U5094 ( .A1(n5876), .A2(n5873), .ZN(n7532) );
  NOR2_X1 U5095 ( .A1(n10213), .A2(n10484), .ZN(n10214) );
  NAND2_X1 U5096 ( .A1(n5201), .A2(n5200), .ZN(n7669) );
  NAND2_X1 U5097 ( .A1(n6131), .A2(n6130), .ZN(n10298) );
  NOR2_X1 U5098 ( .A1(n10486), .A2(n10485), .ZN(n10484) );
  INV_X1 U5099 ( .A(n7542), .ZN(n10414) );
  AND2_X1 U5100 ( .A1(n5181), .A2(n5180), .ZN(n7542) );
  INV_X1 U5101 ( .A(n4381), .ZN(n7055) );
  NAND2_X1 U5102 ( .A1(n6127), .A2(n6126), .ZN(n7786) );
  NAND2_X2 U5103 ( .A1(n7065), .A2(n7018), .ZN(n9157) );
  XNOR2_X1 U5104 ( .A(n5216), .B(n5214), .ZN(n6734) );
  AND4_X1 U5105 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n8455)
         );
  AND4_X1 U5106 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n7876)
         );
  INV_X1 U5107 ( .A(n7301), .ZN(n9648) );
  INV_X1 U5108 ( .A(n7517), .ZN(n8609) );
  CLKBUF_X1 U5109 ( .A(n5289), .Z(n4389) );
  AND4_X2 U5110 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n9364)
         );
  AND4_X1 U5111 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n7301)
         );
  NAND2_X1 U5112 ( .A1(n5196), .A2(n5195), .ZN(n5277) );
  NAND2_X1 U5113 ( .A1(n5176), .A2(n5175), .ZN(n5196) );
  NAND3_X1 U5114 ( .A1(n6816), .A2(n5720), .A3(n7609), .ZN(n5059) );
  CLKBUF_X1 U5115 ( .A(n5720), .Z(n5983) );
  INV_X1 U5116 ( .A(n5137), .ZN(n4394) );
  XNOR2_X1 U5117 ( .A(n6283), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9740) );
  INV_X1 U5118 ( .A(n5851), .ZN(n7609) );
  INV_X1 U5119 ( .A(n6396), .ZN(n9550) );
  NAND2_X1 U5120 ( .A1(n6029), .A2(n6030), .ZN(n8186) );
  XNOR2_X1 U5121 ( .A(n6432), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6438) );
  AND2_X1 U5122 ( .A1(n5033), .A2(n5032), .ZN(n5035) );
  MUX2_X1 U5123 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6028), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n6029) );
  INV_X2 U5124 ( .A(n6085), .ZN(n6284) );
  XNOR2_X1 U5125 ( .A(n6388), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6396) );
  CLKBUF_X1 U5126 ( .A(n6848), .Z(n10184) );
  NAND2_X1 U5127 ( .A1(n5050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5051) );
  OAI21_X1 U5128 ( .B1(n6282), .B2(n4404), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6388) );
  NAND2_X1 U5129 ( .A1(n5029), .A2(n5027), .ZN(n5032) );
  NAND2_X1 U5130 ( .A1(n4598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U5131 ( .A1(n4607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5132 ( .A1(n5219), .A2(n5218), .ZN(n5273) );
  NAND2_X2 U5133 ( .A1(n5026), .A2(n5025), .ZN(n5042) );
  NAND2_X2 U5134 ( .A1(n4391), .A2(P1_U3084), .ZN(n10186) );
  NAND3_X1 U5135 ( .A1(n5047), .A2(n5046), .A3(n4606), .ZN(n4607) );
  AND2_X1 U5136 ( .A1(n6003), .A2(n4565), .ZN(n4567) );
  AND3_X1 U5137 ( .A1(n5999), .A2(n5998), .A3(n5997), .ZN(n6189) );
  NOR3_X1 U5138 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .A3(
        P1_IR_REG_12__SCAN_IN), .ZN(n6000) );
  INV_X1 U5139 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6231) );
  NOR2_X1 U5140 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6001) );
  INV_X1 U5141 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U5142 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5997) );
  NOR2_X1 U5143 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5998) );
  NOR2_X1 U5144 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5999) );
  INV_X1 U5145 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6265) );
  INV_X1 U5146 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6254) );
  INV_X1 U5147 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4788) );
  INV_X1 U5148 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5044) );
  INV_X1 U5149 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5698) );
  NOR2_X1 U5150 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4616) );
  NOR2_X1 U5151 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4615) );
  INV_X1 U5152 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8644) );
  INV_X4 U5153 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U5154 ( .A1(n4985), .A2(n4647), .ZN(n4492) );
  XNOR2_X1 U5155 ( .A(n8609), .B(n7311), .ZN(n4381) );
  OAI21_X1 U5156 ( .B1(n7051), .B2(n4381), .A(n7313), .ZN(n8928) );
  NAND2_X1 U5157 ( .A1(n7050), .A2(n4381), .ZN(n7313) );
  NAND2_X2 U5158 ( .A1(n4817), .A2(n4397), .ZN(n5137) );
  NAND2_X2 U5159 ( .A1(n5043), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5160 ( .A1(n4379), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5066) );
  INV_X1 U5161 ( .A(n4382), .ZN(n8670) );
  OAI21_X2 U5162 ( .B1(n8705), .B2(n8694), .A(n4654), .ZN(n4382) );
  NAND2_X2 U5163 ( .A1(n8707), .A2(n8706), .ZN(n8705) );
  NOR2_X2 U5164 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4385) );
  NOR2_X2 U5165 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4383) );
  NOR2_X2 U5166 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4384) );
  AND3_X2 U5167 ( .A1(n4385), .A2(n4384), .A3(n4383), .ZN(n5017) );
  AND4_X4 U5168 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n5754)
         );
  NAND3_X1 U5169 ( .A1(n6054), .A2(n4916), .A3(n6055), .ZN(n9363) );
  OAI221_X1 U5170 ( .B1(n6634), .B2(keyinput108), .C1(n5040), .C2(keyinput63), 
        .A(n6633), .ZN(n6637) );
  AND4_X2 U5171 ( .A1(n5039), .A2(n5038), .A3(n5036), .A4(n5037), .ZN(n10380)
         );
  NOR2_X2 U5172 ( .A1(n8651), .A2(n8652), .ZN(n8650) );
  OAI211_X1 U5173 ( .C1(n5434), .C2(n4664), .A(n4661), .B(n4660), .ZN(n6975)
         );
  NAND2_X1 U5174 ( .A1(n5623), .A2(n5622), .ZN(n8976) );
  OAI21_X1 U5175 ( .B1(n5618), .B2(n4785), .A(n5617), .ZN(n5636) );
  INV_X1 U5176 ( .A(n5313), .ZN(n5289) );
  NAND2_X2 U5177 ( .A1(n7279), .A2(n7018), .ZN(n7022) );
  OR4_X2 U5178 ( .A1(n8669), .A2(n10418), .A3(n8656), .A4(n8657), .ZN(n8364)
         );
  AND2_X2 U5179 ( .A1(n8158), .A2(n9040), .ZN(n8175) );
  NAND2_X2 U5180 ( .A1(n6085), .A2(n6727), .ZN(n9409) );
  NAND2_X1 U5181 ( .A1(n5177), .A2(n6730), .ZN(n5121) );
  OAI222_X1 U5182 ( .A1(n4369), .A2(n8367), .B1(n9101), .B2(n8369), .C1(n8368), 
        .C2(n8378), .ZN(P2_U3328) );
  AND2_X2 U5183 ( .A1(n8381), .A2(n8367), .ZN(n5129) );
  NAND2_X1 U5184 ( .A1(n5852), .A2(n5853), .ZN(n7046) );
  AND2_X1 U5185 ( .A1(n4896), .A2(n4895), .ZN(n8962) );
  NOR2_X2 U5186 ( .A1(n6009), .A2(n6008), .ZN(n6426) );
  AND2_X2 U5187 ( .A1(n5034), .A2(n5035), .ZN(n5127) );
  INV_X2 U5188 ( .A(n5128), .ZN(n5593) );
  AND2_X2 U5189 ( .A1(n5034), .A2(n8381), .ZN(n5128) );
  AOI211_X1 U5190 ( .C1(n5930), .C2(n5929), .A(n5928), .B(n5927), .ZN(n5935)
         );
  AND2_X4 U5191 ( .A1(n7630), .A2(n7279), .ZN(n8237) );
  INV_X2 U5192 ( .A(n5034), .ZN(n8367) );
  OAI21_X4 U5193 ( .B1(n8705), .B2(n4653), .A(n4651), .ZN(n8669) );
  INV_X1 U5194 ( .A(n5137), .ZN(n4395) );
  INV_X2 U5195 ( .A(n8927), .ZN(n7311) );
  INV_X2 U5196 ( .A(n6120), .ZN(n6213) );
  OAI21_X2 U5197 ( .B1(n8340), .B2(n4991), .A(n4990), .ZN(n8858) );
  BUF_X8 U5198 ( .A(n5249), .Z(n4397) );
  AND2_X1 U5199 ( .A1(n5035), .A2(n8367), .ZN(n4398) );
  INV_X1 U5200 ( .A(n4690), .ZN(n4682) );
  INV_X1 U5201 ( .A(n8676), .ZN(n5828) );
  INV_X1 U5202 ( .A(n5597), .ZN(n5589) );
  INV_X1 U5203 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5023) );
  AND4_X1 U5204 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n6682), .ZN(n5021)
         );
  NOR2_X1 U5205 ( .A1(n9757), .A2(n4921), .ZN(n4920) );
  NAND2_X1 U5206 ( .A1(n9779), .A2(n6422), .ZN(n4921) );
  AOI21_X1 U5207 ( .B1(n4670), .B2(n4668), .A(n4667), .ZN(n4666) );
  INV_X1 U5208 ( .A(n5401), .ZN(n4668) );
  NAND2_X1 U5209 ( .A1(n4659), .A2(n4433), .ZN(n5356) );
  INV_X1 U5210 ( .A(n5353), .ZN(n4658) );
  AND2_X1 U5211 ( .A1(n5604), .A2(n5603), .ZN(n8538) );
  NAND2_X1 U5212 ( .A1(n8743), .A2(n5775), .ZN(n8725) );
  OR2_X1 U5213 ( .A1(n9046), .A2(n8600), .ZN(n8147) );
  INV_X1 U5214 ( .A(n9527), .ZN(n4862) );
  NOR2_X1 U5215 ( .A1(n4623), .A2(n4417), .ZN(n4621) );
  AOI21_X1 U5216 ( .B1(n4641), .B2(n4646), .A(n4439), .ZN(n4639) );
  INV_X1 U5217 ( .A(n6008), .ZN(n4565) );
  AOI21_X1 U5218 ( .B1(n4795), .B2(n8150), .A(n5905), .ZN(n4793) );
  INV_X1 U5219 ( .A(n5901), .ZN(n4795) );
  INV_X1 U5220 ( .A(n5917), .ZN(n4814) );
  NAND2_X1 U5221 ( .A1(n4558), .A2(n4557), .ZN(n4556) );
  NOR2_X1 U5222 ( .A1(n9491), .A2(n9540), .ZN(n4557) );
  NAND2_X1 U5223 ( .A1(n9494), .A2(n9962), .ZN(n4558) );
  INV_X1 U5224 ( .A(n5958), .ZN(n5960) );
  NAND2_X1 U5225 ( .A1(n9780), .A2(n9529), .ZN(n4564) );
  NAND2_X1 U5226 ( .A1(n8695), .A2(n4530), .ZN(n5776) );
  INV_X1 U5227 ( .A(n9526), .ZN(n4561) );
  NAND2_X1 U5228 ( .A1(n7075), .A2(n7161), .ZN(n9366) );
  OR2_X1 U5229 ( .A1(n5787), .A2(SI_29_), .ZN(n4752) );
  NAND2_X1 U5230 ( .A1(n5358), .A2(n6667), .ZN(n5376) );
  NOR2_X1 U5231 ( .A1(n8037), .A2(n4954), .ZN(n4953) );
  INV_X1 U5232 ( .A(n5270), .ZN(n4954) );
  NAND2_X1 U5233 ( .A1(n5126), .A2(n7512), .ZN(n4948) );
  AND2_X1 U5234 ( .A1(n4690), .A2(n5823), .ZN(n4687) );
  OR2_X1 U5235 ( .A1(n8992), .A2(n8794), .ZN(n5933) );
  INV_X1 U5236 ( .A(n5927), .ZN(n5919) );
  OR2_X1 U5237 ( .A1(n9035), .A2(n8335), .ZN(n5906) );
  NOR2_X1 U5238 ( .A1(n4677), .A2(n8127), .ZN(n4676) );
  INV_X1 U5239 ( .A(n5895), .ZN(n4677) );
  NAND2_X1 U5240 ( .A1(n5058), .A2(n8640), .ZN(n6816) );
  AND2_X1 U5241 ( .A1(n5048), .A2(n4960), .ZN(n4959) );
  INV_X1 U5242 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4960) );
  INV_X1 U5243 ( .A(n4607), .ZN(n5052) );
  NAND2_X1 U5244 ( .A1(n4571), .A2(n4569), .ZN(n8268) );
  INV_X1 U5245 ( .A(n8192), .ZN(n4587) );
  INV_X1 U5246 ( .A(n8186), .ZN(n6033) );
  NAND2_X1 U5247 ( .A1(n9584), .A2(n7825), .ZN(n6141) );
  INV_X1 U5248 ( .A(n9836), .ZN(n9833) );
  AND2_X1 U5249 ( .A1(n9550), .A2(n9615), .ZN(n7023) );
  NAND2_X1 U5250 ( .A1(n9629), .A2(n9615), .ZN(n7065) );
  INV_X1 U5251 ( .A(n6096), .ZN(n6003) );
  INV_X1 U5252 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6002) );
  NOR2_X1 U5253 ( .A1(n5635), .A2(n4784), .ZN(n4783) );
  INV_X1 U5254 ( .A(n5617), .ZN(n4784) );
  NAND2_X1 U5255 ( .A1(n5513), .A2(n6523), .ZN(n5534) );
  NAND2_X1 U5256 ( .A1(n5433), .A2(n5401), .ZN(n4671) );
  NAND2_X1 U5257 ( .A1(n5398), .A2(n5397), .ZN(n5401) );
  INV_X1 U5258 ( .A(SI_15_), .ZN(n5397) );
  AOI21_X1 U5259 ( .B1(n4405), .B2(n4759), .A(n4446), .ZN(n4754) );
  AOI21_X1 U5260 ( .B1(n5009), .B2(n4758), .A(n4757), .ZN(n4756) );
  INV_X1 U5261 ( .A(n5376), .ZN(n4757) );
  INV_X1 U5262 ( .A(n5355), .ZN(n4758) );
  INV_X1 U5263 ( .A(n5009), .ZN(n4759) );
  NAND2_X1 U5264 ( .A1(n5355), .A2(n5332), .ZN(n5353) );
  INV_X1 U5265 ( .A(n4932), .ZN(n4931) );
  OAI21_X1 U5266 ( .B1(n8572), .B2(n4933), .A(n4939), .ZN(n4932) );
  NAND2_X1 U5267 ( .A1(n5652), .A2(n5653), .ZN(n4939) );
  NAND2_X1 U5268 ( .A1(n8466), .A2(n8469), .ZN(n4933) );
  AND2_X1 U5269 ( .A1(n5530), .A2(n5509), .ZN(n4958) );
  INV_X1 U5270 ( .A(n4948), .ZN(n4945) );
  OAI21_X1 U5271 ( .B1(n8413), .B2(n4948), .A(n7514), .ZN(n4947) );
  AND2_X1 U5272 ( .A1(n5742), .A2(n7266), .ZN(n5740) );
  AND2_X1 U5273 ( .A1(n5545), .A2(n5544), .ZN(n8536) );
  NAND2_X1 U5274 ( .A1(n7098), .A2(n7099), .ZN(n7190) );
  NAND2_X1 U5275 ( .A1(n8355), .A2(n8686), .ZN(n4653) );
  NAND2_X1 U5276 ( .A1(n8355), .A2(n4652), .ZN(n4651) );
  NOR2_X1 U5277 ( .A1(n8505), .A2(n8406), .ZN(n4533) );
  NAND2_X1 U5278 ( .A1(n4492), .A2(n8351), .ZN(n8731) );
  AND2_X1 U5279 ( .A1(n4984), .A2(n8740), .ZN(n4647) );
  NAND2_X1 U5280 ( .A1(n8755), .A2(n4694), .ZN(n8743) );
  AND2_X1 U5281 ( .A1(n4648), .A2(n5847), .ZN(n4694) );
  INV_X1 U5282 ( .A(n8147), .ZN(n4998) );
  INV_X1 U5283 ( .A(n8795), .ZN(n8908) );
  OR2_X1 U5284 ( .A1(n5989), .A2(n5983), .ZN(n10398) );
  NAND2_X1 U5285 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5027), .ZN(n5030) );
  NAND2_X1 U5286 ( .A1(n9629), .A2(n6393), .ZN(n7031) );
  AND2_X1 U5287 ( .A1(n9549), .A2(n6392), .ZN(n4545) );
  MUX2_X1 U5288 ( .A(n9579), .B(n9539), .S(n9540), .Z(n9546) );
  NAND2_X1 U5289 ( .A1(n9579), .A2(n9576), .ZN(n9543) );
  INV_X1 U5290 ( .A(n6079), .ZN(n6355) );
  NAND2_X1 U5291 ( .A1(n8366), .A2(n8186), .ZN(n6120) );
  AND2_X1 U5292 ( .A1(n8366), .A2(n6033), .ZN(n6077) );
  NAND2_X1 U5293 ( .A1(n9798), .A2(n4860), .ZN(n4859) );
  AND2_X1 U5294 ( .A1(n6418), .A2(n6417), .ZN(n9763) );
  INV_X1 U5295 ( .A(n6353), .ZN(n6352) );
  OAI21_X1 U5296 ( .B1(n4399), .B2(n6295), .A(n4831), .ZN(n4624) );
  INV_X1 U5297 ( .A(n4832), .ZN(n4831) );
  OAI21_X1 U5298 ( .B1(n4833), .B2(n4403), .A(n4838), .ZN(n4832) );
  NOR2_X1 U5299 ( .A1(n9884), .A2(n4875), .ZN(n4874) );
  INV_X1 U5300 ( .A(n9516), .ZN(n4875) );
  NAND2_X1 U5301 ( .A1(n9907), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U5302 ( .A1(n4846), .A2(n6253), .ZN(n4844) );
  NAND2_X1 U5303 ( .A1(n9952), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U5304 ( .A1(n6235), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U5305 ( .A1(n4448), .A2(n7953), .ZN(n4852) );
  NAND2_X1 U5306 ( .A1(n7721), .A2(n4426), .ZN(n4851) );
  INV_X1 U5307 ( .A(n9583), .ZN(n4549) );
  OR2_X1 U5308 ( .A1(n7031), .A2(n10180), .ZN(n10014) );
  OR2_X1 U5309 ( .A1(n9540), .A2(n6396), .ZN(n10133) );
  NAND2_X1 U5310 ( .A1(n6438), .A2(n6437), .ZN(n7279) );
  NOR2_X1 U5311 ( .A1(n8166), .A2(n7952), .ZN(n6437) );
  NAND2_X1 U5312 ( .A1(n6011), .A2(n6013), .ZN(n4857) );
  NAND2_X1 U5313 ( .A1(n6030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5314 ( .A1(n8470), .A2(n4935), .ZN(n4934) );
  NOR2_X1 U5315 ( .A1(n8572), .A2(n4936), .ZN(n4935) );
  AOI21_X1 U5316 ( .B1(n4927), .B2(n4406), .A(n5729), .ZN(n4923) );
  NAND2_X1 U5317 ( .A1(n7492), .A2(n7493), .ZN(n7491) );
  INV_X1 U5318 ( .A(n9097), .ZN(n4819) );
  OAI22_X1 U5319 ( .A1(n9210), .A2(n4737), .B1(n4739), .B2(n9107), .ZN(n9165)
         );
  NAND2_X1 U5320 ( .A1(n4738), .A2(n4741), .ZN(n4737) );
  INV_X1 U5321 ( .A(n9211), .ZN(n4738) );
  NAND2_X1 U5322 ( .A1(n9165), .A2(n9164), .ZN(n9175) );
  OAI21_X1 U5323 ( .B1(n10065), .B2(n10021), .A(n4509), .ZN(n4508) );
  NAND2_X1 U5324 ( .A1(n4414), .A2(n4798), .ZN(n4797) );
  INV_X1 U5325 ( .A(n5893), .ZN(n4801) );
  NAND2_X1 U5326 ( .A1(n4483), .A2(n4425), .ZN(n4791) );
  NAND2_X1 U5327 ( .A1(n5879), .A2(n5878), .ZN(n4483) );
  OR2_X1 U5328 ( .A1(n9436), .A2(n9530), .ZN(n4553) );
  AOI21_X1 U5329 ( .B1(n7778), .B2(n9439), .A(n4412), .ZN(n9436) );
  NAND2_X1 U5330 ( .A1(n5936), .A2(n4400), .ZN(n4825) );
  OAI21_X1 U5331 ( .B1(n5918), .B2(n5923), .A(n5922), .ZN(n5920) );
  NOR2_X1 U5332 ( .A1(n4807), .A2(n4806), .ZN(n4805) );
  OR2_X1 U5333 ( .A1(n5939), .A2(n4822), .ZN(n4821) );
  AND2_X1 U5334 ( .A1(n5940), .A2(n5976), .ZN(n4822) );
  NAND2_X1 U5335 ( .A1(n9494), .A2(n9493), .ZN(n4713) );
  OAI21_X1 U5336 ( .B1(n4713), .B2(n10119), .A(n4712), .ZN(n4711) );
  NOR2_X1 U5337 ( .A1(n9495), .A2(n9530), .ZN(n4712) );
  NAND2_X1 U5338 ( .A1(n9823), .A2(n9417), .ZN(n9425) );
  AND2_X1 U5339 ( .A1(n8695), .A2(n5829), .ZN(n5950) );
  AND2_X1 U5340 ( .A1(n5771), .A2(n8597), .ZN(n5927) );
  NAND2_X1 U5341 ( .A1(n8607), .A2(n7570), .ZN(n5871) );
  AOI21_X1 U5342 ( .B1(n4781), .B2(n4779), .A(n4778), .ZN(n4777) );
  INV_X1 U5343 ( .A(n5654), .ZN(n4778) );
  INV_X1 U5344 ( .A(n4783), .ZN(n4779) );
  INV_X1 U5345 ( .A(n4781), .ZN(n4780) );
  INV_X1 U5346 ( .A(n4768), .ZN(n4767) );
  OAI21_X1 U5347 ( .B1(n4770), .B2(n4769), .A(n5480), .ZN(n4768) );
  INV_X1 U5348 ( .A(n5479), .ZN(n5480) );
  INV_X1 U5349 ( .A(n5453), .ZN(n4769) );
  INV_X1 U5350 ( .A(n5342), .ZN(n5341) );
  NOR4_X1 U5351 ( .A1(n8706), .A2(n5842), .A3(n8740), .A4(n8730), .ZN(n5843)
         );
  INV_X1 U5352 ( .A(n7478), .ZN(n4703) );
  NOR2_X1 U5353 ( .A1(n7456), .A2(n4705), .ZN(n4704) );
  INV_X1 U5354 ( .A(n7452), .ZN(n4705) );
  INV_X1 U5355 ( .A(n4374), .ZN(n4531) );
  NAND2_X1 U5356 ( .A1(n5420), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U5357 ( .A1(n5000), .A2(n8181), .ZN(n4995) );
  NAND2_X1 U5358 ( .A1(n5988), .A2(n7609), .ZN(n5720) );
  INV_X1 U5359 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4606) );
  NOR2_X2 U5360 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4617) );
  INV_X1 U5361 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5094) );
  OR2_X1 U5362 ( .A1(n10108), .A2(n9925), .ZN(n6295) );
  NAND2_X1 U5363 ( .A1(n4525), .A2(n4524), .ZN(n9898) );
  INV_X1 U5364 ( .A(n9915), .ZN(n4524) );
  NOR2_X1 U5365 ( .A1(n10113), .A2(n10119), .ZN(n4919) );
  INV_X1 U5366 ( .A(n9450), .ZN(n4869) );
  NAND2_X1 U5367 ( .A1(n6020), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6162) );
  INV_X1 U5368 ( .A(n6149), .ZN(n6020) );
  NAND2_X1 U5369 ( .A1(n7778), .A2(n9373), .ZN(n4881) );
  AND2_X1 U5370 ( .A1(n6421), .A2(n10286), .ZN(n4914) );
  NAND2_X1 U5371 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  NAND2_X1 U5372 ( .A1(n7614), .A2(n7820), .ZN(n7617) );
  OR2_X1 U5373 ( .A1(n6085), .A2(n6070), .ZN(n6071) );
  NAND2_X1 U5374 ( .A1(n4751), .A2(n4753), .ZN(n4749) );
  AND2_X1 U5375 ( .A1(n6005), .A2(n6004), .ZN(n6010) );
  AOI21_X1 U5376 ( .B1(n4785), .B2(n4783), .A(n4782), .ZN(n4781) );
  INV_X1 U5377 ( .A(n5634), .ZN(n4782) );
  NAND2_X1 U5378 ( .A1(n5634), .A2(n5621), .ZN(n5635) );
  INV_X1 U5379 ( .A(n5614), .ZN(n4785) );
  INV_X1 U5380 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U5381 ( .A1(n6384), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U5382 ( .A1(n4745), .A2(n4744), .ZN(n6384) );
  AOI21_X1 U5383 ( .B1(n4404), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4744) );
  XNOR2_X1 U5384 ( .A(n5549), .B(SI_21_), .ZN(n5548) );
  AND2_X1 U5385 ( .A1(n5534), .A2(n5515), .ZN(n5532) );
  NOR2_X1 U5386 ( .A1(n5454), .A2(n4667), .ZN(n4770) );
  NAND2_X1 U5387 ( .A1(n4666), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5388 ( .A1(n4669), .A2(n5454), .ZN(n4663) );
  AND2_X1 U5389 ( .A1(n5449), .A2(n5406), .ZN(n5011) );
  NAND2_X1 U5390 ( .A1(n5401), .A2(n5400), .ZN(n5433) );
  NAND2_X1 U5391 ( .A1(n5330), .A2(n5329), .ZN(n5355) );
  AND2_X1 U5392 ( .A1(n5376), .A2(n5360), .ZN(n5009) );
  NOR2_X1 U5393 ( .A1(n5327), .A2(n4657), .ZN(n4656) );
  INV_X1 U5394 ( .A(n5299), .ZN(n4657) );
  NOR2_X1 U5395 ( .A1(n4529), .A2(n4527), .ZN(n4526) );
  INV_X1 U5396 ( .A(n5392), .ZN(n4952) );
  OR2_X1 U5397 ( .A1(n5388), .A2(n4952), .ZN(n4951) );
  INV_X1 U5398 ( .A(n5447), .ZN(n4950) );
  NAND2_X1 U5399 ( .A1(n7863), .A2(n7862), .ZN(n7861) );
  NAND2_X1 U5400 ( .A1(n5341), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5365) );
  AOI21_X1 U5401 ( .B1(n4593), .B2(n4953), .A(n4445), .ZN(n4592) );
  INV_X1 U5402 ( .A(n7862), .ZN(n4593) );
  INV_X1 U5403 ( .A(n4953), .ZN(n4594) );
  OR2_X1 U5404 ( .A1(n5472), .A2(n5471), .ZN(n5474) );
  NAND2_X1 U5405 ( .A1(n5459), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5490) );
  AOI21_X1 U5406 ( .B1(n4681), .B2(n4683), .A(n4684), .ZN(n4679) );
  AND4_X1 U5407 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n8335)
         );
  NAND2_X1 U5408 ( .A1(n7190), .A2(n7189), .ZN(n7120) );
  NAND2_X1 U5409 ( .A1(n7142), .A2(n7141), .ZN(n7239) );
  OR2_X1 U5410 ( .A1(n7259), .A2(n7258), .ZN(n7412) );
  INV_X1 U5411 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n4699) );
  AOI21_X1 U5412 ( .B1(n8621), .B2(n8613), .A(n8612), .ZN(n10358) );
  NAND2_X1 U5413 ( .A1(n8718), .A2(n4964), .ZN(n8651) );
  NOR2_X1 U5414 ( .A1(n8662), .A2(n4965), .ZN(n4964) );
  INV_X1 U5415 ( .A(n4966), .ZN(n4965) );
  AOI21_X1 U5416 ( .B1(n8686), .B2(n4655), .A(n4438), .ZN(n4654) );
  INV_X1 U5417 ( .A(n8353), .ZN(n4655) );
  AND2_X1 U5418 ( .A1(n5682), .A2(n5681), .ZN(n8699) );
  OR2_X1 U5419 ( .A1(n5741), .A2(n5733), .ZN(n5682) );
  NAND2_X1 U5420 ( .A1(n8718), .A2(n8692), .ZN(n8689) );
  NAND2_X1 U5421 ( .A1(n5644), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5673) );
  AOI21_X1 U5422 ( .B1(n4986), .B2(n8771), .A(n4437), .ZN(n4984) );
  OR2_X1 U5423 ( .A1(n8992), .A2(n8758), .ZN(n8350) );
  AND2_X1 U5424 ( .A1(n8766), .A2(n8350), .ZN(n4986) );
  NAND2_X1 U5425 ( .A1(n4905), .A2(n5933), .ZN(n4904) );
  NAND2_X1 U5426 ( .A1(n4906), .A2(n5933), .ZN(n4903) );
  NAND2_X1 U5427 ( .A1(n8771), .A2(n5931), .ZN(n4906) );
  NOR2_X1 U5428 ( .A1(n8788), .A2(n5773), .ZN(n8772) );
  AOI21_X1 U5429 ( .B1(n5772), .B2(n8348), .A(n4407), .ZN(n4975) );
  AOI21_X1 U5430 ( .B1(n4992), .B2(n4435), .A(n4440), .ZN(n4990) );
  INV_X1 U5431 ( .A(n4992), .ZN(n4991) );
  AND2_X1 U5432 ( .A1(n8870), .A2(n8341), .ZN(n4992) );
  NAND2_X1 U5433 ( .A1(n8340), .A2(n8339), .ZN(n8886) );
  NAND2_X1 U5434 ( .A1(n4902), .A2(n5760), .ZN(n4900) );
  NAND2_X1 U5435 ( .A1(n4675), .A2(n4674), .ZN(n4899) );
  AND2_X1 U5436 ( .A1(n4456), .A2(n5896), .ZN(n4674) );
  NAND2_X1 U5437 ( .A1(n5001), .A2(n5000), .ZN(n4999) );
  INV_X1 U5438 ( .A(n8149), .ZN(n5001) );
  NAND2_X1 U5439 ( .A1(n7527), .A2(n4978), .ZN(n4981) );
  NOR2_X1 U5440 ( .A1(n7576), .A2(n4982), .ZN(n4978) );
  OR2_X1 U5441 ( .A1(n6992), .A2(n5739), .ZN(n8795) );
  NOR2_X1 U5442 ( .A1(n9102), .A2(n5707), .ZN(n10364) );
  AND2_X1 U5443 ( .A1(n8168), .A2(n5706), .ZN(n5707) );
  AND3_X2 U5444 ( .A1(n5026), .A2(n5025), .A3(n4423), .ZN(n5029) );
  INV_X1 U5445 ( .A(n5045), .ZN(n5046) );
  OR2_X1 U5446 ( .A1(n5092), .A2(n9088), .ZN(n5139) );
  INV_X1 U5447 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5448 ( .B1(n7692), .B2(n7691), .A(n7377), .ZN(n4730) );
  AND2_X1 U5449 ( .A1(n9192), .A2(n4724), .ZN(n4723) );
  NAND2_X1 U5450 ( .A1(n9269), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5451 ( .A1(n7733), .A2(n7614), .ZN(n7027) );
  NAND2_X1 U5452 ( .A1(n8268), .A2(n8267), .ZN(n9266) );
  NAND2_X1 U5453 ( .A1(n9266), .A2(n9267), .ZN(n9265) );
  INV_X1 U5454 ( .A(n8187), .ZN(n4584) );
  INV_X1 U5455 ( .A(n4586), .ZN(n4585) );
  INV_X1 U5456 ( .A(n9199), .ZN(n4581) );
  OR2_X1 U5457 ( .A1(n7285), .A2(n7034), .ZN(n7037) );
  NAND2_X1 U5458 ( .A1(n7071), .A2(n4873), .ZN(n7072) );
  NAND2_X1 U5459 ( .A1(n7070), .A2(n7069), .ZN(n7163) );
  OAI21_X1 U5460 ( .B1(n7022), .B2(n7161), .A(n4746), .ZN(n7162) );
  INV_X1 U5461 ( .A(n9925), .ZN(n9508) );
  INV_X1 U5462 ( .A(n6120), .ZN(n4547) );
  AND2_X1 U5463 ( .A1(n9681), .A2(n6859), .ZN(n6948) );
  AOI21_X1 U5464 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n10233) );
  OR2_X1 U5465 ( .A1(n6907), .A2(n6908), .ZN(n6969) );
  AOI21_X1 U5466 ( .B1(n9798), .B2(n9603), .A(n4862), .ZN(n4487) );
  NAND2_X1 U5467 ( .A1(n4638), .A2(n4637), .ZN(n9788) );
  AND2_X1 U5468 ( .A1(n6349), .A2(n6348), .ZN(n9799) );
  OR2_X1 U5469 ( .A1(n9212), .A2(n6355), .ZN(n6349) );
  OR2_X1 U5470 ( .A1(n10089), .A2(n9867), .ZN(n9347) );
  NAND2_X1 U5471 ( .A1(n4522), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6342) );
  INV_X1 U5472 ( .A(n4836), .ZN(n4830) );
  INV_X1 U5473 ( .A(n9899), .ZN(n4834) );
  NOR2_X1 U5474 ( .A1(n4837), .A2(n6308), .ZN(n4836) );
  INV_X1 U5475 ( .A(n5006), .ZN(n4837) );
  OR2_X1 U5476 ( .A1(n9909), .A2(n9508), .ZN(n5006) );
  AND2_X1 U5477 ( .A1(n6307), .A2(n6306), .ZN(n9917) );
  INV_X1 U5478 ( .A(n10108), .ZN(n9909) );
  OR2_X1 U5479 ( .A1(n9929), .A2(n9918), .ZN(n5005) );
  INV_X1 U5480 ( .A(n6252), .ZN(n4847) );
  AND2_X1 U5481 ( .A1(n9922), .A2(n9921), .ZN(n9943) );
  NAND2_X1 U5482 ( .A1(n4496), .A2(n9450), .ZN(n4866) );
  NOR2_X1 U5483 ( .A1(n10128), .A2(n4909), .ZN(n4907) );
  CLKBUF_X1 U5484 ( .A(n9994), .Z(n4496) );
  AOI21_X1 U5485 ( .B1(n6218), .B2(n4645), .A(n4430), .ZN(n4644) );
  INV_X1 U5486 ( .A(n6206), .ZN(n4645) );
  INV_X1 U5487 ( .A(n6218), .ZN(n4646) );
  NOR2_X1 U5488 ( .A1(n9595), .A2(n4850), .ZN(n4849) );
  INV_X1 U5489 ( .A(n4852), .ZN(n4850) );
  AND4_X1 U5490 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n10013)
         );
  NOR2_X1 U5491 ( .A1(n4402), .A2(n4626), .ZN(n4625) );
  NAND2_X1 U5492 ( .A1(n6155), .A2(n5012), .ZN(n4626) );
  INV_X1 U5493 ( .A(n6141), .ZN(n6128) );
  NAND3_X1 U5494 ( .A1(n4715), .A2(n9581), .A3(n4714), .ZN(n8010) );
  INV_X1 U5495 ( .A(n10016), .ZN(n9938) );
  INV_X1 U5496 ( .A(n10012), .ZN(n9981) );
  INV_X1 U5497 ( .A(n7023), .ZN(n9623) );
  OR2_X1 U5498 ( .A1(n6760), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U5499 ( .A1(n9404), .A2(n9403), .ZN(n9407) );
  NAND2_X1 U5500 ( .A1(n9098), .A2(n6350), .ZN(n4473) );
  AND2_X1 U5501 ( .A1(n6395), .A2(n6394), .ZN(n10311) );
  OR2_X1 U5502 ( .A1(n7818), .A2(n6396), .ZN(n10320) );
  INV_X1 U5503 ( .A(n6015), .ZN(n6012) );
  INV_X1 U5504 ( .A(n4857), .ZN(n4855) );
  NAND2_X1 U5505 ( .A1(n4420), .A2(n6426), .ZN(n6440) );
  NAND2_X1 U5506 ( .A1(n6386), .A2(n6385), .ZN(n6389) );
  NOR2_X1 U5507 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10474), .ZN(n10207) );
  OAI21_X1 U5508 ( .B1(n10487), .B2(n10490), .A(n10211), .ZN(n10212) );
  AND4_X1 U5509 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n8458)
         );
  OR2_X1 U5510 ( .A1(n5500), .A2(n8423), .ZN(n5478) );
  NAND2_X1 U5511 ( .A1(n4934), .A2(n4925), .ZN(n4924) );
  NOR2_X1 U5512 ( .A1(n4928), .A2(n4938), .ZN(n4925) );
  NAND2_X1 U5513 ( .A1(n4937), .A2(n8382), .ZN(n4926) );
  AND2_X1 U5514 ( .A1(n5747), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8464) );
  INV_X1 U5515 ( .A(n8471), .ZN(n4611) );
  AND2_X1 U5516 ( .A1(n4387), .A2(n8590), .ZN(n4609) );
  AND4_X1 U5517 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n8481)
         );
  OR2_X1 U5518 ( .A1(n8573), .A2(n8793), .ZN(n8565) );
  AND2_X1 U5519 ( .A1(n7269), .A2(n7268), .ZN(n8564) );
  NAND2_X1 U5520 ( .A1(n7390), .A2(n5165), .ZN(n4596) );
  NOR2_X2 U5521 ( .A1(n5728), .A2(n5727), .ZN(n8583) );
  INV_X1 U5522 ( .A(n5740), .ZN(n5728) );
  INV_X1 U5523 ( .A(n8583), .ZN(n8579) );
  INV_X1 U5524 ( .A(n8570), .ZN(n8590) );
  AOI21_X1 U5525 ( .B1(n8639), .B2(n10355), .A(n10354), .ZN(n4709) );
  OAI21_X1 U5526 ( .B1(n8643), .B2(n8644), .A(n8642), .ZN(n4707) );
  NAND2_X1 U5527 ( .A1(n4898), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U5528 ( .A1(n8693), .A2(n8680), .ZN(n4897) );
  NOR2_X1 U5529 ( .A1(n8679), .A2(n8868), .ZN(n4898) );
  NAND2_X1 U5530 ( .A1(n8684), .A2(n8686), .ZN(n8685) );
  NAND2_X1 U5531 ( .A1(n8705), .A2(n8353), .ZN(n8684) );
  NOR2_X1 U5532 ( .A1(n8713), .A2(n8712), .ZN(n8715) );
  AND2_X1 U5533 ( .A1(n5645), .A2(n5627), .ZN(n8734) );
  INV_X1 U5534 ( .A(n8932), .ZN(n8944) );
  NAND2_X2 U5535 ( .A1(n7325), .A2(n8877), .ZN(n8945) );
  INV_X1 U5536 ( .A(n8361), .ZN(n4535) );
  INV_X1 U5537 ( .A(n8666), .ZN(n4534) );
  NAND2_X1 U5538 ( .A1(n4575), .A2(n4578), .ZN(n9124) );
  NAND2_X1 U5539 ( .A1(n9279), .A2(n9276), .ZN(n4578) );
  NAND2_X1 U5540 ( .A1(n4579), .A2(n9277), .ZN(n4575) );
  INV_X1 U5541 ( .A(n8069), .ZN(n4732) );
  AND2_X1 U5542 ( .A1(n9170), .A2(n4491), .ZN(n4490) );
  AND2_X1 U5543 ( .A1(n9169), .A2(n9311), .ZN(n4491) );
  AND2_X1 U5544 ( .A1(n6319), .A2(n6318), .ZN(n9886) );
  OR2_X1 U5545 ( .A1(n9795), .A2(n6355), .ZN(n6360) );
  AOI22_X2 U5546 ( .A1(n9257), .A2(n9256), .B1(n8305), .B2(n8304), .ZN(n9210)
         );
  AND2_X1 U5547 ( .A1(n6263), .A2(n6262), .ZN(n9962) );
  OR2_X1 U5548 ( .A1(n7035), .A2(n9662), .ZN(n9320) );
  NAND2_X1 U5549 ( .A1(n7289), .A2(n7288), .ZN(n9305) );
  NOR2_X1 U5550 ( .A1(n8315), .A2(n4740), .ZN(n4739) );
  INV_X1 U5551 ( .A(n4742), .ZN(n4740) );
  NAND2_X1 U5552 ( .A1(n10072), .A2(n9338), .ZN(n8321) );
  AND2_X1 U5553 ( .A1(n8094), .A2(n10299), .ZN(n9338) );
  INV_X1 U5554 ( .A(n9311), .ZN(n9340) );
  OAI211_X1 U5555 ( .C1(n4546), .C2(n9622), .A(n4544), .B(n9621), .ZN(n4543)
         );
  NAND2_X1 U5556 ( .A1(n4546), .A2(n4429), .ZN(n4544) );
  INV_X1 U5557 ( .A(n6392), .ZN(n9629) );
  OR2_X1 U5558 ( .A1(n6229), .A2(n6228), .ZN(n9637) );
  OR2_X1 U5559 ( .A1(n6120), .A2(n6119), .ZN(n6121) );
  OAI21_X1 U5560 ( .B1(n10244), .B2(n9744), .A(n9743), .ZN(n4502) );
  NAND2_X1 U5561 ( .A1(n4859), .A2(n4858), .ZN(n6419) );
  AOI21_X1 U5562 ( .B1(n4860), .B2(n4862), .A(n6416), .ZN(n4858) );
  INV_X1 U5563 ( .A(n9990), .ZN(n10034) );
  OR2_X1 U5564 ( .A1(n10133), .A2(n7036), .ZN(n9999) );
  NOR2_X1 U5565 ( .A1(n4857), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4856) );
  NOR2_X1 U5566 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  NOR2_X1 U5567 ( .A1(n4804), .A2(n4803), .ZN(n4802) );
  INV_X1 U5568 ( .A(n8125), .ZN(n4803) );
  INV_X1 U5569 ( .A(n4802), .ZN(n4798) );
  NAND2_X1 U5570 ( .A1(n4435), .A2(n4811), .ZN(n4810) );
  INV_X1 U5571 ( .A(n5911), .ZN(n4811) );
  INV_X1 U5572 ( .A(n5908), .ZN(n4484) );
  NAND2_X1 U5573 ( .A1(n9440), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5574 ( .A1(n4826), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U5575 ( .A1(n4711), .A2(n4556), .ZN(n4555) );
  INV_X1 U5576 ( .A(n4713), .ZN(n9496) );
  NOR4_X1 U5577 ( .A1(n5831), .A2(n7350), .A3(n7321), .A4(n5833), .ZN(n5834)
         );
  AOI21_X1 U5578 ( .B1(n5964), .B2(n8699), .A(n8657), .ZN(n5967) );
  INV_X1 U5579 ( .A(n7806), .ZN(n4888) );
  INV_X1 U5580 ( .A(n5880), .ZN(n4889) );
  INV_X1 U5581 ( .A(n4890), .ZN(n4517) );
  OR2_X1 U5582 ( .A1(n5223), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5337) );
  NOR2_X1 U5583 ( .A1(n4573), .A2(n4441), .ZN(n4570) );
  INV_X1 U5584 ( .A(n8250), .ZN(n4577) );
  NAND2_X1 U5585 ( .A1(n10050), .A2(n9576), .ZN(n4772) );
  NOR2_X1 U5586 ( .A1(n10050), .A2(n10053), .ZN(n4721) );
  NAND2_X1 U5587 ( .A1(n4720), .A2(n9542), .ZN(n4719) );
  NAND2_X1 U5588 ( .A1(n10050), .A2(n9530), .ZN(n4720) );
  AND2_X1 U5589 ( .A1(n4559), .A2(n9536), .ZN(n4518) );
  NAND2_X1 U5590 ( .A1(n5619), .A2(n6646), .ZN(n5634) );
  NOR2_X1 U5591 ( .A1(n4763), .A2(n4762), .ZN(n4761) );
  INV_X1 U5592 ( .A(n5534), .ZN(n4762) );
  INV_X1 U5593 ( .A(n5548), .ZN(n4763) );
  NAND2_X1 U5594 ( .A1(n5484), .A2(n5483), .ZN(n5510) );
  INV_X1 U5595 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5280) );
  INV_X1 U5596 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5597 ( .A1(n4397), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4505) );
  INV_X1 U5598 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U5599 ( .A1(n4397), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5600 ( .A1(n4396), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4515) );
  NOR2_X1 U5601 ( .A1(n7588), .A2(n4956), .ZN(n4955) );
  INV_X1 U5602 ( .A(n5193), .ZN(n4956) );
  NOR2_X1 U5603 ( .A1(n8522), .A2(n8454), .ZN(n4540) );
  INV_X1 U5604 ( .A(n5182), .ZN(n4528) );
  AND2_X1 U5605 ( .A1(n5341), .A2(n4539), .ZN(n5420) );
  AND2_X1 U5606 ( .A1(n4411), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5607 ( .A1(n4686), .A2(n4685), .ZN(n4684) );
  NAND2_X1 U5608 ( .A1(n5823), .A2(n4689), .ZN(n4685) );
  INV_X1 U5609 ( .A(n5975), .ZN(n4686) );
  INV_X1 U5610 ( .A(n4688), .ZN(n4683) );
  INV_X1 U5611 ( .A(n5778), .ZN(n5779) );
  NOR2_X1 U5612 ( .A1(n8959), .A2(n8964), .ZN(n4966) );
  INV_X1 U5613 ( .A(n4654), .ZN(n4652) );
  AND2_X1 U5614 ( .A1(n5624), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U5615 ( .A1(n8987), .A2(n8992), .ZN(n4963) );
  NOR2_X1 U5616 ( .A1(n8432), .A2(n4537), .ZN(n4536) );
  NOR2_X1 U5617 ( .A1(n8851), .A2(n8837), .ZN(n8815) );
  NAND2_X1 U5618 ( .A1(n8357), .A2(n4971), .ZN(n4970) );
  AND2_X1 U5619 ( .A1(n5990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4961) );
  NOR2_X1 U5620 ( .A1(n9024), .A2(n9030), .ZN(n4971) );
  NAND2_X1 U5621 ( .A1(n7804), .A2(n5758), .ZN(n8128) );
  OAI211_X1 U5622 ( .C1(n7578), .C2(n4673), .A(n4672), .B(n7921), .ZN(n7804)
         );
  INV_X1 U5623 ( .A(n4887), .ZN(n4673) );
  NAND2_X1 U5624 ( .A1(n4887), .A2(n4517), .ZN(n4672) );
  AOI21_X1 U5625 ( .B1(n4890), .B2(n4889), .A(n4888), .ZN(n4887) );
  INV_X1 U5626 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5227) );
  OR2_X1 U5627 ( .A1(n5228), .A2(n5227), .ZN(n5259) );
  NAND2_X1 U5628 ( .A1(n4892), .A2(n5880), .ZN(n4891) );
  NAND2_X1 U5629 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5147) );
  NAND2_X1 U5630 ( .A1(n7352), .A2(n5753), .ZN(n5852) );
  NAND2_X1 U5631 ( .A1(n5754), .A2(n10391), .ZN(n5853) );
  NAND2_X1 U5632 ( .A1(n5752), .A2(n8938), .ZN(n6810) );
  NOR2_X1 U5633 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5092) );
  INV_X1 U5634 ( .A(n9267), .ZN(n4725) );
  NAND2_X1 U5635 ( .A1(n8051), .A2(n8050), .ZN(n8088) );
  NAND2_X1 U5636 ( .A1(n9609), .A2(n10043), .ZN(n9579) );
  INV_X1 U5637 ( .A(n6362), .ZN(n4854) );
  NOR2_X1 U5638 ( .A1(n6312), .A2(n6311), .ZN(n4522) );
  NAND2_X1 U5639 ( .A1(n9876), .A2(n9866), .ZN(n4838) );
  NOR2_X1 U5640 ( .A1(n6273), .A2(n6024), .ZN(n4521) );
  AND2_X1 U5641 ( .A1(n6023), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6235) );
  NOR2_X1 U5642 ( .A1(n4642), .A2(n6230), .ZN(n4641) );
  INV_X1 U5643 ( .A(n4644), .ZN(n4642) );
  NOR2_X1 U5644 ( .A1(n6211), .A2(n9280), .ZN(n4520) );
  NOR2_X1 U5645 ( .A1(n10141), .A2(n8206), .ZN(n4911) );
  NAND2_X1 U5646 ( .A1(n4519), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6172) );
  INV_X1 U5647 ( .A(n6162), .ZN(n4519) );
  AND3_X1 U5648 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5649 ( .A1(n6139), .A2(n7853), .ZN(n9557) );
  NAND2_X1 U5650 ( .A1(n9645), .A2(n6421), .ZN(n9374) );
  INV_X1 U5651 ( .A(n4412), .ZN(n4716) );
  NAND2_X1 U5652 ( .A1(n4547), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6081) );
  INV_X1 U5653 ( .A(SI_13_), .ZN(n6667) );
  AOI21_X1 U5654 ( .B1(n4777), .B2(n4780), .A(n4774), .ZN(n4773) );
  NAND2_X1 U5655 ( .A1(n5618), .A2(n4777), .ZN(n4775) );
  INV_X1 U5656 ( .A(n5656), .ZN(n4774) );
  AND2_X1 U5657 ( .A1(n5687), .A2(n5660), .ZN(n5685) );
  AND2_X1 U5658 ( .A1(n5585), .A2(n5580), .ZN(n5583) );
  NAND2_X1 U5659 ( .A1(n5572), .A2(n5555), .ZN(n5573) );
  AOI21_X1 U5660 ( .B1(n4767), .B2(n4769), .A(n4443), .ZN(n4765) );
  XNOR2_X1 U5661 ( .A(n5324), .B(SI_11_), .ZN(n5323) );
  NOR2_X2 U5662 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6052) );
  NAND2_X1 U5663 ( .A1(n8518), .A2(n5388), .ZN(n8393) );
  AOI21_X1 U5664 ( .B1(n5569), .B2(n4941), .A(n4409), .ZN(n4940) );
  INV_X1 U5665 ( .A(n5569), .ZN(n4942) );
  XNOR2_X1 U5666 ( .A(n5643), .B(n8938), .ZN(n5071) );
  AOI21_X1 U5667 ( .B1(n4592), .B2(n4594), .A(n4591), .ZN(n4590) );
  INV_X1 U5668 ( .A(n8545), .ZN(n4591) );
  NAND2_X1 U5669 ( .A1(n8393), .A2(n5392), .ZN(n8474) );
  NAND2_X1 U5670 ( .A1(n4604), .A2(n4603), .ZN(n7512) );
  INV_X1 U5671 ( .A(n5144), .ZN(n4604) );
  INV_X1 U5672 ( .A(n7044), .ZN(n6811) );
  NAND2_X1 U5673 ( .A1(n5459), .A2(n4536), .ZN(n5518) );
  NAND2_X1 U5674 ( .A1(n5341), .A2(n4540), .ZN(n5381) );
  OR2_X1 U5675 ( .A1(n5311), .A2(n5310), .ZN(n5342) );
  NAND2_X1 U5676 ( .A1(n5258), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5311) );
  INV_X1 U5677 ( .A(n5259), .ZN(n5258) );
  NAND2_X1 U5678 ( .A1(n5145), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5182) );
  INV_X1 U5679 ( .A(n5147), .ZN(n5145) );
  NAND2_X1 U5680 ( .A1(n4528), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U5681 ( .A1(n5341), .A2(n4411), .ZN(n5426) );
  AND2_X1 U5682 ( .A1(n5983), .A2(n6816), .ZN(n4816) );
  XNOR2_X1 U5683 ( .A(n4493), .B(n8640), .ZN(n5845) );
  INV_X1 U5684 ( .A(n5974), .ZN(n4494) );
  NOR2_X1 U5685 ( .A1(n5975), .A2(n8657), .ZN(n4495) );
  AND3_X1 U5686 ( .A1(n5463), .A2(n5462), .A3(n5461), .ZN(n8488) );
  AND3_X1 U5687 ( .A1(n5424), .A2(n5423), .A3(n5422), .ZN(n8487) );
  AND4_X1 U5688 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n8153)
         );
  NAND2_X1 U5689 ( .A1(n7123), .A2(n7122), .ZN(n7237) );
  NAND2_X1 U5690 ( .A1(n7144), .A2(n7143), .ZN(n7206) );
  AOI21_X1 U5691 ( .B1(n4704), .B2(n7414), .A(n4703), .ZN(n4702) );
  NAND2_X1 U5692 ( .A1(n7453), .A2(n4704), .ZN(n7480) );
  OAI21_X1 U5693 ( .B1(n7657), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7654), .ZN(
        n7704) );
  OR2_X1 U5694 ( .A1(n10352), .A2(n8614), .ZN(n4472) );
  NAND2_X1 U5695 ( .A1(n10348), .A2(n4696), .ZN(n8628) );
  OR2_X1 U5696 ( .A1(n10352), .A2(n8622), .ZN(n4696) );
  NAND2_X1 U5697 ( .A1(n8615), .A2(n4413), .ZN(n8633) );
  NOR2_X1 U5698 ( .A1(n8959), .A2(n8329), .ZN(n8656) );
  NAND2_X1 U5699 ( .A1(n8718), .A2(n4966), .ZN(n8671) );
  OR2_X1 U5700 ( .A1(n4375), .A2(n4532), .ZN(n8353) );
  NAND2_X1 U5701 ( .A1(n8724), .A2(n4432), .ZN(n8709) );
  NAND2_X1 U5702 ( .A1(n8796), .A2(n4418), .ZN(n8749) );
  AND2_X1 U5703 ( .A1(n8796), .A2(n4963), .ZN(n8760) );
  OR2_X1 U5704 ( .A1(n5558), .A2(n8535), .ZN(n5597) );
  AND2_X1 U5705 ( .A1(n8796), .A2(n8779), .ZN(n8777) );
  OR2_X1 U5706 ( .A1(n5538), .A2(n8444), .ZN(n5558) );
  AND2_X1 U5707 ( .A1(n5565), .A2(n5564), .ZN(n8794) );
  CLKBUF_X1 U5708 ( .A(n8808), .Z(n8809) );
  OR2_X1 U5709 ( .A1(n8809), .A2(n5772), .ZN(n8811) );
  AND2_X1 U5710 ( .A1(n5517), .A2(n5516), .ZN(n5771) );
  NOR2_X1 U5711 ( .A1(n8804), .A2(n4807), .ZN(n4693) );
  OR2_X1 U5712 ( .A1(n8916), .A2(n4967), .ZN(n8851) );
  NAND2_X1 U5713 ( .A1(n4968), .A2(n8857), .ZN(n4967) );
  INV_X1 U5714 ( .A(n4970), .ZN(n4968) );
  NOR2_X1 U5715 ( .A1(n8916), .A2(n4969), .ZN(n8893) );
  INV_X1 U5716 ( .A(n4971), .ZN(n4969) );
  NOR2_X2 U5717 ( .A1(n5014), .A2(n9046), .ZN(n8158) );
  AND2_X1 U5718 ( .A1(n4675), .A2(n5896), .ZN(n7993) );
  NAND2_X1 U5719 ( .A1(n7993), .A2(n8148), .ZN(n7992) );
  NAND2_X1 U5720 ( .A1(n8128), .A2(n5889), .ZN(n8131) );
  NOR2_X2 U5721 ( .A1(n7813), .A2(n9061), .ZN(n8137) );
  INV_X1 U5722 ( .A(n7921), .ZN(n7805) );
  NAND2_X1 U5723 ( .A1(n7839), .A2(n7592), .ZN(n4983) );
  NAND3_X1 U5724 ( .A1(n4981), .A2(n7575), .A3(n7579), .ZN(n4980) );
  NAND2_X1 U5725 ( .A1(n4980), .A2(n4977), .ZN(n7802) );
  NOR2_X1 U5726 ( .A1(n4979), .A2(n7677), .ZN(n4977) );
  INV_X1 U5727 ( .A(n4983), .ZN(n4979) );
  AND2_X1 U5728 ( .A1(n4891), .A2(n5881), .ZN(n7678) );
  NAND2_X1 U5729 ( .A1(n5819), .A2(n6732), .ZN(n4829) );
  AND2_X1 U5730 ( .A1(n5859), .A2(n5856), .ZN(n4691) );
  NAND2_X1 U5731 ( .A1(n7054), .A2(n7055), .ZN(n4692) );
  NAND2_X1 U5732 ( .A1(n7353), .A2(n7352), .ZN(n7355) );
  NAND4_X1 U5733 ( .A1(n5831), .A2(n6809), .A3(n5853), .A4(n5852), .ZN(n7348)
         );
  CLKBUF_X1 U5734 ( .A(n7046), .Z(n7350) );
  NAND2_X1 U5735 ( .A1(n8657), .A2(n8356), .ZN(n8362) );
  INV_X1 U5736 ( .A(n7570), .ZN(n10408) );
  OR2_X1 U5737 ( .A1(n5983), .A2(n5832), .ZN(n10400) );
  INV_X1 U5738 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5739 ( .A1(n4976), .A2(n5990), .ZN(n5731) );
  INV_X1 U5740 ( .A(n5042), .ZN(n4976) );
  NAND2_X1 U5741 ( .A1(n5042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U5742 ( .A1(n5692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5049) );
  OR3_X1 U5743 ( .A1(n5409), .A2(P2_IR_REG_15__SCAN_IN), .A3(n5408), .ZN(n5411) );
  INV_X1 U5744 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5745 ( .A1(n4957), .A2(n5092), .ZN(n5158) );
  AND2_X1 U5746 ( .A1(n4617), .A2(n5094), .ZN(n4957) );
  NAND2_X1 U5747 ( .A1(n7753), .A2(n7752), .ZN(n8051) );
  INV_X1 U5748 ( .A(n4735), .ZN(n4734) );
  INV_X1 U5749 ( .A(n8050), .ZN(n4736) );
  NAND2_X1 U5750 ( .A1(n6021), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6200) );
  INV_X1 U5751 ( .A(n6183), .ZN(n6021) );
  NAND2_X1 U5752 ( .A1(n6022), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6211) );
  INV_X1 U5753 ( .A(n6200), .ZN(n6022) );
  NAND2_X1 U5754 ( .A1(n4728), .A2(n7693), .ZN(n7746) );
  NAND2_X1 U5755 ( .A1(n7378), .A2(n4729), .ZN(n4728) );
  XNOR2_X1 U5756 ( .A(n7380), .B(n9157), .ZN(n7692) );
  NAND2_X1 U5757 ( .A1(n9286), .A2(n9288), .ZN(n9287) );
  NAND2_X1 U5758 ( .A1(n8289), .A2(n8290), .ZN(n9286) );
  INV_X1 U5759 ( .A(n8289), .ZN(n8292) );
  AND2_X1 U5760 ( .A1(n9626), .A2(n7282), .ZN(n7074) );
  OR2_X1 U5761 ( .A1(n8310), .A2(n8309), .ZN(n4742) );
  AND2_X1 U5762 ( .A1(n6851), .A2(n6850), .ZN(n6982) );
  INV_X1 U5763 ( .A(n6111), .ZN(n6219) );
  AND2_X1 U5764 ( .A1(n6946), .A2(n6862), .ZN(n6923) );
  OR2_X1 U5765 ( .A1(n6191), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6142) );
  OR2_X1 U5766 ( .A1(n6157), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6168) );
  OR2_X1 U5767 ( .A1(n10233), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U5768 ( .A1(n9701), .A2(n9700), .ZN(n9699) );
  AOI21_X1 U5769 ( .B1(n9699), .B2(n6884), .A(n6883), .ZN(n6913) );
  OAI21_X1 U5770 ( .B1(n6913), .B2(n6912), .A(n6911), .ZN(n6962) );
  INV_X1 U5771 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9280) );
  OAI21_X1 U5772 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n7641), .A(n7637), .ZN(
        n7762) );
  INV_X1 U5773 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U5774 ( .A1(n4637), .A2(n4401), .ZN(n4635) );
  NAND2_X1 U5775 ( .A1(n4634), .A2(n4401), .ZN(n4633) );
  NAND2_X1 U5776 ( .A1(n4636), .A2(n4853), .ZN(n4634) );
  NOR2_X1 U5777 ( .A1(n9780), .A2(n4854), .ZN(n4853) );
  NAND2_X1 U5778 ( .A1(n4637), .A2(n9806), .ZN(n4636) );
  NAND2_X1 U5779 ( .A1(n9797), .A2(n9527), .ZN(n4861) );
  OR3_X1 U5780 ( .A1(n6342), .A2(n9259), .A3(n6341), .ZN(n6353) );
  INV_X1 U5781 ( .A(n4884), .ZN(n4883) );
  NAND2_X1 U5782 ( .A1(n9850), .A2(n9849), .ZN(n4886) );
  NAND2_X1 U5783 ( .A1(n4886), .A2(n4884), .ZN(n9822) );
  INV_X1 U5784 ( .A(n4522), .ZN(n6322) );
  INV_X1 U5785 ( .A(n9633), .ZN(n9852) );
  NOR2_X2 U5786 ( .A1(n9856), .A2(n10089), .ZN(n9844) );
  OR2_X1 U5787 ( .A1(n6302), .A2(n9194), .ZN(n6312) );
  NAND2_X1 U5788 ( .A1(n6025), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6302) );
  INV_X1 U5789 ( .A(n6300), .ZN(n6025) );
  NAND2_X1 U5790 ( .A1(n4521), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U5791 ( .A1(n9909), .A2(n4919), .ZN(n4918) );
  INV_X1 U5792 ( .A(n4521), .ZN(n6288) );
  NOR2_X1 U5793 ( .A1(n9964), .A2(n4917), .ZN(n9928) );
  INV_X1 U5794 ( .A(n4919), .ZN(n4917) );
  INV_X1 U5795 ( .A(n4871), .ZN(n4870) );
  OR2_X1 U5796 ( .A1(n9952), .A2(n9975), .ZN(n9977) );
  OAI21_X1 U5797 ( .B1(n4496), .B2(n9993), .A(n9450), .ZN(n9973) );
  NAND2_X1 U5798 ( .A1(n4520), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6247) );
  INV_X1 U5799 ( .A(n4520), .ZN(n6225) );
  NAND2_X1 U5800 ( .A1(n7958), .A2(n4911), .ZN(n5008) );
  NAND2_X1 U5801 ( .A1(n7958), .A2(n10146), .ZN(n10018) );
  INV_X1 U5802 ( .A(n8029), .ZN(n4480) );
  NAND2_X1 U5803 ( .A1(n7721), .A2(n9471), .ZN(n7956) );
  AND4_X1 U5804 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n8073)
         );
  NAND2_X1 U5805 ( .A1(n6103), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U5806 ( .A1(n6019), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6149) );
  INV_X1 U5807 ( .A(n6133), .ZN(n6019) );
  INV_X1 U5808 ( .A(n10298), .ZN(n4915) );
  NAND2_X1 U5809 ( .A1(n4881), .A2(n6409), .ZN(n7890) );
  INV_X1 U5810 ( .A(n4880), .ZN(n4879) );
  NAND2_X1 U5811 ( .A1(n4914), .A2(n8013), .ZN(n7899) );
  NAND2_X1 U5812 ( .A1(n8013), .A2(n10286), .ZN(n7830) );
  NAND2_X1 U5813 ( .A1(n4717), .A2(n4716), .ZN(n9437) );
  INV_X1 U5814 ( .A(n7778), .ZN(n4717) );
  NAND2_X1 U5815 ( .A1(n7084), .A2(n9369), .ZN(n9554) );
  NAND2_X1 U5816 ( .A1(n7612), .A2(n6407), .ZN(n9368) );
  NAND2_X1 U5817 ( .A1(n9368), .A2(n6074), .ZN(n7084) );
  NAND2_X1 U5818 ( .A1(n4547), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U5819 ( .A1(n4547), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6050) );
  OR2_X1 U5820 ( .A1(n7626), .A2(n7625), .ZN(n7633) );
  INV_X1 U5821 ( .A(n7786), .ZN(n10286) );
  INV_X1 U5822 ( .A(n10320), .ZN(n10307) );
  INV_X1 U5823 ( .A(n4482), .ZN(n4481) );
  OAI21_X1 U5824 ( .B1(n9409), .B2(n6769), .A(n6071), .ZN(n4482) );
  OR2_X1 U5825 ( .A1(n6454), .A2(n7626), .ZN(n7368) );
  OAI211_X1 U5826 ( .C1(P1_B_REG_SCAN_IN), .C2(n7952), .A(n6438), .B(n6435), 
        .ZN(n6760) );
  XNOR2_X1 U5827 ( .A(n5818), .B(n5817), .ZN(n9408) );
  NAND2_X1 U5828 ( .A1(n4748), .A2(n4747), .ZN(n5796) );
  NAND2_X1 U5829 ( .A1(n4750), .A2(SI_29_), .ZN(n4747) );
  XNOR2_X1 U5830 ( .A(n5784), .B(n5783), .ZN(n9091) );
  XNOR2_X1 U5831 ( .A(n6016), .B(n6011), .ZN(n6848) );
  NAND2_X1 U5832 ( .A1(n6015), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  AND2_X1 U5833 ( .A1(n6426), .A2(n6429), .ZN(n4599) );
  INV_X1 U5834 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U5835 ( .A1(n5535), .A2(n5534), .ZN(n5547) );
  NAND2_X1 U5836 ( .A1(n4766), .A2(n5453), .ZN(n5481) );
  NAND2_X1 U5837 ( .A1(n5450), .A2(n4770), .ZN(n4766) );
  NAND2_X1 U5838 ( .A1(n4670), .A2(n5464), .ZN(n4664) );
  OAI21_X1 U5839 ( .B1(n5464), .B2(n4666), .A(n4662), .ZN(n4661) );
  OAI21_X1 U5840 ( .B1(n5434), .B2(n5433), .A(n5401), .ZN(n5448) );
  OAI21_X1 U5841 ( .B1(n5356), .B2(n4759), .A(n4756), .ZN(n5396) );
  NAND2_X1 U5842 ( .A1(n5356), .A2(n5355), .ZN(n5375) );
  XNOR2_X1 U5843 ( .A(n5354), .B(n5353), .ZN(n6772) );
  OR2_X1 U5844 ( .A1(n6168), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U5845 ( .A(n6087), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6856) );
  OR2_X1 U5846 ( .A1(n8720), .A2(n5733), .ZN(n5651) );
  AND2_X1 U5847 ( .A1(n8405), .A2(n4478), .ZN(n8496) );
  INV_X1 U5848 ( .A(n8404), .ZN(n4478) );
  AND2_X1 U5849 ( .A1(n5596), .A2(n5595), .ZN(n8499) );
  OR2_X1 U5850 ( .A1(n8746), .A2(n5733), .ZN(n5596) );
  XNOR2_X1 U5851 ( .A(n5608), .B(n5606), .ZN(n8405) );
  NAND2_X1 U5852 ( .A1(n7861), .A2(n5270), .ZN(n8038) );
  NAND2_X1 U5853 ( .A1(n5122), .A2(n8413), .ZN(n8415) );
  NAND2_X1 U5854 ( .A1(n7273), .A2(n7274), .ZN(n7272) );
  NAND2_X1 U5855 ( .A1(n5546), .A2(n8439), .ZN(n8441) );
  NAND2_X1 U5856 ( .A1(n4946), .A2(n4944), .ZN(n7389) );
  INV_X1 U5857 ( .A(n4947), .ZN(n4946) );
  AOI21_X1 U5858 ( .B1(n4419), .B2(n4952), .A(n4950), .ZN(n4949) );
  NAND2_X1 U5859 ( .A1(n8415), .A2(n5126), .ZN(n7513) );
  NAND2_X1 U5860 ( .A1(n8437), .A2(n5509), .ZN(n8513) );
  INV_X1 U5861 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8522) );
  OAI21_X1 U5862 ( .B1(n7863), .B2(n4594), .A(n4592), .ZN(n8544) );
  NAND2_X1 U5863 ( .A1(n7272), .A2(n5074), .ZN(n7564) );
  AND3_X1 U5864 ( .A1(n5477), .A2(n5476), .A3(n5475), .ZN(n8566) );
  NAND2_X1 U5865 ( .A1(n4930), .A2(n8469), .ZN(n8571) );
  AND3_X1 U5866 ( .A1(n5802), .A2(n5801), .A3(n5800), .ZN(n8646) );
  NAND2_X1 U5867 ( .A1(n5668), .A2(n5667), .ZN(n8595) );
  INV_X1 U5868 ( .A(n8499), .ZN(n8757) );
  INV_X1 U5869 ( .A(n8509), .ZN(n8848) );
  INV_X1 U5870 ( .A(n8488), .ZN(n8598) );
  INV_X2 U5871 ( .A(P2_U3966), .ZN(n8610) );
  NAND2_X1 U5872 ( .A1(n7107), .A2(n7106), .ZN(n7110) );
  INV_X1 U5873 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10203) );
  AOI21_X1 U5874 ( .B1(n7224), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7220), .ZN(
        n7421) );
  AOI22_X1 U5875 ( .A1(n7254), .A2(n7253), .B1(n7255), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7404) );
  OR2_X1 U5876 ( .A1(n7415), .A2(n7414), .ZN(n7453) );
  NOR2_X1 U5877 ( .A1(n7405), .A2(n7406), .ZN(n7462) );
  NAND2_X1 U5878 ( .A1(n7453), .A2(n7452), .ZN(n7455) );
  NAND2_X1 U5879 ( .A1(n7661), .A2(n4700), .ZN(n7662) );
  OR2_X1 U5880 ( .A1(n7713), .A2(n7712), .ZN(n8620) );
  NAND2_X1 U5881 ( .A1(n10351), .A2(n10350), .ZN(n10348) );
  NAND2_X1 U5882 ( .A1(n8620), .A2(n4697), .ZN(n10351) );
  NAND2_X1 U5883 ( .A1(n4698), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4697) );
  INV_X1 U5884 ( .A(n8621), .ZN(n4698) );
  AND2_X1 U5885 ( .A1(n7000), .A2(n6999), .ZN(n10354) );
  XNOR2_X1 U5886 ( .A(n8628), .B(n4695), .ZN(n8623) );
  INV_X1 U5887 ( .A(n8952), .ZN(n8645) );
  NAND2_X1 U5888 ( .A1(n8331), .A2(n8330), .ZN(n8666) );
  AOI21_X1 U5889 ( .B1(n8329), .B2(n8907), .A(n8328), .ZN(n8330) );
  NAND2_X1 U5890 ( .A1(n8325), .A2(n8902), .ZN(n8331) );
  AND2_X1 U5891 ( .A1(n8728), .A2(n8727), .ZN(n8981) );
  NAND2_X1 U5892 ( .A1(n8755), .A2(n5847), .ZN(n8741) );
  NAND2_X1 U5893 ( .A1(n4985), .A2(n4984), .ZN(n8739) );
  NAND2_X1 U5894 ( .A1(n4987), .A2(n4986), .ZN(n8765) );
  AND2_X1 U5895 ( .A1(n8776), .A2(n8775), .ZN(n8995) );
  OR2_X1 U5896 ( .A1(n8788), .A2(n4906), .ZN(n8770) );
  NAND2_X1 U5897 ( .A1(n8886), .A2(n4992), .ZN(n8865) );
  AOI21_X1 U5898 ( .B1(n4997), .B2(n8148), .A(n4996), .ZN(n4993) );
  NAND2_X1 U5899 ( .A1(n8149), .A2(n4997), .ZN(n4994) );
  AND2_X1 U5900 ( .A1(n8174), .A2(n8173), .ZN(n9038) );
  NAND2_X1 U5901 ( .A1(n4999), .A2(n4997), .ZN(n8182) );
  NAND2_X1 U5902 ( .A1(n4999), .A2(n8147), .ZN(n8151) );
  NAND2_X1 U5903 ( .A1(n4981), .A2(n7575), .ZN(n7671) );
  CLKBUF_X1 U5904 ( .A(n7050), .Z(n7051) );
  OAI21_X1 U5905 ( .B1(n8973), .B2(n10418), .A(n8972), .ZN(n8974) );
  OR2_X1 U5906 ( .A1(n9013), .A2(n9012), .ZN(n9077) );
  AND2_X2 U5907 ( .A1(n7014), .A2(n7317), .ZN(n10433) );
  AND2_X1 U5908 ( .A1(n5987), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10379) );
  INV_X1 U5909 ( .A(n10373), .ZN(n10376) );
  NAND2_X1 U5910 ( .A1(n5701), .A2(n5042), .ZN(n9102) );
  NOR2_X1 U5911 ( .A1(n5987), .A2(n4369), .ZN(n7798) );
  INV_X1 U5912 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7509) );
  INV_X1 U5913 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5055) );
  INV_X1 U5914 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7308) );
  NAND2_X1 U5915 ( .A1(n5047), .A2(n5046), .ZN(n5455) );
  INV_X1 U5916 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6976) );
  INV_X1 U5917 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6828) );
  INV_X1 U5918 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6800) );
  INV_X1 U5919 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6794) );
  INV_X1 U5920 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6775) );
  INV_X1 U5921 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6749) );
  XNOR2_X1 U5922 ( .A(n5119), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7131) );
  XNOR2_X1 U5923 ( .A(n4710), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U5924 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4710) );
  AND4_X1 U5925 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n8054)
         );
  NAND2_X1 U5926 ( .A1(n4726), .A2(n7744), .ZN(n4612) );
  NAND2_X1 U5927 ( .A1(n9265), .A2(n9269), .ZN(n9191) );
  INV_X1 U5928 ( .A(n9638), .ZN(n9996) );
  AND3_X1 U5929 ( .A1(n6240), .A2(n6239), .A3(n6238), .ZN(n9974) );
  AND2_X1 U5930 ( .A1(n6329), .A2(n6328), .ZN(n9867) );
  NAND2_X1 U5931 ( .A1(n7378), .A2(n7377), .ZN(n7694) );
  NAND2_X1 U5932 ( .A1(n4582), .A2(n4580), .ZN(n8211) );
  NAND2_X1 U5933 ( .A1(n4588), .A2(n8192), .ZN(n9302) );
  NAND2_X1 U5934 ( .A1(n8188), .A2(n8187), .ZN(n4588) );
  AND2_X1 U5935 ( .A1(n7074), .A2(n9662), .ZN(n9322) );
  INV_X1 U5936 ( .A(n9320), .ZN(n9334) );
  INV_X1 U5937 ( .A(n9646), .ZN(n7855) );
  AND3_X1 U5938 ( .A1(n6832), .A2(n6831), .A3(n6830), .ZN(n9749) );
  INV_X1 U5939 ( .A(n9799), .ZN(n9824) );
  NAND2_X1 U5940 ( .A1(n6077), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U5941 ( .A1(n4547), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6042) );
  OR2_X1 U5942 ( .A1(n9679), .A2(n9678), .ZN(n9681) );
  AND2_X1 U5943 ( .A1(n6969), .A2(n6968), .ZN(n6972) );
  OR2_X1 U5944 ( .A1(P1_U3083), .A2(n6866), .ZN(n10244) );
  XOR2_X1 U5945 ( .A(n7769), .B(n7762), .Z(n7765) );
  XNOR2_X1 U5946 ( .A(n9746), .B(n10043), .ZN(n10045) );
  AND2_X1 U5947 ( .A1(n6377), .A2(n6398), .ZN(n9166) );
  INV_X1 U5948 ( .A(n9782), .ZN(n9783) );
  XNOR2_X1 U5949 ( .A(n4487), .B(n9780), .ZN(n9784) );
  AOI22_X1 U5950 ( .A1(n9781), .A2(n9938), .B1(n9936), .B2(n6361), .ZN(n9782)
         );
  NAND2_X1 U5951 ( .A1(n9788), .A2(n6362), .ZN(n9775) );
  AND2_X1 U5952 ( .A1(n4638), .A2(n4422), .ZN(n9789) );
  INV_X1 U5953 ( .A(n10079), .ZN(n9819) );
  NAND2_X1 U5954 ( .A1(n7950), .A2(n4620), .ZN(n6331) );
  OAI21_X1 U5955 ( .B1(n9907), .B2(n4399), .A(n4623), .ZN(n9855) );
  NAND2_X1 U5956 ( .A1(n9901), .A2(n9516), .ZN(n9883) );
  NAND2_X1 U5957 ( .A1(n4835), .A2(n4833), .ZN(n9873) );
  NAND2_X1 U5958 ( .A1(n6296), .A2(n4836), .ZN(n4835) );
  NAND2_X1 U5959 ( .A1(n6296), .A2(n5006), .ZN(n9889) );
  AND2_X1 U5960 ( .A1(n9927), .A2(n4465), .ZN(n4843) );
  AND2_X1 U5961 ( .A1(n4844), .A2(n4465), .ZN(n4841) );
  AND2_X1 U5962 ( .A1(n4848), .A2(n4846), .ZN(n9941) );
  NAND2_X1 U5963 ( .A1(n4848), .A2(n6252), .ZN(n9942) );
  OR2_X1 U5964 ( .A1(n9952), .A2(n6253), .ZN(n4848) );
  NAND2_X1 U5965 ( .A1(n4866), .A2(n4871), .ZN(n9958) );
  NAND2_X1 U5966 ( .A1(n4643), .A2(n4644), .ZN(n9992) );
  OR2_X1 U5967 ( .A1(n7912), .A2(n4646), .ZN(n4643) );
  NAND2_X1 U5968 ( .A1(n4876), .A2(n9478), .ZN(n10009) );
  NAND2_X1 U5969 ( .A1(n7912), .A2(n6206), .ZN(n10006) );
  NAND2_X1 U5970 ( .A1(n4851), .A2(n4852), .ZN(n7914) );
  NOR2_X1 U5971 ( .A1(n4402), .A2(n4629), .ZN(n4627) );
  NAND2_X1 U5972 ( .A1(n7787), .A2(n6128), .ZN(n7897) );
  XNOR2_X1 U5973 ( .A(n7778), .B(n9587), .ZN(n7779) );
  NAND2_X1 U5974 ( .A1(n10036), .A2(n7627), .ZN(n10024) );
  OR2_X1 U5975 ( .A1(n9409), .A2(n6771), .ZN(n6054) );
  NAND2_X1 U5976 ( .A1(n6284), .A2(n6988), .ZN(n4916) );
  NOR2_X1 U5977 ( .A1(n10021), .A2(n7819), .ZN(n9990) );
  INV_X1 U5978 ( .A(n10024), .ZN(n10032) );
  NAND2_X1 U5979 ( .A1(n4513), .A2(n10325), .ZN(n4512) );
  NOR2_X1 U5980 ( .A1(n7368), .A2(n7367), .ZN(n10272) );
  INV_X1 U5981 ( .A(n10272), .ZN(n10326) );
  AND2_X1 U5982 ( .A1(n7279), .A2(n6442), .ZN(n7286) );
  NAND2_X1 U5983 ( .A1(n7286), .A2(n6760), .ZN(n10255) );
  NAND2_X1 U5984 ( .A1(n6012), .A2(n4855), .ZN(n6027) );
  CLKBUF_X1 U5985 ( .A(n6397), .Z(n10180) );
  INV_X1 U5986 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U5987 ( .A1(n6389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6391) );
  INV_X1 U5988 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7599) );
  INV_X1 U5989 ( .A(n6393), .ZN(n9611) );
  INV_X1 U5990 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7310) );
  INV_X1 U5991 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6991) );
  INV_X1 U5992 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6796) );
  INV_X1 U5993 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U5994 ( .A1(n10210), .A2(n10209), .ZN(n10490) );
  NOR2_X1 U5995 ( .A1(n10216), .A2(n10481), .ZN(n10472) );
  AOI21_X1 U5996 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10470), .ZN(n10469) );
  NOR2_X1 U5997 ( .A1(n10469), .A2(n10468), .ZN(n10467) );
  AOI21_X1 U5998 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10467), .ZN(n10466) );
  OAI21_X1 U5999 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10464), .ZN(n10462) );
  OAI21_X1 U6000 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10458), .ZN(n10456) );
  NAND2_X1 U6001 ( .A1(n7491), .A2(n5193), .ZN(n7589) );
  OAI211_X1 U6002 ( .C1(n4934), .C2(n4926), .A(n4924), .B(n4408), .ZN(n5751)
         );
  NAND2_X1 U6003 ( .A1(n4610), .A2(n4608), .ZN(P2_U3227) );
  NOR2_X1 U6004 ( .A1(n8472), .A2(n4609), .ZN(n4608) );
  AOI21_X1 U6005 ( .B1(n4708), .B2(n8640), .A(n4707), .ZN(n4706) );
  INV_X1 U6006 ( .A(n4893), .ZN(n8683) );
  AOI21_X1 U6007 ( .B1(n8960), .B2(n8944), .A(n8682), .ZN(n4894) );
  AOI211_X1 U6008 ( .C1(n8965), .C2(n8944), .A(n8703), .B(n8702), .ZN(n8704)
         );
  NAND2_X1 U6009 ( .A1(n10441), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U6010 ( .A1(n8365), .A2(n10444), .ZN(n4650) );
  NAND2_X1 U6011 ( .A1(n9175), .A2(n4490), .ZN(n9174) );
  NAND2_X1 U6012 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  INV_X1 U6013 ( .A(n4502), .ZN(n4501) );
  OR2_X1 U6014 ( .A1(n9741), .A2(n9615), .ZN(n4503) );
  OR2_X1 U6015 ( .A1(n9742), .A2(n9740), .ZN(n4500) );
  INV_X1 U6016 ( .A(n4508), .ZN(n9773) );
  INV_X2 U6017 ( .A(n4400), .ZN(n5976) );
  OR2_X1 U6018 ( .A1(n4830), .A2(n4403), .ZN(n4399) );
  NOR2_X1 U6019 ( .A1(n5058), .A2(n5846), .ZN(n4400) );
  INV_X1 U6020 ( .A(n8790), .ZN(n4905) );
  XNOR2_X1 U6021 ( .A(n6391), .B(n6390), .ZN(n6392) );
  NAND2_X1 U6022 ( .A1(n9779), .A2(n9800), .ZN(n4401) );
  AND2_X1 U6023 ( .A1(n7895), .A2(n6410), .ZN(n4402) );
  AND2_X1 U6024 ( .A1(n4377), .A2(n4839), .ZN(n4403) );
  OR2_X1 U6025 ( .A1(n6281), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4404) );
  INV_X1 U6026 ( .A(n5922), .ZN(n4807) );
  AND2_X1 U6027 ( .A1(n4756), .A2(n5393), .ZN(n4405) );
  INV_X1 U6028 ( .A(n4396), .ZN(n4489) );
  AND2_X1 U6029 ( .A1(n4929), .A2(n5726), .ZN(n4406) );
  NOR2_X1 U6030 ( .A1(n9000), .A2(n8773), .ZN(n4407) );
  AND2_X1 U6031 ( .A1(n4449), .A2(n4923), .ZN(n4408) );
  AND2_X1 U6032 ( .A1(n8530), .A2(n8532), .ZN(n4409) );
  AND3_X1 U6033 ( .A1(n9438), .A2(n9440), .A3(n9439), .ZN(n4410) );
  INV_X1 U6034 ( .A(n4387), .ZN(n4962) );
  AND2_X1 U6035 ( .A1(n5762), .A2(n5761), .ZN(n8905) );
  AND2_X1 U6036 ( .A1(n4540), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U6037 ( .A1(n4628), .A2(n4625), .ZN(n7873) );
  NAND2_X1 U6038 ( .A1(n7992), .A2(n4901), .ZN(n8146) );
  INV_X1 U6039 ( .A(n5754), .ZN(n5753) );
  AND2_X1 U6040 ( .A1(n9646), .A2(n10286), .ZN(n4412) );
  INV_X1 U6041 ( .A(n9276), .ZN(n4574) );
  AND2_X1 U6042 ( .A1(n10356), .A2(n4472), .ZN(n4413) );
  NAND2_X1 U6043 ( .A1(n6392), .A2(n9740), .ZN(n9540) );
  AND2_X1 U6044 ( .A1(n4799), .A2(n5894), .ZN(n4414) );
  INV_X2 U6045 ( .A(n8237), .ZN(n8217) );
  NAND2_X1 U6046 ( .A1(n4605), .A2(n4949), .ZN(n8422) );
  NAND2_X1 U6047 ( .A1(n4640), .A2(n4639), .ZN(n9952) );
  INV_X1 U6048 ( .A(n7018), .ZN(n7630) );
  NAND4_X1 U6049 ( .A1(n9522), .A2(n9521), .A3(n9520), .A4(n9519), .ZN(n4415)
         );
  AND2_X1 U6050 ( .A1(n6265), .A2(n6254), .ZN(n4416) );
  INV_X1 U6051 ( .A(n5129), .ZN(n5313) );
  AND2_X1 U6052 ( .A1(n9864), .A2(n9426), .ZN(n4417) );
  AND2_X1 U6053 ( .A1(n4963), .A2(n8748), .ZN(n4418) );
  XNOR2_X1 U6054 ( .A(n5451), .B(SI_17_), .ZN(n5464) );
  INV_X1 U6055 ( .A(n5464), .ZN(n5454) );
  INV_X1 U6056 ( .A(n8469), .ZN(n4936) );
  AND2_X1 U6057 ( .A1(n5441), .A2(n4951), .ZN(n4419) );
  AND2_X1 U6058 ( .A1(n5933), .A2(n5932), .ZN(n8771) );
  INV_X1 U6059 ( .A(n8771), .ZN(n4988) );
  NAND2_X1 U6060 ( .A1(n8811), .A2(n8348), .ZN(n8787) );
  AND3_X1 U6061 ( .A1(n4372), .A2(n6111), .A3(n6428), .ZN(n4420) );
  INV_X1 U6062 ( .A(n8333), .ZN(n4485) );
  INV_X1 U6063 ( .A(n5969), .ZN(n4689) );
  OR3_X1 U6064 ( .A1(n4936), .A2(n8466), .A3(n8579), .ZN(n4421) );
  INV_X1 U6065 ( .A(n8825), .ZN(n4806) );
  INV_X1 U6066 ( .A(n9433), .ZN(n4872) );
  NAND2_X1 U6067 ( .A1(n9815), .A2(n4920), .ZN(n9760) );
  NOR2_X1 U6068 ( .A1(n8916), .A2(n4970), .ZN(n8850) );
  NOR2_X1 U6069 ( .A1(n8789), .A2(n8790), .ZN(n8788) );
  NAND2_X1 U6070 ( .A1(n5770), .A2(n4693), .ZN(n8805) );
  AND2_X1 U6071 ( .A1(n5662), .A2(n5661), .ZN(n8692) );
  INV_X1 U6072 ( .A(n8766), .ZN(n4826) );
  NAND2_X1 U6073 ( .A1(n5770), .A2(n5922), .ZN(n8803) );
  NAND2_X1 U6074 ( .A1(n9819), .A2(n9799), .ZN(n4422) );
  INV_X1 U6075 ( .A(n8382), .ZN(n4929) );
  AND2_X1 U6076 ( .A1(n5990), .A2(n4820), .ZN(n4423) );
  NAND2_X1 U6077 ( .A1(n6053), .A2(n6066), .ZN(n6849) );
  AND2_X1 U6078 ( .A1(n6038), .A2(n6037), .ZN(n9866) );
  INV_X1 U6079 ( .A(n9866), .ZN(n4839) );
  AND2_X1 U6080 ( .A1(n4987), .A2(n8350), .ZN(n4424) );
  INV_X1 U6081 ( .A(n5726), .ZN(n4938) );
  NOR2_X1 U6082 ( .A1(n5877), .A2(n7579), .ZN(n4425) );
  AND2_X1 U6083 ( .A1(n9456), .A2(n9454), .ZN(n9588) );
  INV_X1 U6084 ( .A(n9588), .ZN(n6410) );
  AND2_X1 U6085 ( .A1(n7953), .A2(n9471), .ZN(n4426) );
  OR2_X1 U6086 ( .A1(n10051), .A2(n9540), .ZN(n4427) );
  NAND2_X1 U6087 ( .A1(n5828), .A2(n5956), .ZN(n8686) );
  XNOR2_X1 U6088 ( .A(n5394), .B(SI_14_), .ZN(n5393) );
  INV_X1 U6089 ( .A(n5730), .ZN(n4937) );
  AND2_X1 U6090 ( .A1(n4886), .A2(n9347), .ZN(n4428) );
  INV_X1 U6091 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9088) );
  AND2_X1 U6092 ( .A1(n9606), .A2(n4545), .ZN(n4429) );
  INV_X1 U6093 ( .A(n4928), .ZN(n4927) );
  OAI21_X1 U6094 ( .B1(n4931), .B2(n4929), .A(n4442), .ZN(n4928) );
  AND2_X1 U6095 ( .A1(n10141), .A2(n9638), .ZN(n4430) );
  NAND2_X1 U6096 ( .A1(n9220), .A2(n9224), .ZN(n4431) );
  AND2_X1 U6097 ( .A1(n8710), .A2(n8711), .ZN(n4432) );
  AND2_X1 U6098 ( .A1(n4658), .A2(n5326), .ZN(n4433) );
  INV_X1 U6099 ( .A(n8181), .ZN(n4996) );
  INV_X1 U6100 ( .A(n8127), .ZN(n5889) );
  AND2_X1 U6101 ( .A1(n4418), .A2(n4962), .ZN(n4434) );
  INV_X1 U6102 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6013) );
  AND2_X1 U6103 ( .A1(n5830), .A2(n8845), .ZN(n4435) );
  OR2_X1 U6104 ( .A1(n6282), .A2(n6281), .ZN(n4436) );
  AND2_X1 U6105 ( .A1(n8987), .A2(n8774), .ZN(n4437) );
  AND2_X1 U6106 ( .A1(n8692), .A2(n8354), .ZN(n4438) );
  NOR2_X1 U6107 ( .A1(n10136), .A2(n9637), .ZN(n4439) );
  NOR2_X1 U6108 ( .A1(n9020), .A2(n8888), .ZN(n4440) );
  INV_X1 U6109 ( .A(n4972), .ZN(n8915) );
  NOR2_X1 U6110 ( .A1(n8916), .A2(n9030), .ZN(n4972) );
  NOR2_X1 U6111 ( .A1(n9792), .A2(n10067), .ZN(n4922) );
  INV_X1 U6112 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U6113 ( .A1(n5404), .A2(n5403), .ZN(n5449) );
  INV_X1 U6114 ( .A(n5449), .ZN(n4667) );
  AND2_X1 U6115 ( .A1(n4577), .A2(n4574), .ZN(n4441) );
  NAND2_X1 U6116 ( .A1(n5671), .A2(n5670), .ZN(n4442) );
  INV_X1 U6117 ( .A(n9107), .ZN(n4741) );
  INV_X1 U6118 ( .A(n4909), .ZN(n4908) );
  NAND2_X1 U6119 ( .A1(n4910), .A2(n4911), .ZN(n4909) );
  INV_X1 U6120 ( .A(n10380), .ZN(n4973) );
  AND2_X1 U6121 ( .A1(n5482), .A2(SI_18_), .ZN(n4443) );
  INV_X1 U6122 ( .A(n6308), .ZN(n4840) );
  AND2_X1 U6123 ( .A1(n10103), .A2(n9635), .ZN(n6308) );
  INV_X1 U6124 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6382) );
  AND4_X1 U6125 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n7839)
         );
  AND2_X1 U6126 ( .A1(n5651), .A2(n5650), .ZN(n8698) );
  INV_X1 U6127 ( .A(n8698), .ZN(n4532) );
  AND2_X1 U6128 ( .A1(n8200), .A2(n9299), .ZN(n4444) );
  AND2_X1 U6129 ( .A1(n5297), .A2(n5296), .ZN(n4445) );
  AND2_X1 U6130 ( .A1(n5395), .A2(SI_14_), .ZN(n4446) );
  NAND2_X1 U6131 ( .A1(n8437), .A2(n4958), .ZN(n8438) );
  AND2_X1 U6132 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n4820), .ZN(n4447) );
  NAND2_X1 U6133 ( .A1(n7955), .A2(n7954), .ZN(n4448) );
  INV_X1 U6134 ( .A(n4670), .ZN(n4669) );
  AND2_X1 U6135 ( .A1(n4671), .A2(n5011), .ZN(n4670) );
  AND2_X1 U6136 ( .A1(n9797), .A2(n4422), .ZN(n4637) );
  OR2_X1 U6137 ( .A1(n4927), .A2(n5730), .ZN(n4449) );
  INV_X1 U6138 ( .A(n4902), .ZN(n4901) );
  NAND2_X1 U6139 ( .A1(n8150), .A2(n5899), .ZN(n4902) );
  AND3_X1 U6140 ( .A1(n8677), .A2(n8694), .A3(n5843), .ZN(n4450) );
  AND2_X1 U6141 ( .A1(n4666), .A2(n5454), .ZN(n4451) );
  OR2_X1 U6142 ( .A1(n8261), .A2(n8260), .ZN(n4452) );
  AND3_X1 U6143 ( .A1(n10399), .A2(n7311), .A3(n7352), .ZN(n4453) );
  AND2_X1 U6144 ( .A1(n6412), .A2(n9478), .ZN(n4454) );
  AND2_X1 U6145 ( .A1(n6010), .A2(n6011), .ZN(n4455) );
  AND4_X1 U6146 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n7615)
         );
  NAND2_X1 U6147 ( .A1(n5775), .A2(n5774), .ZN(n8740) );
  INV_X1 U6148 ( .A(n8740), .ZN(n4648) );
  NAND2_X1 U6149 ( .A1(n7855), .A2(n7786), .ZN(n9439) );
  AND2_X1 U6150 ( .A1(n5760), .A2(n8148), .ZN(n4456) );
  AND2_X1 U6151 ( .A1(n9538), .A2(n9537), .ZN(n4457) );
  INV_X1 U6152 ( .A(n7853), .ZN(n6421) );
  AND2_X1 U6153 ( .A1(n9603), .A2(n9525), .ZN(n4458) );
  AND2_X1 U6154 ( .A1(n9269), .A2(n8267), .ZN(n4459) );
  AND2_X1 U6155 ( .A1(n4552), .A2(n4550), .ZN(n4460) );
  NAND2_X1 U6156 ( .A1(n7615), .A2(n7987), .ZN(n9369) );
  AND2_X1 U6157 ( .A1(n6128), .A2(n6410), .ZN(n4461) );
  OR2_X1 U6158 ( .A1(n4576), .A2(n4574), .ZN(n4462) );
  OR2_X1 U6159 ( .A1(n8363), .A2(n8362), .ZN(n4463) );
  AND2_X2 U6160 ( .A1(n7014), .A2(n7013), .ZN(n10444) );
  INV_X1 U6161 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4516) );
  AND2_X1 U6162 ( .A1(n6387), .A2(n6389), .ZN(n6393) );
  INV_X1 U6163 ( .A(n8439), .ZN(n4941) );
  NAND2_X1 U6164 ( .A1(n4891), .A2(n4890), .ZN(n7676) );
  OR2_X1 U6165 ( .A1(n9964), .A2(n10119), .ZN(n4464) );
  INV_X1 U6166 ( .A(n8681), .ZN(n4895) );
  INV_X1 U6167 ( .A(n9461), .ZN(n4507) );
  NAND2_X1 U6168 ( .A1(n4994), .A2(n4993), .ZN(n8332) );
  NAND2_X1 U6169 ( .A1(n4733), .A2(n4731), .ZN(n8188) );
  NAND2_X1 U6170 ( .A1(n4692), .A2(n5856), .ZN(n7320) );
  OR2_X1 U6171 ( .A1(n10119), .A2(n6264), .ZN(n4465) );
  AOI21_X1 U6172 ( .B1(n8734), .B2(n4393), .A(n5630), .ZN(n8502) );
  AND2_X1 U6173 ( .A1(n4628), .A2(n4627), .ZN(n7872) );
  INV_X1 U6174 ( .A(n8148), .ZN(n5000) );
  NAND2_X1 U6175 ( .A1(n4980), .A2(n4983), .ZN(n7672) );
  INV_X1 U6176 ( .A(n9563), .ZN(n4551) );
  INV_X1 U6177 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4527) );
  NAND2_X1 U6178 ( .A1(n7958), .A2(n4908), .ZN(n4912) );
  INV_X1 U6179 ( .A(n9492), .ZN(n4864) );
  INV_X1 U6180 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U6181 ( .A1(n8886), .A2(n8341), .ZN(n4466) );
  NAND2_X1 U6182 ( .A1(n6427), .A2(n6426), .ZN(n4467) );
  INV_X1 U6183 ( .A(n5012), .ZN(n4629) );
  INV_X1 U6184 ( .A(n4751), .ZN(n4750) );
  NAND2_X1 U6185 ( .A1(n4752), .A2(n5806), .ZN(n4751) );
  AND2_X1 U6186 ( .A1(n4536), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4468) );
  AND2_X1 U6187 ( .A1(n4845), .A2(n4841), .ZN(n4469) );
  AND2_X1 U6188 ( .A1(n7992), .A2(n5899), .ZN(n4470) );
  INV_X1 U6189 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5425) );
  INV_X1 U6190 ( .A(n5752), .ZN(n7336) );
  INV_X1 U6191 ( .A(n8077), .ZN(n4479) );
  INV_X1 U6192 ( .A(n7521), .ZN(n4603) );
  INV_X1 U6193 ( .A(n10136), .ZN(n4910) );
  AND2_X1 U6194 ( .A1(n10311), .A2(n10133), .ZN(n10144) );
  INV_X1 U6195 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4820) );
  AND2_X1 U6196 ( .A1(n7536), .A2(n7570), .ZN(n7537) );
  NAND2_X1 U6197 ( .A1(n5831), .A2(n6809), .ZN(n7347) );
  INV_X1 U6198 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4537) );
  INV_X1 U6199 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4538) );
  NAND2_X1 U6200 ( .A1(n8646), .A2(n5851), .ZN(n4471) );
  INV_X1 U6201 ( .A(n8627), .ZN(n4695) );
  INV_X1 U6202 ( .A(n9740), .ZN(n9615) );
  AOI21_X1 U6203 ( .B1(n10055), .B2(n10019), .A(n9772), .ZN(n4509) );
  NOR2_X2 U6204 ( .A1(n7633), .A2(n9740), .ZN(n10019) );
  OAI211_X2 U6205 ( .C1(n9850), .C2(n4883), .A(n4882), .B(n6415), .ZN(n9810)
         );
  OAI21_X1 U6206 ( .B1(n8641), .B2(n8640), .A(n4706), .ZN(P2_U3264) );
  OAI21_X1 U6207 ( .B1(n8638), .B2(n8637), .A(n4709), .ZN(n4708) );
  NAND2_X1 U6208 ( .A1(n5169), .A2(SI_4_), .ZN(n5166) );
  NOR2_X1 U6209 ( .A1(n4718), .A2(n4474), .ZN(n9544) );
  NOR2_X1 U6210 ( .A1(n9541), .A2(n4427), .ZN(n4474) );
  INV_X1 U6211 ( .A(n8377), .ZN(n4513) );
  NAND2_X1 U6212 ( .A1(n4632), .A2(n4631), .ZN(n10062) );
  AOI21_X1 U6213 ( .B1(n4771), .B2(n9579), .A(n4457), .ZN(n9539) );
  NAND2_X4 U6214 ( .A1(n5059), .A2(n7318), .ZN(n5643) );
  NAND2_X1 U6215 ( .A1(n4477), .A2(n4475), .ZN(n8508) );
  NAND2_X1 U6216 ( .A1(n4476), .A2(n5610), .ZN(n4475) );
  INV_X1 U6217 ( .A(n8501), .ZN(n4476) );
  OAI22_X1 U6218 ( .A1(n8501), .A2(n8579), .B1(n8499), .B2(n8559), .ZN(n4477)
         );
  NAND2_X1 U6219 ( .A1(n8518), .A2(n4419), .ZN(n4605) );
  OR2_X1 U6220 ( .A1(n8370), .A2(n6423), .ZN(n6424) );
  XNOR2_X1 U6221 ( .A(n5091), .B(n5090), .ZN(n6768) );
  AOI21_X2 U6222 ( .B1(n8022), .B2(n9441), .A(n4507), .ZN(n5003) );
  NAND2_X1 U6223 ( .A1(n4865), .A2(n4863), .ZN(n9935) );
  INV_X1 U6224 ( .A(n7161), .ZN(n7987) );
  NAND3_X1 U6225 ( .A1(n7040), .A2(n7161), .A3(n6406), .ZN(n7973) );
  AND2_X2 U6226 ( .A1(n4618), .A2(n4481), .ZN(n7161) );
  NAND2_X1 U6227 ( .A1(n10007), .A2(n9380), .ZN(n9994) );
  NAND2_X1 U6228 ( .A1(n9369), .A2(n6408), .ZN(n4714) );
  OAI211_X1 U6229 ( .C1(n4458), .C2(n4564), .A(n9534), .B(n9533), .ZN(n4559)
         );
  NOR2_X1 U6230 ( .A1(n4563), .A2(n4564), .ZN(n4562) );
  AOI21_X1 U6231 ( .B1(n9541), .B2(n4721), .A(n4719), .ZN(n4718) );
  NAND2_X1 U6232 ( .A1(n5991), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5043) );
  INV_X1 U6233 ( .A(n5026), .ZN(n5697) );
  AND2_X2 U6234 ( .A1(n5022), .A2(n5021), .ZN(n5026) );
  MUX2_X1 U6235 ( .A(n7806), .B(n5883), .S(n5976), .Z(n5884) );
  NAND2_X1 U6236 ( .A1(n4797), .A2(n4801), .ZN(n4796) );
  AOI21_X1 U6237 ( .B1(n4827), .B2(n4823), .A(n4821), .ZN(n5945) );
  NAND3_X1 U6238 ( .A1(n4794), .A2(n4793), .A3(n4792), .ZN(n4486) );
  OAI21_X1 U6239 ( .B1(n5924), .B2(n5923), .A(n4805), .ZN(n5926) );
  NAND2_X1 U6240 ( .A1(n4665), .A2(n4670), .ZN(n5450) );
  NAND2_X1 U6241 ( .A1(n5533), .A2(n5532), .ZN(n5535) );
  NAND2_X1 U6242 ( .A1(n4760), .A2(n5551), .ZN(n5574) );
  XNOR2_X1 U6243 ( .A(n5136), .B(n5109), .ZN(n5135) );
  NAND2_X1 U6244 ( .A1(n4488), .A2(n4515), .ZN(n5136) );
  NAND2_X1 U6245 ( .A1(n4489), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4488) );
  MUX2_X1 U6246 ( .A(n5952), .B(n5951), .S(n5976), .Z(n5953) );
  MUX2_X1 U6247 ( .A(n9421), .B(n9420), .S(n9540), .Z(n9526) );
  NOR2_X1 U6248 ( .A1(n9541), .A2(n4772), .ZN(n4771) );
  INV_X1 U6249 ( .A(n9827), .ZN(n4885) );
  NAND2_X1 U6250 ( .A1(n5948), .A2(n8711), .ZN(n4530) );
  NAND2_X2 U6251 ( .A1(n6331), .A2(n6330), .ZN(n9836) );
  NAND2_X1 U6252 ( .A1(n8249), .A2(n4371), .ZN(n4573) );
  NAND2_X1 U6253 ( .A1(n4722), .A2(n4723), .ZN(n9190) );
  NAND2_X1 U6254 ( .A1(n4601), .A2(n8315), .ZN(n4600) );
  NAND2_X1 U6255 ( .A1(n8912), .A2(n8914), .ZN(n8913) );
  NAND3_X1 U6256 ( .A1(n4450), .A2(n4495), .A3(n4494), .ZN(n4493) );
  NAND2_X1 U6257 ( .A1(n4884), .A2(n9840), .ZN(n4882) );
  NAND2_X1 U6258 ( .A1(n4764), .A2(n4765), .ZN(n5512) );
  NAND2_X1 U6259 ( .A1(n5584), .A2(n5583), .ZN(n5586) );
  AOI21_X1 U6260 ( .B1(n9605), .B2(n6419), .A(n9763), .ZN(n6420) );
  AOI21_X1 U6261 ( .B1(n10154), .B2(n10344), .A(n6457), .ZN(n6718) );
  MUX2_X1 U6262 ( .A(n5898), .B(n5897), .S(n5976), .Z(n5902) );
  AOI21_X1 U6263 ( .B1(n5938), .B2(n5937), .A(n4824), .ZN(n4823) );
  NAND3_X1 U6264 ( .A1(n4796), .A2(n8150), .A3(n4800), .ZN(n4794) );
  NAND2_X2 U6265 ( .A1(n9881), .A2(n9431), .ZN(n9861) );
  NAND2_X1 U6266 ( .A1(n4876), .A2(n4454), .ZN(n10007) );
  NAND2_X1 U6267 ( .A1(n4497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U6268 ( .A1(n7907), .A2(n9444), .ZN(n4876) );
  NAND2_X1 U6269 ( .A1(n9557), .A2(n4412), .ZN(n9561) );
  NAND4_X1 U6270 ( .A1(n4372), .A2(n6111), .A3(n6426), .A4(n4455), .ZN(n4497)
         );
  NAND2_X1 U6271 ( .A1(n4871), .A2(n4869), .ZN(n4868) );
  NAND2_X1 U6272 ( .A1(n4498), .A2(n7798), .ZN(n5996) );
  OAI211_X1 U6273 ( .C1(n5985), .C2(n5984), .A(n4815), .B(n5986), .ZN(n4498)
         );
  NAND2_X1 U6274 ( .A1(n4499), .A2(n5954), .ZN(n4504) );
  NAND2_X1 U6275 ( .A1(n5946), .A2(n5947), .ZN(n4499) );
  NAND2_X1 U6276 ( .A1(n4828), .A2(n5976), .ZN(n4827) );
  AOI211_X1 U6277 ( .C1(n5973), .C2(n5972), .A(n5971), .B(n5970), .ZN(n5981)
         );
  NOR2_X1 U6278 ( .A1(n8110), .A2(n8109), .ZN(n9725) );
  NAND3_X1 U6279 ( .A1(n4503), .A2(n4501), .A3(n4500), .ZN(P1_U3260) );
  NAND2_X1 U6280 ( .A1(n5134), .A2(n5135), .ZN(n5168) );
  NAND2_X1 U6281 ( .A1(n5116), .A2(n5115), .ZN(n5134) );
  NAND2_X1 U6282 ( .A1(n7802), .A2(n7801), .ZN(n8001) );
  NAND2_X1 U6283 ( .A1(n4504), .A2(n8694), .ZN(n4790) );
  INV_X1 U6284 ( .A(n5776), .ZN(n5952) );
  OAI21_X2 U6285 ( .B1(n5512), .B2(n5511), .A(n5510), .ZN(n5533) );
  NAND3_X1 U6286 ( .A1(n5245), .A2(n5242), .A3(n5243), .ZN(n5274) );
  OAI21_X1 U6287 ( .B1(n4397), .B2(n4506), .A(n4505), .ZN(n5238) );
  NAND2_X1 U6288 ( .A1(n6425), .A2(n4512), .ZN(n10154) );
  AOI21_X2 U6289 ( .B1(n9287), .B2(n9289), .A(n8298), .ZN(n9133) );
  OAI21_X2 U6290 ( .B1(n9133), .B2(n9135), .A(n9132), .ZN(n9257) );
  NAND2_X1 U6291 ( .A1(n4743), .A2(n4742), .ZN(n4601) );
  AOI21_X1 U6292 ( .B1(n4602), .B2(n4600), .A(n8322), .ZN(n8323) );
  OAI21_X1 U6293 ( .B1(n4397), .B2(n4511), .A(n4510), .ZN(n5174) );
  AOI21_X2 U6294 ( .B1(n5042), .B2(n4961), .A(n4447), .ZN(n4818) );
  NAND2_X1 U6295 ( .A1(n8358), .A2(n8651), .ZN(n8664) );
  NAND2_X1 U6296 ( .A1(n9890), .A2(n9894), .ZN(n9891) );
  AND2_X2 U6297 ( .A1(n4453), .A2(n7353), .ZN(n7536) );
  NOR2_X4 U6298 ( .A1(n8817), .A2(n9000), .ZN(n8796) );
  NAND2_X1 U6299 ( .A1(n4650), .A2(n4649), .ZN(P2_U3549) );
  INV_X1 U6300 ( .A(n4922), .ZN(n9776) );
  INV_X1 U6301 ( .A(n6768), .ZN(n4619) );
  NAND2_X1 U6302 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  NAND4_X1 U6303 ( .A1(n4535), .A2(n4463), .A3(n8364), .A4(n4534), .ZN(n8365)
         );
  NAND2_X1 U6304 ( .A1(n5168), .A2(n4514), .ZN(n5173) );
  AND2_X1 U6305 ( .A1(n5166), .A2(n5167), .ZN(n4514) );
  NAND2_X1 U6306 ( .A1(n8903), .A2(n5762), .ZN(n8844) );
  NAND2_X1 U6307 ( .A1(n4543), .A2(n4541), .ZN(n9631) );
  AOI21_X2 U6308 ( .B1(n4560), .B2(n4415), .A(n4518), .ZN(n9541) );
  INV_X1 U6309 ( .A(n5884), .ZN(n4804) );
  NAND2_X1 U6310 ( .A1(n4802), .A2(n5885), .ZN(n4799) );
  NAND2_X1 U6311 ( .A1(n5984), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U6312 ( .A1(n4813), .A2(n8914), .ZN(n4812) );
  NAND2_X1 U6313 ( .A1(n4814), .A2(n4808), .ZN(n5924) );
  OAI21_X1 U6314 ( .B1(n5935), .B2(n5934), .A(n5933), .ZN(n4828) );
  NAND4_X2 U6315 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n9646)
         );
  NAND2_X2 U6316 ( .A1(n9861), .A2(n9864), .ZN(n9850) );
  INV_X1 U6317 ( .A(n9373), .ZN(n4878) );
  OAI21_X1 U6318 ( .B1(n9798), .B2(n4862), .A(n4860), .ZN(n6418) );
  INV_X1 U6319 ( .A(n9914), .ZN(n4525) );
  NAND2_X1 U6320 ( .A1(n4790), .A2(n5961), .ZN(n5964) );
  NAND2_X2 U6321 ( .A1(n9898), .A2(n6413), .ZN(n9901) );
  NOR2_X1 U6322 ( .A1(n10070), .A2(n10021), .ZN(n9785) );
  AND2_X1 U6323 ( .A1(n9561), .A2(n9374), .ZN(n6409) );
  NAND2_X1 U6324 ( .A1(n4528), .A2(n4526), .ZN(n5228) );
  INV_X1 U6325 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U6326 ( .A1(n5589), .A2(n4533), .ZN(n5626) );
  NAND2_X1 U6327 ( .A1(n5589), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5599) );
  INV_X1 U6328 ( .A(n5626), .ZN(n5624) );
  NAND2_X1 U6329 ( .A1(n5459), .A2(n4468), .ZN(n5538) );
  NAND2_X2 U6330 ( .A1(n4548), .A2(n9555), .ZN(n7778) );
  NAND3_X1 U6331 ( .A1(n4549), .A2(n8010), .A3(n9558), .ZN(n4548) );
  NAND3_X1 U6332 ( .A1(n4554), .A2(n4553), .A3(n4410), .ZN(n4552) );
  NAND3_X1 U6333 ( .A1(n4554), .A2(n9438), .A3(n4553), .ZN(n9455) );
  OR2_X1 U6334 ( .A1(n9437), .A2(n9540), .ZN(n4554) );
  NAND2_X1 U6335 ( .A1(n4555), .A2(n9497), .ZN(n9511) );
  AND2_X1 U6336 ( .A1(n4562), .A2(n4561), .ZN(n4560) );
  INV_X1 U6337 ( .A(n9536), .ZN(n4563) );
  NAND2_X1 U6338 ( .A1(n6010), .A2(n6002), .ZN(n4568) );
  NAND4_X1 U6339 ( .A1(n4566), .A2(n4567), .A3(n4372), .A4(n4856), .ZN(n6030)
         );
  NAND3_X1 U6340 ( .A1(n4566), .A2(n4567), .A3(n4372), .ZN(n6015) );
  AND2_X2 U6341 ( .A1(n6003), .A2(n6002), .ZN(n6111) );
  NAND2_X1 U6342 ( .A1(n4572), .A2(n9279), .ZN(n4571) );
  NAND2_X1 U6343 ( .A1(n4462), .A2(n4573), .ZN(n4572) );
  OAI21_X1 U6344 ( .B1(n9279), .B2(n4570), .A(n4572), .ZN(n9144) );
  NOR2_X1 U6345 ( .A1(n4570), .A2(n4452), .ZN(n4569) );
  INV_X1 U6346 ( .A(n8249), .ZN(n4576) );
  OR2_X1 U6347 ( .A1(n9279), .A2(n9276), .ZN(n4579) );
  INV_X4 U6348 ( .A(n7022), .ZN(n9159) );
  NAND2_X1 U6349 ( .A1(n8188), .A2(n4583), .ZN(n4582) );
  OAI21_X1 U6350 ( .B1(n8188), .B2(n4585), .A(n4583), .ZN(n9201) );
  AOI21_X1 U6351 ( .B1(n4583), .B2(n4585), .A(n4581), .ZN(n4580) );
  NAND2_X1 U6352 ( .A1(n7863), .A2(n4592), .ZN(n4589) );
  NAND2_X1 U6353 ( .A1(n4589), .A2(n4590), .ZN(n5322) );
  NAND2_X1 U6354 ( .A1(n4947), .A2(n5165), .ZN(n4597) );
  NAND3_X1 U6355 ( .A1(n4597), .A2(n4596), .A3(n4595), .ZN(n7492) );
  NAND3_X1 U6356 ( .A1(n4945), .A2(n5165), .A3(n4943), .ZN(n4595) );
  NAND2_X1 U6357 ( .A1(n4945), .A2(n4943), .ZN(n4944) );
  NAND2_X1 U6358 ( .A1(n4599), .A2(n4420), .ZN(n4598) );
  AND2_X2 U6359 ( .A1(n4372), .A2(n6111), .ZN(n6427) );
  XNOR2_X2 U6360 ( .A(n5057), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8640) );
  MUX2_X1 U6361 ( .A(n4421), .B(n4611), .S(n8470), .Z(n4610) );
  NAND3_X1 U6362 ( .A1(n5612), .A2(n5613), .A3(n5611), .ZN(n8470) );
  NAND3_X1 U6363 ( .A1(n4613), .A2(n7846), .A3(n4612), .ZN(n7751) );
  NAND3_X1 U6364 ( .A1(n7378), .A2(n4729), .A3(n7744), .ZN(n4613) );
  AND4_X2 U6365 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n5198)
         );
  INV_X2 U6366 ( .A(n6065), .ZN(n4620) );
  NOR3_X1 U6367 ( .A1(n4622), .A2(n4621), .A3(n5007), .ZN(n9841) );
  NAND2_X1 U6368 ( .A1(n7787), .A2(n4461), .ZN(n4628) );
  OR2_X1 U6369 ( .A1(n9805), .A2(n4635), .ZN(n4630) );
  NAND2_X1 U6370 ( .A1(n9805), .A2(n9807), .ZN(n4638) );
  NAND2_X1 U6371 ( .A1(n4630), .A2(n4633), .ZN(n6381) );
  AOI21_X1 U6372 ( .B1(n4633), .B2(n4635), .A(n9534), .ZN(n4631) );
  NAND2_X1 U6373 ( .A1(n9805), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U6374 ( .A1(n7912), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U6375 ( .A1(n5300), .A2(n5299), .ZN(n5328) );
  NAND2_X1 U6376 ( .A1(n4659), .A2(n5326), .ZN(n5354) );
  NAND2_X1 U6377 ( .A1(n5356), .A2(n4405), .ZN(n4755) );
  NAND2_X1 U6378 ( .A1(n5434), .A2(n4451), .ZN(n4660) );
  NAND2_X1 U6379 ( .A1(n5434), .A2(n5401), .ZN(n4665) );
  NAND2_X1 U6380 ( .A1(n5757), .A2(n5876), .ZN(n7578) );
  NAND2_X1 U6381 ( .A1(n8128), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U6382 ( .A1(n4678), .A2(n4679), .ZN(n5824) );
  NAND2_X1 U6383 ( .A1(n8678), .A2(n4680), .ZN(n4678) );
  NAND2_X1 U6384 ( .A1(n8678), .A2(n5782), .ZN(n8324) );
  NAND2_X1 U6385 ( .A1(n4692), .A2(n4691), .ZN(n7546) );
  INV_X4 U6386 ( .A(n4817), .ZN(n5487) );
  NAND2_X1 U6387 ( .A1(n4376), .A2(n6727), .ZN(n5108) );
  NAND2_X1 U6388 ( .A1(n7660), .A2(n7705), .ZN(n4700) );
  NAND3_X1 U6389 ( .A1(n7661), .A2(n4700), .A3(n4699), .ZN(n7710) );
  NAND2_X1 U6390 ( .A1(n7710), .A2(n4700), .ZN(n7713) );
  NAND2_X1 U6391 ( .A1(n4701), .A2(n4702), .ZN(n7476) );
  NAND2_X1 U6392 ( .A1(n7415), .A2(n4704), .ZN(n4701) );
  MUX2_X1 U6393 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8947), .S(n7108), .Z(n7107)
         );
  AOI21_X1 U6394 ( .B1(n9489), .B2(n9490), .A(n9488), .ZN(n9494) );
  NAND3_X1 U6395 ( .A1(n7612), .A2(n6407), .A3(n9369), .ZN(n4715) );
  NOR2_X1 U6396 ( .A1(n7614), .A2(n7040), .ZN(n7613) );
  INV_X1 U6397 ( .A(n7820), .ZN(n7040) );
  MUX2_X1 U6398 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10190), .S(n6085), .Z(n7820)
         );
  NAND2_X2 U6399 ( .A1(n6397), .A2(n6848), .ZN(n6085) );
  NAND2_X1 U6400 ( .A1(n8268), .A2(n4459), .ZN(n4722) );
  OR2_X1 U6401 ( .A1(n7745), .A2(n4727), .ZN(n4726) );
  INV_X1 U6402 ( .A(n7693), .ZN(n4727) );
  NAND2_X1 U6403 ( .A1(n7753), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6404 ( .A1(n6282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U6405 ( .A1(n8237), .A2(n7075), .ZN(n4746) );
  NAND2_X1 U6406 ( .A1(n5788), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U6407 ( .A1(n5787), .A2(SI_29_), .ZN(n4753) );
  NAND2_X1 U6408 ( .A1(n5535), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6409 ( .A1(n5450), .A2(n4767), .ZN(n4764) );
  NAND2_X1 U6410 ( .A1(n5618), .A2(n4783), .ZN(n4776) );
  NAND2_X4 U6411 ( .A1(n4787), .A2(n4786), .ZN(n5249) );
  NAND3_X2 U6412 ( .A1(n5040), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4786) );
  INV_X1 U6413 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U6414 ( .A1(n5279), .A2(n5278), .ZN(n5298) );
  NAND2_X2 U6415 ( .A1(n5586), .A2(n5585), .ZN(n5618) );
  NAND2_X1 U6416 ( .A1(n5784), .A2(n5783), .ZN(n5788) );
  NAND2_X1 U6417 ( .A1(n5688), .A2(n5687), .ZN(n5784) );
  OAI21_X1 U6418 ( .B1(n5277), .B2(n5276), .A(n5275), .ZN(n5279) );
  OAI21_X2 U6419 ( .B1(n5574), .B2(n5573), .A(n5572), .ZN(n5584) );
  NAND2_X1 U6420 ( .A1(n5686), .A2(n5685), .ZN(n5688) );
  NAND4_X1 U6421 ( .A1(n4791), .A2(n4414), .A3(n8150), .A4(n4800), .ZN(n4792)
         );
  INV_X1 U6422 ( .A(n5902), .ZN(n4800) );
  NOR2_X1 U6423 ( .A1(n5914), .A2(n8870), .ZN(n4809) );
  NOR2_X1 U6424 ( .A1(n5487), .A2(n4819), .ZN(n7004) );
  MUX2_X1 U6425 ( .A(n9103), .B(P2_IR_REG_0__SCAN_IN), .S(n5487), .Z(n10381)
         );
  OAI22_X1 U6426 ( .A1(n8621), .A2(n4376), .B1(n5137), .B2(n6828), .ZN(n5415)
         );
  OAI22_X1 U6427 ( .A1(n10352), .A2(n4817), .B1(n5137), .B2(n6976), .ZN(n5468)
         );
  OAI21_X1 U6428 ( .B1(n10363), .B2(n6992), .A(n4817), .ZN(n6784) );
  NAND2_X1 U6429 ( .A1(n7005), .A2(n4376), .ZN(n6997) );
  NAND2_X1 U6430 ( .A1(n9374), .A2(n9557), .ZN(n9584) );
  INV_X1 U6431 ( .A(n6139), .ZN(n9645) );
  NAND2_X1 U6432 ( .A1(n4834), .A2(n4840), .ZN(n4833) );
  NAND2_X1 U6433 ( .A1(n4851), .A2(n4849), .ZN(n7912) );
  NAND2_X1 U6434 ( .A1(n9994), .A2(n4867), .ZN(n4865) );
  AOI21_X2 U6435 ( .B1(n9993), .B2(n9450), .A(n4872), .ZN(n4871) );
  NAND2_X1 U6436 ( .A1(n9159), .A2(n4386), .ZN(n4873) );
  NAND2_X2 U6437 ( .A1(n9901), .A2(n4874), .ZN(n9881) );
  NAND2_X1 U6438 ( .A1(n6409), .A2(n9588), .ZN(n4880) );
  NAND3_X1 U6439 ( .A1(n6409), .A2(n9588), .A3(n4878), .ZN(n4877) );
  NAND2_X1 U6440 ( .A1(n4881), .A2(n4879), .ZN(n7892) );
  INV_X1 U6441 ( .A(n7578), .ZN(n4892) );
  NAND2_X1 U6442 ( .A1(n4899), .A2(n4900), .ZN(n8172) );
  OAI21_X2 U6443 ( .B1(n8789), .B2(n4904), .A(n4903), .ZN(n8756) );
  AND2_X2 U6444 ( .A1(n7958), .A2(n4907), .ZN(n9982) );
  INV_X1 U6445 ( .A(n4912), .ZN(n9998) );
  NAND2_X1 U6446 ( .A1(n4913), .A2(n8013), .ZN(n7900) );
  AND2_X1 U6447 ( .A1(n4914), .A2(n4915), .ZN(n4913) );
  NOR2_X2 U6448 ( .A1(n7973), .A2(n7972), .ZN(n10265) );
  NOR2_X2 U6449 ( .A1(n9964), .A2(n4918), .ZN(n9890) );
  INV_X1 U6450 ( .A(n9760), .ZN(n9745) );
  NAND2_X1 U6451 ( .A1(n9815), .A2(n6422), .ZN(n9792) );
  NAND2_X1 U6452 ( .A1(n4934), .A2(n4931), .ZN(n8383) );
  OR2_X1 U6453 ( .A1(n8470), .A2(n8466), .ZN(n4930) );
  OAI21_X2 U6454 ( .B1(n5546), .B2(n4942), .A(n4940), .ZN(n5608) );
  INV_X1 U6455 ( .A(n5122), .ZN(n4943) );
  NAND2_X1 U6456 ( .A1(n7491), .A2(n4955), .ZN(n5213) );
  NAND3_X1 U6457 ( .A1(n7272), .A2(n5074), .A3(n5102), .ZN(n7561) );
  NAND2_X1 U6458 ( .A1(n5052), .A2(n5048), .ZN(n5050) );
  NAND2_X1 U6459 ( .A1(n5052), .A2(n4959), .ZN(n5692) );
  NAND2_X2 U6460 ( .A1(n8796), .A2(n4434), .ZN(n8732) );
  NAND3_X1 U6461 ( .A1(n7353), .A2(n7352), .A3(n7311), .ZN(n7327) );
  NAND3_X1 U6462 ( .A1(n7046), .A2(n7045), .A3(n7044), .ZN(n7049) );
  NAND2_X1 U6463 ( .A1(n4973), .A2(n10381), .ZN(n7044) );
  NAND2_X2 U6464 ( .A1(n7336), .A2(n7270), .ZN(n6809) );
  NAND2_X1 U6465 ( .A1(n8808), .A2(n8348), .ZN(n4974) );
  NAND2_X1 U6466 ( .A1(n7527), .A2(n7526), .ZN(n7577) );
  INV_X1 U6467 ( .A(n7526), .ZN(n4982) );
  NAND2_X1 U6468 ( .A1(n4989), .A2(n4988), .ZN(n4987) );
  INV_X1 U6469 ( .A(n8784), .ZN(n4989) );
  NOR2_X2 U6470 ( .A1(n8150), .A2(n4998), .ZN(n4997) );
  INV_X1 U6471 ( .A(n9407), .ZN(n9753) );
  NAND2_X2 U6472 ( .A1(n9572), .A2(n9393), .ZN(n9827) );
  AOI21_X1 U6473 ( .B1(n5815), .B2(n5814), .A(n5813), .ZN(n5818) );
  INV_X1 U6474 ( .A(n8815), .ZN(n8834) );
  CLKBUF_X1 U6475 ( .A(n7907), .Z(n7961) );
  XNOR2_X1 U6476 ( .A(n8650), .B(n8645), .ZN(n8954) );
  CLKBUF_X1 U6477 ( .A(n7804), .Z(n8126) );
  AND4_X4 U6478 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n7571)
         );
  INV_X1 U6479 ( .A(n6080), .ZN(n6091) );
  OAI211_X2 U6480 ( .C1(n5137), .C2(n4516), .A(n5121), .B(n5120), .ZN(n8927)
         );
  XNOR2_X1 U6481 ( .A(n5636), .B(n5635), .ZN(n8165) );
  XNOR2_X2 U6482 ( .A(n5064), .B(n5063), .ZN(n6770) );
  NOR2_X1 U6483 ( .A1(n8375), .A2(n6424), .ZN(n6425) );
  NAND2_X1 U6484 ( .A1(n6032), .A2(n8186), .ZN(n6080) );
  XNOR2_X1 U6485 ( .A(n5049), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5058) );
  NAND2_X2 U6486 ( .A1(n9647), .A2(n8015), .ZN(n9555) );
  AND2_X1 U6487 ( .A1(n5198), .A2(n5024), .ZN(n5025) );
  INV_X1 U6488 ( .A(n5223), .ZN(n5047) );
  NOR2_X1 U6489 ( .A1(n5608), .A2(n5607), .ZN(n8495) );
  INV_X1 U6490 ( .A(n5058), .ZN(n5988) );
  INV_X1 U6491 ( .A(n5799), .ZN(n5307) );
  INV_X4 U6492 ( .A(n5593), .ZN(n5663) );
  NAND2_X2 U6493 ( .A1(n7633), .A2(n9999), .ZN(n10036) );
  OR2_X1 U6494 ( .A1(n5826), .A2(n6815), .ZN(n5004) );
  OR2_X1 U6495 ( .A1(n6992), .A2(n6999), .ZN(n8793) );
  INV_X1 U6496 ( .A(n8804), .ZN(n5772) );
  AND2_X1 U6497 ( .A1(n6817), .A2(n6816), .ZN(n8868) );
  INV_X1 U6498 ( .A(n9962), .ZN(n6264) );
  INV_X1 U6499 ( .A(n8699), .ZN(n8329) );
  AND2_X1 U6500 ( .A1(n9860), .A2(n9886), .ZN(n5007) );
  INV_X1 U6501 ( .A(n9215), .ZN(n6361) );
  AND2_X1 U6502 ( .A1(n5299), .A2(n5284), .ZN(n5010) );
  OR2_X1 U6503 ( .A1(n9644), .A2(n10298), .ZN(n5012) );
  AND2_X1 U6504 ( .A1(n5956), .A2(n5950), .ZN(n5013) );
  INV_X1 U6505 ( .A(n6032), .ZN(n8366) );
  INV_X1 U6506 ( .A(n8692), .ZN(n8964) );
  OR2_X2 U6507 ( .A1(n8138), .A2(n9052), .ZN(n5014) );
  INV_X1 U6508 ( .A(n5963), .ZN(n5959) );
  NOR2_X1 U6509 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  INV_X1 U6510 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5015) );
  AND2_X1 U6511 ( .A1(n8652), .A2(n8327), .ZN(n5970) );
  INV_X1 U6512 ( .A(n9364), .ZN(n6057) );
  NOR2_X1 U6513 ( .A1(n4806), .A2(n5763), .ZN(n5764) );
  INV_X1 U6514 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6383) );
  INV_X1 U6515 ( .A(n10010), .ZN(n6412) );
  INV_X1 U6516 ( .A(n9884), .ZN(n6414) );
  NAND2_X1 U6517 ( .A1(n4416), .A2(n6280), .ZN(n6281) );
  INV_X1 U6518 ( .A(n7563), .ZN(n5102) );
  INV_X1 U6519 ( .A(n8514), .ZN(n5530) );
  INV_X1 U6520 ( .A(n8595), .ZN(n8354) );
  INV_X1 U6521 ( .A(n10418), .ZN(n8356) );
  AND3_X1 U6522 ( .A1(n5698), .A2(n5044), .A3(n5023), .ZN(n5024) );
  INV_X1 U6523 ( .A(n6247), .ZN(n6023) );
  INV_X1 U6524 ( .A(n9363), .ZN(n6406) );
  INV_X1 U6525 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6872) );
  AND2_X1 U6526 ( .A1(n9757), .A2(n10299), .ZN(n6423) );
  NAND2_X1 U6527 ( .A1(n9648), .A2(n10267), .ZN(n9371) );
  INV_X1 U6528 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6385) );
  INV_X1 U6529 ( .A(SI_20_), .ZN(n6523) );
  INV_X1 U6530 ( .A(n5323), .ZN(n5327) );
  OR2_X1 U6531 ( .A1(n8497), .A2(n8500), .ZN(n5611) );
  NOR2_X1 U6532 ( .A1(n8647), .A2(n8327), .ZN(n8328) );
  AND2_X1 U6533 ( .A1(n4375), .A2(n10423), .ZN(n8970) );
  OR2_X1 U6534 ( .A1(n5692), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n5693) );
  INV_X1 U6535 ( .A(n7755), .ZN(n7752) );
  INV_X1 U6536 ( .A(n8290), .ZN(n8291) );
  NAND2_X1 U6537 ( .A1(n7068), .A2(n7067), .ZN(n7166) );
  AND2_X1 U6538 ( .A1(n9124), .A2(n9220), .ZN(n9239) );
  INV_X1 U6539 ( .A(n8019), .ZN(n8015) );
  AND2_X1 U6540 ( .A1(n7286), .A2(n7033), .ZN(n6453) );
  NAND2_X1 U6541 ( .A1(n5553), .A2(n5552), .ZN(n5572) );
  AND2_X1 U6542 ( .A1(n7501), .A2(n5060), .ZN(n7274) );
  NAND2_X1 U6543 ( .A1(n5322), .A2(n5321), .ZN(n8452) );
  INV_X1 U6544 ( .A(n10363), .ZN(n7266) );
  OR2_X1 U6545 ( .A1(n8573), .A2(n8795), .ZN(n8537) );
  INV_X1 U6546 ( .A(n4393), .ZN(n5733) );
  INV_X1 U6547 ( .A(n5939), .ZN(n5774) );
  INV_X1 U6548 ( .A(n8905), .ZN(n8914) );
  AND2_X1 U6549 ( .A1(n10364), .A2(n10375), .ZN(n5708) );
  NOR2_X1 U6550 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  INV_X1 U6551 ( .A(n10398), .ZN(n10423) );
  NAND2_X1 U6552 ( .A1(n5693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5719) );
  AND2_X1 U6553 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  NAND2_X1 U6554 ( .A1(n7028), .A2(n7021), .ZN(n7068) );
  OR2_X1 U6555 ( .A1(n7031), .A2(n7023), .ZN(n7280) );
  INV_X1 U6556 ( .A(n9637), .ZN(n10015) );
  INV_X1 U6557 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6456) );
  AND2_X1 U6558 ( .A1(n9442), .A2(n9460), .ZN(n9595) );
  AND2_X1 U6559 ( .A1(n6405), .A2(n9548), .ZN(n10012) );
  OR2_X1 U6560 ( .A1(n7031), .A2(n9662), .ZN(n10016) );
  AND2_X1 U6561 ( .A1(n5656), .A2(n5640), .ZN(n5654) );
  XNOR2_X1 U6562 ( .A(n5482), .B(SI_18_), .ZN(n5479) );
  OR2_X1 U6563 ( .A1(n7983), .A2(n5718), .ZN(n6719) );
  NAND2_X1 U6564 ( .A1(n7266), .A2(n5721), .ZN(n8877) );
  AND2_X1 U6565 ( .A1(n5496), .A2(n5495), .ZN(n8509) );
  INV_X1 U6566 ( .A(n8637), .ZN(n10349) );
  AND2_X1 U6567 ( .A1(n7005), .A2(n7004), .ZN(n10355) );
  INV_X1 U6568 ( .A(n8793), .ZN(n8907) );
  INV_X1 U6569 ( .A(n8868), .ZN(n8902) );
  AND2_X1 U6570 ( .A1(n8945), .A2(n7324), .ZN(n8939) );
  NOR2_X1 U6571 ( .A1(n10374), .A2(n5708), .ZN(n7013) );
  AND2_X1 U6572 ( .A1(n8890), .A2(n10429), .ZN(n10418) );
  NOR2_X1 U6573 ( .A1(n6808), .A2(n6807), .ZN(n7014) );
  NAND2_X1 U6574 ( .A1(n6719), .A2(n10379), .ZN(n10363) );
  INV_X1 U6575 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5990) );
  AND2_X1 U6576 ( .A1(n6404), .A2(n6403), .ZN(n10051) );
  AND2_X1 U6577 ( .A1(n6279), .A2(n6278), .ZN(n9918) );
  INV_X1 U6578 ( .A(n10180), .ZN(n9662) );
  INV_X1 U6579 ( .A(n9735), .ZN(n10235) );
  INV_X1 U6580 ( .A(n10228), .ZN(n9733) );
  INV_X1 U6581 ( .A(n10239), .ZN(n9716) );
  INV_X1 U6582 ( .A(n10014), .ZN(n9936) );
  INV_X1 U6583 ( .A(n10028), .ZN(n10041) );
  NOR2_X1 U6584 ( .A1(n10344), .A2(n6456), .ZN(n6457) );
  NAND2_X1 U6585 ( .A1(n6455), .A2(n10172), .ZN(n7623) );
  INV_X1 U6586 ( .A(n10144), .ZN(n10325) );
  INV_X1 U6587 ( .A(n7623), .ZN(n7367) );
  INV_X1 U6588 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6429) );
  AND2_X1 U6589 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10206), .ZN(n10474) );
  INV_X1 U6590 ( .A(n8643), .ZN(n10347) );
  INV_X1 U6591 ( .A(n5749), .ZN(n5750) );
  INV_X1 U6592 ( .A(n8982), .ZN(n8748) );
  AND2_X1 U6593 ( .A1(n5722), .A2(n8877), .ZN(n8570) );
  AND2_X1 U6594 ( .A1(n5738), .A2(n5737), .ZN(n7511) );
  INV_X1 U6595 ( .A(n8538), .ZN(n8774) );
  INV_X1 U6596 ( .A(n10355), .ZN(n7719) );
  INV_X1 U6597 ( .A(n10354), .ZN(n8626) );
  INV_X1 U6598 ( .A(n8939), .ZN(n8920) );
  AND2_X1 U6599 ( .A1(n8911), .A2(n8910), .ZN(n9033) );
  NAND2_X1 U6600 ( .A1(n8945), .A2(n7319), .ZN(n8860) );
  INV_X1 U6601 ( .A(n10444), .ZN(n10441) );
  INV_X1 U6602 ( .A(n10433), .ZN(n10431) );
  NOR2_X1 U6603 ( .A1(n10364), .A2(n10363), .ZN(n10373) );
  AND2_X1 U6604 ( .A1(n7983), .A2(n9102), .ZN(n10374) );
  XNOR2_X1 U6605 ( .A(n5696), .B(n5695), .ZN(n7983) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7611) );
  INV_X1 U6607 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6782) );
  CLKBUF_X1 U6608 ( .A(n8378), .Z(n9099) );
  INV_X1 U6609 ( .A(n9305), .ZN(n9336) );
  INV_X1 U6610 ( .A(n9338), .ZN(n9298) );
  INV_X1 U6611 ( .A(n10051), .ZN(n10053) );
  INV_X1 U6612 ( .A(n9867), .ZN(n9825) );
  OR2_X1 U6613 ( .A1(n9734), .A2(n9662), .ZN(n10239) );
  OR2_X1 U6614 ( .A1(n9734), .A2(n10180), .ZN(n10228) );
  OR3_X1 U6615 ( .A1(n9655), .A2(n9652), .A3(n10180), .ZN(n9735) );
  INV_X1 U6616 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U6617 ( .A1(n10036), .A2(n7791), .ZN(n10028) );
  INV_X2 U6618 ( .A(n10341), .ZN(n10344) );
  OR2_X1 U6619 ( .A1(n7368), .A2(n7623), .ZN(n10341) );
  INV_X1 U6620 ( .A(n10326), .ZN(n10328) );
  INV_X1 U6621 ( .A(n10255), .ZN(n10254) );
  XNOR2_X1 U6622 ( .A(n6430), .B(n6429), .ZN(n7952) );
  INV_X1 U6623 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7490) );
  INV_X1 U6624 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6798) );
  INV_X1 U6625 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U6626 ( .B1(n10203), .B2(n6536), .A(n10202), .ZN(n10495) );
  NOR2_X1 U6627 ( .A1(n10472), .A2(n10471), .ZN(n10470) );
  OAI21_X1 U6628 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10461), .ZN(n10459) );
  AND2_X1 U6629 ( .A1(n6993), .A2(n10379), .ZN(P2_U3966) );
  INV_X2 U6630 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5407) );
  INV_X2 U6631 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5335) );
  INV_X2 U6632 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5467) );
  AND4_X2 U6633 ( .A1(n5407), .A2(n5335), .A3(n5015), .A4(n5467), .ZN(n5016)
         );
  NAND2_X1 U6634 ( .A1(n5017), .A2(n5016), .ZN(n5045) );
  INV_X1 U6635 ( .A(n5045), .ZN(n5022) );
  NOR2_X1 U6636 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5020) );
  NOR2_X1 U6637 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5019) );
  NOR2_X1 U6638 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5018) );
  INV_X2 U6639 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6682) );
  XNOR2_X2 U6640 ( .A(n5028), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5034) );
  OAI21_X1 U6641 ( .B1(n5029), .B2(n9088), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5031) );
  NAND2_X1 U6642 ( .A1(n5031), .A2(n5030), .ZN(n5033) );
  AND2_X4 U6643 ( .A1(n5035), .A2(n8367), .ZN(n5799) );
  NAND2_X1 U6644 ( .A1(n5799), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5039) );
  INV_X1 U6645 ( .A(n5035), .ZN(n8381) );
  NAND2_X1 U6646 ( .A1(n5128), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5038) );
  NAND2_X1 U6647 ( .A1(n5129), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6648 ( .A1(n5127), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5036) );
  INV_X2 U6649 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6650 ( .A1(n6727), .A2(SI_0_), .ZN(n5041) );
  XNOR2_X1 U6651 ( .A(n5041), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9103) );
  INV_X1 U6652 ( .A(n10381), .ZN(n7500) );
  NAND2_X1 U6653 ( .A1(n5198), .A2(n5044), .ZN(n5223) );
  NOR2_X1 U6654 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5048) );
  INV_X1 U6655 ( .A(n5720), .ZN(n10382) );
  INV_X1 U6656 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6657 ( .A1(n5057), .A2(n5053), .ZN(n5054) );
  NAND2_X1 U6658 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5056) );
  XNOR2_X2 U6659 ( .A(n5056), .B(n5055), .ZN(n7507) );
  AND2_X2 U6660 ( .A1(n10382), .A2(n5989), .ZN(n5826) );
  NAND2_X1 U6661 ( .A1(n6811), .A2(n5525), .ZN(n7501) );
  NAND2_X1 U6662 ( .A1(n7507), .A2(n5851), .ZN(n7318) );
  OR2_X1 U6663 ( .A1(n5643), .A2(n10381), .ZN(n5060) );
  AND2_X1 U6664 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6665 ( .A1(n4391), .A2(n5083), .ZN(n6045) );
  AND2_X1 U6666 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6667 ( .A1(n6727), .A2(n5079), .ZN(n5061) );
  NAND2_X1 U6668 ( .A1(n6045), .A2(n5061), .ZN(n5062) );
  INV_X1 U6669 ( .A(SI_1_), .ZN(n6478) );
  XNOR2_X1 U6670 ( .A(n5062), .B(n6478), .ZN(n5064) );
  MUX2_X1 U6671 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4391), .Z(n5063) );
  NAND2_X1 U6672 ( .A1(n5487), .A2(n7108), .ZN(n5065) );
  OAI211_X2 U6673 ( .C1(n5108), .C2(n6770), .A(n5066), .B(n5065), .ZN(n8938)
         );
  NAND2_X1 U6674 ( .A1(n4398), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6675 ( .A1(n5127), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6676 ( .A1(n5128), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6677 ( .A1(n5129), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5067) );
  AND4_X2 U6678 ( .A1(n5070), .A2(n5069), .A3(n5068), .A4(n5067), .ZN(n5752)
         );
  CLKBUF_X1 U6679 ( .A(n5752), .Z(n7560) );
  OR2_X1 U6680 ( .A1(n7560), .A2(n5826), .ZN(n5073) );
  XNOR2_X1 U6681 ( .A(n5071), .B(n5073), .ZN(n7273) );
  INV_X1 U6682 ( .A(n5071), .ZN(n5072) );
  NAND2_X1 U6683 ( .A1(n5073), .A2(n5072), .ZN(n5074) );
  NAND2_X1 U6684 ( .A1(n4398), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6685 ( .A1(n5129), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6686 ( .A1(n5127), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6687 ( .A1(n5128), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U6688 ( .A1(n5754), .A2(n5826), .ZN(n5098) );
  INV_X1 U6689 ( .A(n5079), .ZN(n5080) );
  NOR2_X1 U6690 ( .A1(n5080), .A2(n6478), .ZN(n5082) );
  INV_X1 U6691 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6754) );
  AOI21_X1 U6692 ( .B1(n6478), .B2(n5080), .A(n6754), .ZN(n5081) );
  OAI21_X1 U6693 ( .B1(n5082), .B2(n5081), .A(n4489), .ZN(n5089) );
  INV_X1 U6694 ( .A(n5083), .ZN(n5086) );
  INV_X1 U6695 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U6696 ( .A1(n5086), .A2(n6771), .ZN(n5084) );
  NAND2_X1 U6697 ( .A1(n5084), .A2(SI_1_), .ZN(n5085) );
  OAI21_X1 U6698 ( .B1(n5086), .B2(n6771), .A(n5085), .ZN(n5087) );
  NAND2_X1 U6699 ( .A1(n4391), .A2(n5087), .ZN(n5088) );
  NAND2_X1 U6700 ( .A1(n5089), .A2(n5088), .ZN(n5113) );
  INV_X1 U6701 ( .A(SI_2_), .ZN(n5110) );
  XNOR2_X1 U6702 ( .A(n5113), .B(n5110), .ZN(n5091) );
  MUX2_X1 U6703 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4392), .Z(n5090) );
  NAND2_X1 U6704 ( .A1(n4379), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5097) );
  INV_X1 U6705 ( .A(n5139), .ZN(n5093) );
  NAND2_X1 U6706 ( .A1(n5093), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6707 ( .A1(n5139), .A2(n5094), .ZN(n5118) );
  AND2_X1 U6708 ( .A1(n5095), .A2(n5118), .ZN(n7182) );
  NAND2_X1 U6709 ( .A1(n5487), .A2(n7182), .ZN(n5096) );
  OAI211_X2 U6710 ( .C1(n5108), .C2(n6768), .A(n5097), .B(n5096), .ZN(n10391)
         );
  XNOR2_X1 U6711 ( .A(n5643), .B(n10391), .ZN(n5099) );
  NAND2_X1 U6712 ( .A1(n5098), .A2(n5099), .ZN(n5103) );
  INV_X1 U6713 ( .A(n5098), .ZN(n5100) );
  INV_X1 U6714 ( .A(n5099), .ZN(n8412) );
  NAND2_X1 U6715 ( .A1(n5100), .A2(n8412), .ZN(n5101) );
  NAND2_X1 U6716 ( .A1(n5103), .A2(n5101), .ZN(n7563) );
  NAND2_X1 U6717 ( .A1(n7561), .A2(n5103), .ZN(n5122) );
  NAND2_X1 U6718 ( .A1(n5799), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6719 ( .A1(n5129), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6720 ( .A1(n5128), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6721 ( .A1(n5127), .A2(n8930), .ZN(n5104) );
  AND4_X2 U6722 ( .A1(n5107), .A2(n5106), .A3(n5105), .A4(n5104), .ZN(n7517)
         );
  OR2_X1 U6723 ( .A1(n7517), .A2(n5826), .ZN(n5123) );
  INV_X2 U6724 ( .A(n5108), .ZN(n5177) );
  INV_X1 U6725 ( .A(SI_3_), .ZN(n5109) );
  INV_X1 U6726 ( .A(n5135), .ZN(n5117) );
  INV_X1 U6727 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U6728 ( .A1(n4392), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5111) );
  OAI211_X1 U6729 ( .C1(n4397), .C2(n6752), .A(n5111), .B(n5110), .ZN(n5112)
         );
  NAND2_X1 U6730 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  INV_X1 U6731 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6769) );
  NAND2_X1 U6732 ( .A1(n4397), .A2(n6769), .ZN(n5114) );
  OAI211_X1 U6733 ( .C1(n4392), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5114), .B(
        SI_2_), .ZN(n5115) );
  XNOR2_X1 U6734 ( .A(n5134), .B(n5117), .ZN(n6730) );
  NAND2_X1 U6735 ( .A1(n5118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6736 ( .A1(n5487), .A2(n7131), .ZN(n5120) );
  XNOR2_X1 U6737 ( .A(n5643), .B(n8927), .ZN(n5124) );
  XNOR2_X1 U6738 ( .A(n5123), .B(n5124), .ZN(n8413) );
  INV_X1 U6739 ( .A(n5123), .ZN(n5125) );
  NAND2_X1 U6740 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  NAND2_X1 U6741 ( .A1(n5799), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5133) );
  OAI21_X1 U6742 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5147), .ZN(n7329) );
  INV_X1 U6743 ( .A(n7329), .ZN(n7520) );
  NAND2_X1 U6744 ( .A1(n4393), .A2(n7520), .ZN(n5132) );
  NAND2_X1 U6745 ( .A1(n5663), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U6746 ( .A1(n5289), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5130) );
  AND4_X2 U6747 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n7525)
         );
  OR2_X1 U6748 ( .A1(n7525), .A2(n5826), .ZN(n5144) );
  NAND2_X1 U6749 ( .A1(n5136), .A2(SI_3_), .ZN(n5167) );
  NAND2_X1 U6750 ( .A1(n5168), .A2(n5167), .ZN(n5155) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4396), .Z(n5169) );
  XNOR2_X1 U6752 ( .A(n5169), .B(SI_4_), .ZN(n5153) );
  XNOR2_X1 U6753 ( .A(n5155), .B(n5153), .ZN(n6725) );
  NAND2_X1 U6754 ( .A1(n6725), .A2(n5177), .ZN(n5143) );
  OAI21_X1 U6755 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(P2_IR_REG_3__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6756 ( .A1(n5139), .A2(n5138), .ZN(n5141) );
  INV_X1 U6757 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5140) );
  XNOR2_X1 U6758 ( .A(n5141), .B(n5140), .ZN(n7195) );
  AOI22_X1 U6759 ( .A1(n4394), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n5487), .B2(
        n7195), .ZN(n5142) );
  NAND2_X1 U6760 ( .A1(n5143), .A2(n5142), .ZN(n7331) );
  INV_X2 U6761 ( .A(n7331), .ZN(n10399) );
  XNOR2_X1 U6762 ( .A(n5643), .B(n10399), .ZN(n7521) );
  NAND2_X1 U6763 ( .A1(n5144), .A2(n7521), .ZN(n7514) );
  NAND2_X1 U6764 ( .A1(n5799), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5152) );
  INV_X1 U6765 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6766 ( .A1(n5147), .A2(n5146), .ZN(n5148) );
  AND2_X1 U6767 ( .A1(n5182), .A2(n5148), .ZN(n7391) );
  NAND2_X1 U6768 ( .A1(n4393), .A2(n7391), .ZN(n5151) );
  NAND2_X1 U6769 ( .A1(n5663), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6770 ( .A1(n5289), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5149) );
  OR2_X1 U6771 ( .A1(n7571), .A2(n5826), .ZN(n5161) );
  INV_X1 U6772 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6773 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6774 ( .A1(n5156), .A2(n5166), .ZN(n5157) );
  XNOR2_X1 U6775 ( .A(n5174), .B(SI_5_), .ZN(n5171) );
  XNOR2_X1 U6776 ( .A(n5157), .B(n5171), .ZN(n6732) );
  NAND2_X1 U6777 ( .A1(n5158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5159) );
  XNOR2_X1 U6778 ( .A(n5159), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7150) );
  AOI22_X1 U6779 ( .A1(n4394), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5487), .B2(
        n7150), .ZN(n5160) );
  XNOR2_X1 U6780 ( .A(n5643), .B(n7570), .ZN(n5162) );
  XNOR2_X1 U6781 ( .A(n5161), .B(n5162), .ZN(n7390) );
  INV_X1 U6782 ( .A(n5161), .ZN(n5164) );
  INV_X1 U6783 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6784 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NOR2_X1 U6785 ( .A1(n5169), .A2(SI_4_), .ZN(n5170) );
  NOR2_X1 U6786 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  NAND2_X1 U6787 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
  NAND2_X1 U6788 ( .A1(n5174), .A2(SI_5_), .ZN(n5175) );
  MUX2_X1 U6789 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4391), .Z(n5197) );
  XNOR2_X1 U6790 ( .A(n5197), .B(SI_6_), .ZN(n5194) );
  XNOR2_X1 U6791 ( .A(n5196), .B(n5194), .ZN(n6723) );
  NAND2_X1 U6792 ( .A1(n6723), .A2(n5819), .ZN(n5181) );
  OR2_X1 U6793 ( .A1(n5158), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6794 ( .A1(n5178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6795 ( .A(n5179), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7242) );
  AOI22_X1 U6796 ( .A1(n4394), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5487), .B2(
        n7242), .ZN(n5180) );
  XNOR2_X1 U6797 ( .A(n10414), .B(n5643), .ZN(n5188) );
  NAND2_X1 U6798 ( .A1(n5799), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6799 ( .A1(n5182), .A2(n4527), .ZN(n5183) );
  AND2_X1 U6800 ( .A1(n5202), .A2(n5183), .ZN(n7540) );
  NAND2_X1 U6801 ( .A1(n4393), .A2(n7540), .ZN(n5186) );
  NAND2_X1 U6802 ( .A1(n5289), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6803 ( .A1(n5663), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5184) );
  NAND4_X1 U6804 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n8606)
         );
  AND2_X1 U6805 ( .A1(n5525), .A2(n8606), .ZN(n5189) );
  NAND2_X1 U6806 ( .A1(n5188), .A2(n5189), .ZN(n5192) );
  INV_X1 U6807 ( .A(n5188), .ZN(n5191) );
  INV_X1 U6808 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6809 ( .A1(n5191), .A2(n5190), .ZN(n5193) );
  AND2_X1 U6810 ( .A1(n5192), .A2(n5193), .ZN(n7493) );
  INV_X1 U6811 ( .A(n5194), .ZN(n5195) );
  NAND2_X1 U6812 ( .A1(n5197), .A2(SI_6_), .ZN(n5240) );
  NAND2_X1 U6813 ( .A1(n5277), .A2(n5240), .ZN(n5216) );
  XNOR2_X1 U6814 ( .A(n5238), .B(SI_7_), .ZN(n5214) );
  NAND2_X1 U6815 ( .A1(n6734), .A2(n5819), .ZN(n5201) );
  OR2_X1 U6816 ( .A1(n5198), .A2(n9088), .ZN(n5199) );
  XNOR2_X1 U6817 ( .A(n5199), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7210) );
  AOI22_X1 U6818 ( .A1(n4394), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5487), .B2(
        n7210), .ZN(n5200) );
  XNOR2_X1 U6819 ( .A(n7669), .B(n5683), .ZN(n5209) );
  NAND2_X1 U6820 ( .A1(n5799), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6821 ( .A1(n5202), .A2(n4529), .ZN(n5203) );
  AND2_X1 U6822 ( .A1(n5228), .A2(n5203), .ZN(n7595) );
  NAND2_X1 U6823 ( .A1(n4393), .A2(n7595), .ZN(n5206) );
  NAND2_X1 U6824 ( .A1(n5289), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6825 ( .A1(n5663), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5204) );
  OR2_X1 U6826 ( .A1(n7839), .A2(n5826), .ZN(n5208) );
  XNOR2_X1 U6827 ( .A(n5209), .B(n5208), .ZN(n7588) );
  INV_X1 U6828 ( .A(n5208), .ZN(n5211) );
  INV_X1 U6829 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6830 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6831 ( .A1(n5213), .A2(n5212), .ZN(n7835) );
  INV_X1 U6832 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6833 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6834 ( .A1(n5238), .A2(SI_7_), .ZN(n5242) );
  NAND2_X1 U6835 ( .A1(n5217), .A2(n5242), .ZN(n5222) );
  INV_X1 U6836 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6751) );
  INV_X1 U6837 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6737) );
  MUX2_X1 U6838 ( .A(n6751), .B(n6737), .S(n4396), .Z(n5219) );
  INV_X1 U6839 ( .A(SI_8_), .ZN(n5218) );
  INV_X1 U6840 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6841 ( .A1(n5220), .A2(SI_8_), .ZN(n5221) );
  NAND2_X1 U6842 ( .A1(n5273), .A2(n5221), .ZN(n5244) );
  XNOR2_X1 U6843 ( .A(n5222), .B(n5244), .ZN(n6736) );
  NAND2_X1 U6844 ( .A1(n6736), .A2(n5819), .ZN(n5226) );
  NAND2_X1 U6845 ( .A1(n5223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5224) );
  XNOR2_X1 U6846 ( .A(n5224), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7224) );
  AOI22_X1 U6847 ( .A1(n4394), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5487), .B2(
        n7224), .ZN(n5225) );
  XNOR2_X1 U6848 ( .A(n4523), .B(n5643), .ZN(n5236) );
  NAND2_X1 U6849 ( .A1(n5799), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6850 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  AND2_X1 U6851 ( .A1(n5259), .A2(n5229), .ZN(n7685) );
  NAND2_X1 U6852 ( .A1(n4393), .A2(n7685), .ZN(n5232) );
  NAND2_X1 U6853 ( .A1(n5289), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6854 ( .A1(n5128), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6855 ( .A1(n5525), .A2(n8604), .ZN(n5234) );
  XNOR2_X1 U6856 ( .A(n5236), .B(n5234), .ZN(n7836) );
  INV_X1 U6857 ( .A(n5234), .ZN(n5235) );
  AND2_X1 U6858 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  INV_X1 U6859 ( .A(n5238), .ZN(n5239) );
  INV_X1 U6860 ( .A(SI_7_), .ZN(n6477) );
  NAND2_X1 U6861 ( .A1(n5239), .A2(n6477), .ZN(n5271) );
  INV_X1 U6862 ( .A(n5271), .ZN(n5247) );
  INV_X1 U6863 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U6864 ( .A1(n5241), .A2(n5271), .ZN(n5243) );
  INV_X1 U6865 ( .A(n5244), .ZN(n5245) );
  INV_X1 U6866 ( .A(n5274), .ZN(n5246) );
  OAI21_X1 U6867 ( .B1(n5277), .B2(n5247), .A(n5246), .ZN(n5248) );
  NAND2_X1 U6868 ( .A1(n5248), .A2(n5273), .ZN(n5255) );
  INV_X1 U6869 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6757) );
  INV_X1 U6870 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6765) );
  MUX2_X1 U6871 ( .A(n6757), .B(n6765), .S(n4397), .Z(n5251) );
  INV_X1 U6872 ( .A(SI_9_), .ZN(n5250) );
  NAND2_X1 U6873 ( .A1(n5251), .A2(n5250), .ZN(n5278) );
  INV_X1 U6874 ( .A(n5251), .ZN(n5252) );
  NAND2_X1 U6875 ( .A1(n5252), .A2(SI_9_), .ZN(n5253) );
  NAND2_X1 U6876 ( .A1(n5278), .A2(n5253), .ZN(n5272) );
  INV_X1 U6877 ( .A(n5272), .ZN(n5254) );
  XNOR2_X1 U6878 ( .A(n5255), .B(n5254), .ZN(n6756) );
  NAND2_X1 U6879 ( .A1(n6756), .A2(n5819), .ZN(n5257) );
  NAND2_X1 U6880 ( .A1(n5337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6881 ( .A(n5285), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7424) );
  AOI22_X1 U6882 ( .A1(n4394), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5487), .B2(
        n7424), .ZN(n5256) );
  XNOR2_X1 U6883 ( .A(n9061), .B(n5683), .ZN(n5265) );
  NAND2_X1 U6884 ( .A1(n5799), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5264) );
  INV_X1 U6885 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U6886 ( .A1(n5259), .A2(n6599), .ZN(n5260) );
  AND2_X1 U6887 ( .A1(n5311), .A2(n5260), .ZN(n7814) );
  NAND2_X1 U6888 ( .A1(n4393), .A2(n7814), .ZN(n5263) );
  NAND2_X1 U6889 ( .A1(n5663), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6890 ( .A1(n4390), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5261) );
  AND4_X2 U6891 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n8132)
         );
  OR2_X1 U6892 ( .A1(n8132), .A2(n5826), .ZN(n5266) );
  NAND2_X1 U6893 ( .A1(n5265), .A2(n5266), .ZN(n5270) );
  INV_X1 U6894 ( .A(n5265), .ZN(n5268) );
  INV_X1 U6895 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6896 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  AND2_X1 U6897 ( .A1(n5270), .A2(n5269), .ZN(n7862) );
  NAND2_X1 U6898 ( .A1(n5271), .A2(n5273), .ZN(n5276) );
  AOI21_X1 U6899 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5275) );
  MUX2_X1 U6900 ( .A(n5280), .B(n6767), .S(n4392), .Z(n5282) );
  INV_X1 U6901 ( .A(SI_10_), .ZN(n5281) );
  NAND2_X1 U6902 ( .A1(n5282), .A2(n5281), .ZN(n5299) );
  INV_X1 U6903 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6904 ( .A1(n5283), .A2(SI_10_), .ZN(n5284) );
  XNOR2_X1 U6905 ( .A(n5298), .B(n5010), .ZN(n6738) );
  NAND2_X1 U6906 ( .A1(n6738), .A2(n5819), .ZN(n5288) );
  NAND2_X1 U6907 ( .A1(n5285), .A2(n5335), .ZN(n5286) );
  NAND2_X1 U6908 ( .A1(n5286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6909 ( .A(n5302), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7255) );
  AOI22_X1 U6910 ( .A1(n7255), .A2(n5487), .B1(n4394), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5287) );
  XNOR2_X1 U6911 ( .A(n8142), .B(n5643), .ZN(n5294) );
  NAND2_X1 U6912 ( .A1(n5799), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5293) );
  XNOR2_X1 U6913 ( .A(n5311), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U6914 ( .A1(n4393), .A2(n8040), .ZN(n5292) );
  NAND2_X1 U6915 ( .A1(n5663), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6916 ( .A1(n5289), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5290) );
  NAND4_X1 U6917 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n8602)
         );
  NAND2_X1 U6918 ( .A1(n5525), .A2(n8602), .ZN(n5295) );
  XNOR2_X1 U6919 ( .A(n5294), .B(n5295), .ZN(n8037) );
  INV_X1 U6920 ( .A(n5294), .ZN(n5297) );
  INV_X1 U6921 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6922 ( .A1(n5298), .A2(n5010), .ZN(n5300) );
  INV_X1 U6923 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5301) );
  MUX2_X1 U6924 ( .A(n6749), .B(n5301), .S(n4397), .Z(n5324) );
  NAND2_X1 U6925 ( .A1(n6746), .A2(n5819), .ZN(n5306) );
  INV_X1 U6926 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6927 ( .A1(n5302), .A2(n5334), .ZN(n5303) );
  NAND2_X1 U6928 ( .A1(n5303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5304) );
  XNOR2_X1 U6929 ( .A(n5304), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7410) );
  AOI22_X1 U6930 ( .A1(n7410), .A2(n5487), .B1(n4394), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6931 ( .A(n9052), .B(n5683), .ZN(n5318) );
  NAND2_X1 U6932 ( .A1(n5799), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5317) );
  INV_X1 U6933 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5309) );
  INV_X1 U6934 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5308) );
  OAI21_X1 U6935 ( .B1(n5311), .B2(n5309), .A(n5308), .ZN(n5312) );
  NAND2_X1 U6936 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5310) );
  AND2_X1 U6937 ( .A1(n5312), .A2(n5342), .ZN(n8551) );
  NAND2_X1 U6938 ( .A1(n4393), .A2(n8551), .ZN(n5316) );
  NAND2_X1 U6939 ( .A1(n4390), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6940 ( .A1(n5663), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U6941 ( .A1(n8455), .A2(n5826), .ZN(n5319) );
  XNOR2_X1 U6942 ( .A(n5318), .B(n5319), .ZN(n8545) );
  INV_X1 U6943 ( .A(n5318), .ZN(n5320) );
  NAND2_X1 U6944 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  INV_X1 U6945 ( .A(n5324), .ZN(n5325) );
  NAND2_X1 U6946 ( .A1(n5325), .A2(SI_11_), .ZN(n5326) );
  MUX2_X1 U6947 ( .A(n6775), .B(n6773), .S(n4391), .Z(n5330) );
  INV_X1 U6948 ( .A(SI_12_), .ZN(n5329) );
  INV_X1 U6949 ( .A(n5330), .ZN(n5331) );
  NAND2_X1 U6950 ( .A1(n5331), .A2(SI_12_), .ZN(n5332) );
  NAND2_X1 U6951 ( .A1(n6772), .A2(n5177), .ZN(n5340) );
  INV_X1 U6952 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5333) );
  NAND3_X1 U6953 ( .A1(n5335), .A2(n5334), .A3(n5333), .ZN(n5336) );
  NOR2_X1 U6954 ( .A1(n5337), .A2(n5336), .ZN(n5362) );
  OR2_X1 U6955 ( .A1(n5362), .A2(n9088), .ZN(n5338) );
  XNOR2_X1 U6956 ( .A(n5338), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7451) );
  AOI22_X1 U6957 ( .A1(n7451), .A2(n5487), .B1(n4394), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U6958 ( .A(n9046), .B(n5683), .ZN(n5348) );
  NAND2_X1 U6959 ( .A1(n5799), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5347) );
  INV_X1 U6960 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U6961 ( .A1(n5342), .A2(n8454), .ZN(n5343) );
  AND2_X1 U6962 ( .A1(n5365), .A2(n5343), .ZN(n8456) );
  NAND2_X1 U6963 ( .A1(n4393), .A2(n8456), .ZN(n5346) );
  NAND2_X1 U6964 ( .A1(n4389), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6965 ( .A1(n5663), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6966 ( .A1(n8153), .A2(n5826), .ZN(n5349) );
  NAND2_X1 U6967 ( .A1(n5348), .A2(n5349), .ZN(n8450) );
  NAND2_X1 U6968 ( .A1(n8452), .A2(n8450), .ZN(n5352) );
  INV_X1 U6969 ( .A(n5348), .ZN(n5351) );
  INV_X1 U6970 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6971 ( .A1(n5351), .A2(n5350), .ZN(n8451) );
  NAND2_X1 U6972 ( .A1(n5352), .A2(n8451), .ZN(n8519) );
  INV_X1 U6973 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5357) );
  MUX2_X1 U6974 ( .A(n6782), .B(n5357), .S(n4391), .Z(n5358) );
  INV_X1 U6975 ( .A(n5358), .ZN(n5359) );
  NAND2_X1 U6976 ( .A1(n5359), .A2(SI_13_), .ZN(n5360) );
  NAND2_X1 U6977 ( .A1(n6779), .A2(n5177), .ZN(n5364) );
  INV_X1 U6978 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6979 ( .A1(n5362), .A2(n5361), .ZN(n5409) );
  NAND2_X1 U6980 ( .A1(n5409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U6981 ( .A(n5377), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7458) );
  AOI22_X1 U6982 ( .A1(n7458), .A2(n5487), .B1(n4379), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5363) );
  XNOR2_X1 U6983 ( .A(n8180), .B(n5643), .ZN(n5371) );
  NAND2_X1 U6984 ( .A1(n5799), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6985 ( .A1(n5365), .A2(n8522), .ZN(n5366) );
  AND2_X1 U6986 ( .A1(n5381), .A2(n5366), .ZN(n8525) );
  NAND2_X1 U6987 ( .A1(n4393), .A2(n8525), .ZN(n5369) );
  NAND2_X1 U6988 ( .A1(n4389), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6989 ( .A1(n5663), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5367) );
  NOR2_X1 U6990 ( .A1(n8458), .A2(n5826), .ZN(n5372) );
  NAND2_X1 U6991 ( .A1(n5371), .A2(n5372), .ZN(n5387) );
  INV_X1 U6992 ( .A(n5371), .ZN(n8390) );
  INV_X1 U6993 ( .A(n5372), .ZN(n5373) );
  NAND2_X1 U6994 ( .A1(n8390), .A2(n5373), .ZN(n5374) );
  AND2_X1 U6995 ( .A1(n5387), .A2(n5374), .ZN(n8520) );
  NAND2_X1 U6996 ( .A1(n8519), .A2(n8520), .ZN(n8518) );
  MUX2_X1 U6997 ( .A(n6794), .B(n6796), .S(n4392), .Z(n5394) );
  XNOR2_X1 U6998 ( .A(n5396), .B(n5393), .ZN(n6793) );
  NAND2_X1 U6999 ( .A1(n6793), .A2(n5177), .ZN(n5380) );
  NAND2_X1 U7000 ( .A1(n5377), .A2(n5407), .ZN(n5378) );
  NAND2_X1 U7001 ( .A1(n5378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U7002 ( .A(n5436), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7657) );
  AOI22_X1 U7003 ( .A1(n7657), .A2(n5487), .B1(n4379), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5379) );
  XNOR2_X1 U7004 ( .A(n9035), .B(n5683), .ZN(n5391) );
  NAND2_X1 U7005 ( .A1(n5799), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U7006 ( .A1(n5381), .A2(n8394), .ZN(n5382) );
  AND2_X1 U7007 ( .A1(n5426), .A2(n5382), .ZN(n8395) );
  NAND2_X1 U7008 ( .A1(n4393), .A2(n8395), .ZN(n5385) );
  NAND2_X1 U7009 ( .A1(n4389), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U7010 ( .A1(n5663), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5383) );
  NOR2_X1 U7011 ( .A1(n8335), .A2(n5826), .ZN(n5389) );
  XNOR2_X1 U7012 ( .A(n5391), .B(n5389), .ZN(n8402) );
  AND2_X1 U7013 ( .A1(n8402), .A2(n5387), .ZN(n5388) );
  INV_X1 U7014 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U7015 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  INV_X1 U7016 ( .A(n5394), .ZN(n5395) );
  MUX2_X1 U7017 ( .A(n6800), .B(n6798), .S(n4397), .Z(n5398) );
  INV_X1 U7018 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U7019 ( .A1(n5399), .A2(SI_15_), .ZN(n5400) );
  INV_X1 U7020 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5402) );
  MUX2_X1 U7021 ( .A(n6828), .B(n5402), .S(n4397), .Z(n5404) );
  INV_X1 U7022 ( .A(SI_16_), .ZN(n5403) );
  INV_X1 U7023 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U7024 ( .A1(n5405), .A2(SI_16_), .ZN(n5406) );
  NAND2_X1 U7025 ( .A1(n6802), .A2(n5177), .ZN(n5417) );
  INV_X1 U7026 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U7027 ( .A1(n5407), .A2(n5435), .ZN(n5408) );
  NAND2_X1 U7028 ( .A1(n5411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5410) );
  INV_X1 U7029 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5412) );
  MUX2_X1 U7030 ( .A(n5410), .B(P2_IR_REG_31__SCAN_IN), .S(n5412), .Z(n5414)
         );
  INV_X1 U7031 ( .A(n5411), .ZN(n5413) );
  NAND2_X1 U7032 ( .A1(n5413), .A2(n5412), .ZN(n5465) );
  NAND2_X1 U7033 ( .A1(n5414), .A2(n5465), .ZN(n8621) );
  INV_X1 U7034 ( .A(n5415), .ZN(n5416) );
  XNOR2_X1 U7035 ( .A(n9024), .B(n5643), .ZN(n8477) );
  NAND2_X1 U7036 ( .A1(n5799), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U7037 ( .A1(n4389), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5418) );
  AND2_X1 U7038 ( .A1(n5419), .A2(n5418), .ZN(n5424) );
  INV_X1 U7039 ( .A(n5420), .ZN(n5428) );
  INV_X1 U7040 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U7041 ( .A1(n5428), .A2(n8480), .ZN(n5421) );
  NAND2_X1 U7042 ( .A1(n5472), .A2(n5421), .ZN(n8894) );
  OR2_X1 U7043 ( .A1(n5733), .A2(n8894), .ZN(n5423) );
  NAND2_X1 U7044 ( .A1(n5663), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5422) );
  NOR2_X1 U7045 ( .A1(n8487), .A2(n5826), .ZN(n5442) );
  NAND2_X1 U7046 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  AND2_X1 U7047 ( .A1(n5428), .A2(n5427), .ZN(n8917) );
  NAND2_X1 U7048 ( .A1(n8917), .A2(n4393), .ZN(n5432) );
  NAND2_X1 U7049 ( .A1(n5799), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7050 ( .A1(n4389), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7051 ( .A1(n5663), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5429) );
  NOR2_X1 U7052 ( .A1(n8481), .A2(n5826), .ZN(n5443) );
  XNOR2_X1 U7053 ( .A(n5434), .B(n5433), .ZN(n6797) );
  NAND2_X1 U7054 ( .A1(n6797), .A2(n5177), .ZN(n5440) );
  NAND2_X1 U7055 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NAND2_X1 U7056 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U7057 ( .A(n5438), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7666) );
  AOI22_X1 U7058 ( .A1(n7666), .A2(n5487), .B1(n4394), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U7059 ( .A(n9030), .B(n5643), .ZN(n8473) );
  AOI22_X1 U7060 ( .A1(n8477), .A2(n5442), .B1(n5443), .B2(n8473), .ZN(n5441)
         );
  INV_X1 U7061 ( .A(n8477), .ZN(n5446) );
  OAI21_X1 U7062 ( .B1(n8473), .B2(n5443), .A(n5442), .ZN(n5445) );
  INV_X1 U7063 ( .A(n8473), .ZN(n8475) );
  INV_X1 U7064 ( .A(n5442), .ZN(n8476) );
  INV_X1 U7065 ( .A(n5443), .ZN(n8582) );
  AND2_X1 U7066 ( .A1(n8476), .A2(n8582), .ZN(n5444) );
  AOI22_X1 U7067 ( .A1(n5446), .A2(n5445), .B1(n8475), .B2(n5444), .ZN(n5447)
         );
  MUX2_X1 U7068 ( .A(n6976), .B(n6991), .S(n4397), .Z(n5451) );
  INV_X1 U7069 ( .A(n5451), .ZN(n5452) );
  NAND2_X1 U7070 ( .A1(n5452), .A2(SI_17_), .ZN(n5453) );
  MUX2_X1 U7071 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4392), .Z(n5482) );
  XNOR2_X1 U7072 ( .A(n5481), .B(n5479), .ZN(n7091) );
  NAND2_X1 U7073 ( .A1(n7091), .A2(n5177), .ZN(n5458) );
  NAND2_X1 U7074 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  XNOR2_X1 U7075 ( .A(n5456), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8627) );
  AOI22_X1 U7076 ( .A1(n4395), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5487), .B2(
        n8627), .ZN(n5457) );
  XNOR2_X1 U7077 ( .A(n9014), .B(n5683), .ZN(n5497) );
  INV_X1 U7078 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5471) );
  INV_X1 U7079 ( .A(n5474), .ZN(n5459) );
  NAND2_X1 U7080 ( .A1(n5474), .A2(n4537), .ZN(n5460) );
  NAND2_X1 U7081 ( .A1(n5490), .A2(n5460), .ZN(n8854) );
  OR2_X1 U7082 ( .A1(n8854), .A2(n5733), .ZN(n5463) );
  AOI22_X1 U7083 ( .A1(n5799), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n4389), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7084 ( .A1(n5663), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7085 ( .A1(n8598), .A2(n5525), .ZN(n5498) );
  AND2_X1 U7086 ( .A1(n5497), .A2(n5498), .ZN(n5500) );
  NAND2_X1 U7087 ( .A1(n6975), .A2(n5819), .ZN(n5470) );
  NAND2_X1 U7088 ( .A1(n5465), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5466) );
  XNOR2_X1 U7089 ( .A(n5467), .B(n5466), .ZN(n10352) );
  INV_X1 U7090 ( .A(n5468), .ZN(n5469) );
  XNOR2_X1 U7091 ( .A(n9020), .B(n5683), .ZN(n8560) );
  NAND2_X1 U7092 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  AND2_X1 U7093 ( .A1(n5474), .A2(n5473), .ZN(n8486) );
  NAND2_X1 U7094 ( .A1(n8486), .A2(n4393), .ZN(n5477) );
  AOI22_X1 U7095 ( .A1(n5799), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n4389), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7096 ( .A1(n5663), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5475) );
  OR2_X1 U7097 ( .A1(n8566), .A2(n5826), .ZN(n5501) );
  AND2_X1 U7098 ( .A1(n8560), .A2(n5501), .ZN(n8423) );
  MUX2_X1 U7099 ( .A(n7308), .B(n7310), .S(n4397), .Z(n5484) );
  INV_X1 U7100 ( .A(SI_19_), .ZN(n5483) );
  INV_X1 U7101 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U7102 ( .A1(n5485), .A2(SI_19_), .ZN(n5486) );
  NAND2_X1 U7103 ( .A1(n5510), .A2(n5486), .ZN(n5511) );
  XNOR2_X1 U7104 ( .A(n5512), .B(n5511), .ZN(n7307) );
  NAND2_X1 U7105 ( .A1(n7307), .A2(n5819), .ZN(n5489) );
  AOI22_X1 U7106 ( .A1(n8640), .A2(n5487), .B1(n4395), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5488) );
  XNOR2_X1 U7107 ( .A(n8837), .B(n5683), .ZN(n5508) );
  INV_X1 U7108 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U7109 ( .A1(n5490), .A2(n8432), .ZN(n5491) );
  AND2_X1 U7110 ( .A1(n5518), .A2(n5491), .ZN(n8836) );
  NAND2_X1 U7111 ( .A1(n8836), .A2(n4393), .ZN(n5496) );
  INV_X1 U7112 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U7113 ( .A1(n5799), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7114 ( .A1(n5663), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7115 ( .C1(n5313), .C2(n6565), .A(n5493), .B(n5492), .ZN(n5494)
         );
  INV_X1 U7116 ( .A(n5494), .ZN(n5495) );
  NOR2_X1 U7117 ( .A1(n8509), .A2(n5826), .ZN(n5506) );
  XNOR2_X1 U7118 ( .A(n5508), .B(n5506), .ZN(n8429) );
  INV_X1 U7119 ( .A(n5497), .ZN(n8427) );
  INV_X1 U7120 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7121 ( .A1(n8427), .A2(n5499), .ZN(n8424) );
  INV_X1 U7122 ( .A(n5500), .ZN(n8425) );
  INV_X1 U7123 ( .A(n8560), .ZN(n5503) );
  INV_X1 U7124 ( .A(n5501), .ZN(n5502) );
  AND2_X1 U7125 ( .A1(n5503), .A2(n5502), .ZN(n8426) );
  NAND2_X1 U7126 ( .A1(n8425), .A2(n8426), .ZN(n5504) );
  AND3_X1 U7127 ( .A1(n8429), .A2(n8424), .A3(n5504), .ZN(n5505) );
  INV_X1 U7128 ( .A(n5506), .ZN(n5507) );
  NAND2_X1 U7129 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  MUX2_X1 U7130 ( .A(n7509), .B(n7490), .S(n4391), .Z(n5513) );
  INV_X1 U7131 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7132 ( .A1(n5514), .A2(SI_20_), .ZN(n5515) );
  XNOR2_X1 U7133 ( .A(n5533), .B(n5532), .ZN(n7489) );
  NAND2_X1 U7134 ( .A1(n7489), .A2(n5819), .ZN(n5517) );
  NAND2_X1 U7135 ( .A1(n4395), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5516) );
  XNOR2_X1 U7136 ( .A(n5771), .B(n5683), .ZN(n5526) );
  NAND2_X1 U7137 ( .A1(n5518), .A2(n4538), .ZN(n5519) );
  NAND2_X1 U7138 ( .A1(n5538), .A2(n5519), .ZN(n8812) );
  OR2_X1 U7139 ( .A1(n8812), .A2(n5733), .ZN(n5524) );
  INV_X1 U7140 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7141 ( .A1(n4389), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7142 ( .A1(n5663), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5520) );
  OAI211_X1 U7143 ( .C1(n5307), .C2(n6601), .A(n5521), .B(n5520), .ZN(n5522)
         );
  INV_X1 U7144 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U7145 ( .A1(n5524), .A2(n5523), .ZN(n8597) );
  AND2_X1 U7146 ( .A1(n8597), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U7147 ( .A1(n5526), .A2(n5527), .ZN(n5531) );
  INV_X1 U7148 ( .A(n5526), .ZN(n8440) );
  INV_X1 U7149 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U7150 ( .A1(n8440), .A2(n5528), .ZN(n5529) );
  NAND2_X1 U7151 ( .A1(n5531), .A2(n5529), .ZN(n8514) );
  NAND2_X1 U7152 ( .A1(n8438), .A2(n5531), .ZN(n5546) );
  MUX2_X1 U7153 ( .A(n7611), .B(n7599), .S(n4397), .Z(n5549) );
  XNOR2_X1 U7154 ( .A(n5547), .B(n5548), .ZN(n7598) );
  NAND2_X1 U7155 ( .A1(n7598), .A2(n5819), .ZN(n5537) );
  NAND2_X1 U7156 ( .A1(n4395), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5536) );
  XNOR2_X1 U7157 ( .A(n9000), .B(n5683), .ZN(n5566) );
  INV_X1 U7158 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U7159 ( .A1(n5538), .A2(n8444), .ZN(n5539) );
  AND2_X1 U7160 ( .A1(n5558), .A2(n5539), .ZN(n8798) );
  NAND2_X1 U7161 ( .A1(n8798), .A2(n4393), .ZN(n5545) );
  INV_X1 U7162 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7163 ( .A1(n5799), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7164 ( .A1(n4389), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7165 ( .C1(n5542), .C2(n5593), .A(n5541), .B(n5540), .ZN(n5543)
         );
  INV_X1 U7166 ( .A(n5543), .ZN(n5544) );
  NOR2_X1 U7167 ( .A1(n8536), .A2(n5826), .ZN(n5567) );
  XNOR2_X1 U7168 ( .A(n5566), .B(n5567), .ZN(n8439) );
  INV_X1 U7169 ( .A(n5549), .ZN(n5550) );
  NAND2_X1 U7170 ( .A1(n5550), .A2(SI_21_), .ZN(n5551) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7653) );
  INV_X1 U7172 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7650) );
  MUX2_X1 U7173 ( .A(n7653), .B(n7650), .S(n4391), .Z(n5553) );
  INV_X1 U7174 ( .A(SI_22_), .ZN(n5552) );
  INV_X1 U7175 ( .A(n5553), .ZN(n5554) );
  NAND2_X1 U7176 ( .A1(n5554), .A2(SI_22_), .ZN(n5555) );
  XNOR2_X1 U7177 ( .A(n5574), .B(n5573), .ZN(n7649) );
  NAND2_X1 U7178 ( .A1(n7649), .A2(n5819), .ZN(n5557) );
  NAND2_X1 U7179 ( .A1(n4395), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5556) );
  XNOR2_X1 U7180 ( .A(n8992), .B(n5643), .ZN(n5570) );
  INV_X1 U7181 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U7182 ( .A1(n5558), .A2(n8535), .ZN(n5559) );
  NAND2_X1 U7183 ( .A1(n5597), .A2(n5559), .ZN(n8780) );
  INV_X1 U7184 ( .A(n8780), .ZN(n5560) );
  NAND2_X1 U7185 ( .A1(n5560), .A2(n4393), .ZN(n5565) );
  INV_X1 U7186 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8781) );
  NAND2_X1 U7187 ( .A1(n5799), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7188 ( .A1(n4390), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5561) );
  OAI211_X1 U7189 ( .C1(n8781), .C2(n5593), .A(n5562), .B(n5561), .ZN(n5563)
         );
  INV_X1 U7190 ( .A(n5563), .ZN(n5564) );
  NOR2_X1 U7191 ( .A1(n8794), .A2(n5826), .ZN(n5571) );
  INV_X1 U7192 ( .A(n5566), .ZN(n5568) );
  AND2_X1 U7193 ( .A1(n5568), .A2(n5567), .ZN(n8528) );
  AOI21_X1 U7194 ( .B1(n5570), .B2(n5571), .A(n8528), .ZN(n5569) );
  INV_X1 U7195 ( .A(n5570), .ZN(n8530) );
  INV_X1 U7196 ( .A(n5571), .ZN(n8532) );
  INV_X1 U7197 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5576) );
  INV_X1 U7198 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5575) );
  MUX2_X1 U7199 ( .A(n5576), .B(n5575), .S(n4392), .Z(n5578) );
  INV_X1 U7200 ( .A(SI_23_), .ZN(n5577) );
  NAND2_X1 U7201 ( .A1(n5578), .A2(n5577), .ZN(n5585) );
  INV_X1 U7202 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7203 ( .A1(n5579), .A2(SI_23_), .ZN(n5580) );
  XNOR2_X1 U7204 ( .A(n5584), .B(n5583), .ZN(n7795) );
  NAND2_X1 U7205 ( .A1(n7795), .A2(n5819), .ZN(n5582) );
  NAND2_X1 U7206 ( .A1(n4395), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5581) );
  XNOR2_X1 U7207 ( .A(n8987), .B(n5643), .ZN(n5606) );
  INV_X1 U7208 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7981) );
  INV_X1 U7209 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7951) );
  MUX2_X1 U7210 ( .A(n7981), .B(n7951), .S(n4392), .Z(n5615) );
  XNOR2_X1 U7211 ( .A(n5615), .B(SI_24_), .ZN(n5614) );
  NAND2_X1 U7212 ( .A1(n7950), .A2(n5177), .ZN(n5588) );
  NAND2_X1 U7213 ( .A1(n4395), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5587) );
  XNOR2_X1 U7214 ( .A(n8982), .B(n5683), .ZN(n8497) );
  INV_X1 U7215 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U7216 ( .A1(n5599), .A2(n8505), .ZN(n5590) );
  NAND2_X1 U7217 ( .A1(n5626), .A2(n5590), .ZN(n8746) );
  INV_X1 U7218 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U7219 ( .A1(n5799), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7220 ( .A1(n4389), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7221 ( .C1(n8745), .C2(n5593), .A(n5592), .B(n5591), .ZN(n5594)
         );
  INV_X1 U7222 ( .A(n5594), .ZN(n5595) );
  INV_X1 U7223 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U7224 ( .A1(n5597), .A2(n8406), .ZN(n5598) );
  AND2_X1 U7225 ( .A1(n5599), .A2(n5598), .ZN(n8762) );
  NAND2_X1 U7226 ( .A1(n8762), .A2(n4393), .ZN(n5604) );
  INV_X1 U7227 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U7228 ( .A1(n4389), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7229 ( .A1(n5663), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U7230 ( .C1(n5307), .C2(n6658), .A(n5601), .B(n5600), .ZN(n5602)
         );
  INV_X1 U7231 ( .A(n5602), .ZN(n5603) );
  OR2_X1 U7232 ( .A1(n8538), .A2(n5826), .ZN(n8404) );
  AOI21_X1 U7233 ( .B1(n8497), .B2(n8499), .A(n8404), .ZN(n5605) );
  NAND2_X1 U7234 ( .A1(n8405), .A2(n5605), .ZN(n5613) );
  NOR2_X1 U7235 ( .A1(n8499), .A2(n5826), .ZN(n5610) );
  INV_X1 U7236 ( .A(n8497), .ZN(n5609) );
  INV_X1 U7237 ( .A(n5606), .ZN(n5607) );
  OAI21_X1 U7238 ( .B1(n5610), .B2(n5609), .A(n8495), .ZN(n5612) );
  INV_X1 U7239 ( .A(n5610), .ZN(n8500) );
  INV_X1 U7240 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U7241 ( .A1(n5616), .A2(SI_24_), .ZN(n5617) );
  INV_X1 U7242 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8170) );
  INV_X1 U7243 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8167) );
  MUX2_X1 U7244 ( .A(n8170), .B(n8167), .S(n4397), .Z(n5619) );
  INV_X1 U7245 ( .A(SI_25_), .ZN(n6646) );
  INV_X1 U7246 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7247 ( .A1(n5620), .A2(SI_25_), .ZN(n5621) );
  NAND2_X1 U7248 ( .A1(n8165), .A2(n5819), .ZN(n5623) );
  NAND2_X1 U7249 ( .A1(n4395), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5622) );
  XNOR2_X1 U7250 ( .A(n4387), .B(n5643), .ZN(n8467) );
  INV_X1 U7251 ( .A(n5644), .ZN(n5645) );
  INV_X1 U7252 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7253 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  INV_X1 U7254 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U7255 ( .A1(n5799), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7256 ( .A1(n5663), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5628) );
  OAI211_X1 U7257 ( .C1(n5313), .C2(n6607), .A(n5629), .B(n5628), .ZN(n5630)
         );
  NOR2_X1 U7258 ( .A1(n8502), .A2(n5826), .ZN(n5631) );
  AND2_X1 U7259 ( .A1(n8467), .A2(n5631), .ZN(n8466) );
  INV_X1 U7260 ( .A(n8467), .ZN(n5633) );
  INV_X1 U7261 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7262 ( .A1(n5633), .A2(n5632), .ZN(n8469) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9100) );
  MUX2_X1 U7264 ( .A(n9100), .B(n10187), .S(n4397), .Z(n5638) );
  INV_X1 U7265 ( .A(SI_26_), .ZN(n5637) );
  NAND2_X1 U7266 ( .A1(n5638), .A2(n5637), .ZN(n5656) );
  INV_X1 U7267 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7268 ( .A1(n5639), .A2(SI_26_), .ZN(n5640) );
  XNOR2_X2 U7269 ( .A(n5655), .B(n5654), .ZN(n9098) );
  NAND2_X1 U7270 ( .A1(n4395), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5641) );
  XNOR2_X1 U7271 ( .A(n4375), .B(n5643), .ZN(n5652) );
  INV_X1 U7272 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U7273 ( .A1(n5645), .A2(n8574), .ZN(n5646) );
  NAND2_X1 U7274 ( .A1(n5673), .A2(n5646), .ZN(n8720) );
  INV_X1 U7275 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7276 ( .A1(n5663), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7277 ( .A1(n4390), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5647) );
  OAI211_X1 U7278 ( .C1(n5307), .C2(n6498), .A(n5648), .B(n5647), .ZN(n5649)
         );
  INV_X1 U7279 ( .A(n5649), .ZN(n5650) );
  NOR2_X1 U7280 ( .A1(n8698), .A2(n5826), .ZN(n5653) );
  XNOR2_X1 U7281 ( .A(n5652), .B(n5653), .ZN(n8572) );
  INV_X1 U7282 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9096) );
  INV_X1 U7283 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10183) );
  MUX2_X1 U7284 ( .A(n9096), .B(n10183), .S(n4397), .Z(n5658) );
  INV_X1 U7285 ( .A(SI_27_), .ZN(n5657) );
  NAND2_X1 U7286 ( .A1(n5658), .A2(n5657), .ZN(n5687) );
  INV_X1 U7287 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7288 ( .A1(n5659), .A2(SI_27_), .ZN(n5660) );
  NAND2_X1 U7289 ( .A1(n9095), .A2(n5177), .ZN(n5662) );
  NAND2_X1 U7290 ( .A1(n4395), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U7291 ( .A(n8692), .B(n5683), .ZN(n5671) );
  XNOR2_X1 U7292 ( .A(n5673), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U7293 ( .A1(n8690), .A2(n4393), .ZN(n5668) );
  INV_X1 U7294 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7295 ( .A1(n5663), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7296 ( .A1(n4389), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5664) );
  OAI211_X1 U7297 ( .C1(n5307), .C2(n6657), .A(n5665), .B(n5664), .ZN(n5666)
         );
  INV_X1 U7298 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7299 ( .A1(n8595), .A2(n5525), .ZN(n5669) );
  XNOR2_X1 U7300 ( .A(n5671), .B(n5669), .ZN(n8382) );
  INV_X1 U7301 ( .A(n5669), .ZN(n5670) );
  INV_X1 U7302 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8385) );
  INV_X1 U7303 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5672) );
  OAI21_X1 U7304 ( .B1(n5673), .B2(n8385), .A(n5672), .ZN(n5676) );
  INV_X1 U7305 ( .A(n5673), .ZN(n5675) );
  AND2_X1 U7306 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5674) );
  NAND2_X1 U7307 ( .A1(n5675), .A2(n5674), .ZN(n8660) );
  NAND2_X1 U7308 ( .A1(n5676), .A2(n8660), .ZN(n5741) );
  INV_X1 U7309 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7310 ( .A1(n5799), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7311 ( .A1(n4390), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5677) );
  OAI211_X1 U7312 ( .C1(n5679), .C2(n5593), .A(n5678), .B(n5677), .ZN(n5680)
         );
  INV_X1 U7313 ( .A(n5680), .ZN(n5681) );
  OR2_X1 U7314 ( .A1(n8699), .A2(n5826), .ZN(n5684) );
  XNOR2_X1 U7315 ( .A(n5684), .B(n5683), .ZN(n5725) );
  INV_X1 U7316 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5689) );
  INV_X1 U7317 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10179) );
  MUX2_X1 U7318 ( .A(n5689), .B(n10179), .S(n4391), .Z(n5786) );
  XNOR2_X1 U7319 ( .A(n5786), .B(SI_28_), .ZN(n5783) );
  NAND2_X1 U7320 ( .A1(n9091), .A2(n5819), .ZN(n5691) );
  NAND2_X1 U7321 ( .A1(n4395), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5690) );
  INV_X1 U7322 ( .A(n8959), .ZN(n8675) );
  NAND2_X1 U7323 ( .A1(n5719), .A2(n6682), .ZN(n5694) );
  NAND2_X1 U7324 ( .A1(n5694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5696) );
  INV_X1 U7325 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5695) );
  OR2_X1 U7326 ( .A1(n5223), .A2(n5697), .ZN(n5702) );
  INV_X1 U7327 ( .A(n5702), .ZN(n5699) );
  NAND2_X1 U7328 ( .A1(n5699), .A2(n5698), .ZN(n5704) );
  NAND2_X1 U7329 ( .A1(n5704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5700) );
  MUX2_X1 U7330 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5700), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5701) );
  NAND2_X1 U7331 ( .A1(n5702), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5703) );
  MUX2_X1 U7332 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5703), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5705) );
  NAND2_X1 U7333 ( .A1(n5705), .A2(n5704), .ZN(n8168) );
  INV_X1 U7334 ( .A(P2_B_REG_SCAN_IN), .ZN(n8326) );
  XOR2_X1 U7335 ( .A(n7983), .B(n8326), .Z(n5706) );
  INV_X1 U7336 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10375) );
  INV_X1 U7337 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10377) );
  AND2_X1 U7338 ( .A1(n9102), .A2(n8168), .ZN(n10378) );
  AOI21_X1 U7339 ( .B1(n10364), .B2(n10377), .A(n10378), .ZN(n6807) );
  NOR4_X1 U7340 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5712) );
  NOR4_X1 U7341 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5711) );
  NOR4_X1 U7342 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5710) );
  NOR4_X1 U7343 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5709) );
  NAND4_X1 U7344 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n5717)
         );
  NOR2_X1 U7345 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .ZN(
        n6482) );
  NOR4_X1 U7346 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5715) );
  NOR4_X1 U7347 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5714) );
  NOR4_X1 U7348 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5713) );
  NAND4_X1 U7349 ( .A1(n6482), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(n5716)
         );
  OAI21_X1 U7350 ( .B1(n5717), .B2(n5716), .A(n10364), .ZN(n6806) );
  AND2_X1 U7351 ( .A1(n6807), .A2(n6806), .ZN(n7315) );
  AND2_X1 U7352 ( .A1(n7013), .A2(n7315), .ZN(n5742) );
  OR2_X1 U7353 ( .A1(n8168), .A2(n9102), .ZN(n5718) );
  XNOR2_X1 U7354 ( .A(n5719), .B(n6682), .ZN(n5987) );
  NOR2_X1 U7355 ( .A1(n5983), .A2(n7507), .ZN(n7324) );
  NAND2_X1 U7356 ( .A1(n5740), .A2(n7324), .ZN(n5722) );
  INV_X1 U7357 ( .A(n7507), .ZN(n5832) );
  NAND2_X1 U7358 ( .A1(n10424), .A2(n8640), .ZN(n6805) );
  INV_X1 U7359 ( .A(n6805), .ZN(n5721) );
  NOR3_X1 U7360 ( .A1(n8675), .A2(n5725), .A3(n8590), .ZN(n5723) );
  AOI21_X1 U7361 ( .B1(n5725), .B2(n8675), .A(n5723), .ZN(n5730) );
  NAND3_X1 U7362 ( .A1(n8959), .A2(n5725), .A3(n8570), .ZN(n5724) );
  OAI21_X1 U7363 ( .B1(n8959), .B2(n5725), .A(n5724), .ZN(n5726) );
  NAND2_X1 U7364 ( .A1(n5058), .A2(n5851), .ZN(n6992) );
  NAND2_X1 U7365 ( .A1(n10398), .A2(n6992), .ZN(n5727) );
  AOI21_X1 U7366 ( .B1(n8959), .B2(n8590), .A(n8583), .ZN(n5729) );
  NAND2_X1 U7367 ( .A1(n5731), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5732) );
  XNOR2_X1 U7368 ( .A(n5732), .B(n4820), .ZN(n6999) );
  OR2_X1 U7369 ( .A1(n8660), .A2(n5733), .ZN(n5738) );
  INV_X1 U7370 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U7371 ( .A1(n5799), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7372 ( .A1(n4390), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7373 ( .C1(n8659), .C2(n5593), .A(n5735), .B(n5734), .ZN(n5736)
         );
  INV_X1 U7374 ( .A(n5736), .ZN(n5737) );
  INV_X1 U7375 ( .A(n6999), .ZN(n5739) );
  OAI22_X1 U7376 ( .A1(n8354), .A2(n8793), .B1(n7511), .B2(n8795), .ZN(n8681)
         );
  NAND2_X1 U7377 ( .A1(n5740), .A2(n5989), .ZN(n8573) );
  INV_X1 U7378 ( .A(n5741), .ZN(n8673) );
  INV_X1 U7379 ( .A(n5742), .ZN(n5746) );
  NAND2_X1 U7380 ( .A1(n5746), .A2(n10398), .ZN(n5745) );
  NOR2_X1 U7381 ( .A1(n5989), .A2(n6992), .ZN(n6804) );
  INV_X1 U7382 ( .A(n6804), .ZN(n5743) );
  AND3_X1 U7383 ( .A1(n6719), .A2(n5743), .A3(n5987), .ZN(n5744) );
  NAND2_X1 U7384 ( .A1(n5745), .A2(n5744), .ZN(n7265) );
  AND2_X1 U7385 ( .A1(n5746), .A2(n7324), .ZN(n7267) );
  OR2_X1 U7386 ( .A1(n7265), .A2(n7267), .ZN(n5747) );
  AOI22_X1 U7387 ( .A1(n8673), .A2(n8464), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        n4369), .ZN(n5748) );
  OAI21_X1 U7388 ( .B1(n4895), .B2(n8573), .A(n5748), .ZN(n5749) );
  NAND2_X1 U7389 ( .A1(n5751), .A2(n5750), .ZN(P2_U3222) );
  NAND2_X1 U7390 ( .A1(n7348), .A2(n5853), .ZN(n7054) );
  NAND2_X1 U7391 ( .A1(n7517), .A2(n8927), .ZN(n5856) );
  NAND2_X1 U7392 ( .A1(n7525), .A2(n7331), .ZN(n5859) );
  INV_X1 U7393 ( .A(n7525), .ZN(n8608) );
  NAND2_X1 U7394 ( .A1(n8608), .A2(n10399), .ZN(n7547) );
  NAND2_X1 U7395 ( .A1(n7547), .A2(n5871), .ZN(n5869) );
  INV_X1 U7396 ( .A(n5869), .ZN(n5755) );
  NAND2_X1 U7397 ( .A1(n7546), .A2(n5755), .ZN(n5756) );
  NAND2_X1 U7398 ( .A1(n7571), .A2(n10408), .ZN(n5861) );
  NAND2_X1 U7399 ( .A1(n5756), .A2(n5861), .ZN(n7531) );
  NOR2_X1 U7400 ( .A1(n8606), .A2(n7542), .ZN(n5863) );
  INV_X1 U7401 ( .A(n5863), .ZN(n5876) );
  NAND2_X1 U7402 ( .A1(n8606), .A2(n7542), .ZN(n5873) );
  NAND2_X1 U7403 ( .A1(n7531), .A2(n7532), .ZN(n5757) );
  NAND2_X1 U7404 ( .A1(n7839), .A2(n7669), .ZN(n5880) );
  INV_X1 U7405 ( .A(n7669), .ZN(n7592) );
  INV_X1 U7406 ( .A(n7839), .ZN(n8605) );
  NAND2_X1 U7407 ( .A1(n7592), .A2(n8605), .ZN(n5881) );
  XNOR2_X1 U7408 ( .A(n10422), .B(n8604), .ZN(n7677) );
  INV_X1 U7409 ( .A(n8604), .ZN(n7866) );
  NAND2_X1 U7410 ( .A1(n10422), .A2(n7866), .ZN(n7806) );
  NOR2_X1 U7411 ( .A1(n9061), .A2(n8132), .ZN(n5886) );
  INV_X1 U7412 ( .A(n5886), .ZN(n5890) );
  NAND2_X1 U7413 ( .A1(n9061), .A2(n8132), .ZN(n8125) );
  INV_X1 U7414 ( .A(n8142), .ZN(n9056) );
  INV_X1 U7415 ( .A(n8602), .ZN(n7922) );
  NAND2_X1 U7416 ( .A1(n9056), .A2(n7922), .ZN(n5888) );
  NAND2_X1 U7417 ( .A1(n5888), .A2(n8125), .ZN(n5887) );
  INV_X1 U7418 ( .A(n5887), .ZN(n5758) );
  AND2_X1 U7419 ( .A1(n8142), .A2(n8602), .ZN(n8127) );
  NAND2_X1 U7420 ( .A1(n9052), .A2(n8455), .ZN(n5896) );
  NAND2_X1 U7421 ( .A1(n9046), .A2(n8153), .ZN(n5900) );
  NOR2_X1 U7422 ( .A1(n8180), .A2(n8458), .ZN(n5903) );
  INV_X1 U7423 ( .A(n5903), .ZN(n5759) );
  AND2_X2 U7424 ( .A1(n5759), .A2(n5760), .ZN(n8150) );
  NAND2_X1 U7425 ( .A1(n9035), .A2(n8335), .ZN(n5907) );
  NAND2_X1 U7426 ( .A1(n5906), .A2(n5907), .ZN(n8333) );
  NAND2_X1 U7427 ( .A1(n8172), .A2(n4485), .ZN(n8171) );
  NAND2_X1 U7428 ( .A1(n8171), .A2(n5906), .ZN(n8904) );
  NOR2_X1 U7429 ( .A1(n9030), .A2(n8481), .ZN(n5909) );
  INV_X1 U7430 ( .A(n5909), .ZN(n5762) );
  AND2_X1 U7431 ( .A1(n9030), .A2(n8481), .ZN(n5910) );
  INV_X1 U7432 ( .A(n5910), .ZN(n5761) );
  NAND2_X1 U7433 ( .A1(n8904), .A2(n8905), .ZN(n8903) );
  NAND2_X1 U7434 ( .A1(n9014), .A2(n8488), .ZN(n8825) );
  NAND2_X1 U7435 ( .A1(n9020), .A2(n8566), .ZN(n5915) );
  NAND2_X1 U7436 ( .A1(n9024), .A2(n8487), .ZN(n8845) );
  AND2_X1 U7437 ( .A1(n5915), .A2(n8845), .ZN(n8824) );
  INV_X1 U7438 ( .A(n8824), .ZN(n5763) );
  NAND2_X1 U7439 ( .A1(n8844), .A2(n5764), .ZN(n5769) );
  NOR2_X1 U7440 ( .A1(n9014), .A2(n8488), .ZN(n5923) );
  INV_X1 U7441 ( .A(n5923), .ZN(n5765) );
  INV_X1 U7442 ( .A(n9020), .ZN(n8357) );
  NAND2_X1 U7443 ( .A1(n5830), .A2(n8566), .ZN(n5766) );
  INV_X1 U7444 ( .A(n5830), .ZN(n5913) );
  INV_X1 U7445 ( .A(n8566), .ZN(n8888) );
  AOI22_X1 U7446 ( .A1(n8357), .A2(n5766), .B1(n5913), .B2(n8888), .ZN(n5767)
         );
  NAND2_X1 U7447 ( .A1(n8859), .A2(n5767), .ZN(n8823) );
  OR2_X1 U7448 ( .A1(n8837), .A2(n8509), .ZN(n5925) );
  NAND2_X1 U7449 ( .A1(n8837), .A2(n8509), .ZN(n5922) );
  NAND2_X1 U7450 ( .A1(n5925), .A2(n5922), .ZN(n8833) );
  AOI21_X1 U7451 ( .B1(n8825), .B2(n8823), .A(n8833), .ZN(n5768) );
  NAND2_X1 U7452 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  INV_X1 U7453 ( .A(n8597), .ZN(n8792) );
  NAND2_X1 U7454 ( .A1(n9004), .A2(n8792), .ZN(n5929) );
  NAND2_X1 U7455 ( .A1(n5919), .A2(n5929), .ZN(n8804) );
  XNOR2_X1 U7456 ( .A(n9000), .B(n8536), .ZN(n8790) );
  NAND2_X1 U7457 ( .A1(n9000), .A2(n8536), .ZN(n5931) );
  INV_X1 U7458 ( .A(n5931), .ZN(n5773) );
  NAND2_X1 U7459 ( .A1(n8992), .A2(n8794), .ZN(n5932) );
  OR2_X1 U7460 ( .A1(n8987), .A2(n8538), .ZN(n5941) );
  NAND2_X1 U7461 ( .A1(n8987), .A2(n8538), .ZN(n5847) );
  NAND2_X1 U7462 ( .A1(n5941), .A2(n5847), .ZN(n8766) );
  NAND2_X1 U7463 ( .A1(n4387), .A2(n8502), .ZN(n5829) );
  NAND2_X1 U7464 ( .A1(n8725), .A2(n5013), .ZN(n5780) );
  INV_X1 U7465 ( .A(n5956), .ZN(n5777) );
  OAI21_X1 U7466 ( .B1(n5777), .B2(n5776), .A(n5828), .ZN(n5778) );
  NAND2_X1 U7467 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  INV_X1 U7468 ( .A(n5955), .ZN(n5782) );
  NAND2_X1 U7469 ( .A1(n8959), .A2(n8699), .ZN(n5963) );
  NAND2_X1 U7470 ( .A1(n5781), .A2(n8677), .ZN(n8678) );
  INV_X1 U7471 ( .A(SI_28_), .ZN(n5785) );
  NAND2_X1 U7472 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  INV_X1 U7473 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8379) );
  INV_X1 U7474 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9343) );
  MUX2_X1 U7475 ( .A(n8379), .B(n9343), .S(n4397), .Z(n5808) );
  XNOR2_X1 U7476 ( .A(n5808), .B(SI_29_), .ZN(n5789) );
  NAND2_X1 U7477 ( .A1(n9342), .A2(n5819), .ZN(n5791) );
  NAND2_X1 U7478 ( .A1(n4395), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5790) );
  INV_X1 U7479 ( .A(n5968), .ZN(n5962) );
  NAND2_X1 U7480 ( .A1(n8662), .A2(n7511), .ZN(n5969) );
  INV_X1 U7481 ( .A(SI_29_), .ZN(n5809) );
  INV_X1 U7482 ( .A(n5808), .ZN(n5806) );
  MUX2_X1 U7483 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4392), .Z(n5792) );
  NAND2_X1 U7484 ( .A1(n5792), .A2(SI_30_), .ZN(n5810) );
  INV_X1 U7485 ( .A(n5792), .ZN(n5794) );
  INV_X1 U7486 ( .A(SI_30_), .ZN(n5793) );
  NAND2_X1 U7487 ( .A1(n5794), .A2(n5793), .ZN(n5811) );
  NAND2_X1 U7488 ( .A1(n5810), .A2(n5811), .ZN(n5795) );
  NAND2_X1 U7489 ( .A1(n9401), .A2(n5819), .ZN(n5798) );
  NAND2_X1 U7490 ( .A1(n4395), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7491 ( .A1(n5799), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7492 ( .A1(n4390), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7493 ( .A1(n5663), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7494 ( .A1(n5799), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7495 ( .A1(n5663), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7496 ( .A1(n4389), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5803) );
  AND3_X1 U7497 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n8327) );
  NOR2_X1 U7498 ( .A1(n8652), .A2(n8327), .ZN(n5971) );
  INV_X1 U7499 ( .A(n5971), .ZN(n5823) );
  INV_X1 U7500 ( .A(n5970), .ZN(n5822) );
  NAND2_X1 U7501 ( .A1(n5806), .A2(SI_29_), .ZN(n5807) );
  AND2_X1 U7502 ( .A1(n5810), .A2(n5807), .ZN(n5814) );
  NAND3_X1 U7503 ( .A1(n5810), .A2(n5809), .A3(n5808), .ZN(n5812) );
  NAND2_X1 U7504 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  MUX2_X1 U7505 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4397), .Z(n5816) );
  XNOR2_X1 U7506 ( .A(n5816), .B(SI_31_), .ZN(n5817) );
  NAND2_X1 U7507 ( .A1(n9408), .A2(n5819), .ZN(n5821) );
  NAND2_X1 U7508 ( .A1(n4395), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5820) );
  OR2_X1 U7509 ( .A1(n8952), .A2(n8646), .ZN(n5977) );
  NAND2_X1 U7510 ( .A1(n5822), .A2(n5977), .ZN(n5975) );
  NAND2_X1 U7511 ( .A1(n8952), .A2(n8646), .ZN(n5978) );
  NAND2_X1 U7512 ( .A1(n5824), .A2(n5978), .ZN(n5825) );
  XNOR2_X1 U7513 ( .A(n5825), .B(n8640), .ZN(n5827) );
  AND2_X1 U7514 ( .A1(n5832), .A2(n5851), .ZN(n6815) );
  NAND2_X1 U7515 ( .A1(n5827), .A2(n5004), .ZN(n5986) );
  NAND2_X1 U7516 ( .A1(n5823), .A2(n5978), .ZN(n5974) );
  INV_X1 U7517 ( .A(n8686), .ZN(n8694) );
  NAND2_X1 U7518 ( .A1(n5859), .A2(n7547), .ZN(n7321) );
  NAND2_X1 U7519 ( .A1(n4973), .A2(n7500), .ZN(n10385) );
  NAND3_X1 U7520 ( .A1(n10385), .A2(n6809), .A3(n5832), .ZN(n5833) );
  XNOR2_X1 U7521 ( .A(n8607), .B(n10408), .ZN(n7549) );
  NAND4_X1 U7522 ( .A1(n5834), .A2(n7532), .A3(n7055), .A4(n7549), .ZN(n5835)
         );
  NAND2_X1 U7523 ( .A1(n5880), .A2(n5881), .ZN(n7579) );
  NAND2_X1 U7524 ( .A1(n5889), .A2(n5888), .ZN(n8124) );
  NOR4_X1 U7525 ( .A1(n5835), .A2(n7579), .A3(n7805), .A4(n8124), .ZN(n5836)
         );
  AND2_X2 U7526 ( .A1(n5895), .A2(n5896), .ZN(n7999) );
  NAND4_X1 U7527 ( .A1(n5836), .A2(n8148), .A3(n7999), .A4(n7677), .ZN(n5838)
         );
  INV_X1 U7528 ( .A(n8150), .ZN(n5837) );
  NOR4_X1 U7529 ( .A1(n8914), .A2(n5838), .A3(n8333), .A4(n5837), .ZN(n5839)
         );
  XNOR2_X1 U7530 ( .A(n9020), .B(n8566), .ZN(n8870) );
  INV_X1 U7531 ( .A(n8870), .ZN(n8864) );
  NAND4_X1 U7532 ( .A1(n8859), .A2(n4435), .A3(n5839), .A4(n8864), .ZN(n5840)
         );
  NOR4_X1 U7533 ( .A1(n4988), .A2(n8833), .A3(n8804), .A4(n5840), .ZN(n5841)
         );
  NAND3_X1 U7534 ( .A1(n5841), .A2(n4826), .A3(n4905), .ZN(n5842) );
  INV_X1 U7535 ( .A(n6816), .ZN(n5844) );
  AOI22_X1 U7536 ( .A1(n5845), .A2(n7609), .B1(n5844), .B2(n7507), .ZN(n5985)
         );
  NAND2_X1 U7537 ( .A1(n5851), .A2(n8640), .ZN(n5846) );
  INV_X1 U7538 ( .A(n5847), .ZN(n5940) );
  INV_X1 U7539 ( .A(n5933), .ZN(n5848) );
  NOR2_X1 U7540 ( .A1(n9000), .A2(n8536), .ZN(n5928) );
  NOR3_X1 U7541 ( .A1(n5848), .A2(n5928), .A3(n5976), .ZN(n5938) );
  INV_X1 U7542 ( .A(n6810), .ZN(n5850) );
  INV_X1 U7543 ( .A(n5853), .ZN(n5849) );
  AOI211_X1 U7544 ( .C1(n10385), .C2(n6809), .A(n5850), .B(n5849), .ZN(n5868)
         );
  NAND2_X1 U7545 ( .A1(n5852), .A2(n4400), .ZN(n5867) );
  AOI21_X1 U7546 ( .B1(n5851), .B2(n10385), .A(n5831), .ZN(n5855) );
  NAND2_X1 U7547 ( .A1(n6809), .A2(n5852), .ZN(n5854) );
  OAI211_X1 U7548 ( .C1(n5855), .C2(n5854), .A(n5976), .B(n5853), .ZN(n5858)
         );
  NAND2_X1 U7549 ( .A1(n5859), .A2(n5856), .ZN(n5857) );
  AOI22_X1 U7550 ( .A1(n5858), .A2(n7055), .B1(n5976), .B2(n5857), .ZN(n5865)
         );
  NAND2_X1 U7551 ( .A1(n5859), .A2(n5861), .ZN(n5860) );
  INV_X1 U7552 ( .A(n5861), .ZN(n5862) );
  OAI21_X1 U7553 ( .B1(n5863), .B2(n5862), .A(n5976), .ZN(n5864) );
  OAI211_X1 U7554 ( .C1(n5868), .C2(n5867), .A(n5866), .B(n5873), .ZN(n5879)
         );
  AOI21_X1 U7555 ( .B1(n7311), .B2(n8609), .A(n5869), .ZN(n5870) );
  AOI21_X1 U7556 ( .B1(n5872), .B2(n5871), .A(n5870), .ZN(n5875) );
  INV_X1 U7557 ( .A(n5873), .ZN(n5874) );
  OAI21_X1 U7558 ( .B1(n5875), .B2(n5874), .A(n4400), .ZN(n5878) );
  NOR2_X1 U7559 ( .A1(n5876), .A2(n5976), .ZN(n5877) );
  MUX2_X1 U7560 ( .A(n5881), .B(n5880), .S(n5976), .Z(n5882) );
  NAND2_X1 U7561 ( .A1(n7677), .A2(n5882), .ZN(n5885) );
  INV_X1 U7562 ( .A(n10422), .ZN(n7845) );
  NAND2_X1 U7563 ( .A1(n7845), .A2(n8604), .ZN(n5883) );
  AOI211_X1 U7564 ( .C1(n5976), .C2(n5887), .A(n5886), .B(n8127), .ZN(n5894)
         );
  NAND2_X1 U7565 ( .A1(n5896), .A2(n5888), .ZN(n5892) );
  INV_X1 U7566 ( .A(n5888), .ZN(n8130) );
  OAI211_X1 U7567 ( .C1(n8130), .C2(n5890), .A(n5895), .B(n5889), .ZN(n5891)
         );
  MUX2_X1 U7568 ( .A(n5892), .B(n5891), .S(n5976), .Z(n5893) );
  NAND2_X1 U7569 ( .A1(n5899), .A2(n5895), .ZN(n5898) );
  NAND2_X1 U7570 ( .A1(n5900), .A2(n5896), .ZN(n5897) );
  MUX2_X1 U7571 ( .A(n5900), .B(n5899), .S(n5976), .Z(n5901) );
  MUX2_X1 U7572 ( .A(n5904), .B(n5903), .S(n5976), .Z(n5905) );
  MUX2_X1 U7573 ( .A(n5907), .B(n5906), .S(n5976), .Z(n5908) );
  MUX2_X1 U7574 ( .A(n5910), .B(n5909), .S(n5976), .Z(n5911) );
  INV_X1 U7575 ( .A(n8845), .ZN(n5912) );
  MUX2_X1 U7576 ( .A(n5913), .B(n5912), .S(n5976), .Z(n5914) );
  NAND2_X1 U7577 ( .A1(n8825), .A2(n5915), .ZN(n5916) );
  NOR2_X1 U7578 ( .A1(n9020), .A2(n8566), .ZN(n8846) );
  MUX2_X1 U7579 ( .A(n5916), .B(n8846), .S(n5976), .Z(n5917) );
  INV_X1 U7580 ( .A(n5924), .ZN(n5918) );
  NAND3_X1 U7581 ( .A1(n5920), .A2(n5925), .A3(n5919), .ZN(n5921) );
  NAND3_X1 U7582 ( .A1(n5921), .A2(n5929), .A3(n5931), .ZN(n5937) );
  INV_X1 U7583 ( .A(n5932), .ZN(n5936) );
  NAND2_X1 U7584 ( .A1(n5926), .A2(n5925), .ZN(n5930) );
  NAND2_X1 U7585 ( .A1(n5932), .A2(n5931), .ZN(n5934) );
  INV_X1 U7586 ( .A(n5941), .ZN(n5942) );
  NOR2_X1 U7587 ( .A1(n5944), .A2(n5942), .ZN(n5943) );
  OAI22_X1 U7588 ( .A1(n5945), .A2(n5944), .B1(n5943), .B2(n5976), .ZN(n5946)
         );
  INV_X1 U7589 ( .A(n5948), .ZN(n5949) );
  NOR2_X1 U7590 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  INV_X1 U7591 ( .A(n5953), .ZN(n5954) );
  NOR2_X1 U7592 ( .A1(n5955), .A2(n8676), .ZN(n5957) );
  MUX2_X1 U7593 ( .A(n5957), .B(n5956), .S(n5976), .Z(n5958) );
  NOR2_X1 U7594 ( .A1(n5962), .A2(n5976), .ZN(n5966) );
  OAI211_X1 U7595 ( .C1(n4400), .C2(n8959), .A(n5964), .B(n5963), .ZN(n5965)
         );
  OAI21_X1 U7596 ( .B1(n5967), .B2(n5966), .A(n5965), .ZN(n5973) );
  MUX2_X1 U7597 ( .A(n5969), .B(n5968), .S(n5976), .Z(n5972) );
  MUX2_X1 U7598 ( .A(n5975), .B(n5974), .S(n5976), .Z(n5980) );
  MUX2_X1 U7599 ( .A(n5978), .B(n5977), .S(n5976), .Z(n5979) );
  OAI21_X1 U7600 ( .B1(n5981), .B2(n5980), .A(n5979), .ZN(n5982) );
  INV_X1 U7601 ( .A(n5989), .ZN(n5992) );
  XNOR2_X1 U7602 ( .A(n5991), .B(n5990), .ZN(n9097) );
  NOR4_X1 U7603 ( .A1(n10363), .A2(n5992), .A3(n8793), .A4(n9097), .ZN(n5993)
         );
  AOI211_X1 U7604 ( .C1(n7798), .C2(n5988), .A(n8326), .B(n5993), .ZN(n5994)
         );
  INV_X1 U7605 ( .A(n5994), .ZN(n5995) );
  NAND2_X1 U7606 ( .A1(n5996), .A2(n5995), .ZN(P2_U3244) );
  NAND2_X1 U7607 ( .A1(n6052), .A2(n6001), .ZN(n6096) );
  NOR2_X1 U7608 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6005) );
  NOR2_X1 U7609 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6004) );
  NOR2_X1 U7610 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n6006) );
  NAND2_X1 U7611 ( .A1(n4416), .A2(n6006), .ZN(n6009) );
  NAND4_X1 U7612 ( .A1(n6007), .A2(n6232), .A3(n6383), .A4(n6231), .ZN(n6008)
         );
  INV_X1 U7613 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7614 ( .A1(n6085), .A2(n4391), .ZN(n6065) );
  NAND2_X1 U7615 ( .A1(n7598), .A2(n4620), .ZN(n6018) );
  OR2_X1 U7616 ( .A1(n9409), .A2(n7599), .ZN(n6017) );
  NAND2_X1 U7617 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n6024) );
  INV_X1 U7618 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U7619 ( .A1(n6302), .A2(n9194), .ZN(n6026) );
  NAND2_X1 U7620 ( .A1(n6312), .A2(n6026), .ZN(n9877) );
  NAND2_X1 U7621 ( .A1(n6027), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6028) );
  AND2_X4 U7622 ( .A1(n6033), .A2(n6032), .ZN(n6079) );
  OR2_X1 U7623 ( .A1(n9877), .A2(n6355), .ZN(n6038) );
  INV_X1 U7624 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U7625 ( .A1(n6829), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7626 ( .A1(n6213), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6034) );
  OAI211_X1 U7627 ( .C1(n6080), .C2(n9878), .A(n6035), .B(n6034), .ZN(n6036)
         );
  INV_X1 U7628 ( .A(n6036), .ZN(n6037) );
  NAND2_X1 U7629 ( .A1(n6091), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7630 ( .A1(n6079), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7631 ( .A1(n4397), .A2(SI_0_), .ZN(n6044) );
  INV_X1 U7632 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7633 ( .A1(n6044), .A2(n6043), .ZN(n6046) );
  AND2_X1 U7634 ( .A1(n6046), .A2(n6045), .ZN(n10190) );
  NAND2_X1 U7635 ( .A1(n6077), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7636 ( .A1(n6091), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7637 ( .A1(n6079), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7638 ( .A1(n7617), .A2(n9364), .ZN(n6056) );
  NAND2_X1 U7639 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6051) );
  MUX2_X1 U7640 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6051), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n6053) );
  INV_X1 U7641 ( .A(n6052), .ZN(n6066) );
  NAND2_X1 U7642 ( .A1(n6056), .A2(n4386), .ZN(n6060) );
  INV_X1 U7643 ( .A(n7617), .ZN(n6058) );
  NAND2_X1 U7644 ( .A1(n6058), .A2(n6057), .ZN(n6059) );
  NAND2_X1 U7645 ( .A1(n6060), .A2(n6059), .ZN(n6072) );
  NAND2_X1 U7646 ( .A1(n6077), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7647 ( .A1(n6079), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7648 ( .A1(n6091), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7649 ( .A1(n6066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6068) );
  INV_X1 U7650 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6067) );
  OR2_X1 U7651 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NAND2_X1 U7652 ( .A1(n6068), .A2(n6067), .ZN(n6086) );
  AND2_X1 U7653 ( .A1(n6069), .A2(n6086), .ZN(n9671) );
  INV_X1 U7654 ( .A(n9671), .ZN(n6070) );
  NAND2_X1 U7655 ( .A1(n7615), .A2(n7161), .ZN(n6073) );
  NAND2_X1 U7656 ( .A1(n6072), .A2(n6073), .ZN(n6076) );
  NAND2_X1 U7657 ( .A1(n9369), .A2(n9366), .ZN(n6408) );
  INV_X1 U7658 ( .A(n6408), .ZN(n6074) );
  NAND2_X1 U7659 ( .A1(n6076), .A2(n6075), .ZN(n7967) );
  NAND2_X1 U7660 ( .A1(n6077), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6084) );
  INV_X1 U7661 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7662 ( .A1(n6079), .A2(n6078), .ZN(n6083) );
  NAND2_X1 U7663 ( .A1(n6091), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6082) );
  INV_X1 U7664 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U7665 ( .A1(n4620), .A2(n6730), .ZN(n6089) );
  NAND2_X1 U7666 ( .A1(n6086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7667 ( .A1(n6284), .A2(n6856), .ZN(n6088) );
  NAND2_X1 U7668 ( .A1(n7301), .A2(n7972), .ZN(n9558) );
  OAI22_X1 U7669 ( .A1(n7967), .A2(n9581), .B1(n7972), .B2(n9648), .ZN(n8009)
         );
  NAND2_X1 U7670 ( .A1(n6829), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6095) );
  INV_X1 U7671 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6090) );
  XNOR2_X1 U7672 ( .A(n6090), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U7673 ( .A1(n6079), .A2(n8016), .ZN(n6094) );
  NAND2_X1 U7674 ( .A1(n6091), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7675 ( .A1(n6213), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6092) );
  AND4_X2 U7676 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n7780)
         );
  NAND2_X1 U7677 ( .A1(n6096), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6097) );
  MUX2_X1 U7678 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6097), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6098) );
  AND2_X1 U7679 ( .A1(n6219), .A2(n6098), .ZN(n9690) );
  AOI22_X1 U7680 ( .A1(n6371), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6284), .B2(
        n9690), .ZN(n6100) );
  NAND2_X1 U7681 ( .A1(n6725), .A2(n4620), .ZN(n6099) );
  NAND2_X1 U7682 ( .A1(n6100), .A2(n6099), .ZN(n8019) );
  NAND2_X1 U7683 ( .A1(n7780), .A2(n8019), .ZN(n9556) );
  NAND2_X1 U7684 ( .A1(n8009), .A2(n9583), .ZN(n6102) );
  NAND2_X1 U7685 ( .A1(n7780), .A2(n8015), .ZN(n6101) );
  NAND2_X1 U7686 ( .A1(n6102), .A2(n6101), .ZN(n7787) );
  NAND2_X1 U7687 ( .A1(n6829), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6109) );
  INV_X1 U7688 ( .A(n6103), .ZN(n6118) );
  INV_X1 U7689 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7690 ( .A1(n6118), .A2(n6104), .ZN(n6105) );
  AND2_X1 U7691 ( .A1(n6133), .A2(n6105), .ZN(n7858) );
  NAND2_X1 U7692 ( .A1(n6079), .A2(n7858), .ZN(n6108) );
  NAND2_X1 U7693 ( .A1(n6787), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7694 ( .A1(n6213), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7695 ( .A1(n6723), .A2(n4620), .ZN(n6114) );
  INV_X1 U7696 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7697 ( .A1(n6111), .A2(n6110), .ZN(n6191) );
  NAND2_X1 U7698 ( .A1(n6191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6112) );
  XNOR2_X1 U7699 ( .A(n6112), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6863) );
  AOI22_X1 U7700 ( .A1(n6371), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6284), .B2(
        n6863), .ZN(n6113) );
  NAND2_X1 U7701 ( .A1(n6114), .A2(n6113), .ZN(n7853) );
  NAND2_X1 U7702 ( .A1(n6829), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6124) );
  INV_X1 U7703 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7704 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6115) );
  NAND2_X1 U7705 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  AND2_X1 U7706 ( .A1(n6118), .A2(n6117), .ZN(n7781) );
  NAND2_X1 U7707 ( .A1(n6079), .A2(n7781), .ZN(n6123) );
  NAND2_X1 U7708 ( .A1(n6787), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6122) );
  INV_X1 U7709 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7710 ( .A1(n6732), .A2(n4620), .ZN(n6127) );
  NAND2_X1 U7711 ( .A1(n6219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7712 ( .A(n6125), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6861) );
  AOI22_X1 U7713 ( .A1(n6371), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6284), .B2(
        n6861), .ZN(n6126) );
  NAND2_X1 U7714 ( .A1(n9646), .A2(n7786), .ZN(n7825) );
  NAND2_X1 U7715 ( .A1(n6734), .A2(n6350), .ZN(n6131) );
  NAND2_X1 U7716 ( .A1(n6142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7717 ( .A(n6129), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U7718 ( .A1(n6371), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6284), .B2(
        n6891), .ZN(n6130) );
  NAND2_X1 U7719 ( .A1(n6829), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6138) );
  INV_X1 U7720 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7721 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  AND2_X1 U7722 ( .A1(n6149), .A2(n6134), .ZN(n7902) );
  NAND2_X1 U7723 ( .A1(n6079), .A2(n7902), .ZN(n6137) );
  NAND2_X1 U7724 ( .A1(n6787), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7725 ( .A1(n6213), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7726 ( .A1(n10298), .A2(n7876), .ZN(n9456) );
  NAND2_X1 U7727 ( .A1(n9439), .A2(n4716), .ZN(n7788) );
  NAND2_X1 U7728 ( .A1(n6139), .A2(n6421), .ZN(n6140) );
  OAI21_X1 U7729 ( .B1(n6141), .B2(n7788), .A(n6140), .ZN(n7895) );
  INV_X1 U7730 ( .A(n7876), .ZN(n9644) );
  NAND2_X1 U7731 ( .A1(n6736), .A2(n6350), .ZN(n6147) );
  INV_X1 U7732 ( .A(n6142), .ZN(n6144) );
  INV_X1 U7733 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7734 ( .A1(n6144), .A2(n6143), .ZN(n6157) );
  NAND2_X1 U7735 ( .A1(n6157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7736 ( .A(n6145), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U7737 ( .A1(n4388), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6284), .B2(
        n10231), .ZN(n6146) );
  NAND2_X1 U7738 ( .A1(n6147), .A2(n6146), .ZN(n9177) );
  NAND2_X1 U7739 ( .A1(n6829), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6154) );
  INV_X1 U7740 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7741 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  AND2_X1 U7742 ( .A1(n6162), .A2(n6150), .ZN(n9184) );
  NAND2_X1 U7743 ( .A1(n6079), .A2(n9184), .ZN(n6153) );
  NAND2_X1 U7744 ( .A1(n6787), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7745 ( .A1(n6213), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6151) );
  OR2_X1 U7746 ( .A1(n9177), .A2(n8054), .ZN(n9457) );
  NAND2_X1 U7747 ( .A1(n9177), .A2(n8054), .ZN(n9462) );
  AND2_X1 U7748 ( .A1(n9457), .A2(n9462), .ZN(n9590) );
  INV_X1 U7749 ( .A(n9590), .ZN(n6155) );
  INV_X1 U7750 ( .A(n8054), .ZN(n9643) );
  NAND2_X1 U7751 ( .A1(n9177), .A2(n9643), .ZN(n6156) );
  NAND2_X1 U7752 ( .A1(n7873), .A2(n6156), .ZN(n8028) );
  NAND2_X1 U7753 ( .A1(n6756), .A2(n6350), .ZN(n6160) );
  NAND2_X1 U7754 ( .A1(n6168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6158) );
  XNOR2_X1 U7755 ( .A(n6158), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9696) );
  AOI22_X1 U7756 ( .A1(n4388), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9696), .B2(
        n6284), .ZN(n6159) );
  NAND2_X1 U7757 ( .A1(n6160), .A2(n6159), .ZN(n8093) );
  NAND2_X1 U7758 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  AND2_X1 U7759 ( .A1(n6172), .A2(n6163), .ZN(n8095) );
  NAND2_X1 U7760 ( .A1(n6079), .A2(n8095), .ZN(n6167) );
  NAND2_X1 U7761 ( .A1(n6829), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7762 ( .A1(n6787), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7763 ( .A1(n6213), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6164) );
  NAND4_X1 U7764 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n9642)
         );
  OR2_X1 U7765 ( .A1(n8093), .A2(n9642), .ZN(n8023) );
  AND2_X1 U7766 ( .A1(n8093), .A2(n9642), .ZN(n8024) );
  AOI21_X2 U7767 ( .B1(n8028), .B2(n8023), .A(n8024), .ZN(n7721) );
  NAND2_X1 U7768 ( .A1(n6738), .A2(n6350), .ZN(n6171) );
  NAND2_X1 U7769 ( .A1(n6178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U7770 ( .A(n6169), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U7771 ( .A1(n6903), .A2(n6284), .B1(n4388), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7772 ( .A1(n6171), .A2(n6170), .ZN(n8077) );
  NAND2_X1 U7773 ( .A1(n6172), .A2(n6872), .ZN(n6173) );
  AND2_X1 U7774 ( .A1(n6183), .A2(n6173), .ZN(n8078) );
  NAND2_X1 U7775 ( .A1(n6079), .A2(n8078), .ZN(n6177) );
  NAND2_X1 U7776 ( .A1(n6829), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7777 ( .A1(n6787), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7778 ( .A1(n6213), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7779 ( .A1(n8077), .A2(n8073), .ZN(n9466) );
  NAND2_X1 U7780 ( .A1(n8077), .A2(n8073), .ZN(n9459) );
  NAND2_X1 U7781 ( .A1(n9466), .A2(n9459), .ZN(n9471) );
  INV_X1 U7782 ( .A(n8073), .ZN(n9641) );
  OR2_X1 U7783 ( .A1(n8077), .A2(n9641), .ZN(n7955) );
  NAND2_X1 U7784 ( .A1(n6746), .A2(n6350), .ZN(n6181) );
  OAI21_X1 U7785 ( .B1(n6178), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7786 ( .A(n6179), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7787 ( .A1(n6967), .A2(n6284), .B1(n4388), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6180) );
  INV_X1 U7788 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7789 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  AND2_X1 U7790 ( .A1(n6200), .A2(n6184), .ZN(n10030) );
  NAND2_X1 U7791 ( .A1(n6079), .A2(n10030), .ZN(n6188) );
  NAND2_X1 U7792 ( .A1(n6829), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7793 ( .A1(n6787), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7794 ( .A1(n6213), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6185) );
  NAND4_X1 U7795 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n9640)
         );
  OR2_X1 U7796 ( .A1(n10031), .A2(n9640), .ZN(n7954) );
  NAND2_X1 U7797 ( .A1(n10031), .A2(n9640), .ZN(n7953) );
  NAND2_X1 U7798 ( .A1(n6772), .A2(n6350), .ZN(n6198) );
  INV_X1 U7799 ( .A(n6189), .ZN(n6190) );
  OR2_X1 U7800 ( .A1(n6191), .A2(n6190), .ZN(n6193) );
  NAND2_X1 U7801 ( .A1(n6193), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6192) );
  MUX2_X1 U7802 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6192), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6196) );
  INV_X1 U7803 ( .A(n6193), .ZN(n6195) );
  INV_X1 U7804 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7805 ( .A1(n6195), .A2(n6194), .ZN(n6207) );
  NAND2_X1 U7806 ( .A1(n6196), .A2(n6207), .ZN(n6970) );
  INV_X1 U7807 ( .A(n6970), .ZN(n7433) );
  AOI22_X1 U7808 ( .A1(n4388), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6284), .B2(
        n7433), .ZN(n6197) );
  NAND2_X1 U7809 ( .A1(n6198), .A2(n6197), .ZN(n8206) );
  NAND2_X1 U7810 ( .A1(n6829), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6205) );
  INV_X1 U7811 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7812 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  AND2_X1 U7813 ( .A1(n6211), .A2(n6201), .ZN(n9207) );
  NAND2_X1 U7814 ( .A1(n6079), .A2(n9207), .ZN(n6204) );
  NAND2_X1 U7815 ( .A1(n6787), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7816 ( .A1(n6213), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7817 ( .A1(n8206), .A2(n10013), .ZN(n9442) );
  NAND2_X1 U7818 ( .A1(n8206), .A2(n10013), .ZN(n9460) );
  INV_X1 U7819 ( .A(n10013), .ZN(n9639) );
  NAND2_X1 U7820 ( .A1(n8206), .A2(n9639), .ZN(n6206) );
  NAND2_X1 U7821 ( .A1(n6779), .A2(n6350), .ZN(n6210) );
  NAND2_X1 U7822 ( .A1(n6207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6208) );
  XNOR2_X1 U7823 ( .A(n6208), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9715) );
  AOI22_X1 U7824 ( .A1(n4388), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6284), .B2(
        n9715), .ZN(n6209) );
  NAND2_X1 U7825 ( .A1(n6829), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7826 ( .A1(n6211), .A2(n9280), .ZN(n6212) );
  AND2_X1 U7827 ( .A1(n6225), .A2(n6212), .ZN(n10020) );
  NAND2_X1 U7828 ( .A1(n6079), .A2(n10020), .ZN(n6216) );
  INV_X2 U7829 ( .A(n6080), .ZN(n6787) );
  NAND2_X1 U7830 ( .A1(n6787), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7831 ( .A1(n6213), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6214) );
  NAND4_X1 U7832 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n9638)
         );
  OR2_X1 U7833 ( .A1(n10141), .A2(n9638), .ZN(n6218) );
  NAND2_X1 U7834 ( .A1(n6793), .A2(n6350), .ZN(n6223) );
  INV_X1 U7835 ( .A(n6427), .ZN(n6220) );
  NAND2_X1 U7836 ( .A1(n6220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6221) );
  XNOR2_X1 U7837 ( .A(n6221), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7641) );
  AOI22_X1 U7838 ( .A1(n4388), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6284), .B2(
        n7641), .ZN(n6222) );
  INV_X1 U7839 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7840 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U7841 ( .A1(n6247), .A2(n6226), .ZN(n10000) );
  INV_X1 U7842 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6227) );
  OAI22_X1 U7843 ( .A1(n10000), .A2(n6355), .B1(n6120), .B2(n6227), .ZN(n6229)
         );
  INV_X1 U7844 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6643) );
  INV_X1 U7845 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10001) );
  OAI22_X1 U7846 ( .A1(n6401), .A2(n6643), .B1(n6080), .B2(n10001), .ZN(n6228)
         );
  AND2_X1 U7847 ( .A1(n10136), .A2(n9637), .ZN(n6230) );
  NAND2_X1 U7848 ( .A1(n6802), .A2(n6350), .ZN(n6234) );
  NAND2_X1 U7849 ( .A1(n6241), .A2(n6232), .ZN(n6282) );
  NAND2_X1 U7850 ( .A1(n6282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6255) );
  XNOR2_X1 U7851 ( .A(n6255), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7941) );
  AOI22_X1 U7852 ( .A1(n4388), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6284), .B2(
        n7941), .ZN(n6233) );
  INV_X1 U7853 ( .A(n6235), .ZN(n6249) );
  INV_X1 U7854 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7855 ( .A1(n6249), .A2(n6236), .ZN(n6237) );
  NAND2_X1 U7856 ( .A1(n6273), .A2(n6237), .ZN(n9966) );
  OR2_X1 U7857 ( .A1(n9966), .A2(n6355), .ZN(n6240) );
  AOI22_X1 U7858 ( .A1(n6829), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6787), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7859 ( .A1(n6213), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6238) );
  OR2_X1 U7860 ( .A1(n10125), .A2(n9974), .ZN(n9487) );
  NAND2_X1 U7861 ( .A1(n10125), .A2(n9974), .ZN(n9492) );
  NAND2_X1 U7862 ( .A1(n9487), .A2(n9492), .ZN(n9955) );
  NAND2_X1 U7863 ( .A1(n6797), .A2(n6350), .ZN(n6245) );
  INV_X1 U7864 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U7865 ( .A1(n6242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6243) );
  XNOR2_X1 U7866 ( .A(n6243), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7769) );
  AOI22_X1 U7867 ( .A1(n4388), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6284), .B2(
        n7769), .ZN(n6244) );
  INV_X1 U7868 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7869 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  NAND2_X1 U7870 ( .A1(n6249), .A2(n6248), .ZN(n9983) );
  AOI22_X1 U7871 ( .A1(n6213), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n6787), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7872 ( .A1(n6829), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6250) );
  OAI211_X1 U7873 ( .C1(n9983), .C2(n6355), .A(n6251), .B(n6250), .ZN(n9636)
         );
  INV_X1 U7874 ( .A(n9636), .ZN(n9997) );
  OR2_X1 U7875 ( .A1(n10128), .A2(n9997), .ZN(n9957) );
  NAND2_X1 U7876 ( .A1(n9957), .A2(n9433), .ZN(n9972) );
  NAND2_X1 U7877 ( .A1(n9955), .A2(n9972), .ZN(n6253) );
  AND2_X1 U7878 ( .A1(n10128), .A2(n9636), .ZN(n9953) );
  INV_X1 U7879 ( .A(n9974), .ZN(n9937) );
  AOI22_X1 U7880 ( .A1(n9955), .A2(n9953), .B1(n9937), .B2(n10125), .ZN(n6252)
         );
  NAND2_X1 U7881 ( .A1(n6975), .A2(n6350), .ZN(n6258) );
  NAND2_X1 U7882 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  NAND2_X1 U7883 ( .A1(n6256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6266) );
  XNOR2_X1 U7884 ( .A(n6266), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8112) );
  AOI22_X1 U7885 ( .A1(n8112), .A2(n6284), .B1(n4388), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7886 ( .A(n6273), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U7887 ( .A1(n9945), .A2(n6079), .ZN(n6263) );
  INV_X1 U7888 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8104) );
  NAND2_X1 U7889 ( .A1(n6787), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7890 ( .A1(n6213), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7891 ( .C1(n8104), .C2(n6401), .A(n6260), .B(n6259), .ZN(n6261)
         );
  INV_X1 U7892 ( .A(n6261), .ZN(n6262) );
  OR2_X1 U7893 ( .A1(n10119), .A2(n9962), .ZN(n9922) );
  NAND2_X1 U7894 ( .A1(n10119), .A2(n9962), .ZN(n9921) );
  INV_X1 U7895 ( .A(n10119), .ZN(n9948) );
  NAND2_X1 U7896 ( .A1(n7091), .A2(n6350), .ZN(n6271) );
  NAND2_X1 U7897 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  NAND2_X1 U7898 ( .A1(n6267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6268) );
  XNOR2_X1 U7899 ( .A(n6268), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9728) );
  INV_X1 U7900 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7252) );
  NOR2_X1 U7901 ( .A1(n9409), .A2(n7252), .ZN(n6269) );
  AOI21_X1 U7902 ( .B1(n9728), .B2(n6284), .A(n6269), .ZN(n6270) );
  INV_X1 U7903 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7938) );
  INV_X1 U7904 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7905 ( .B1(n6273), .B2(n7938), .A(n6272), .ZN(n6274) );
  NAND2_X1 U7906 ( .A1(n6274), .A2(n6288), .ZN(n9930) );
  OR2_X1 U7907 ( .A1(n9930), .A2(n6355), .ZN(n6279) );
  INV_X1 U7908 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U7909 ( .A1(n6829), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7910 ( .A1(n6787), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6275) );
  OAI211_X1 U7911 ( .C1(n6560), .C2(n6120), .A(n6276), .B(n6275), .ZN(n6277)
         );
  INV_X1 U7912 ( .A(n6277), .ZN(n6278) );
  OR2_X1 U7913 ( .A1(n10113), .A2(n9918), .ZN(n9502) );
  NAND2_X1 U7914 ( .A1(n10113), .A2(n9918), .ZN(n9510) );
  NAND2_X1 U7915 ( .A1(n9502), .A2(n9510), .ZN(n9927) );
  INV_X1 U7916 ( .A(n10113), .ZN(n9929) );
  NAND2_X1 U7917 ( .A1(n10111), .A2(n5005), .ZN(n9907) );
  NAND2_X1 U7918 ( .A1(n7307), .A2(n4620), .ZN(n6286) );
  NAND2_X1 U7919 ( .A1(n4436), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6283) );
  AOI22_X1 U7920 ( .A1(n4388), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9740), .B2(
        n6284), .ZN(n6285) );
  INV_X1 U7921 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7922 ( .A1(n6288), .A2(n6287), .ZN(n6289) );
  NAND2_X1 U7923 ( .A1(n6300), .A2(n6289), .ZN(n9910) );
  OR2_X1 U7924 ( .A1(n9910), .A2(n6355), .ZN(n6294) );
  INV_X1 U7925 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U7926 ( .A1(n6787), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7927 ( .A1(n6213), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6290) );
  OAI211_X1 U7928 ( .C1(n9726), .C2(n6401), .A(n6291), .B(n6290), .ZN(n6292)
         );
  INV_X1 U7929 ( .A(n6292), .ZN(n6293) );
  NAND2_X1 U7930 ( .A1(n6294), .A2(n6293), .ZN(n9925) );
  NAND2_X1 U7931 ( .A1(n7489), .A2(n4620), .ZN(n6298) );
  NAND2_X1 U7932 ( .A1(n4388), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6297) );
  INV_X1 U7933 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7934 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NAND2_X1 U7935 ( .A1(n6302), .A2(n6301), .ZN(n9895) );
  OR2_X1 U7936 ( .A1(n9895), .A2(n6355), .ZN(n6307) );
  INV_X1 U7937 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U7938 ( .A1(n6787), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7939 ( .A1(n6213), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6303) );
  OAI211_X1 U7940 ( .C1(n6558), .C2(n6401), .A(n6304), .B(n6303), .ZN(n6305)
         );
  INV_X1 U7941 ( .A(n6305), .ZN(n6306) );
  NAND2_X1 U7942 ( .A1(n10103), .A2(n9917), .ZN(n9514) );
  INV_X1 U7943 ( .A(n9917), .ZN(n9635) );
  NAND2_X1 U7944 ( .A1(n7649), .A2(n4620), .ZN(n6310) );
  NAND2_X1 U7945 ( .A1(n4388), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6309) );
  INV_X1 U7946 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7947 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  AND2_X1 U7948 ( .A1(n6322), .A2(n6313), .ZN(n9858) );
  NAND2_X1 U7949 ( .A1(n9858), .A2(n6079), .ZN(n6319) );
  INV_X1 U7950 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7951 ( .A1(n6213), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7952 ( .A1(n6787), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6314) );
  OAI211_X1 U7953 ( .C1(n6401), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6317)
         );
  INV_X1 U7954 ( .A(n6317), .ZN(n6318) );
  NAND2_X1 U7955 ( .A1(n10092), .A2(n9886), .ZN(n9426) );
  INV_X1 U7956 ( .A(n10092), .ZN(n9860) );
  NAND2_X1 U7957 ( .A1(n7795), .A2(n4620), .ZN(n6321) );
  NAND2_X1 U7958 ( .A1(n4388), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6320) );
  INV_X1 U7959 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U7960 ( .A1(n6322), .A2(n9137), .ZN(n6323) );
  NAND2_X1 U7961 ( .A1(n6342), .A2(n6323), .ZN(n9847) );
  OR2_X1 U7962 ( .A1(n9847), .A2(n6355), .ZN(n6329) );
  INV_X1 U7963 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7964 ( .A1(n6213), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7965 ( .A1(n6787), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6324) );
  OAI211_X1 U7966 ( .C1(n6401), .C2(n6326), .A(n6325), .B(n6324), .ZN(n6327)
         );
  INV_X1 U7967 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U7968 ( .A1(n10089), .A2(n9867), .ZN(n9551) );
  NAND2_X1 U7969 ( .A1(n9347), .A2(n9551), .ZN(n9840) );
  NAND2_X1 U7970 ( .A1(n9841), .A2(n9840), .ZN(n9839) );
  NAND2_X1 U7971 ( .A1(n10089), .A2(n9825), .ZN(n9422) );
  NAND2_X1 U7972 ( .A1(n9839), .A2(n9422), .ZN(n9828) );
  NAND2_X1 U7973 ( .A1(n4388), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6330) );
  XNOR2_X1 U7974 ( .A(n6342), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9829) );
  NAND2_X1 U7975 ( .A1(n9829), .A2(n6079), .ZN(n6336) );
  INV_X1 U7976 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U7977 ( .A1(n6829), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7978 ( .A1(n6213), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6332) );
  OAI211_X1 U7979 ( .C1(n6080), .C2(n9830), .A(n6333), .B(n6332), .ZN(n6334)
         );
  INV_X1 U7980 ( .A(n6334), .ZN(n6335) );
  NAND2_X1 U7981 ( .A1(n6336), .A2(n6335), .ZN(n9633) );
  OR2_X1 U7982 ( .A1(n9836), .A2(n9633), .ZN(n6338) );
  AND2_X1 U7983 ( .A1(n9836), .A2(n9633), .ZN(n6337) );
  AOI21_X2 U7984 ( .B1(n9828), .B2(n6338), .A(n6337), .ZN(n9805) );
  NAND2_X1 U7985 ( .A1(n8165), .A2(n4620), .ZN(n6340) );
  NAND2_X1 U7986 ( .A1(n4388), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6339) );
  NAND2_X2 U7987 ( .A1(n6340), .A2(n6339), .ZN(n10079) );
  INV_X1 U7988 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9259) );
  INV_X1 U7989 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7990 ( .B1(n6342), .B2(n9259), .A(n6341), .ZN(n6343) );
  NAND2_X1 U7991 ( .A1(n6343), .A2(n6353), .ZN(n9212) );
  INV_X1 U7992 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7993 ( .A1(n6787), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U7994 ( .A1(n6213), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6344) );
  OAI211_X1 U7995 ( .C1(n6401), .C2(n6346), .A(n6345), .B(n6344), .ZN(n6347)
         );
  INV_X1 U7996 ( .A(n6347), .ZN(n6348) );
  OR2_X2 U7997 ( .A1(n10079), .A2(n9799), .ZN(n9524) );
  NAND2_X1 U7998 ( .A1(n10079), .A2(n9799), .ZN(n9523) );
  NAND2_X1 U7999 ( .A1(n9524), .A2(n9523), .ZN(n9807) );
  OR2_X1 U8000 ( .A1(n9409), .A2(n10187), .ZN(n6351) );
  INV_X1 U8001 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U8002 ( .A1(n6353), .A2(n8316), .ZN(n6354) );
  NAND2_X1 U8003 ( .A1(n6376), .A2(n6354), .ZN(n9795) );
  INV_X1 U8004 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8005 ( .A1(n6213), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U8006 ( .A1(n6787), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6356) );
  OAI211_X1 U8007 ( .C1(n6401), .C2(n6510), .A(n6357), .B(n6356), .ZN(n6358)
         );
  INV_X1 U8008 ( .A(n6358), .ZN(n6359) );
  NAND2_X1 U8009 ( .A1(n10072), .A2(n9215), .ZN(n9528) );
  INV_X1 U8010 ( .A(n10072), .ZN(n6422) );
  NAND2_X1 U8011 ( .A1(n10072), .A2(n6361), .ZN(n6362) );
  NAND2_X1 U8012 ( .A1(n9095), .A2(n4620), .ZN(n6364) );
  NAND2_X1 U8013 ( .A1(n4388), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6363) );
  XNOR2_X1 U8014 ( .A(n6376), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U8015 ( .A1(n9777), .A2(n6079), .ZN(n6370) );
  INV_X1 U8016 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U8017 ( .A1(n6787), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8018 ( .A1(n6213), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6365) );
  OAI211_X1 U8019 ( .C1(n6367), .C2(n6401), .A(n6366), .B(n6365), .ZN(n6368)
         );
  INV_X1 U8020 ( .A(n6368), .ZN(n6369) );
  AND2_X2 U8021 ( .A1(n6370), .A2(n6369), .ZN(n9800) );
  NAND2_X1 U8022 ( .A1(n10067), .A2(n9800), .ZN(n9532) );
  INV_X1 U8023 ( .A(n10067), .ZN(n9779) );
  NAND2_X1 U8024 ( .A1(n9091), .A2(n4620), .ZN(n6373) );
  NAND2_X1 U8025 ( .A1(n4388), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6372) );
  INV_X1 U8026 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9118) );
  INV_X1 U8027 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6374) );
  OAI21_X1 U8028 ( .B1(n6376), .B2(n9118), .A(n6374), .ZN(n6377) );
  NAND2_X1 U8029 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6375) );
  NAND2_X1 U8030 ( .A1(n6787), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8031 ( .A1(n6213), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6378) );
  OAI211_X1 U8032 ( .C1(n6401), .C2(n6456), .A(n6379), .B(n6378), .ZN(n6380)
         );
  AOI21_X2 U8033 ( .B1(n9166), .B2(n6079), .A(n6380), .ZN(n9769) );
  NAND2_X1 U8034 ( .A1(n9757), .A2(n9769), .ZN(n9764) );
  OAI21_X1 U8035 ( .B1(n6381), .B2(n9605), .A(n10062), .ZN(n8377) );
  OR2_X1 U8036 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  INV_X1 U8037 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6390) );
  OR2_X1 U8038 ( .A1(n7630), .A2(n7065), .ZN(n6395) );
  NAND3_X1 U8039 ( .A1(n6392), .A2(n6393), .A3(n7023), .ZN(n6394) );
  INV_X1 U8040 ( .A(n6398), .ZN(n9761) );
  NAND2_X1 U8041 ( .A1(n9761), .A2(n6079), .ZN(n6404) );
  INV_X1 U8042 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8043 ( .A1(n6787), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U8044 ( .A1(n6213), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6399) );
  OAI211_X1 U8045 ( .C1(n6401), .C2(n6654), .A(n6400), .B(n6399), .ZN(n6402)
         );
  INV_X1 U8046 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U8047 ( .A1(n9629), .A2(n9740), .ZN(n6405) );
  OR2_X1 U8048 ( .A1(n9611), .A2(n9550), .ZN(n9548) );
  XNOR2_X2 U8049 ( .A(n6406), .B(n9364), .ZN(n7081) );
  NAND2_X1 U8050 ( .A1(n7081), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U8051 ( .A1(n9364), .A2(n4386), .ZN(n6407) );
  AND2_X1 U8052 ( .A1(n9439), .A2(n9557), .ZN(n9373) );
  AND2_X1 U8053 ( .A1(n9462), .A2(n9454), .ZN(n9440) );
  INV_X1 U8054 ( .A(n9642), .ZN(n8061) );
  OR2_X1 U8055 ( .A1(n8093), .A2(n8061), .ZN(n9469) );
  AND2_X1 U8056 ( .A1(n9457), .A2(n9469), .ZN(n9441) );
  NAND2_X1 U8057 ( .A1(n8093), .A2(n8061), .ZN(n9461) );
  INV_X1 U8058 ( .A(n9471), .ZN(n6411) );
  NAND2_X1 U8059 ( .A1(n5003), .A2(n6411), .ZN(n7723) );
  NAND2_X1 U8060 ( .A1(n7723), .A2(n9466), .ZN(n7907) );
  INV_X1 U8061 ( .A(n9640), .ZN(n8196) );
  NAND2_X1 U8062 ( .A1(n10031), .A2(n8196), .ZN(n9472) );
  AND2_X1 U8063 ( .A1(n9460), .A2(n9472), .ZN(n9444) );
  OR2_X1 U8064 ( .A1(n10031), .A2(n8196), .ZN(n7908) );
  NAND2_X1 U8065 ( .A1(n9442), .A2(n7908), .ZN(n9468) );
  NAND2_X1 U8066 ( .A1(n9468), .A2(n9460), .ZN(n9478) );
  OR2_X1 U8067 ( .A1(n10141), .A2(n9996), .ZN(n9382) );
  NAND2_X1 U8068 ( .A1(n10141), .A2(n9996), .ZN(n9380) );
  NAND2_X1 U8069 ( .A1(n9382), .A2(n9380), .ZN(n10010) );
  XNOR2_X1 U8070 ( .A(n10136), .B(n10015), .ZN(n9993) );
  OR2_X1 U8071 ( .A1(n10136), .A2(n10015), .ZN(n9450) );
  AND2_X1 U8072 ( .A1(n9487), .A2(n9957), .ZN(n9435) );
  NAND2_X1 U8073 ( .A1(n9510), .A2(n9921), .ZN(n9491) );
  NAND2_X1 U8074 ( .A1(n9502), .A2(n9922), .ZN(n9495) );
  NAND2_X1 U8075 ( .A1(n9495), .A2(n9510), .ZN(n9355) );
  OAI21_X1 U8076 ( .B1(n9935), .B2(n9491), .A(n9355), .ZN(n9914) );
  XNOR2_X1 U8077 ( .A(n10108), .B(n9508), .ZN(n9915) );
  AND2_X1 U8078 ( .A1(n10108), .A2(n9508), .ZN(n9900) );
  NOR2_X1 U8079 ( .A1(n9899), .A2(n9900), .ZN(n6413) );
  XNOR2_X1 U8080 ( .A(n4377), .B(n9866), .ZN(n9884) );
  NAND2_X1 U8081 ( .A1(n4377), .A2(n9866), .ZN(n9862) );
  AND2_X1 U8082 ( .A1(n9426), .A2(n9862), .ZN(n9431) );
  INV_X1 U8083 ( .A(n9840), .ZN(n9849) );
  NAND2_X1 U8084 ( .A1(n9836), .A2(n9852), .ZN(n9393) );
  INV_X1 U8085 ( .A(n9393), .ZN(n9808) );
  NAND2_X2 U8086 ( .A1(n9810), .A2(n9524), .ZN(n9798) );
  INV_X1 U8087 ( .A(n9531), .ZN(n6416) );
  NOR2_X1 U8088 ( .A1(n9605), .A2(n6416), .ZN(n6417) );
  OAI222_X1 U8089 ( .A1(n10014), .A2(n9800), .B1(n10016), .B2(n10051), .C1(
        n10012), .C2(n6420), .ZN(n8375) );
  NOR2_X2 U8090 ( .A1(n7900), .A2(n9177), .ZN(n8031) );
  INV_X1 U8091 ( .A(n8093), .ZN(n8030) );
  NAND2_X1 U8092 ( .A1(n8031), .A2(n8030), .ZN(n8029) );
  NOR2_X4 U8093 ( .A1(n5002), .A2(n10031), .ZN(n7958) );
  INV_X1 U8094 ( .A(n8206), .ZN(n10146) );
  INV_X1 U8095 ( .A(n10128), .ZN(n9986) );
  INV_X1 U8096 ( .A(n10125), .ZN(n9965) );
  INV_X1 U8097 ( .A(n10103), .ZN(n9894) );
  OR2_X2 U8098 ( .A1(n9891), .A2(n4377), .ZN(n9874) );
  OR2_X2 U8099 ( .A1(n9874), .A2(n10092), .ZN(n9856) );
  AND2_X2 U8100 ( .A1(n9814), .A2(n9819), .ZN(n9815) );
  NAND2_X1 U8101 ( .A1(n6392), .A2(n9611), .ZN(n7818) );
  AOI211_X1 U8102 ( .C1(n9757), .C2(n9776), .A(n10320), .B(n9745), .ZN(n8370)
         );
  INV_X1 U8103 ( .A(n7818), .ZN(n7042) );
  AND2_X2 U8104 ( .A1(n7042), .A2(n9623), .ZN(n10299) );
  NAND2_X1 U8105 ( .A1(n6440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U8106 ( .A1(n6434), .A2(n6433), .ZN(n6431) );
  NAND2_X1 U8107 ( .A1(n6431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6432) );
  XNOR2_X1 U8108 ( .A(n6434), .B(n6433), .ZN(n8166) );
  NAND3_X1 U8109 ( .A1(n8166), .A2(P1_B_REG_SCAN_IN), .A3(n7952), .ZN(n6435)
         );
  OR2_X1 U8110 ( .A1(n6760), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6436) );
  INV_X1 U8111 ( .A(n6438), .ZN(n10188) );
  NAND2_X1 U8112 ( .A1(n10188), .A2(n8166), .ZN(n6761) );
  NAND2_X1 U8113 ( .A1(n6436), .A2(n6761), .ZN(n7032) );
  OAI21_X1 U8114 ( .B1(n10133), .B2(n6393), .A(n7032), .ZN(n6454) );
  NAND2_X1 U8115 ( .A1(n4467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6439) );
  MUX2_X1 U8116 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6439), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6441) );
  NAND2_X1 U8117 ( .A1(n6441), .A2(n6440), .ZN(n7796) );
  AND2_X1 U8118 ( .A1(n7796), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6442) );
  NOR2_X1 U8119 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .ZN(
        n6488) );
  NOR4_X1 U8120 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6445) );
  NOR4_X1 U8121 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6444) );
  NOR4_X1 U8122 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6443) );
  NAND4_X1 U8123 ( .A1(n6488), .A2(n6445), .A3(n6444), .A4(n6443), .ZN(n6451)
         );
  NOR4_X1 U8124 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6449) );
  NOR4_X1 U8125 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6448) );
  NOR4_X1 U8126 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6447) );
  NOR4_X1 U8127 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6446) );
  NAND4_X1 U8128 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n6450)
         );
  NOR2_X1 U8129 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  OR2_X1 U8130 ( .A1(n6760), .A2(n6452), .ZN(n7033) );
  NAND2_X1 U8131 ( .A1(n7280), .A2(n6453), .ZN(n7626) );
  NAND2_X1 U8132 ( .A1(n10188), .A2(n7952), .ZN(n10172) );
  INV_X1 U8133 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6458) );
  NAND4_X1 U8134 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .A3(
        n6682), .A4(n6458), .ZN(n6463) );
  AND2_X1 U8135 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7106) );
  NAND3_X1 U8136 ( .A1(n7106), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .ZN(n6462) );
  NAND4_X1 U8137 ( .A1(SI_27_), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_REG2_REG_20__SCAN_IN), .ZN(n6461) );
  INV_X1 U8138 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6459) );
  INV_X1 U8139 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6536) );
  NAND4_X1 U8140 ( .A1(n6459), .A2(n6536), .A3(P2_REG1_REG_31__SCAN_IN), .A4(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n6460) );
  NOR4_X1 U8141 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n6466)
         );
  INV_X1 U8142 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10369) );
  INV_X1 U8143 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9650) );
  AND4_X1 U8144 ( .A1(n9650), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_2__SCAN_IN), .A4(P1_REG2_REG_28__SCAN_IN), .ZN(n6465) );
  INV_X1 U8145 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7581) );
  NOR4_X1 U8146 ( .A1(n6976), .A2(n7581), .A3(P2_IR_REG_6__SCAN_IN), .A4(
        P2_IR_REG_5__SCAN_IN), .ZN(n6464) );
  NAND4_X1 U8147 ( .A1(n6466), .A2(n10369), .A3(n6465), .A4(n6464), .ZN(n6486)
         );
  INV_X1 U8148 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10245) );
  NAND4_X1 U8149 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(n10245), .ZN(n6485) );
  INV_X1 U8150 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10173) );
  NOR4_X1 U8151 ( .A1(n7938), .A2(n10173), .A3(P1_IR_REG_20__SCAN_IN), .A4(
        P1_REG1_REG_29__SCAN_IN), .ZN(n6481) );
  AND2_X1 U8152 ( .A1(n4369), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8618) );
  INV_X1 U8153 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6618) );
  NAND4_X1 U8154 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P2_DATAO_REG_26__SCAN_IN), 
        .A3(P2_REG0_REG_25__SCAN_IN), .A4(n6618), .ZN(n6470) );
  INV_X1 U8155 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6609) );
  NAND4_X1 U8156 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(P2_REG1_REG_15__SCAN_IN), 
        .A3(n6609), .A4(n6658), .ZN(n6469) );
  NAND4_X1 U8157 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(P2_REG0_REG_4__SCAN_IN), 
        .A3(P2_ADDR_REG_11__SCAN_IN), .A4(n8454), .ZN(n6468) );
  NAND4_X1 U8158 ( .A1(SI_8_), .A2(P1_REG3_REG_15__SCAN_IN), .A3(
        P1_REG1_REG_20__SCAN_IN), .A4(n6796), .ZN(n6467) );
  OR4_X1 U8159 ( .A1(n6470), .A2(n6469), .A3(n6468), .A4(n6467), .ZN(n6476) );
  NAND4_X1 U8160 ( .A1(SI_13_), .A2(P2_REG3_REG_9__SCAN_IN), .A3(
        P2_REG0_REG_5__SCAN_IN), .A4(n9137), .ZN(n6472) );
  INV_X1 U8161 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7608) );
  NAND4_X1 U8162 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .A3(P2_B_REG_SCAN_IN), .A4(n7608), .ZN(n6471) );
  NOR2_X1 U8163 ( .A1(n6472), .A2(n6471), .ZN(n6474) );
  INV_X1 U8164 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6836) );
  NOR4_X1 U8165 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(P2_REG0_REG_11__SCAN_IN), 
        .A3(n6510), .A4(n8574), .ZN(n6473) );
  INV_X1 U8166 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10434) );
  NAND4_X1 U8167 ( .A1(n6474), .A2(n6836), .A3(n6473), .A4(
        P2_REG1_REG_0__SCAN_IN), .ZN(n6475) );
  NOR4_X1 U8168 ( .A1(n10248), .A2(P1_IR_REG_19__SCAN_IN), .A3(n6476), .A4(
        n6475), .ZN(n6480) );
  AND4_X1 U8169 ( .A1(n6773), .A2(n6478), .A3(n6477), .A4(SI_3_), .ZN(n6479)
         );
  NAND4_X1 U8170 ( .A1(n6481), .A2(n8618), .A3(n6480), .A4(n6479), .ZN(n6484)
         );
  INV_X1 U8171 ( .A(n6482), .ZN(n6483) );
  NOR4_X1 U8172 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6490)
         );
  NAND4_X1 U8173 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_REG1_REG_13__SCAN_IN), 
        .A3(P2_REG3_REG_16__SCAN_IN), .A4(P2_REG2_REG_22__SCAN_IN), .ZN(n6487)
         );
  NOR3_X1 U8174 ( .A1(SI_20_), .A2(n7252), .A3(n6487), .ZN(n6489) );
  NOR2_X1 U8175 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .ZN(n10488) );
  AND4_X1 U8176 ( .A1(n6490), .A2(n6489), .A3(n10488), .A4(n6488), .ZN(n6497)
         );
  INV_X1 U8177 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10247) );
  NAND4_X1 U8178 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_REG1_REG_6__SCAN_IN), 
        .A3(P1_REG0_REG_4__SCAN_IN), .A4(n10247), .ZN(n6494) );
  INV_X1 U8179 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6517) );
  NAND4_X1 U8180 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P2_REG2_REG_27__SCAN_IN), 
        .A3(SI_31_), .A4(n6517), .ZN(n6493) );
  INV_X1 U8181 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6567) );
  NAND4_X1 U8182 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P2_REG1_REG_20__SCAN_IN), 
        .A3(P2_REG2_REG_14__SCAN_IN), .A4(n6567), .ZN(n6492) );
  NAND4_X1 U8183 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(P1_REG2_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_12__SCAN_IN), .A4(P2_REG1_REG_6__SCAN_IN), .ZN(n6491)
         );
  NOR4_X1 U8184 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n6496)
         );
  NOR4_X1 U8185 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .A3(P1_ADDR_REG_14__SCAN_IN), .A4(P1_ADDR_REG_13__SCAN_IN), .ZN(n6495)
         );
  NAND3_X1 U8186 ( .A1(n6497), .A2(n6496), .A3(n6495), .ZN(n6508) );
  INV_X1 U8187 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6902) );
  NAND4_X1 U8188 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), 
        .A3(n6902), .A4(n6565), .ZN(n6502) );
  INV_X1 U8189 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8622) );
  NAND4_X1 U8190 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(n8622), .ZN(n6501) );
  INV_X1 U8191 ( .A(SI_11_), .ZN(n6648) );
  NAND4_X1 U8192 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(P2_REG0_REG_9__SCAN_IN), 
        .A3(n6648), .A4(n6498), .ZN(n6500) );
  NAND4_X1 U8193 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P2_REG0_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_11__SCAN_IN), .A4(n6646), .ZN(n6499) );
  NOR4_X1 U8194 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n6505)
         );
  INV_X1 U8195 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10372) );
  INV_X1 U8196 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6634) );
  NOR4_X1 U8197 ( .A1(P2_RD_REG_SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .A3(
        n10372), .A4(n6634), .ZN(n6504) );
  INV_X1 U8198 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10367) );
  NOR4_X1 U8199 ( .A1(SI_4_), .A2(P1_REG0_REG_31__SCAN_IN), .A3(n7599), .A4(
        n10367), .ZN(n6503) );
  NAND3_X1 U8200 ( .A1(n6505), .A2(n6504), .A3(n6503), .ZN(n6507) );
  INV_X1 U8201 ( .A(keyinput39), .ZN(n6506) );
  OAI21_X1 U8202 ( .B1(n6508), .B2(n6507), .A(n6506), .ZN(n6716) );
  AOI22_X1 U8203 ( .A1(n10001), .A2(keyinput69), .B1(n6510), .B2(keyinput93), 
        .ZN(n6509) );
  OAI221_X1 U8204 ( .B1(n10001), .B2(keyinput69), .C1(n6510), .C2(keyinput93), 
        .A(n6509), .ZN(n6521) );
  INV_X1 U8205 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6512) );
  AOI22_X1 U8206 ( .A1(n6512), .A2(keyinput61), .B1(n8574), .B2(keyinput90), 
        .ZN(n6511) );
  OAI221_X1 U8207 ( .B1(n6512), .B2(keyinput61), .C1(n8574), .C2(keyinput90), 
        .A(n6511), .ZN(n6520) );
  INV_X1 U8208 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U8209 ( .A1(n6514), .A2(keyinput16), .B1(P1_U3084), .B2(keyinput33), 
        .ZN(n6513) );
  OAI221_X1 U8210 ( .B1(n6514), .B2(keyinput16), .C1(P1_U3084), .C2(keyinput33), .A(n6513), .ZN(n6519) );
  INV_X1 U8211 ( .A(SI_31_), .ZN(n6516) );
  AOI22_X1 U8212 ( .A1(n6517), .A2(keyinput126), .B1(keyinput18), .B2(n6516), 
        .ZN(n6515) );
  OAI221_X1 U8213 ( .B1(n6517), .B2(keyinput126), .C1(n6516), .C2(keyinput18), 
        .A(n6515), .ZN(n6518) );
  NOR4_X1 U8214 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n6533)
         );
  AOI22_X1 U8215 ( .A1(n6523), .A2(keyinput110), .B1(keyinput46), .B2(n6976), 
        .ZN(n6522) );
  OAI221_X1 U8216 ( .B1(n6523), .B2(keyinput110), .C1(n6976), .C2(keyinput46), 
        .A(n6522), .ZN(n6531) );
  INV_X1 U8217 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U8218 ( .A1(n10246), .A2(keyinput87), .B1(n7252), .B2(keyinput65), 
        .ZN(n6524) );
  OAI221_X1 U8219 ( .B1(n10246), .B2(keyinput87), .C1(n7252), .C2(keyinput65), 
        .A(n6524), .ZN(n6530) );
  AOI22_X1 U8220 ( .A1(P2_U3152), .A2(keyinput82), .B1(keyinput99), .B2(n8781), 
        .ZN(n6525) );
  OAI221_X1 U8221 ( .B1(n4369), .B2(keyinput82), .C1(n8781), .C2(keyinput99), 
        .A(n6525), .ZN(n6529) );
  INV_X1 U8222 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6527) );
  AOI22_X1 U8223 ( .A1(n6527), .A2(keyinput100), .B1(keyinput35), .B2(n8480), 
        .ZN(n6526) );
  OAI221_X1 U8224 ( .B1(n6527), .B2(keyinput100), .C1(n8480), .C2(keyinput35), 
        .A(n6526), .ZN(n6528) );
  NOR4_X1 U8225 ( .A1(n6531), .A2(n6530), .A3(n6529), .A4(n6528), .ZN(n6532)
         );
  NAND2_X1 U8226 ( .A1(n6533), .A2(n6532), .ZN(n6715) );
  INV_X1 U8227 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10251) );
  INV_X1 U8228 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n6535) );
  AOI22_X1 U8229 ( .A1(n10251), .A2(keyinput28), .B1(keyinput112), .B2(n6535), 
        .ZN(n6534) );
  OAI221_X1 U8230 ( .B1(n10251), .B2(keyinput28), .C1(n6535), .C2(keyinput112), 
        .A(n6534), .ZN(n6542) );
  XNOR2_X1 U8231 ( .A(SI_8_), .B(keyinput72), .ZN(n6540) );
  XNOR2_X1 U8232 ( .A(SI_27_), .B(keyinput105), .ZN(n6539) );
  XNOR2_X1 U8233 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput7), .ZN(n6538) );
  NAND2_X1 U8234 ( .A1(n6536), .A2(keyinput11), .ZN(n6537) );
  NAND4_X1 U8235 ( .A1(n6540), .A2(n6539), .A3(n6538), .A4(n6537), .ZN(n6541)
         );
  NOR2_X1 U8236 ( .A1(n6542), .A2(n6541), .ZN(n6554) );
  XNOR2_X1 U8237 ( .A(SI_4_), .B(keyinput70), .ZN(n6546) );
  XNOR2_X1 U8238 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput60), .ZN(n6545) );
  XNOR2_X1 U8239 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput78), .ZN(n6544) );
  XNOR2_X1 U8240 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput15), .ZN(n6543) );
  NAND4_X1 U8241 ( .A1(n6546), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(n6552)
         );
  XNOR2_X1 U8242 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput85), .ZN(n6550) );
  XNOR2_X1 U8243 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput30), .ZN(n6549) );
  XNOR2_X1 U8244 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput117), .ZN(n6548) );
  XNOR2_X1 U8245 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput101), .ZN(n6547)
         );
  NAND4_X1 U8246 ( .A1(n6550), .A2(n6549), .A3(n6548), .A4(n6547), .ZN(n6551)
         );
  NOR2_X1 U8247 ( .A1(n6552), .A2(n6551), .ZN(n6553) );
  AND2_X1 U8248 ( .A1(n6554), .A2(n6553), .ZN(n6596) );
  INV_X1 U8249 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6556) );
  INV_X1 U8250 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U8251 ( .A1(n6556), .A2(keyinput6), .B1(keyinput12), .B2(n10439), 
        .ZN(n6555) );
  OAI221_X1 U8252 ( .B1(n6556), .B2(keyinput6), .C1(n10439), .C2(keyinput12), 
        .A(n6555), .ZN(n6563) );
  INV_X1 U8253 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U8254 ( .A1(n10366), .A2(keyinput97), .B1(n6558), .B2(keyinput96), 
        .ZN(n6557) );
  OAI221_X1 U8255 ( .B1(n10366), .B2(keyinput97), .C1(n6558), .C2(keyinput96), 
        .A(n6557), .ZN(n6562) );
  NAND2_X1 U8256 ( .A1(n6560), .A2(keyinput127), .ZN(n6559) );
  OAI221_X1 U8257 ( .B1(n6536), .B2(keyinput11), .C1(n6560), .C2(keyinput127), 
        .A(n6559), .ZN(n6561) );
  NOR3_X1 U8258 ( .A1(n6563), .A2(n6562), .A3(n6561), .ZN(n6595) );
  AOI22_X1 U8259 ( .A1(n6902), .A2(keyinput120), .B1(keyinput37), .B2(n6565), 
        .ZN(n6564) );
  OAI221_X1 U8260 ( .B1(n6902), .B2(keyinput120), .C1(n6565), .C2(keyinput37), 
        .A(n6564), .ZN(n6570) );
  INV_X1 U8261 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7475) );
  AOI22_X1 U8262 ( .A1(n7475), .A2(keyinput27), .B1(n6567), .B2(keyinput98), 
        .ZN(n6566) );
  OAI221_X1 U8263 ( .B1(n7475), .B2(keyinput27), .C1(n6567), .C2(keyinput98), 
        .A(n6566), .ZN(n6569) );
  INV_X1 U8264 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10249) );
  XNOR2_X1 U8265 ( .A(n10249), .B(keyinput80), .ZN(n6568) );
  NOR3_X1 U8266 ( .A1(n6570), .A2(n6569), .A3(n6568), .ZN(n6594) );
  XNOR2_X1 U8267 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput21), .ZN(n6574) );
  XNOR2_X1 U8268 ( .A(P2_REG0_REG_18__SCAN_IN), .B(keyinput26), .ZN(n6573) );
  XNOR2_X1 U8269 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput125), .ZN(n6572) );
  XNOR2_X1 U8270 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput114), .ZN(n6571) );
  NAND4_X1 U8271 ( .A1(n6574), .A2(n6573), .A3(n6572), .A4(n6571), .ZN(n6580)
         );
  XNOR2_X1 U8272 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput84), .ZN(n6578) );
  XNOR2_X1 U8273 ( .A(SI_7_), .B(keyinput111), .ZN(n6577) );
  XNOR2_X1 U8274 ( .A(SI_1_), .B(keyinput86), .ZN(n6576) );
  XNOR2_X1 U8275 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput102), .ZN(n6575) );
  NAND4_X1 U8276 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6579)
         );
  NOR2_X1 U8277 ( .A1(n6580), .A2(n6579), .ZN(n6592) );
  XNOR2_X1 U8278 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput52), .ZN(n6584) );
  XNOR2_X1 U8279 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput79), .ZN(n6583) );
  XNOR2_X1 U8280 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput22), .ZN(n6582) );
  XNOR2_X1 U8281 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput45), .ZN(n6581) );
  NAND4_X1 U8282 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n6590)
         );
  XNOR2_X1 U8283 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput2), .ZN(n6588) );
  XNOR2_X1 U8284 ( .A(SI_3_), .B(keyinput3), .ZN(n6587) );
  XNOR2_X1 U8285 ( .A(P2_REG1_REG_31__SCAN_IN), .B(keyinput1), .ZN(n6586) );
  XNOR2_X1 U8286 ( .A(keyinput77), .B(P1_D_REG_21__SCAN_IN), .ZN(n6585) );
  NAND4_X1 U8287 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6589)
         );
  NOR2_X1 U8288 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  AND2_X1 U8289 ( .A1(n6592), .A2(n6591), .ZN(n6593) );
  NAND4_X1 U8290 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6628)
         );
  INV_X1 U8291 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7445) );
  AOI22_X1 U8292 ( .A1(n7581), .A2(keyinput103), .B1(keyinput58), .B2(n7445), 
        .ZN(n6597) );
  OAI221_X1 U8293 ( .B1(n7581), .B2(keyinput103), .C1(n7445), .C2(keyinput58), 
        .A(n6597), .ZN(n6604) );
  AOI22_X1 U8294 ( .A1(n9137), .A2(keyinput57), .B1(keyinput106), .B2(n6599), 
        .ZN(n6598) );
  OAI221_X1 U8295 ( .B1(n9137), .B2(keyinput57), .C1(n6599), .C2(keyinput106), 
        .A(n6598), .ZN(n6603) );
  AOI22_X1 U8296 ( .A1(n7308), .A2(keyinput10), .B1(keyinput74), .B2(n6601), 
        .ZN(n6600) );
  OAI221_X1 U8297 ( .B1(n7308), .B2(keyinput10), .C1(n6601), .C2(keyinput74), 
        .A(n6600), .ZN(n6602) );
  NOR3_X1 U8298 ( .A1(n6604), .A2(n6603), .A3(n6602), .ZN(n6626) );
  INV_X1 U8299 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U8300 ( .A1(n6836), .A2(keyinput88), .B1(keyinput62), .B2(n9712), 
        .ZN(n6605) );
  OAI221_X1 U8301 ( .B1(n6836), .B2(keyinput88), .C1(n9712), .C2(keyinput62), 
        .A(n6605), .ZN(n6612) );
  AOI22_X1 U8302 ( .A1(n10187), .A2(keyinput13), .B1(keyinput104), .B2(n6607), 
        .ZN(n6606) );
  OAI221_X1 U8303 ( .B1(n10187), .B2(keyinput13), .C1(n6607), .C2(keyinput104), 
        .A(n6606), .ZN(n6611) );
  INV_X1 U8304 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7706) );
  AOI22_X1 U8305 ( .A1(n7706), .A2(keyinput48), .B1(n6609), .B2(keyinput44), 
        .ZN(n6608) );
  OAI221_X1 U8306 ( .B1(n7706), .B2(keyinput48), .C1(n6609), .C2(keyinput44), 
        .A(n6608), .ZN(n6610) );
  NOR3_X1 U8307 ( .A1(n6612), .A2(n6611), .A3(n6610), .ZN(n6625) );
  INV_X1 U8308 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U8309 ( .A1(n6116), .A2(keyinput14), .B1(keyinput83), .B2(n10197), 
        .ZN(n6613) );
  OAI221_X1 U8310 ( .B1(n6116), .B2(keyinput14), .C1(n10197), .C2(keyinput83), 
        .A(n6613), .ZN(n6616) );
  AOI22_X1 U8311 ( .A1(n8316), .A2(keyinput47), .B1(keyinput31), .B2(n10367), 
        .ZN(n6614) );
  OAI221_X1 U8312 ( .B1(n8316), .B2(keyinput47), .C1(n10367), .C2(keyinput31), 
        .A(n6614), .ZN(n6615) );
  NOR2_X1 U8313 ( .A1(n6616), .A2(n6615), .ZN(n6624) );
  AOI22_X1 U8314 ( .A1(n6618), .A2(keyinput42), .B1(keyinput0), .B2(n10434), 
        .ZN(n6617) );
  OAI221_X1 U8315 ( .B1(n6618), .B2(keyinput42), .C1(n10434), .C2(keyinput0), 
        .A(n6617), .ZN(n6622) );
  INV_X1 U8316 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U8317 ( .A1(n6620), .A2(keyinput71), .B1(keyinput118), .B2(n10203), 
        .ZN(n6619) );
  OAI221_X1 U8318 ( .B1(n6620), .B2(keyinput71), .C1(n10203), .C2(keyinput118), 
        .A(n6619), .ZN(n6621) );
  NOR2_X1 U8319 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  NAND4_X1 U8320 ( .A1(n6626), .A2(n6625), .A3(n6624), .A4(n6623), .ZN(n6627)
         );
  NOR2_X1 U8321 ( .A1(n6628), .A2(n6627), .ZN(n6713) );
  INV_X1 U8322 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6630) );
  INV_X1 U8323 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U8324 ( .A1(n6630), .A2(keyinput55), .B1(n10253), .B2(keyinput5), 
        .ZN(n6629) );
  OAI221_X1 U8325 ( .B1(n6630), .B2(keyinput55), .C1(n10253), .C2(keyinput5), 
        .A(n6629), .ZN(n6639) );
  INV_X1 U8326 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6632) );
  INV_X1 U8327 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U8328 ( .A1(n6632), .A2(keyinput109), .B1(keyinput91), .B2(n10479), 
        .ZN(n6631) );
  OAI221_X1 U8329 ( .B1(n6632), .B2(keyinput109), .C1(n10479), .C2(keyinput91), 
        .A(n6631), .ZN(n6638) );
  AOI22_X1 U8330 ( .A1(n6634), .A2(keyinput108), .B1(n5040), .B2(keyinput63), 
        .ZN(n6633) );
  AOI22_X1 U8331 ( .A1(n10372), .A2(keyinput9), .B1(keyinput64), .B2(n8622), 
        .ZN(n6635) );
  OAI221_X1 U8332 ( .B1(n10372), .B2(keyinput9), .C1(n8622), .C2(keyinput64), 
        .A(n6635), .ZN(n6636) );
  NOR4_X1 U8333 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6712)
         );
  INV_X1 U8334 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6641) );
  INV_X1 U8335 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U8336 ( .A1(n6641), .A2(keyinput113), .B1(keyinput41), .B2(n10215), 
        .ZN(n6640) );
  OAI221_X1 U8337 ( .B1(n6641), .B2(keyinput113), .C1(n10215), .C2(keyinput41), 
        .A(n6640), .ZN(n6652) );
  INV_X1 U8338 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7401) );
  AOI22_X1 U8339 ( .A1(n6643), .A2(keyinput115), .B1(keyinput17), .B2(n7401), 
        .ZN(n6642) );
  OAI221_X1 U8340 ( .B1(n6643), .B2(keyinput115), .C1(n7401), .C2(keyinput17), 
        .A(n6642), .ZN(n6651) );
  INV_X1 U8341 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U8342 ( .A1(n6646), .A2(keyinput68), .B1(keyinput94), .B2(n6645), 
        .ZN(n6644) );
  OAI221_X1 U8343 ( .B1(n6646), .B2(keyinput68), .C1(n6645), .C2(keyinput94), 
        .A(n6644), .ZN(n6650) );
  AOI22_X1 U8344 ( .A1(n6872), .A2(keyinput121), .B1(n6648), .B2(keyinput116), 
        .ZN(n6647) );
  OAI221_X1 U8345 ( .B1(n6872), .B2(keyinput121), .C1(n6648), .C2(keyinput116), 
        .A(n6647), .ZN(n6649) );
  NOR4_X1 U8346 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6711)
         );
  AOI22_X1 U8347 ( .A1(n6654), .A2(keyinput56), .B1(keyinput54), .B2(n6459), 
        .ZN(n6653) );
  OAI221_X1 U8348 ( .B1(n6654), .B2(keyinput56), .C1(n6459), .C2(keyinput54), 
        .A(n6653), .ZN(n6661) );
  AOI22_X1 U8349 ( .A1(n8454), .A2(keyinput25), .B1(n6796), .B2(keyinput107), 
        .ZN(n6655) );
  OAI221_X1 U8350 ( .B1(n8454), .B2(keyinput25), .C1(n6796), .C2(keyinput107), 
        .A(n6655), .ZN(n6660) );
  AOI22_X1 U8351 ( .A1(n6658), .A2(keyinput24), .B1(n6657), .B2(keyinput59), 
        .ZN(n6656) );
  OAI221_X1 U8352 ( .B1(n6658), .B2(keyinput24), .C1(n6657), .C2(keyinput59), 
        .A(n6656), .ZN(n6659) );
  NOR3_X1 U8353 ( .A1(n6661), .A2(n6660), .A3(n6659), .ZN(n6680) );
  AOI22_X1 U8354 ( .A1(n9830), .A2(keyinput50), .B1(n10245), .B2(keyinput51), 
        .ZN(n6662) );
  OAI221_X1 U8355 ( .B1(n9830), .B2(keyinput50), .C1(n10245), .C2(keyinput51), 
        .A(n6662), .ZN(n6665) );
  INV_X1 U8356 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U8357 ( .A1(n10335), .A2(keyinput49), .B1(n10247), .B2(keyinput92), 
        .ZN(n6663) );
  OAI221_X1 U8358 ( .B1(n10335), .B2(keyinput49), .C1(n10247), .C2(keyinput92), 
        .A(n6663), .ZN(n6664) );
  NOR2_X1 U8359 ( .A1(n6665), .A2(n6664), .ZN(n6679) );
  INV_X1 U8360 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U8361 ( .A1(n6667), .A2(keyinput29), .B1(keyinput81), .B2(n10413), 
        .ZN(n6666) );
  OAI221_X1 U8362 ( .B1(n6667), .B2(keyinput29), .C1(n10413), .C2(keyinput81), 
        .A(n6666), .ZN(n6671) );
  INV_X1 U8363 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6669) );
  AOI22_X1 U8364 ( .A1(n6383), .A2(keyinput40), .B1(keyinput119), .B2(n6669), 
        .ZN(n6668) );
  OAI221_X1 U8365 ( .B1(n6383), .B2(keyinput40), .C1(n6669), .C2(keyinput119), 
        .A(n6668), .ZN(n6670) );
  NOR2_X1 U8366 ( .A1(n6671), .A2(n6670), .ZN(n6678) );
  INV_X1 U8367 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U8368 ( .A1(n7938), .A2(keyinput123), .B1(keyinput67), .B2(n10371), 
        .ZN(n6672) );
  OAI221_X1 U8369 ( .B1(n7938), .B2(keyinput123), .C1(n10371), .C2(keyinput67), 
        .A(n6672), .ZN(n6676) );
  INV_X1 U8370 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6674) );
  INV_X1 U8371 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U8372 ( .A1(n6674), .A2(keyinput36), .B1(keyinput23), .B2(n10368), 
        .ZN(n6673) );
  OAI221_X1 U8373 ( .B1(n6674), .B2(keyinput36), .C1(n10368), .C2(keyinput23), 
        .A(n6673), .ZN(n6675) );
  NOR2_X1 U8374 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  NAND4_X1 U8375 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n6709)
         );
  INV_X1 U8376 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U8377 ( .A1(n6682), .A2(keyinput124), .B1(n10252), .B2(keyinput122), 
        .ZN(n6681) );
  OAI221_X1 U8378 ( .B1(n6682), .B2(keyinput124), .C1(n10252), .C2(keyinput122), .A(n6681), .ZN(n6686) );
  INV_X1 U8379 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6684) );
  INV_X1 U8380 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U8381 ( .A1(n6684), .A2(keyinput53), .B1(n10370), .B2(keyinput32), 
        .ZN(n6683) );
  OAI221_X1 U8382 ( .B1(n6684), .B2(keyinput53), .C1(n10370), .C2(keyinput32), 
        .A(n6683), .ZN(n6685) );
  NOR2_X1 U8383 ( .A1(n6686), .A2(n6685), .ZN(n6707) );
  AOI22_X1 U8384 ( .A1(n7608), .A2(keyinput34), .B1(n8326), .B2(keyinput38), 
        .ZN(n6687) );
  OAI221_X1 U8385 ( .B1(n7608), .B2(keyinput34), .C1(n8326), .C2(keyinput38), 
        .A(n6687), .ZN(n6690) );
  INV_X1 U8386 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7338) );
  INV_X1 U8387 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U8388 ( .A1(n7338), .A2(keyinput8), .B1(n10250), .B2(keyinput76), 
        .ZN(n6688) );
  OAI221_X1 U8389 ( .B1(n7338), .B2(keyinput8), .C1(n10250), .C2(keyinput76), 
        .A(n6688), .ZN(n6689) );
  NOR2_X1 U8390 ( .A1(n6690), .A2(n6689), .ZN(n6706) );
  INV_X1 U8391 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U8392 ( .A1(n10369), .A2(keyinput43), .B1(n6692), .B2(keyinput4), 
        .ZN(n6691) );
  OAI221_X1 U8393 ( .B1(n10369), .B2(keyinput43), .C1(n6692), .C2(keyinput4), 
        .A(n6691), .ZN(n6696) );
  INV_X1 U8394 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10196) );
  INV_X1 U8395 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U8396 ( .A1(n10196), .A2(keyinput75), .B1(n6694), .B2(keyinput66), 
        .ZN(n6693) );
  OAI221_X1 U8397 ( .B1(n10196), .B2(keyinput75), .C1(n6694), .C2(keyinput66), 
        .A(n6693), .ZN(n6695) );
  NOR2_X1 U8398 ( .A1(n6696), .A2(n6695), .ZN(n6705) );
  AOI22_X1 U8399 ( .A1(n9878), .A2(keyinput89), .B1(n6382), .B2(keyinput95), 
        .ZN(n6697) );
  OAI221_X1 U8400 ( .B1(n9878), .B2(keyinput89), .C1(n6382), .C2(keyinput95), 
        .A(n6697), .ZN(n6703) );
  INV_X1 U8401 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10406) );
  XNOR2_X1 U8402 ( .A(keyinput20), .B(n10406), .ZN(n6699) );
  INV_X1 U8403 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10365) );
  XNOR2_X1 U8404 ( .A(keyinput73), .B(n10365), .ZN(n6698) );
  NOR2_X1 U8405 ( .A1(n6699), .A2(n6698), .ZN(n6701) );
  INV_X1 U8406 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10280) );
  XNOR2_X1 U8407 ( .A(keyinput19), .B(P1_REG0_REG_4__SCAN_IN), .ZN(n6700) );
  OAI211_X1 U8408 ( .C1(n10198), .C2(keyinput39), .A(n6701), .B(n6700), .ZN(
        n6702) );
  NOR2_X1 U8409 ( .A1(n6703), .A2(n6702), .ZN(n6704) );
  NAND4_X1 U8410 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6708)
         );
  NOR2_X1 U8411 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND4_X1 U8412 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6714)
         );
  AOI211_X1 U8413 ( .C1(n6716), .C2(n10198), .A(n6715), .B(n6714), .ZN(n6717)
         );
  XNOR2_X1 U8414 ( .A(n6718), .B(n6717), .ZN(P1_U3551) );
  INV_X1 U8415 ( .A(n6719), .ZN(n6993) );
  INV_X1 U8416 ( .A(n7796), .ZN(n6720) );
  NOR2_X1 U8417 ( .A1(n7279), .A2(n6720), .ZN(n6866) );
  AND2_X2 U8418 ( .A1(n6866), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U8419 ( .A1(n7031), .A2(n7279), .ZN(n6721) );
  NAND2_X1 U8420 ( .A1(n6721), .A2(n7796), .ZN(n6847) );
  NAND2_X1 U8421 ( .A1(n6847), .A2(n6085), .ZN(n6722) );
  NAND2_X1 U8422 ( .A1(n6722), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8423 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6724) );
  INV_X1 U8424 ( .A(n6723), .ZN(n6728) );
  INV_X1 U8425 ( .A(n6863), .ZN(n6933) );
  OAI222_X1 U8426 ( .A1(n10182), .A2(n6724), .B1(n10186), .B2(n6728), .C1(
        P1_U3084), .C2(n6933), .ZN(P1_U3347) );
  INV_X1 U8427 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6726) );
  INV_X1 U8428 ( .A(n6725), .ZN(n6758) );
  INV_X1 U8429 ( .A(n9690), .ZN(n6858) );
  OAI222_X1 U8430 ( .A1(n10182), .A2(n6726), .B1(n10186), .B2(n6758), .C1(
        P1_U3084), .C2(n6858), .ZN(P1_U3349) );
  NAND2_X1 U8431 ( .A1(n4397), .A2(n4369), .ZN(n8378) );
  INV_X1 U8432 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6729) );
  NAND2_X1 U8433 ( .A1(n6727), .A2(P2_U3152), .ZN(n9101) );
  INV_X1 U8434 ( .A(n7242), .ZN(n7250) );
  OAI222_X1 U8435 ( .A1(n8378), .A2(n6729), .B1(n9101), .B2(n6728), .C1(
        P2_U3152), .C2(n7250), .ZN(P2_U3352) );
  INV_X1 U8436 ( .A(n6730), .ZN(n6745) );
  INV_X1 U8437 ( .A(n6856), .ZN(n6945) );
  OAI222_X1 U8438 ( .A1(n10182), .A2(n6731), .B1(n10186), .B2(n6745), .C1(
        P1_U3084), .C2(n6945), .ZN(P1_U3350) );
  INV_X1 U8439 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6733) );
  INV_X1 U8440 ( .A(n6732), .ZN(n6741) );
  INV_X1 U8441 ( .A(n6861), .ZN(n6957) );
  OAI222_X1 U8442 ( .A1(n10182), .A2(n6733), .B1(n10186), .B2(n6741), .C1(
        P1_U3084), .C2(n6957), .ZN(P1_U3348) );
  INV_X1 U8443 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6735) );
  INV_X1 U8444 ( .A(n6734), .ZN(n6743) );
  INV_X1 U8445 ( .A(n6891), .ZN(n6867) );
  OAI222_X1 U8446 ( .A1(n10182), .A2(n6735), .B1(n10186), .B2(n6743), .C1(
        P1_U3084), .C2(n6867), .ZN(P1_U3346) );
  INV_X1 U8447 ( .A(n6736), .ZN(n6750) );
  INV_X1 U8448 ( .A(n10231), .ZN(n10238) );
  OAI222_X1 U8449 ( .A1(n10182), .A2(n6737), .B1(n10186), .B2(n6750), .C1(
        P1_U3084), .C2(n10238), .ZN(P1_U3345) );
  INV_X1 U8450 ( .A(n6738), .ZN(n6766) );
  INV_X1 U8451 ( .A(n8378), .ZN(n9093) );
  AOI22_X1 U8452 ( .A1(n7255), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9093), .ZN(n6739) );
  OAI21_X1 U8453 ( .B1(n6766), .B2(n9101), .A(n6739), .ZN(P2_U3348) );
  AOI22_X1 U8454 ( .A1(n7150), .A2(P2_STATE_REG_SCAN_IN), .B1(n9093), .B2(
        P1_DATAO_REG_5__SCAN_IN), .ZN(n6740) );
  OAI21_X1 U8455 ( .B1(n6741), .B2(n9101), .A(n6740), .ZN(P2_U3353) );
  AOI22_X1 U8456 ( .A1(n7210), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9093), .ZN(n6742) );
  OAI21_X1 U8457 ( .B1(n6743), .B2(n9101), .A(n6742), .ZN(P2_U3351) );
  INV_X1 U8458 ( .A(n7131), .ZN(n6744) );
  OAI222_X1 U8459 ( .A1(n9099), .A2(n4516), .B1(n9101), .B2(n6745), .C1(n4369), 
        .C2(n6744), .ZN(P2_U3355) );
  INV_X1 U8460 ( .A(n6746), .ZN(n6748) );
  INV_X1 U8461 ( .A(n10182), .ZN(n10176) );
  AOI22_X1 U8462 ( .A1(n6967), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10176), .ZN(n6747) );
  OAI21_X1 U8463 ( .B1(n6748), .B2(n10186), .A(n6747), .ZN(P1_U3342) );
  CLKBUF_X1 U8464 ( .A(n9101), .Z(n7652) );
  INV_X1 U8465 ( .A(n7410), .ZN(n7402) );
  OAI222_X1 U8466 ( .A1(n8378), .A2(n6749), .B1(n7652), .B2(n6748), .C1(n7402), 
        .C2(n4369), .ZN(P2_U3347) );
  INV_X1 U8467 ( .A(n7224), .ZN(n7219) );
  OAI222_X1 U8468 ( .A1(n9099), .A2(n6751), .B1(n7652), .B2(n6750), .C1(
        P2_U3152), .C2(n7219), .ZN(P2_U3350) );
  INV_X1 U8469 ( .A(n7182), .ZN(n6753) );
  OAI222_X1 U8470 ( .A1(n6753), .A2(P2_U3152), .B1(n7652), .B2(n6768), .C1(
        n6752), .C2(n8378), .ZN(P2_U3356) );
  INV_X1 U8471 ( .A(n7108), .ZN(n6755) );
  OAI222_X1 U8472 ( .A1(n6755), .A2(n4369), .B1(n7652), .B2(n6770), .C1(n6754), 
        .C2(n8378), .ZN(P2_U3357) );
  INV_X1 U8473 ( .A(n6756), .ZN(n6764) );
  INV_X1 U8474 ( .A(n7424), .ZN(n7422) );
  OAI222_X1 U8475 ( .A1(n8378), .A2(n6757), .B1(n7652), .B2(n6764), .C1(n7422), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8476 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6759) );
  INV_X1 U8477 ( .A(n7195), .ZN(n7203) );
  OAI222_X1 U8478 ( .A1(n6759), .A2(n8378), .B1(P2_U3152), .B2(n7203), .C1(
        n7652), .C2(n6758), .ZN(P2_U3354) );
  INV_X1 U8479 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6763) );
  INV_X1 U8480 ( .A(n6761), .ZN(n6762) );
  AOI22_X1 U8481 ( .A1(n10255), .A2(n6763), .B1(n7286), .B2(n6762), .ZN(
        P1_U3441) );
  INV_X1 U8482 ( .A(n9696), .ZN(n6879) );
  OAI222_X1 U8483 ( .A1(n10182), .A2(n6765), .B1(n6879), .B2(P1_U3084), .C1(
        n10186), .C2(n6764), .ZN(P1_U3344) );
  INV_X1 U8484 ( .A(n6903), .ZN(n6881) );
  OAI222_X1 U8485 ( .A1(n10182), .A2(n6767), .B1(n6881), .B2(P1_U3084), .C1(
        n10186), .C2(n6766), .ZN(P1_U3343) );
  OAI222_X1 U8486 ( .A1(n10182), .A2(n6769), .B1(n10186), .B2(n6768), .C1(
        P1_U3084), .C2(n6070), .ZN(P1_U3351) );
  OAI222_X1 U8487 ( .A1(n10182), .A2(n6771), .B1(n10186), .B2(n6770), .C1(
        P1_U3084), .C2(n6849), .ZN(P1_U3352) );
  INV_X1 U8488 ( .A(n6772), .ZN(n6774) );
  OAI222_X1 U8489 ( .A1(n10182), .A2(n6773), .B1(n10186), .B2(n6774), .C1(
        P1_U3084), .C2(n6970), .ZN(P1_U3341) );
  INV_X1 U8490 ( .A(n7451), .ZN(n7407) );
  OAI222_X1 U8491 ( .A1(n8378), .A2(n6775), .B1(n7652), .B2(n6774), .C1(n4369), 
        .C2(n7407), .ZN(P2_U3346) );
  INV_X1 U8492 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6778) );
  INV_X1 U8493 ( .A(n8646), .ZN(n6776) );
  NAND2_X1 U8494 ( .A1(n6776), .A2(P2_U3966), .ZN(n6777) );
  OAI21_X1 U8495 ( .B1(n6778), .B2(P2_U3966), .A(n6777), .ZN(P2_U3583) );
  INV_X1 U8496 ( .A(n6779), .ZN(n6781) );
  AOI22_X1 U8497 ( .A1(n9715), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10176), .ZN(n6780) );
  OAI21_X1 U8498 ( .B1(n6781), .B2(n10186), .A(n6780), .ZN(P1_U3340) );
  INV_X1 U8499 ( .A(n7458), .ZN(n7465) );
  OAI222_X1 U8500 ( .A1(n8378), .A2(n6782), .B1(n7652), .B2(n6781), .C1(n7465), 
        .C2(n4369), .ZN(P2_U3345) );
  INV_X1 U8501 ( .A(n7798), .ZN(n6995) );
  NAND2_X1 U8502 ( .A1(n10363), .A2(n6995), .ZN(n6783) );
  NAND2_X1 U8503 ( .A1(n6784), .A2(n6783), .ZN(n8643) );
  NOR2_X1 U8504 ( .A1(n10347), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8505 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8506 ( .A1(P1_U4006), .A2(n7614), .ZN(n6785) );
  OAI21_X1 U8507 ( .B1(P1_U4006), .B2(n6786), .A(n6785), .ZN(P1_U3555) );
  INV_X1 U8508 ( .A(P1_U4006), .ZN(n6792) );
  NAND2_X1 U8509 ( .A1(n6829), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8510 ( .A1(n6787), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8511 ( .A1(n6213), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6788) );
  AND3_X1 U8512 ( .A1(n6790), .A2(n6789), .A3(n6788), .ZN(n9768) );
  NAND2_X1 U8513 ( .A1(n6792), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6791) );
  OAI21_X1 U8514 ( .B1(n6792), .B2(n9768), .A(n6791), .ZN(P1_U3585) );
  INV_X1 U8515 ( .A(n6793), .ZN(n6795) );
  INV_X1 U8516 ( .A(n7657), .ZN(n7484) );
  OAI222_X1 U8517 ( .A1(n9099), .A2(n6794), .B1(n7652), .B2(n6795), .C1(n7484), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8518 ( .A(n7641), .ZN(n7438) );
  OAI222_X1 U8519 ( .A1(n10182), .A2(n6796), .B1(n7438), .B2(P1_U3084), .C1(
        n10186), .C2(n6795), .ZN(P1_U3339) );
  INV_X1 U8520 ( .A(n6797), .ZN(n6799) );
  INV_X1 U8521 ( .A(n7769), .ZN(n7763) );
  OAI222_X1 U8522 ( .A1(n10182), .A2(n6798), .B1(n10186), .B2(n6799), .C1(
        P1_U3084), .C2(n7763), .ZN(P1_U3338) );
  INV_X1 U8523 ( .A(n7666), .ZN(n7705) );
  OAI222_X1 U8524 ( .A1(n9099), .A2(n6800), .B1(n7652), .B2(n6799), .C1(
        P2_U3152), .C2(n7705), .ZN(P2_U3343) );
  NAND2_X1 U8525 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n8610), .ZN(n6801) );
  OAI21_X1 U8526 ( .B1(n8327), .B2(n8610), .A(n6801), .ZN(P2_U3582) );
  INV_X1 U8527 ( .A(n6802), .ZN(n6827) );
  AOI22_X1 U8528 ( .A1(n7941), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10176), .ZN(n6803) );
  OAI21_X1 U8529 ( .B1(n6827), .B2(n10186), .A(n6803), .ZN(P1_U3337) );
  NOR2_X1 U8530 ( .A1(n10363), .A2(n6804), .ZN(n7316) );
  NAND3_X1 U8531 ( .A1(n6806), .A2(n7316), .A3(n6805), .ZN(n6808) );
  INV_X1 U8532 ( .A(n7013), .ZN(n7317) );
  INV_X1 U8533 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6826) );
  INV_X1 U8534 ( .A(n7045), .ZN(n6812) );
  NOR2_X1 U8535 ( .A1(n6812), .A2(n6811), .ZN(n7345) );
  AOI21_X1 U8536 ( .B1(n6812), .B2(n6811), .A(n7345), .ZN(n8937) );
  XNOR2_X1 U8537 ( .A(n7318), .B(n5058), .ZN(n6813) );
  NAND2_X1 U8538 ( .A1(n6813), .A2(n8874), .ZN(n8890) );
  NAND2_X1 U8539 ( .A1(n7507), .A2(n8640), .ZN(n6814) );
  OR2_X1 U8540 ( .A1(n6814), .A2(n5058), .ZN(n10429) );
  INV_X1 U8541 ( .A(n7335), .ZN(n6820) );
  INV_X1 U8542 ( .A(n6809), .ZN(n6818) );
  INV_X1 U8543 ( .A(n6815), .ZN(n6817) );
  OAI21_X1 U8544 ( .B1(n5831), .B2(n6818), .A(n8902), .ZN(n6819) );
  AOI21_X1 U8545 ( .B1(n6820), .B2(n7045), .A(n6819), .ZN(n6822) );
  OAI22_X1 U8546 ( .A1(n10380), .A2(n8793), .B1(n5754), .B2(n8795), .ZN(n6821)
         );
  NOR2_X1 U8547 ( .A1(n6822), .A2(n6821), .ZN(n8946) );
  NOR2_X2 U8548 ( .A1(n8938), .A2(n10381), .ZN(n7353) );
  AND2_X1 U8549 ( .A1(n8938), .A2(n10381), .ZN(n6823) );
  NOR2_X1 U8550 ( .A1(n7353), .A2(n6823), .ZN(n8943) );
  AOI22_X1 U8551 ( .A1(n8943), .A2(n10424), .B1(n10423), .B2(n8938), .ZN(n6824) );
  OAI211_X1 U8552 ( .C1(n8937), .C2(n10418), .A(n8946), .B(n6824), .ZN(n7015)
         );
  NAND2_X1 U8553 ( .A1(n7015), .A2(n10433), .ZN(n6825) );
  OAI21_X1 U8554 ( .B1(n10433), .B2(n6826), .A(n6825), .ZN(P2_U3454) );
  OAI222_X1 U8555 ( .A1(n8378), .A2(n6828), .B1(n7652), .B2(n6827), .C1(n8621), 
        .C2(n4369), .ZN(P2_U3342) );
  INV_X1 U8556 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8557 ( .A1(n6829), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8558 ( .A1(n6787), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U8559 ( .A1(n6213), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6830) );
  INV_X1 U8560 ( .A(n9749), .ZN(n6833) );
  NAND2_X1 U8561 ( .A1(P1_U4006), .A2(n6833), .ZN(n6834) );
  OAI21_X1 U8562 ( .B1(P1_U4006), .B2(n6835), .A(n6834), .ZN(P1_U3586) );
  MUX2_X1 U8563 ( .A(n6836), .B(P1_REG2_REG_4__SCAN_IN), .S(n9690), .Z(n9685)
         );
  INV_X1 U8564 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6837) );
  XNOR2_X1 U8565 ( .A(n9671), .B(n6837), .ZN(n9674) );
  XNOR2_X1 U8566 ( .A(n6849), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6978) );
  AND2_X1 U8567 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9661) );
  NAND2_X1 U8568 ( .A1(n6978), .A2(n9661), .ZN(n6977) );
  INV_X1 U8569 ( .A(n6849), .ZN(n6988) );
  NAND2_X1 U8570 ( .A1(n6988), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8571 ( .A1(n6977), .A2(n6838), .ZN(n9673) );
  NAND2_X1 U8572 ( .A1(n9674), .A2(n9673), .ZN(n9672) );
  NAND2_X1 U8573 ( .A1(n9671), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U8574 ( .A1(n9672), .A2(n6839), .ZN(n6941) );
  INV_X1 U8575 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6840) );
  XNOR2_X1 U8576 ( .A(n6856), .B(n6840), .ZN(n6942) );
  NAND2_X1 U8577 ( .A1(n6941), .A2(n6942), .ZN(n6940) );
  NAND2_X1 U8578 ( .A1(n6856), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8579 ( .A1(n6940), .A2(n6841), .ZN(n9686) );
  OR2_X1 U8580 ( .A1(n9685), .A2(n9686), .ZN(n9688) );
  NAND2_X1 U8581 ( .A1(n6858), .A2(n6836), .ZN(n6842) );
  AND2_X1 U8582 ( .A1(n9688), .A2(n6842), .ZN(n6953) );
  INV_X1 U8583 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7783) );
  XNOR2_X1 U8584 ( .A(n6861), .B(n7783), .ZN(n6954) );
  NAND2_X1 U8585 ( .A1(n6953), .A2(n6954), .ZN(n6952) );
  NAND2_X1 U8586 ( .A1(n6861), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8587 ( .A1(n6952), .A2(n6843), .ZN(n6929) );
  INV_X1 U8588 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6844) );
  MUX2_X1 U8589 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6844), .S(n6863), .Z(n6930)
         );
  NAND2_X1 U8590 ( .A1(n6929), .A2(n6930), .ZN(n6928) );
  NAND2_X1 U8591 ( .A1(n6863), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8592 ( .A1(n6928), .A2(n6845), .ZN(n6890) );
  XOR2_X1 U8593 ( .A(n6891), .B(P1_REG2_REG_7__SCAN_IN), .Z(n6846) );
  XNOR2_X1 U8594 ( .A(n6890), .B(n6846), .ZN(n6871) );
  NAND2_X1 U8595 ( .A1(n6847), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9655) );
  OR2_X1 U8596 ( .A1(n9655), .A2(n10184), .ZN(n9734) );
  INV_X1 U8597 ( .A(n10184), .ZN(n9652) );
  NAND2_X1 U8598 ( .A1(n6988), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6851) );
  INV_X1 U8599 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U8600 ( .A1(n6849), .A2(n10329), .ZN(n6850) );
  AND2_X1 U8601 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6983) );
  NAND2_X1 U8602 ( .A1(n6982), .A2(n6983), .ZN(n6981) );
  NAND2_X1 U8603 ( .A1(n6981), .A2(n6851), .ZN(n9667) );
  INV_X1 U8604 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6852) );
  XNOR2_X1 U8605 ( .A(n9671), .B(n6852), .ZN(n9666) );
  NAND2_X1 U8606 ( .A1(n9667), .A2(n9666), .ZN(n6854) );
  NAND2_X1 U8607 ( .A1(n9671), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8608 ( .A1(n6854), .A2(n6853), .ZN(n6935) );
  INV_X1 U8609 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6855) );
  MUX2_X1 U8610 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6855), .S(n6856), .Z(n6936)
         );
  NAND2_X1 U8611 ( .A1(n6935), .A2(n6936), .ZN(n6934) );
  NAND2_X1 U8612 ( .A1(n6856), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8613 ( .A1(n6934), .A2(n6857), .ZN(n9679) );
  MUX2_X1 U8614 ( .A(n10332), .B(P1_REG1_REG_4__SCAN_IN), .S(n9690), .Z(n9678)
         );
  NAND2_X1 U8615 ( .A1(n6858), .A2(n10332), .ZN(n6859) );
  INV_X1 U8616 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6860) );
  MUX2_X1 U8617 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6860), .S(n6861), .Z(n6947)
         );
  NAND2_X1 U8618 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  NAND2_X1 U8619 ( .A1(n6861), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6862) );
  MUX2_X1 U8620 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10335), .S(n6863), .Z(n6922)
         );
  NAND2_X1 U8621 ( .A1(n6923), .A2(n6922), .ZN(n6921) );
  OR2_X1 U8622 ( .A1(n6863), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U8623 ( .A1(n6921), .A2(n6864), .ZN(n6877) );
  INV_X1 U8624 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10337) );
  XNOR2_X1 U8625 ( .A(n6891), .B(n10337), .ZN(n6865) );
  XNOR2_X1 U8626 ( .A(n6877), .B(n6865), .ZN(n6869) );
  AND2_X1 U8627 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7756) );
  OAI22_X1 U8628 ( .A1(n10239), .A2(n6867), .B1(n10244), .B2(n10197), .ZN(
        n6868) );
  AOI211_X1 U8629 ( .C1(n10235), .C2(n6869), .A(n7756), .B(n6868), .ZN(n6870)
         );
  OAI21_X1 U8630 ( .B1(n6871), .B2(n10228), .A(n6870), .ZN(P1_U3248) );
  INV_X1 U8631 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6874) );
  NOR2_X1 U8632 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6872), .ZN(n8076) );
  INV_X1 U8633 ( .A(n8076), .ZN(n6873) );
  OAI21_X1 U8634 ( .B1(n10244), .B2(n6874), .A(n6873), .ZN(n6888) );
  NAND2_X1 U8635 ( .A1(n6891), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U8636 ( .A1(n6891), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6875) );
  AOI22_X1 U8637 ( .A1(n6878), .A2(n10231), .B1(n10233), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n9701) );
  INV_X1 U8638 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10342) );
  MUX2_X1 U8639 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10342), .S(n9696), .Z(n9700)
         );
  NAND2_X1 U8640 ( .A1(n6879), .A2(n10342), .ZN(n6884) );
  INV_X1 U8641 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8642 ( .A1(n6881), .A2(n6880), .ZN(n6909) );
  NAND2_X1 U8643 ( .A1(n6903), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U8644 ( .A1(n6909), .A2(n6882), .ZN(n6883) );
  INV_X1 U8645 ( .A(n6913), .ZN(n6886) );
  NAND3_X1 U8646 ( .A1(n9699), .A2(n6884), .A3(n6883), .ZN(n6885) );
  AOI21_X1 U8647 ( .B1(n6886), .B2(n6885), .A(n9735), .ZN(n6887) );
  AOI211_X1 U8648 ( .C1(n9716), .C2(n6903), .A(n6888), .B(n6887), .ZN(n6901)
         );
  OR2_X1 U8649 ( .A1(n6891), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U8650 ( .A1(n6890), .A2(n6889), .ZN(n6893) );
  NAND2_X1 U8651 ( .A1(n6891), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8652 ( .A1(n6893), .A2(n6892), .ZN(n10226) );
  AND2_X1 U8653 ( .A1(n10231), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10223) );
  OR2_X1 U8654 ( .A1(n10226), .A2(n10223), .ZN(n6894) );
  OR2_X1 U8655 ( .A1(n10231), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10227) );
  AND2_X1 U8656 ( .A1(n6894), .A2(n10227), .ZN(n10224) );
  INV_X1 U8657 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6895) );
  XNOR2_X1 U8658 ( .A(n9696), .B(n6895), .ZN(n9698) );
  NAND2_X1 U8659 ( .A1(n10224), .A2(n9698), .ZN(n9697) );
  NAND2_X1 U8660 ( .A1(n9696), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8661 ( .A1(n9697), .A2(n6896), .ZN(n6899) );
  INV_X1 U8662 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6897) );
  XNOR2_X1 U8663 ( .A(n6903), .B(n6897), .ZN(n6898) );
  NAND2_X1 U8664 ( .A1(n6899), .A2(n6898), .ZN(n6905) );
  OAI211_X1 U8665 ( .C1(n6899), .C2(n6898), .A(n6905), .B(n9733), .ZN(n6900)
         );
  NAND2_X1 U8666 ( .A1(n6901), .A2(n6900), .ZN(P1_U3251) );
  MUX2_X1 U8667 ( .A(n6902), .B(P1_REG2_REG_11__SCAN_IN), .S(n6967), .Z(n6908)
         );
  NAND2_X1 U8668 ( .A1(n6903), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8669 ( .A1(n6905), .A2(n6904), .ZN(n6907) );
  INV_X1 U8670 ( .A(n6969), .ZN(n6906) );
  AOI21_X1 U8671 ( .B1(n6908), .B2(n6907), .A(n6906), .ZN(n6920) );
  INV_X1 U8672 ( .A(n6909), .ZN(n6912) );
  OR2_X1 U8673 ( .A1(n6967), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U8674 ( .A1(n6967), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6910) );
  AND2_X1 U8675 ( .A1(n6961), .A2(n6910), .ZN(n6911) );
  INV_X1 U8676 ( .A(n6962), .ZN(n6915) );
  NOR3_X1 U8677 ( .A1(n6913), .A2(n6912), .A3(n6911), .ZN(n6914) );
  OAI21_X1 U8678 ( .B1(n6915), .B2(n6914), .A(n10235), .ZN(n6919) );
  INV_X1 U8679 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8680 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9303) );
  OAI21_X1 U8681 ( .B1(n10244), .B2(n6916), .A(n9303), .ZN(n6917) );
  AOI21_X1 U8682 ( .B1(n6967), .B2(n9716), .A(n6917), .ZN(n6918) );
  OAI211_X1 U8683 ( .C1(n6920), .C2(n10228), .A(n6919), .B(n6918), .ZN(
        P1_U3252) );
  OAI21_X1 U8684 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(n6927) );
  NAND2_X1 U8685 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7854) );
  INV_X1 U8686 ( .A(n7854), .ZN(n6926) );
  INV_X1 U8687 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8688 ( .A1(n10244), .A2(n6924), .ZN(n6925) );
  AOI211_X1 U8689 ( .C1(n10235), .C2(n6927), .A(n6926), .B(n6925), .ZN(n6932)
         );
  OAI211_X1 U8690 ( .C1(n6930), .C2(n6929), .A(n9733), .B(n6928), .ZN(n6931)
         );
  OAI211_X1 U8691 ( .C1(n10239), .C2(n6933), .A(n6932), .B(n6931), .ZN(
        P1_U3247) );
  INV_X1 U8692 ( .A(n10244), .ZN(n9684) );
  OAI21_X1 U8693 ( .B1(n6936), .B2(n6935), .A(n6934), .ZN(n6938) );
  NOR2_X1 U8694 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6078), .ZN(n7291) );
  INV_X1 U8695 ( .A(n7291), .ZN(n6937) );
  OAI21_X1 U8696 ( .B1(n9735), .B2(n6938), .A(n6937), .ZN(n6939) );
  AOI21_X1 U8697 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(n9684), .A(n6939), .ZN(
        n6944) );
  OAI211_X1 U8698 ( .C1(n6942), .C2(n6941), .A(n9733), .B(n6940), .ZN(n6943)
         );
  OAI211_X1 U8699 ( .C1(n10239), .C2(n6945), .A(n6944), .B(n6943), .ZN(
        P1_U3244) );
  OAI21_X1 U8700 ( .B1(n6948), .B2(n6947), .A(n6946), .ZN(n6950) );
  NOR2_X1 U8701 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6116), .ZN(n7700) );
  INV_X1 U8702 ( .A(n7700), .ZN(n6949) );
  OAI21_X1 U8703 ( .B1(n9735), .B2(n6950), .A(n6949), .ZN(n6951) );
  AOI21_X1 U8704 ( .B1(n9684), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6951), .ZN(
        n6956) );
  OAI211_X1 U8705 ( .C1(n6954), .C2(n6953), .A(n9733), .B(n6952), .ZN(n6955)
         );
  OAI211_X1 U8706 ( .C1(n10239), .C2(n6957), .A(n6956), .B(n6955), .ZN(
        P1_U3246) );
  INV_X1 U8707 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6958) );
  NAND2_X1 U8708 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9203) );
  OAI21_X1 U8709 ( .B1(n10244), .B2(n6958), .A(n9203), .ZN(n6966) );
  INV_X1 U8710 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U8711 ( .A1(n6970), .A2(n6959), .ZN(n7439) );
  OAI21_X1 U8712 ( .B1(n6970), .B2(n6959), .A(n7439), .ZN(n6960) );
  AOI21_X1 U8713 ( .B1(n6962), .B2(n6961), .A(n6960), .ZN(n9709) );
  INV_X1 U8714 ( .A(n9709), .ZN(n6964) );
  NAND3_X1 U8715 ( .A1(n6962), .A2(n6961), .A3(n6960), .ZN(n6963) );
  AOI21_X1 U8716 ( .B1(n6964), .B2(n6963), .A(n9735), .ZN(n6965) );
  AOI211_X1 U8717 ( .C1(n9716), .C2(n7433), .A(n6966), .B(n6965), .ZN(n6974)
         );
  OR2_X1 U8718 ( .A1(n6967), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6968) );
  XNOR2_X1 U8719 ( .A(n6970), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8720 ( .A1(n6972), .A2(n6971), .ZN(n7435) );
  OAI211_X1 U8721 ( .C1(n6972), .C2(n6971), .A(n7435), .B(n9733), .ZN(n6973)
         );
  NAND2_X1 U8722 ( .A1(n6974), .A2(n6973), .ZN(P1_U3253) );
  INV_X1 U8723 ( .A(n6975), .ZN(n6990) );
  OAI222_X1 U8724 ( .A1(n8378), .A2(n6976), .B1(n7652), .B2(n6990), .C1(n10352), .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U8725 ( .B1(n6978), .B2(n9661), .A(n6977), .ZN(n6980) );
  INV_X1 U8726 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6979) );
  OAI22_X1 U8727 ( .A1(n10228), .A2(n6980), .B1(n10244), .B2(n6979), .ZN(n6987) );
  INV_X1 U8728 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6985) );
  OAI211_X1 U8729 ( .C1(n6983), .C2(n6982), .A(n10235), .B(n6981), .ZN(n6984)
         );
  OAI21_X1 U8730 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6985), .A(n6984), .ZN(n6986) );
  AOI211_X1 U8731 ( .C1(n9716), .C2(n6988), .A(n6987), .B(n6986), .ZN(n6989)
         );
  INV_X1 U8732 ( .A(n6989), .ZN(P1_U3242) );
  INV_X1 U8733 ( .A(n8112), .ZN(n8103) );
  OAI222_X1 U8734 ( .A1(n10182), .A2(n6991), .B1(n8103), .B2(P1_U3084), .C1(
        n10186), .C2(n6990), .ZN(P1_U3336) );
  INV_X1 U8735 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U8736 ( .A(n7107), .B(n7106), .ZN(n7012) );
  INV_X1 U8737 ( .A(n6992), .ZN(n6996) );
  NOR2_X1 U8738 ( .A1(n6999), .A2(P2_U3152), .ZN(n9092) );
  NAND2_X1 U8739 ( .A1(n6993), .A2(n9092), .ZN(n6994) );
  OAI211_X1 U8740 ( .C1(n10363), .C2(n6996), .A(n6995), .B(n6994), .ZN(n7005)
         );
  NAND2_X1 U8741 ( .A1(n6997), .A2(n8610), .ZN(n7000) );
  NOR2_X1 U8742 ( .A1(n6999), .A2(n9097), .ZN(n6998) );
  NAND2_X1 U8743 ( .A1(n7000), .A2(n6998), .ZN(n8637) );
  INV_X1 U8744 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7001) );
  INV_X1 U8745 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7278) );
  OAI22_X1 U8746 ( .A1(n8643), .A2(n7001), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7278), .ZN(n7010) );
  INV_X1 U8747 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7017) );
  MUX2_X1 U8748 ( .A(n7017), .B(P2_REG1_REG_1__SCAN_IN), .S(n7108), .Z(n7008)
         );
  AND2_X1 U8749 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n7002) );
  INV_X1 U8750 ( .A(n7002), .ZN(n7007) );
  MUX2_X1 U8751 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n7017), .S(n7108), .Z(n7003)
         );
  NAND2_X1 U8752 ( .A1(n7003), .A2(n7002), .ZN(n7176) );
  INV_X1 U8753 ( .A(n7176), .ZN(n7006) );
  AOI211_X1 U8754 ( .C1(n7008), .C2(n7007), .A(n7006), .B(n7719), .ZN(n7009)
         );
  AOI211_X1 U8755 ( .C1(n10354), .C2(n7108), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OAI21_X1 U8756 ( .B1(n7012), .B2(n8637), .A(n7011), .ZN(P2_U3246) );
  NAND2_X1 U8757 ( .A1(n7015), .A2(n10444), .ZN(n7016) );
  OAI21_X1 U8758 ( .B1(n10444), .B2(n7017), .A(n7016), .ZN(P2_U3521) );
  INV_X1 U8759 ( .A(n7279), .ZN(n7025) );
  NAND2_X1 U8760 ( .A1(n8237), .A2(n7614), .ZN(n7020) );
  OR2_X1 U8761 ( .A1(n7279), .A2(n9650), .ZN(n7019) );
  OAI211_X1 U8762 ( .C1(n7022), .C2(n7040), .A(n7020), .B(n7019), .ZN(n7021)
         );
  INV_X1 U8763 ( .A(n7021), .ZN(n7066) );
  NAND2_X1 U8764 ( .A1(n6392), .A2(n7023), .ZN(n7024) );
  AOI22_X1 U8765 ( .A1(n8237), .A2(n7820), .B1(n7025), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U8766 ( .A1(n7027), .A2(n7026), .ZN(n7030) );
  INV_X1 U8767 ( .A(n7030), .ZN(n7028) );
  INV_X1 U8768 ( .A(n7068), .ZN(n7029) );
  AOI21_X1 U8769 ( .B1(n7066), .B2(n7030), .A(n7029), .ZN(n9660) );
  INV_X1 U8770 ( .A(n7031), .ZN(n9547) );
  OR2_X1 U8771 ( .A1(n10299), .A2(n9547), .ZN(n7283) );
  INV_X1 U8772 ( .A(n7032), .ZN(n7624) );
  NAND3_X1 U8773 ( .A1(n7367), .A2(n7624), .A3(n7033), .ZN(n7285) );
  INV_X1 U8774 ( .A(n7286), .ZN(n7034) );
  NOR2_X2 U8775 ( .A1(n7283), .A2(n7037), .ZN(n9311) );
  OR2_X1 U8776 ( .A1(n7018), .A2(n7065), .ZN(n7790) );
  NOR2_X1 U8777 ( .A1(n7790), .A2(n7034), .ZN(n9626) );
  INV_X1 U8778 ( .A(n7285), .ZN(n7282) );
  INV_X1 U8779 ( .A(n7074), .ZN(n7035) );
  NAND2_X1 U8780 ( .A1(n9611), .A2(n7286), .ZN(n7036) );
  NAND2_X1 U8781 ( .A1(n7037), .A2(n9999), .ZN(n8094) );
  NAND2_X1 U8782 ( .A1(n8094), .A2(n7280), .ZN(n7171) );
  AOI22_X1 U8783 ( .A1(n9334), .A2(n6057), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7171), .ZN(n7039) );
  NAND2_X1 U8784 ( .A1(n9338), .A2(n7820), .ZN(n7038) );
  OAI211_X1 U8785 ( .C1(n9660), .C2(n9340), .A(n7039), .B(n7038), .ZN(P1_U3230) );
  INV_X1 U8786 ( .A(n7790), .ZN(n7287) );
  AND2_X1 U8787 ( .A1(n7614), .A2(n7040), .ZN(n9361) );
  NOR2_X1 U8788 ( .A1(n7613), .A2(n9361), .ZN(n9582) );
  OR3_X1 U8789 ( .A1(n7287), .A2(n9582), .A3(n7042), .ZN(n7041) );
  OAI21_X1 U8790 ( .B1(n9364), .B2(n10016), .A(n7041), .ZN(n7821) );
  AOI21_X1 U8791 ( .B1(n7820), .B2(n7042), .A(n7821), .ZN(n7371) );
  NAND2_X1 U8792 ( .A1(n10341), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7043) );
  OAI21_X1 U8793 ( .B1(n7371), .B2(n10341), .A(n7043), .ZN(P1_U3523) );
  INV_X1 U8794 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7064) );
  AND2_X1 U8795 ( .A1(n7560), .A2(n7270), .ZN(n7344) );
  NAND2_X1 U8796 ( .A1(n7046), .A2(n7344), .ZN(n7048) );
  NAND2_X1 U8797 ( .A1(n7352), .A2(n5754), .ZN(n7047) );
  NAND3_X1 U8798 ( .A1(n7049), .A2(n7048), .A3(n7047), .ZN(n7050) );
  INV_X1 U8799 ( .A(n8890), .ZN(n7811) );
  OR2_X1 U8800 ( .A1(n7525), .A2(n8795), .ZN(n7053) );
  OR2_X1 U8801 ( .A1(n5754), .A2(n8793), .ZN(n7052) );
  NAND2_X1 U8802 ( .A1(n7053), .A2(n7052), .ZN(n8418) );
  AOI21_X1 U8803 ( .B1(n8928), .B2(n7811), .A(n8418), .ZN(n7058) );
  XNOR2_X1 U8804 ( .A(n7054), .B(n7055), .ZN(n7056) );
  NAND2_X1 U8805 ( .A1(n7056), .A2(n8902), .ZN(n7057) );
  AND2_X1 U8806 ( .A1(n7058), .A2(n7057), .ZN(n8926) );
  INV_X1 U8807 ( .A(n10429), .ZN(n7061) );
  NAND2_X1 U8808 ( .A1(n7355), .A2(n8927), .ZN(n7059) );
  NAND2_X1 U8809 ( .A1(n7327), .A2(n7059), .ZN(n8931) );
  OAI22_X1 U8810 ( .A1(n8931), .A2(n10400), .B1(n7311), .B2(n10398), .ZN(n7060) );
  AOI21_X1 U8811 ( .B1(n8928), .B2(n7061), .A(n7060), .ZN(n7062) );
  NAND2_X1 U8812 ( .A1(n8926), .A2(n7062), .ZN(n7079) );
  NAND2_X1 U8813 ( .A1(n7079), .A2(n10433), .ZN(n7063) );
  OAI21_X1 U8814 ( .B1(n10433), .B2(n7064), .A(n7063), .ZN(P2_U3460) );
  NAND2_X1 U8815 ( .A1(n7066), .A2(n9157), .ZN(n7067) );
  OR2_X1 U8816 ( .A1(n7299), .A2(n9364), .ZN(n7070) );
  NAND2_X1 U8817 ( .A1(n8237), .A2(n4386), .ZN(n7069) );
  INV_X1 U8818 ( .A(n7163), .ZN(n7167) );
  XNOR2_X1 U8819 ( .A(n7166), .B(n7167), .ZN(n7073) );
  OR2_X1 U8820 ( .A1(n8217), .A2(n9364), .ZN(n7071) );
  XNOR2_X1 U8821 ( .A(n7072), .B(n9157), .ZN(n7164) );
  INV_X1 U8822 ( .A(n7164), .ZN(n7168) );
  XNOR2_X1 U8823 ( .A(n7073), .B(n7168), .ZN(n7078) );
  AND2_X1 U8824 ( .A1(n10299), .A2(n4386), .ZN(n10256) );
  AOI22_X1 U8825 ( .A1(n9322), .A2(n7614), .B1(n10256), .B2(n8094), .ZN(n7077)
         );
  AOI22_X1 U8826 ( .A1(n9334), .A2(n7075), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7171), .ZN(n7076) );
  OAI211_X1 U8827 ( .C1(n7078), .C2(n9340), .A(n7077), .B(n7076), .ZN(P1_U3220) );
  INV_X1 U8828 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U8829 ( .A1(n7079), .A2(n10444), .ZN(n7080) );
  OAI21_X1 U8830 ( .B1(n10444), .B2(n7097), .A(n7080), .ZN(P2_U3523) );
  INV_X1 U8831 ( .A(n10133), .ZN(n10316) );
  NOR2_X1 U8832 ( .A1(n7081), .A2(n7617), .ZN(n7618) );
  AOI21_X1 U8833 ( .B1(n6057), .B2(n4386), .A(n7618), .ZN(n7082) );
  XNOR2_X1 U8834 ( .A(n7082), .B(n6074), .ZN(n7991) );
  INV_X1 U8835 ( .A(n7991), .ZN(n7089) );
  INV_X1 U8836 ( .A(n10299), .ZN(n10285) );
  OAI21_X1 U8837 ( .B1(n7820), .B2(n4386), .A(n7987), .ZN(n7083) );
  NAND2_X1 U8838 ( .A1(n7083), .A2(n7973), .ZN(n7985) );
  OAI22_X1 U8839 ( .A1(n10285), .A2(n7161), .B1(n7985), .B2(n10320), .ZN(n7088) );
  OAI21_X1 U8840 ( .B1(n6074), .B2(n9368), .A(n7084), .ZN(n7086) );
  OAI22_X1 U8841 ( .A1(n7301), .A2(n10016), .B1(n10014), .B2(n9364), .ZN(n7085) );
  AOI21_X1 U8842 ( .B1(n7086), .B2(n9981), .A(n7085), .ZN(n7087) );
  OAI21_X1 U8843 ( .B1(n7991), .B2(n10311), .A(n7087), .ZN(n7988) );
  AOI211_X1 U8844 ( .C1(n10316), .C2(n7089), .A(n7088), .B(n7988), .ZN(n10263)
         );
  NAND2_X1 U8845 ( .A1(n10341), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7090) );
  OAI21_X1 U8846 ( .B1(n10263), .B2(n10341), .A(n7090), .ZN(P1_U3525) );
  INV_X1 U8847 ( .A(n7091), .ZN(n7251) );
  AOI22_X1 U8848 ( .A1(n8627), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9093), .ZN(n7092) );
  OAI21_X1 U8849 ( .B1(n7251), .B2(n9101), .A(n7092), .ZN(P2_U3340) );
  INV_X1 U8850 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8930) );
  OAI22_X1 U8851 ( .A1(n8643), .A2(n10203), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8930), .ZN(n7104) );
  INV_X1 U8852 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7093) );
  MUX2_X1 U8853 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7093), .S(n7182), .Z(n7095)
         );
  NAND2_X1 U8854 ( .A1(n7108), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8855 ( .A1(n7176), .A2(n7175), .ZN(n7094) );
  NAND2_X1 U8856 ( .A1(n7095), .A2(n7094), .ZN(n7179) );
  NAND2_X1 U8857 ( .A1(n7182), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7096) );
  NAND2_X1 U8858 ( .A1(n7179), .A2(n7096), .ZN(n7099) );
  INV_X1 U8859 ( .A(n7099), .ZN(n7102) );
  MUX2_X1 U8860 ( .A(n7097), .B(P2_REG1_REG_3__SCAN_IN), .S(n7131), .Z(n7101)
         );
  MUX2_X1 U8861 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7097), .S(n7131), .Z(n7098)
         );
  INV_X1 U8862 ( .A(n7190), .ZN(n7100) );
  AOI211_X1 U8863 ( .C1(n7102), .C2(n7101), .A(n7100), .B(n7719), .ZN(n7103)
         );
  AOI211_X1 U8864 ( .C1(n10354), .C2(n7131), .A(n7104), .B(n7103), .ZN(n7117)
         );
  INV_X1 U8865 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7105) );
  MUX2_X1 U8866 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7105), .S(n7182), .Z(n7185)
         );
  NAND2_X1 U8867 ( .A1(n7108), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U8868 ( .A1(n7110), .A2(n7109), .ZN(n7184) );
  NAND2_X1 U8869 ( .A1(n7185), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U8870 ( .A1(n7182), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7113) );
  NAND2_X1 U8871 ( .A1(n7183), .A2(n7113), .ZN(n7112) );
  INV_X1 U8872 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8925) );
  MUX2_X1 U8873 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n8925), .S(n7131), .Z(n7111)
         );
  NAND2_X1 U8874 ( .A1(n7112), .A2(n7111), .ZN(n7198) );
  MUX2_X1 U8875 ( .A(n8925), .B(P2_REG2_REG_3__SCAN_IN), .S(n7131), .Z(n7114)
         );
  NAND3_X1 U8876 ( .A1(n7183), .A2(n7114), .A3(n7113), .ZN(n7115) );
  NAND3_X1 U8877 ( .A1(n10349), .A2(n7198), .A3(n7115), .ZN(n7116) );
  NAND2_X1 U8878 ( .A1(n7117), .A2(n7116), .ZN(P2_U3248) );
  INV_X1 U8879 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U8880 ( .A1(n7131), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7189) );
  INV_X1 U8881 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7118) );
  MUX2_X1 U8882 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7118), .S(n7195), .Z(n7119)
         );
  NAND2_X1 U8883 ( .A1(n7120), .A2(n7119), .ZN(n7192) );
  NAND2_X1 U8884 ( .A1(n7195), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7125) );
  NAND2_X1 U8885 ( .A1(n7192), .A2(n7125), .ZN(n7123) );
  INV_X1 U8886 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7121) );
  MUX2_X1 U8887 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7121), .S(n7150), .Z(n7122)
         );
  MUX2_X1 U8888 ( .A(n7121), .B(P2_REG1_REG_5__SCAN_IN), .S(n7150), .Z(n7124)
         );
  NAND3_X1 U8889 ( .A1(n7192), .A2(n7125), .A3(n7124), .ZN(n7126) );
  NAND3_X1 U8890 ( .A1(n10355), .A2(n7237), .A3(n7126), .ZN(n7128) );
  AND2_X1 U8891 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7394) );
  INV_X1 U8892 ( .A(n7394), .ZN(n7127) );
  OAI211_X1 U8893 ( .C1(n7129), .C2(n8643), .A(n7128), .B(n7127), .ZN(n7130)
         );
  AOI21_X1 U8894 ( .B1(n7150), .B2(n10354), .A(n7130), .ZN(n7140) );
  NAND2_X1 U8895 ( .A1(n7131), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7197) );
  NAND2_X1 U8896 ( .A1(n7198), .A2(n7197), .ZN(n7133) );
  INV_X1 U8897 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7323) );
  MUX2_X1 U8898 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7323), .S(n7195), .Z(n7132)
         );
  NAND2_X1 U8899 ( .A1(n7133), .A2(n7132), .ZN(n7200) );
  NAND2_X1 U8900 ( .A1(n7195), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8901 ( .A1(n7200), .A2(n7137), .ZN(n7135) );
  INV_X1 U8902 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7552) );
  MUX2_X1 U8903 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7552), .S(n7150), .Z(n7134)
         );
  NAND2_X1 U8904 ( .A1(n7135), .A2(n7134), .ZN(n7245) );
  MUX2_X1 U8905 ( .A(n7552), .B(P2_REG2_REG_5__SCAN_IN), .S(n7150), .Z(n7136)
         );
  NAND3_X1 U8906 ( .A1(n7200), .A2(n7137), .A3(n7136), .ZN(n7138) );
  NAND3_X1 U8907 ( .A1(n10349), .A2(n7245), .A3(n7138), .ZN(n7139) );
  NAND2_X1 U8908 ( .A1(n7140), .A2(n7139), .ZN(P2_U3250) );
  NAND2_X1 U8909 ( .A1(n7150), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7236) );
  NAND2_X1 U8910 ( .A1(n7237), .A2(n7236), .ZN(n7142) );
  MUX2_X1 U8911 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10439), .S(n7242), .Z(n7141)
         );
  NAND2_X1 U8912 ( .A1(n7242), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U8913 ( .A1(n7239), .A2(n7146), .ZN(n7144) );
  MUX2_X1 U8914 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7608), .S(n7210), .Z(n7143)
         );
  MUX2_X1 U8915 ( .A(n7608), .B(P2_REG1_REG_7__SCAN_IN), .S(n7210), .Z(n7145)
         );
  NAND3_X1 U8916 ( .A1(n7239), .A2(n7146), .A3(n7145), .ZN(n7147) );
  NAND3_X1 U8917 ( .A1(n10355), .A2(n7206), .A3(n7147), .ZN(n7148) );
  NAND2_X1 U8918 ( .A1(n4369), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7590) );
  OAI211_X1 U8919 ( .C1(n10196), .C2(n8643), .A(n7148), .B(n7590), .ZN(n7149)
         );
  AOI21_X1 U8920 ( .B1(n7210), .B2(n10354), .A(n7149), .ZN(n7159) );
  NAND2_X1 U8921 ( .A1(n7150), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U8922 ( .A1(n7245), .A2(n7244), .ZN(n7152) );
  INV_X1 U8923 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7535) );
  MUX2_X1 U8924 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7535), .S(n7242), .Z(n7151)
         );
  NAND2_X1 U8925 ( .A1(n7152), .A2(n7151), .ZN(n7247) );
  NAND2_X1 U8926 ( .A1(n7242), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8927 ( .A1(n7247), .A2(n7156), .ZN(n7154) );
  MUX2_X1 U8928 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7581), .S(n7210), .Z(n7153)
         );
  NAND2_X1 U8929 ( .A1(n7154), .A2(n7153), .ZN(n7215) );
  MUX2_X1 U8930 ( .A(n7581), .B(P2_REG2_REG_7__SCAN_IN), .S(n7210), .Z(n7155)
         );
  NAND3_X1 U8931 ( .A1(n7247), .A2(n7156), .A3(n7155), .ZN(n7157) );
  NAND3_X1 U8932 ( .A1(n10349), .A2(n7215), .A3(n7157), .ZN(n7158) );
  NAND2_X1 U8933 ( .A1(n7159), .A2(n7158), .ZN(P2_U3252) );
  NOR2_X1 U8934 ( .A1(n8217), .A2(n7161), .ZN(n7160) );
  AOI21_X1 U8935 ( .B1(n7733), .B2(n7075), .A(n7160), .ZN(n7296) );
  XNOR2_X1 U8936 ( .A(n7162), .B(n9157), .ZN(n7294) );
  XNOR2_X1 U8937 ( .A(n7296), .B(n7294), .ZN(n7292) );
  NAND2_X1 U8938 ( .A1(n7164), .A2(n7163), .ZN(n7165) );
  NAND2_X1 U8939 ( .A1(n7166), .A2(n7165), .ZN(n7170) );
  NAND2_X1 U8940 ( .A1(n7168), .A2(n7167), .ZN(n7169) );
  NAND2_X1 U8941 ( .A1(n7170), .A2(n7169), .ZN(n7293) );
  XOR2_X1 U8942 ( .A(n7292), .B(n7293), .Z(n7174) );
  AOI22_X1 U8943 ( .A1(n9334), .A2(n9648), .B1(n9322), .B2(n6057), .ZN(n7173)
         );
  AOI22_X1 U8944 ( .A1(n9338), .A2(n7987), .B1(n7171), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7172) );
  OAI211_X1 U8945 ( .C1(n7174), .C2(n9340), .A(n7173), .B(n7172), .ZN(P1_U3235) );
  INV_X1 U8946 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7356) );
  OAI22_X1 U8947 ( .A1(n8643), .A2(n10198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7356), .ZN(n7181) );
  MUX2_X1 U8948 ( .A(n7093), .B(P2_REG1_REG_2__SCAN_IN), .S(n7182), .Z(n7177)
         );
  NAND3_X1 U8949 ( .A1(n7177), .A2(n7176), .A3(n7175), .ZN(n7178) );
  AND3_X1 U8950 ( .A1(n10355), .A2(n7179), .A3(n7178), .ZN(n7180) );
  AOI211_X1 U8951 ( .C1(n10354), .C2(n7182), .A(n7181), .B(n7180), .ZN(n7187)
         );
  OAI211_X1 U8952 ( .C1(n7185), .C2(n7184), .A(n10349), .B(n7183), .ZN(n7186)
         );
  NAND2_X1 U8953 ( .A1(n7187), .A2(n7186), .ZN(P2_U3247) );
  NAND2_X1 U8954 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7516) );
  INV_X1 U8955 ( .A(n7516), .ZN(n7194) );
  MUX2_X1 U8956 ( .A(n7118), .B(P2_REG1_REG_4__SCAN_IN), .S(n7195), .Z(n7188)
         );
  NAND3_X1 U8957 ( .A1(n7190), .A2(n7189), .A3(n7188), .ZN(n7191) );
  AND3_X1 U8958 ( .A1(n10355), .A2(n7192), .A3(n7191), .ZN(n7193) );
  AOI211_X1 U8959 ( .C1(n10347), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7194), .B(
        n7193), .ZN(n7202) );
  MUX2_X1 U8960 ( .A(n7323), .B(P2_REG2_REG_4__SCAN_IN), .S(n7195), .Z(n7196)
         );
  NAND3_X1 U8961 ( .A1(n7198), .A2(n7197), .A3(n7196), .ZN(n7199) );
  NAND3_X1 U8962 ( .A1(n10349), .A2(n7200), .A3(n7199), .ZN(n7201) );
  OAI211_X1 U8963 ( .C1(n7203), .C2(n8626), .A(n7202), .B(n7201), .ZN(P2_U3249) );
  NAND2_X1 U8964 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7840) );
  INV_X1 U8965 ( .A(n7840), .ZN(n7209) );
  NAND2_X1 U8966 ( .A1(n7210), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7205) );
  INV_X1 U8967 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10442) );
  MUX2_X1 U8968 ( .A(n10442), .B(P2_REG1_REG_8__SCAN_IN), .S(n7224), .Z(n7204)
         );
  AOI21_X1 U8969 ( .B1(n7206), .B2(n7205), .A(n7204), .ZN(n7220) );
  AND3_X1 U8970 ( .A1(n7206), .A2(n7205), .A3(n7204), .ZN(n7207) );
  NOR3_X1 U8971 ( .A1(n7719), .A2(n7220), .A3(n7207), .ZN(n7208) );
  AOI211_X1 U8972 ( .C1(n10347), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7209), .B(
        n7208), .ZN(n7218) );
  NAND2_X1 U8973 ( .A1(n7210), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U8974 ( .A1(n7215), .A2(n7214), .ZN(n7212) );
  INV_X1 U8975 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7682) );
  MUX2_X1 U8976 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7682), .S(n7224), .Z(n7211)
         );
  NAND2_X1 U8977 ( .A1(n7212), .A2(n7211), .ZN(n7427) );
  MUX2_X1 U8978 ( .A(n7682), .B(P2_REG2_REG_8__SCAN_IN), .S(n7224), .Z(n7213)
         );
  NAND3_X1 U8979 ( .A1(n7215), .A2(n7214), .A3(n7213), .ZN(n7216) );
  NAND3_X1 U8980 ( .A1(n10349), .A2(n7427), .A3(n7216), .ZN(n7217) );
  OAI211_X1 U8981 ( .C1(n8626), .C2(n7219), .A(n7218), .B(n7217), .ZN(P2_U3253) );
  XNOR2_X1 U8982 ( .A(n7424), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7420) );
  INV_X1 U8983 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7221) );
  OAI22_X1 U8984 ( .A1(n7421), .A2(n7420), .B1(n7422), .B2(n7221), .ZN(n7254)
         );
  XOR2_X1 U8985 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7255), .Z(n7253) );
  XNOR2_X1 U8986 ( .A(n7254), .B(n7253), .ZN(n7234) );
  INV_X1 U8987 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8988 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8041) );
  OAI21_X1 U8989 ( .B1(n8643), .B2(n7222), .A(n8041), .ZN(n7223) );
  AOI21_X1 U8990 ( .B1(n10354), .B2(n7255), .A(n7223), .ZN(n7233) );
  NAND2_X1 U8991 ( .A1(n7224), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8992 ( .A1(n7427), .A2(n7426), .ZN(n7226) );
  INV_X1 U8993 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7812) );
  MUX2_X1 U8994 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7812), .S(n7424), .Z(n7225)
         );
  NAND2_X1 U8995 ( .A1(n7226), .A2(n7225), .ZN(n7429) );
  NAND2_X1 U8996 ( .A1(n7424), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U8997 ( .A1(n7429), .A2(n7230), .ZN(n7228) );
  INV_X1 U8998 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8136) );
  MUX2_X1 U8999 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8136), .S(n7255), .Z(n7227)
         );
  NAND2_X1 U9000 ( .A1(n7228), .A2(n7227), .ZN(n7257) );
  MUX2_X1 U9001 ( .A(n8136), .B(P2_REG2_REG_10__SCAN_IN), .S(n7255), .Z(n7229)
         );
  NAND3_X1 U9002 ( .A1(n7429), .A2(n7230), .A3(n7229), .ZN(n7231) );
  NAND3_X1 U9003 ( .A1(n10349), .A2(n7257), .A3(n7231), .ZN(n7232) );
  OAI211_X1 U9004 ( .C1(n7234), .C2(n7719), .A(n7233), .B(n7232), .ZN(P2_U3255) );
  NAND2_X1 U9005 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n4369), .ZN(n7495) );
  INV_X1 U9006 ( .A(n7495), .ZN(n7241) );
  MUX2_X1 U9007 ( .A(n10439), .B(P2_REG1_REG_6__SCAN_IN), .S(n7242), .Z(n7235)
         );
  NAND3_X1 U9008 ( .A1(n7237), .A2(n7236), .A3(n7235), .ZN(n7238) );
  AND3_X1 U9009 ( .A1(n10355), .A2(n7239), .A3(n7238), .ZN(n7240) );
  AOI211_X1 U9010 ( .C1(n10347), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7241), .B(
        n7240), .ZN(n7249) );
  MUX2_X1 U9011 ( .A(n7535), .B(P2_REG2_REG_6__SCAN_IN), .S(n7242), .Z(n7243)
         );
  NAND3_X1 U9012 ( .A1(n7245), .A2(n7244), .A3(n7243), .ZN(n7246) );
  NAND3_X1 U9013 ( .A1(n10349), .A2(n7247), .A3(n7246), .ZN(n7248) );
  OAI211_X1 U9014 ( .C1(n8626), .C2(n7250), .A(n7249), .B(n7248), .ZN(P2_U3251) );
  INV_X1 U9015 ( .A(n9728), .ZN(n8108) );
  OAI222_X1 U9016 ( .A1(n10182), .A2(n7252), .B1(n10186), .B2(n7251), .C1(
        P1_U3084), .C2(n8108), .ZN(P1_U3335) );
  XNOR2_X1 U9017 ( .A(n7410), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7403) );
  XNOR2_X1 U9018 ( .A(n7404), .B(n7403), .ZN(n7264) );
  NAND2_X1 U9019 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8548) );
  OAI21_X1 U9020 ( .B1(n8643), .B2(n6669), .A(n8548), .ZN(n7262) );
  NAND2_X1 U9021 ( .A1(n7255), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U9022 ( .A1(n7257), .A2(n7256), .ZN(n7259) );
  INV_X1 U9023 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7930) );
  MUX2_X1 U9024 ( .A(n7930), .B(P2_REG2_REG_11__SCAN_IN), .S(n7410), .Z(n7258)
         );
  NAND2_X1 U9025 ( .A1(n7259), .A2(n7258), .ZN(n7260) );
  AOI21_X1 U9026 ( .B1(n7412), .B2(n7260), .A(n8637), .ZN(n7261) );
  AOI211_X1 U9027 ( .C1(n10354), .C2(n7410), .A(n7262), .B(n7261), .ZN(n7263)
         );
  OAI21_X1 U9028 ( .B1(n7264), .B2(n7719), .A(n7263), .ZN(P2_U3256) );
  NAND2_X1 U9029 ( .A1(n7265), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7269) );
  NAND2_X1 U9030 ( .A1(n7267), .A2(n7266), .ZN(n7268) );
  NAND2_X1 U9031 ( .A1(n8564), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7567) );
  INV_X1 U9032 ( .A(n7567), .ZN(n7506) );
  INV_X1 U9033 ( .A(n8565), .ZN(n8587) );
  OAI22_X1 U9034 ( .A1(n7270), .A2(n8570), .B1(n8537), .B2(n5754), .ZN(n7271)
         );
  AOI21_X1 U9035 ( .B1(n8587), .B2(n4973), .A(n7271), .ZN(n7277) );
  OAI21_X1 U9036 ( .B1(n7274), .B2(n7273), .A(n7272), .ZN(n7275) );
  NAND2_X1 U9037 ( .A1(n7275), .A2(n8583), .ZN(n7276) );
  OAI211_X1 U9038 ( .C1(n7506), .C2(n7278), .A(n7277), .B(n7276), .ZN(P2_U3224) );
  AND3_X1 U9039 ( .A1(n7280), .A2(n7279), .A3(n7796), .ZN(n7281) );
  OAI21_X1 U9040 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n7284) );
  NAND2_X1 U9041 ( .A1(n7284), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7289) );
  NOR2_X1 U9042 ( .A1(n7818), .A2(n9550), .ZN(n7627) );
  OAI211_X1 U9043 ( .C1(n7287), .C2(n7627), .A(n7286), .B(n7285), .ZN(n7288)
         );
  OAI22_X1 U9044 ( .A1(n9298), .A2(n10267), .B1(n9320), .B2(n7780), .ZN(n7290)
         );
  AOI211_X1 U9045 ( .C1(n9322), .C2(n7075), .A(n7291), .B(n7290), .ZN(n7306)
         );
  NAND2_X1 U9046 ( .A1(n7293), .A2(n7292), .ZN(n7298) );
  INV_X1 U9047 ( .A(n7294), .ZN(n7295) );
  NAND2_X1 U9048 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  NAND2_X1 U9049 ( .A1(n7298), .A2(n7297), .ZN(n7373) );
  NOR2_X1 U9050 ( .A1(n8217), .A2(n10267), .ZN(n7300) );
  AOI21_X1 U9051 ( .B1(n7733), .B2(n9648), .A(n7300), .ZN(n7376) );
  OR2_X1 U9052 ( .A1(n8217), .A2(n7301), .ZN(n7302) );
  OAI21_X1 U9053 ( .B1(n7022), .B2(n10267), .A(n7302), .ZN(n7303) );
  XNOR2_X1 U9054 ( .A(n7303), .B(n9157), .ZN(n7374) );
  XNOR2_X1 U9055 ( .A(n7376), .B(n7374), .ZN(n7372) );
  XNOR2_X1 U9056 ( .A(n7373), .B(n7372), .ZN(n7304) );
  NAND2_X1 U9057 ( .A1(n7304), .A2(n9311), .ZN(n7305) );
  OAI211_X1 U9058 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9336), .A(n7306), .B(
        n7305), .ZN(P1_U3216) );
  INV_X1 U9059 ( .A(n7307), .ZN(n7309) );
  OAI222_X1 U9060 ( .A1(n8378), .A2(n7308), .B1(n7652), .B2(n7309), .C1(n4369), 
        .C2(n8874), .ZN(P2_U3339) );
  OAI222_X1 U9061 ( .A1(n10182), .A2(n7310), .B1(n10186), .B2(n7309), .C1(
        P1_U3084), .C2(n9615), .ZN(P1_U3334) );
  NAND2_X1 U9062 ( .A1(n7517), .A2(n7311), .ZN(n7312) );
  NAND2_X1 U9063 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  NAND2_X1 U9064 ( .A1(n7314), .A2(n7321), .ZN(n7527) );
  OAI21_X1 U9065 ( .B1(n7314), .B2(n7321), .A(n7527), .ZN(n10405) );
  INV_X1 U9066 ( .A(n10405), .ZN(n7334) );
  NAND3_X1 U9067 ( .A1(n7317), .A2(n7316), .A3(n7315), .ZN(n7325) );
  OR2_X1 U9068 ( .A1(n7318), .A2(n8874), .ZN(n7674) );
  NAND2_X1 U9069 ( .A1(n8890), .A2(n7674), .ZN(n7319) );
  XOR2_X1 U9070 ( .A(n7320), .B(n7321), .Z(n7322) );
  AOI222_X1 U9071 ( .A1(n8902), .A2(n7322), .B1(n8607), .B2(n8908), .C1(n8609), 
        .C2(n8907), .ZN(n10402) );
  MUX2_X1 U9072 ( .A(n7323), .B(n10402), .S(n8945), .Z(n7333) );
  INV_X1 U9073 ( .A(n7325), .ZN(n7326) );
  AND2_X1 U9074 ( .A1(n7326), .A2(n8874), .ZN(n8818) );
  NAND2_X1 U9075 ( .A1(n8818), .A2(n10424), .ZN(n8932) );
  INV_X1 U9076 ( .A(n7327), .ZN(n7328) );
  INV_X1 U9077 ( .A(n7536), .ZN(n7553) );
  OAI21_X1 U9078 ( .B1(n10399), .B2(n7328), .A(n7553), .ZN(n10401) );
  OAI22_X1 U9079 ( .A1(n8932), .A2(n10401), .B1(n7329), .B2(n8877), .ZN(n7330)
         );
  AOI21_X1 U9080 ( .B1(n8939), .B2(n7331), .A(n7330), .ZN(n7332) );
  OAI211_X1 U9081 ( .C1(n7334), .C2(n8860), .A(n7333), .B(n7332), .ZN(P2_U3292) );
  NAND2_X1 U9082 ( .A1(n7335), .A2(n10385), .ZN(n7337) );
  INV_X1 U9083 ( .A(n7337), .ZN(n7343) );
  OAI21_X1 U9084 ( .B1(n8944), .B2(n8939), .A(n10381), .ZN(n7342) );
  INV_X1 U9085 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7505) );
  AOI22_X1 U9086 ( .A1(n7337), .A2(n8902), .B1(n8908), .B2(n7336), .ZN(n10386)
         );
  OAI21_X1 U9087 ( .B1(n7505), .B2(n8877), .A(n10386), .ZN(n7340) );
  NOR2_X1 U9088 ( .A1(n8945), .A2(n7338), .ZN(n7339) );
  AOI21_X1 U9089 ( .B1(n8945), .B2(n7340), .A(n7339), .ZN(n7341) );
  OAI211_X1 U9090 ( .C1(n7343), .C2(n8860), .A(n7342), .B(n7341), .ZN(P2_U3296) );
  NOR2_X1 U9091 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  XNOR2_X1 U9092 ( .A(n7346), .B(n7350), .ZN(n10395) );
  INV_X1 U9093 ( .A(n7348), .ZN(n7349) );
  AOI21_X1 U9094 ( .B1(n7347), .B2(n7350), .A(n7349), .ZN(n7351) );
  OAI222_X1 U9095 ( .A1(n8793), .A2(n7560), .B1(n8795), .B2(n7517), .C1(n8868), 
        .C2(n7351), .ZN(n10390) );
  AOI22_X1 U9096 ( .A1(n10390), .A2(n8945), .B1(n8939), .B2(n10391), .ZN(n7359) );
  OR2_X1 U9097 ( .A1(n7353), .A2(n7352), .ZN(n7354) );
  AND2_X1 U9098 ( .A1(n7355), .A2(n7354), .ZN(n10392) );
  OAI22_X1 U9099 ( .A1(n8945), .A2(n7105), .B1(n7356), .B2(n8877), .ZN(n7357)
         );
  AOI21_X1 U9100 ( .B1(n8944), .B2(n10392), .A(n7357), .ZN(n7358) );
  OAI211_X1 U9101 ( .C1(n10395), .C2(n8860), .A(n7359), .B(n7358), .ZN(
        P2_U3294) );
  INV_X1 U9102 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7366) );
  AOI22_X1 U9103 ( .A1(n10349), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10355), .ZN(n7363) );
  NAND2_X1 U9104 ( .A1(n10355), .A2(n10434), .ZN(n7360) );
  OAI211_X1 U9105 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n8637), .A(n8626), .B(
        n7360), .ZN(n7361) );
  INV_X1 U9106 ( .A(n7361), .ZN(n7362) );
  MUX2_X1 U9107 ( .A(n7363), .B(n7362), .S(P2_IR_REG_0__SCAN_IN), .Z(n7365) );
  NAND2_X1 U9108 ( .A1(n4369), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7364) );
  OAI211_X1 U9109 ( .C1(n8643), .C2(n7366), .A(n7365), .B(n7364), .ZN(P2_U3245) );
  INV_X1 U9110 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7369) );
  OR2_X1 U9111 ( .A1(n10272), .A2(n7369), .ZN(n7370) );
  OAI21_X1 U9112 ( .B1(n7371), .B2(n10326), .A(n7370), .ZN(P1_U3454) );
  NAND2_X1 U9113 ( .A1(n7373), .A2(n7372), .ZN(n7378) );
  INV_X1 U9114 ( .A(n7374), .ZN(n7375) );
  NAND2_X1 U9115 ( .A1(n7376), .A2(n7375), .ZN(n7377) );
  OR2_X1 U9116 ( .A1(n8217), .A2(n7780), .ZN(n7379) );
  OAI21_X1 U9117 ( .B1(n7022), .B2(n8015), .A(n7379), .ZN(n7380) );
  OR2_X1 U9118 ( .A1(n8297), .A2(n7780), .ZN(n7382) );
  NAND2_X1 U9119 ( .A1(n4378), .A2(n8019), .ZN(n7381) );
  XNOR2_X1 U9120 ( .A(n7692), .B(n7691), .ZN(n7383) );
  XNOR2_X1 U9121 ( .A(n7694), .B(n7383), .ZN(n7388) );
  AND2_X1 U9122 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9683) );
  INV_X1 U9123 ( .A(n8094), .ZN(n9264) );
  NAND2_X1 U9124 ( .A1(n10299), .A2(n8019), .ZN(n10274) );
  NOR2_X1 U9125 ( .A1(n9264), .A2(n10274), .ZN(n7384) );
  AOI211_X1 U9126 ( .C1(n9322), .C2(n9648), .A(n9683), .B(n7384), .ZN(n7385)
         );
  OAI21_X1 U9127 ( .B1(n7855), .B2(n9320), .A(n7385), .ZN(n7386) );
  AOI21_X1 U9128 ( .B1(n8016), .B2(n9305), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9129 ( .B1(n7388), .B2(n9340), .A(n7387), .ZN(P1_U3228) );
  XOR2_X1 U9130 ( .A(n7390), .B(n7389), .Z(n7398) );
  INV_X1 U9131 ( .A(n7391), .ZN(n7554) );
  NOR2_X1 U9132 ( .A1(n8564), .A2(n7554), .ZN(n7397) );
  INV_X1 U9133 ( .A(n8573), .ZN(n8510) );
  OR2_X1 U9134 ( .A1(n7525), .A2(n8793), .ZN(n7393) );
  NAND2_X1 U9135 ( .A1(n8606), .A2(n8908), .ZN(n7392) );
  NAND2_X1 U9136 ( .A1(n7393), .A2(n7392), .ZN(n7550) );
  AOI21_X1 U9137 ( .B1(n8510), .B2(n7550), .A(n7394), .ZN(n7395) );
  OAI21_X1 U9138 ( .B1(n7570), .B2(n8570), .A(n7395), .ZN(n7396) );
  AOI211_X1 U9139 ( .C1(n7398), .C2(n8583), .A(n7397), .B(n7396), .ZN(n7399)
         );
  INV_X1 U9140 ( .A(n7399), .ZN(P2_U3229) );
  INV_X1 U9141 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U9142 ( .A1(n7407), .A2(n7400), .ZN(n7457) );
  OAI21_X1 U9143 ( .B1(n7407), .B2(n7400), .A(n7457), .ZN(n7406) );
  OAI22_X1 U9144 ( .A1(n7404), .A2(n7403), .B1(n7402), .B2(n7401), .ZN(n7405)
         );
  AOI21_X1 U9145 ( .B1(n7406), .B2(n7405), .A(n7462), .ZN(n7419) );
  NOR2_X1 U9146 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8454), .ZN(n7409) );
  NOR2_X1 U9147 ( .A1(n8626), .A2(n7407), .ZN(n7408) );
  AOI211_X1 U9148 ( .C1(n10347), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7409), .B(
        n7408), .ZN(n7418) );
  OR2_X1 U9149 ( .A1(n7410), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U9150 ( .A1(n7412), .A2(n7411), .ZN(n7415) );
  INV_X1 U9151 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7413) );
  MUX2_X1 U9152 ( .A(n7413), .B(P2_REG2_REG_12__SCAN_IN), .S(n7451), .Z(n7414)
         );
  AOI21_X1 U9153 ( .B1(n7415), .B2(n7414), .A(n8637), .ZN(n7416) );
  NAND2_X1 U9154 ( .A1(n7416), .A2(n7453), .ZN(n7417) );
  OAI211_X1 U9155 ( .C1(n7419), .C2(n7719), .A(n7418), .B(n7417), .ZN(P2_U3257) );
  XNOR2_X1 U9156 ( .A(n7421), .B(n7420), .ZN(n7432) );
  AND2_X1 U9157 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(n4369), .ZN(n7868) );
  NOR2_X1 U9158 ( .A1(n8626), .A2(n7422), .ZN(n7423) );
  AOI211_X1 U9159 ( .C1(n10347), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7868), .B(
        n7423), .ZN(n7431) );
  MUX2_X1 U9160 ( .A(n7812), .B(P2_REG2_REG_9__SCAN_IN), .S(n7424), .Z(n7425)
         );
  NAND3_X1 U9161 ( .A1(n7427), .A2(n7426), .A3(n7425), .ZN(n7428) );
  NAND3_X1 U9162 ( .A1(n10349), .A2(n7429), .A3(n7428), .ZN(n7430) );
  OAI211_X1 U9163 ( .C1(n7432), .C2(n7719), .A(n7431), .B(n7430), .ZN(P2_U3254) );
  NAND2_X1 U9164 ( .A1(n7433), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U9165 ( .A1(n7435), .A2(n7434), .ZN(n9719) );
  INV_X1 U9166 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7436) );
  XNOR2_X1 U9167 ( .A(n9715), .B(n7436), .ZN(n9718) );
  NAND2_X1 U9168 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U9169 ( .A1(n9715), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9170 ( .A1(n9717), .A2(n7437), .ZN(n7642) );
  XNOR2_X1 U9171 ( .A(n7642), .B(n7438), .ZN(n7640) );
  XNOR2_X1 U9172 ( .A(n7640), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n7449) );
  XOR2_X1 U9173 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7641), .Z(n7443) );
  INV_X1 U9174 ( .A(n7439), .ZN(n9708) );
  OR2_X1 U9175 ( .A1(n9715), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9176 ( .A1(n9715), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7440) );
  AND2_X1 U9177 ( .A1(n7441), .A2(n7440), .ZN(n9707) );
  OAI21_X1 U9178 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(n9706) );
  NAND2_X1 U9179 ( .A1(n9706), .A2(n7441), .ZN(n7442) );
  NAND2_X1 U9180 ( .A1(n7442), .A2(n7443), .ZN(n7637) );
  OAI21_X1 U9181 ( .B1(n7443), .B2(n7442), .A(n7637), .ZN(n7447) );
  NAND2_X1 U9182 ( .A1(n9716), .A2(n7641), .ZN(n7444) );
  NAND2_X1 U9183 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9126) );
  OAI211_X1 U9184 ( .C1(n7445), .C2(n10244), .A(n7444), .B(n9126), .ZN(n7446)
         );
  AOI21_X1 U9185 ( .B1(n7447), .B2(n10235), .A(n7446), .ZN(n7448) );
  OAI21_X1 U9186 ( .B1(n7449), .B2(n10228), .A(n7448), .ZN(P1_U3255) );
  OR2_X1 U9187 ( .A1(n7458), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7478) );
  NAND2_X1 U9188 ( .A1(n7458), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9189 ( .A1(n7478), .A2(n7450), .ZN(n7456) );
  NAND2_X1 U9190 ( .A1(n7451), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7452) );
  INV_X1 U9191 ( .A(n7480), .ZN(n7454) );
  AOI21_X1 U9192 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7470) );
  INV_X1 U9193 ( .A(n7457), .ZN(n7461) );
  OR2_X1 U9194 ( .A1(n7458), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9195 ( .A1(n7458), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7459) );
  AND2_X1 U9196 ( .A1(n7471), .A2(n7459), .ZN(n7460) );
  OAI21_X1 U9197 ( .B1(n7462), .B2(n7461), .A(n7460), .ZN(n7472) );
  INV_X1 U9198 ( .A(n7472), .ZN(n7464) );
  NOR3_X1 U9199 ( .A1(n7462), .A2(n7461), .A3(n7460), .ZN(n7463) );
  OAI21_X1 U9200 ( .B1(n7464), .B2(n7463), .A(n10355), .ZN(n7469) );
  AND2_X1 U9201 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7467) );
  NOR2_X1 U9202 ( .A1(n8626), .A2(n7465), .ZN(n7466) );
  AOI211_X1 U9203 ( .C1(n10347), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n7467), .B(
        n7466), .ZN(n7468) );
  OAI211_X1 U9204 ( .C1(n7470), .C2(n8637), .A(n7469), .B(n7468), .ZN(P2_U3258) );
  XOR2_X1 U9205 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7657), .Z(n7474) );
  NAND2_X1 U9206 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  NAND2_X1 U9207 ( .A1(n7473), .A2(n7474), .ZN(n7654) );
  OAI21_X1 U9208 ( .B1(n7474), .B2(n7473), .A(n7654), .ZN(n7487) );
  MUX2_X1 U9209 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7475), .S(n7657), .Z(n7477)
         );
  NAND2_X1 U9210 ( .A1(n7476), .A2(n7477), .ZN(n7659) );
  INV_X1 U9211 ( .A(n7477), .ZN(n7479) );
  NAND3_X1 U9212 ( .A1(n7480), .A2(n7479), .A3(n7478), .ZN(n7481) );
  AOI21_X1 U9213 ( .B1(n7659), .B2(n7481), .A(n8637), .ZN(n7486) );
  NOR2_X1 U9214 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8394), .ZN(n7482) );
  AOI21_X1 U9215 ( .B1(n10347), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7482), .ZN(
        n7483) );
  OAI21_X1 U9216 ( .B1(n8626), .B2(n7484), .A(n7483), .ZN(n7485) );
  AOI211_X1 U9217 ( .C1(n7487), .C2(n10355), .A(n7486), .B(n7485), .ZN(n7488)
         );
  INV_X1 U9218 ( .A(n7488), .ZN(P2_U3259) );
  INV_X1 U9219 ( .A(n7489), .ZN(n7508) );
  OAI222_X1 U9220 ( .A1(n10186), .A2(n7508), .B1(n9550), .B2(P1_U3084), .C1(
        n7490), .C2(n10182), .ZN(P1_U3333) );
  OAI21_X1 U9221 ( .B1(n7493), .B2(n7492), .A(n7491), .ZN(n7494) );
  NAND2_X1 U9222 ( .A1(n7494), .A2(n8583), .ZN(n7499) );
  INV_X1 U9223 ( .A(n8564), .ZN(n8588) );
  OAI21_X1 U9224 ( .B1(n8570), .B2(n7542), .A(n7495), .ZN(n7497) );
  OAI22_X1 U9225 ( .A1(n7571), .A2(n8565), .B1(n8537), .B2(n7839), .ZN(n7496)
         );
  AOI211_X1 U9226 ( .C1(n7540), .C2(n8588), .A(n7497), .B(n7496), .ZN(n7498)
         );
  NAND2_X1 U9227 ( .A1(n7499), .A2(n7498), .ZN(P2_U3241) );
  INV_X1 U9228 ( .A(n8537), .ZN(n8589) );
  AOI22_X1 U9229 ( .A1(n10381), .A2(n8590), .B1(n8589), .B2(n7336), .ZN(n7504)
         );
  NAND2_X1 U9230 ( .A1(n8583), .A2(n5525), .ZN(n8559) );
  OAI22_X1 U9231 ( .A1(n10380), .A2(n8559), .B1(n8579), .B2(n7500), .ZN(n7502)
         );
  NAND2_X1 U9232 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  OAI211_X1 U9233 ( .C1(n7506), .C2(n7505), .A(n7504), .B(n7503), .ZN(P2_U3234) );
  OAI222_X1 U9234 ( .A1(n8378), .A2(n7509), .B1(n7652), .B2(n7508), .C1(n7507), 
        .C2(n4369), .ZN(P2_U3338) );
  NAND2_X1 U9235 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8610), .ZN(n7510) );
  OAI21_X1 U9236 ( .B1(n7511), .B2(n8610), .A(n7510), .ZN(P2_U3581) );
  NAND2_X1 U9237 ( .A1(n7512), .A2(n7514), .ZN(n7515) );
  MUX2_X1 U9238 ( .A(n7515), .B(n7514), .S(n7513), .Z(n7524) );
  OAI21_X1 U9239 ( .B1(n8570), .B2(n10399), .A(n7516), .ZN(n7519) );
  OAI22_X1 U9240 ( .A1(n7517), .A2(n8565), .B1(n8537), .B2(n7571), .ZN(n7518)
         );
  AOI211_X1 U9241 ( .C1(n7520), .C2(n8588), .A(n7519), .B(n7518), .ZN(n7523)
         );
  INV_X1 U9242 ( .A(n8559), .ZN(n8581) );
  NAND4_X1 U9243 ( .A1(n7513), .A2(n8581), .A3(n4603), .A4(n8608), .ZN(n7522)
         );
  OAI211_X1 U9244 ( .C1(n7524), .C2(n8579), .A(n7523), .B(n7522), .ZN(P2_U3232) );
  NAND2_X1 U9245 ( .A1(n7525), .A2(n10399), .ZN(n7526) );
  INV_X1 U9246 ( .A(n7577), .ZN(n7529) );
  OAI21_X1 U9247 ( .B1(n7577), .B2(n7571), .A(n7570), .ZN(n7528) );
  OAI21_X1 U9248 ( .B1(n7529), .B2(n8607), .A(n7528), .ZN(n7530) );
  XNOR2_X1 U9249 ( .A(n7530), .B(n7532), .ZN(n10419) );
  XNOR2_X1 U9250 ( .A(n7531), .B(n7532), .ZN(n7534) );
  OAI22_X1 U9251 ( .A1(n7571), .A2(n8793), .B1(n7839), .B2(n8795), .ZN(n7533)
         );
  AOI21_X1 U9252 ( .B1(n7534), .B2(n8902), .A(n7533), .ZN(n10417) );
  MUX2_X1 U9253 ( .A(n7535), .B(n10417), .S(n8945), .Z(n7545) );
  INV_X1 U9254 ( .A(n7537), .ZN(n7539) );
  NAND2_X1 U9255 ( .A1(n7537), .A2(n7542), .ZN(n7583) );
  INV_X1 U9256 ( .A(n7583), .ZN(n7538) );
  AOI21_X1 U9257 ( .B1(n10414), .B2(n7539), .A(n7538), .ZN(n10415) );
  INV_X1 U9258 ( .A(n7540), .ZN(n7541) );
  OAI22_X1 U9259 ( .A1(n8920), .A2(n7542), .B1(n8877), .B2(n7541), .ZN(n7543)
         );
  AOI21_X1 U9260 ( .B1(n8944), .B2(n10415), .A(n7543), .ZN(n7544) );
  OAI211_X1 U9261 ( .C1(n10419), .C2(n8860), .A(n7545), .B(n7544), .ZN(
        P2_U3290) );
  XNOR2_X1 U9262 ( .A(n7577), .B(n7549), .ZN(n10411) );
  NAND2_X1 U9263 ( .A1(n7546), .A2(n7547), .ZN(n7548) );
  XOR2_X1 U9264 ( .A(n7549), .B(n7548), .Z(n7551) );
  AOI21_X1 U9265 ( .B1(n7551), .B2(n8902), .A(n7550), .ZN(n10410) );
  MUX2_X1 U9266 ( .A(n10410), .B(n7552), .S(n8924), .Z(n7558) );
  NAND2_X1 U9267 ( .A1(n8945), .A2(n8874), .ZN(n8840) );
  INV_X1 U9268 ( .A(n8840), .ZN(n7556) );
  AOI211_X1 U9269 ( .C1(n10408), .C2(n7553), .A(n10400), .B(n7537), .ZN(n10407) );
  OAI22_X1 U9270 ( .A1(n8920), .A2(n7570), .B1(n8877), .B2(n7554), .ZN(n7555)
         );
  AOI21_X1 U9271 ( .B1(n7556), .B2(n10407), .A(n7555), .ZN(n7557) );
  OAI211_X1 U9272 ( .C1(n8860), .C2(n10411), .A(n7558), .B(n7557), .ZN(
        P2_U3291) );
  AOI22_X1 U9273 ( .A1(n10391), .A2(n8590), .B1(n8589), .B2(n8609), .ZN(n7559)
         );
  OAI21_X1 U9274 ( .B1(n7560), .B2(n8565), .A(n7559), .ZN(n7566) );
  INV_X1 U9275 ( .A(n7561), .ZN(n7562) );
  AOI211_X1 U9276 ( .C1(n7564), .C2(n7563), .A(n8579), .B(n7562), .ZN(n7565)
         );
  AOI211_X1 U9277 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(n7567), .A(n7566), .B(
        n7565), .ZN(n7568) );
  INV_X1 U9278 ( .A(n7568), .ZN(P2_U3239) );
  NAND2_X1 U9279 ( .A1(n7571), .A2(n7570), .ZN(n7569) );
  OAI21_X1 U9280 ( .B1(n8606), .B2(n10414), .A(n7569), .ZN(n7576) );
  INV_X1 U9281 ( .A(n8606), .ZN(n7591) );
  OAI21_X1 U9282 ( .B1(n7571), .B2(n7570), .A(n7591), .ZN(n7572) );
  NAND2_X1 U9283 ( .A1(n7572), .A2(n10414), .ZN(n7574) );
  NAND3_X1 U9284 ( .A1(n8607), .A2(n8606), .A3(n10408), .ZN(n7573) );
  AND2_X1 U9285 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  XNOR2_X1 U9286 ( .A(n7671), .B(n7579), .ZN(n7603) );
  INV_X1 U9287 ( .A(n7579), .ZN(n7670) );
  XNOR2_X1 U9288 ( .A(n7578), .B(n7670), .ZN(n7580) );
  AOI222_X1 U9289 ( .A1(n8902), .A2(n7580), .B1(n8604), .B2(n8908), .C1(n8606), 
        .C2(n8907), .ZN(n7602) );
  MUX2_X1 U9290 ( .A(n7581), .B(n7602), .S(n8945), .Z(n7587) );
  OR2_X2 U9291 ( .A1(n7583), .A2(n7669), .ZN(n7684) );
  INV_X1 U9292 ( .A(n7684), .ZN(n7582) );
  AOI21_X1 U9293 ( .B1(n7669), .B2(n7583), .A(n7582), .ZN(n7600) );
  INV_X1 U9294 ( .A(n7595), .ZN(n7584) );
  OAI22_X1 U9295 ( .A1(n8920), .A2(n7592), .B1(n8877), .B2(n7584), .ZN(n7585)
         );
  AOI21_X1 U9296 ( .B1(n8944), .B2(n7600), .A(n7585), .ZN(n7586) );
  OAI211_X1 U9297 ( .C1(n8860), .C2(n7603), .A(n7587), .B(n7586), .ZN(P2_U3289) );
  XNOR2_X1 U9298 ( .A(n7589), .B(n7588), .ZN(n7597) );
  OAI21_X1 U9299 ( .B1(n8537), .B2(n7866), .A(n7590), .ZN(n7594) );
  OAI22_X1 U9300 ( .A1(n7592), .A2(n8570), .B1(n8565), .B2(n7591), .ZN(n7593)
         );
  AOI211_X1 U9301 ( .C1(n7595), .C2(n8588), .A(n7594), .B(n7593), .ZN(n7596)
         );
  OAI21_X1 U9302 ( .B1(n7597), .B2(n8579), .A(n7596), .ZN(P2_U3215) );
  INV_X1 U9303 ( .A(n7598), .ZN(n7610) );
  OAI222_X1 U9304 ( .A1(n10186), .A2(n7610), .B1(n9611), .B2(P1_U3084), .C1(
        n7599), .C2(n10182), .ZN(P1_U3332) );
  INV_X1 U9305 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7605) );
  AOI22_X1 U9306 ( .A1(n7600), .A2(n10424), .B1(n10423), .B2(n7669), .ZN(n7601) );
  OAI211_X1 U9307 ( .C1(n10418), .C2(n7603), .A(n7602), .B(n7601), .ZN(n7606)
         );
  NAND2_X1 U9308 ( .A1(n7606), .A2(n10433), .ZN(n7604) );
  OAI21_X1 U9309 ( .B1(n10433), .B2(n7605), .A(n7604), .ZN(P2_U3472) );
  NAND2_X1 U9310 ( .A1(n7606), .A2(n10444), .ZN(n7607) );
  OAI21_X1 U9311 ( .B1(n10444), .B2(n7608), .A(n7607), .ZN(P2_U3527) );
  OAI222_X1 U9312 ( .A1(n9099), .A2(n7611), .B1(n7652), .B2(n7610), .C1(n7609), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI21_X1 U9313 ( .B1(n7613), .B2(n7081), .A(n7612), .ZN(n7622) );
  INV_X1 U9314 ( .A(n7614), .ZN(n7616) );
  OAI22_X1 U9315 ( .A1(n7616), .A2(n10014), .B1(n10016), .B2(n7615), .ZN(n7621) );
  AND2_X1 U9316 ( .A1(n7617), .A2(n7081), .ZN(n7619) );
  OR2_X1 U9317 ( .A1(n7619), .A2(n7618), .ZN(n7632) );
  NOR2_X1 U9318 ( .A1(n7632), .A2(n10311), .ZN(n7620) );
  AOI211_X1 U9319 ( .C1(n9981), .C2(n7622), .A(n7621), .B(n7620), .ZN(n10260)
         );
  NAND2_X1 U9320 ( .A1(n7624), .A2(n7623), .ZN(n7625) );
  INV_X1 U9321 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7628) );
  OAI22_X1 U9322 ( .A1(n10036), .A2(n7628), .B1(n6985), .B2(n9999), .ZN(n7629)
         );
  AOI21_X1 U9323 ( .B1(n10032), .B2(n4386), .A(n7629), .ZN(n7636) );
  AND2_X1 U9324 ( .A1(n7630), .A2(n9740), .ZN(n7631) );
  NAND2_X1 U9325 ( .A1(n10036), .A2(n7631), .ZN(n9987) );
  INV_X1 U9326 ( .A(n9987), .ZN(n7978) );
  INV_X1 U9327 ( .A(n7632), .ZN(n10258) );
  XNOR2_X1 U9328 ( .A(n4386), .B(n7820), .ZN(n7634) );
  NOR2_X1 U9329 ( .A1(n10320), .A2(n7634), .ZN(n10257) );
  AOI22_X1 U9330 ( .A1(n7978), .A2(n10258), .B1(n10019), .B2(n10257), .ZN(
        n7635) );
  OAI211_X1 U9331 ( .C1(n10260), .C2(n10021), .A(n7636), .B(n7635), .ZN(
        P1_U3290) );
  XOR2_X1 U9332 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n7765), .Z(n7648) );
  INV_X1 U9333 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9334 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9331) );
  OAI21_X1 U9335 ( .B1(n10244), .B2(n7638), .A(n9331), .ZN(n7639) );
  AOI21_X1 U9336 ( .B1(n7769), .B2(n9716), .A(n7639), .ZN(n7647) );
  NAND2_X1 U9337 ( .A1(n7640), .A2(n10001), .ZN(n7644) );
  OR2_X1 U9338 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  NAND2_X1 U9339 ( .A1(n7644), .A2(n7643), .ZN(n7768) );
  XNOR2_X1 U9340 ( .A(n7768), .B(n7769), .ZN(n7645) );
  NAND2_X1 U9341 ( .A1(n7645), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n7772) );
  OAI211_X1 U9342 ( .C1(n7645), .C2(P1_REG2_REG_15__SCAN_IN), .A(n7772), .B(
        n9733), .ZN(n7646) );
  OAI211_X1 U9343 ( .C1(n7648), .C2(n9735), .A(n7647), .B(n7646), .ZN(P1_U3256) );
  INV_X1 U9344 ( .A(n7649), .ZN(n7651) );
  OAI222_X1 U9345 ( .A1(n10182), .A2(n7650), .B1(n10186), .B2(n7651), .C1(
        P1_U3084), .C2(n6392), .ZN(P1_U3331) );
  OAI222_X1 U9346 ( .A1(n9099), .A2(n7653), .B1(n7652), .B2(n7651), .C1(
        P2_U3152), .C2(n5988), .ZN(P2_U3336) );
  XNOR2_X1 U9347 ( .A(n7704), .B(n7705), .ZN(n7707) );
  XOR2_X1 U9348 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n7707), .Z(n7668) );
  INV_X1 U9349 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U9350 ( .A1(n4369), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7655) );
  OAI21_X1 U9351 ( .B1(n8643), .B2(n7656), .A(n7655), .ZN(n7665) );
  OR2_X1 U9352 ( .A1(n7657), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9353 ( .A1(n7659), .A2(n7658), .ZN(n7660) );
  OR2_X1 U9354 ( .A1(n7660), .A2(n7705), .ZN(n7661) );
  NAND2_X1 U9355 ( .A1(n7662), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7663) );
  AOI21_X1 U9356 ( .B1(n7710), .B2(n7663), .A(n8637), .ZN(n7664) );
  AOI211_X1 U9357 ( .C1(n10354), .C2(n7666), .A(n7665), .B(n7664), .ZN(n7667)
         );
  OAI21_X1 U9358 ( .B1(n7668), .B2(n7719), .A(n7667), .ZN(P2_U3260) );
  NAND2_X1 U9359 ( .A1(n7672), .A2(n7677), .ZN(n7673) );
  NAND2_X1 U9360 ( .A1(n7802), .A2(n7673), .ZN(n10428) );
  INV_X1 U9361 ( .A(n7674), .ZN(n7675) );
  NAND2_X1 U9362 ( .A1(n8945), .A2(n7675), .ZN(n8898) );
  OAI21_X1 U9363 ( .B1(n7678), .B2(n7677), .A(n7676), .ZN(n7681) );
  OAI22_X1 U9364 ( .A1(n7839), .A2(n8793), .B1(n8132), .B2(n8795), .ZN(n7680)
         );
  NOR2_X1 U9365 ( .A1(n10428), .A2(n8890), .ZN(n7679) );
  AOI211_X1 U9366 ( .C1(n8902), .C2(n7681), .A(n7680), .B(n7679), .ZN(n10427)
         );
  MUX2_X1 U9367 ( .A(n7682), .B(n10427), .S(n8945), .Z(n7688) );
  OR2_X2 U9368 ( .A1(n7684), .A2(n4523), .ZN(n7813) );
  INV_X1 U9369 ( .A(n7813), .ZN(n7683) );
  AOI21_X1 U9370 ( .B1(n4523), .B2(n7684), .A(n7683), .ZN(n10425) );
  INV_X1 U9371 ( .A(n7685), .ZN(n7838) );
  OAI22_X1 U9372 ( .A1(n8920), .A2(n7845), .B1(n8877), .B2(n7838), .ZN(n7686)
         );
  AOI21_X1 U9373 ( .B1(n8944), .B2(n10425), .A(n7686), .ZN(n7687) );
  OAI211_X1 U9374 ( .C1(n10428), .C2(n8898), .A(n7688), .B(n7687), .ZN(
        P2_U3288) );
  OR2_X1 U9375 ( .A1(n8297), .A2(n7855), .ZN(n7690) );
  NAND2_X1 U9376 ( .A1(n4378), .A2(n7786), .ZN(n7689) );
  NAND2_X1 U9377 ( .A1(n7690), .A2(n7689), .ZN(n7737) );
  NAND2_X1 U9378 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  NAND2_X1 U9379 ( .A1(n8237), .A2(n9646), .ZN(n7695) );
  OAI21_X1 U9380 ( .B1(n10286), .B2(n7022), .A(n7695), .ZN(n7696) );
  XNOR2_X1 U9381 ( .A(n7696), .B(n9157), .ZN(n7736) );
  OR2_X1 U9382 ( .A1(n7746), .A2(n7736), .ZN(n7848) );
  NAND2_X1 U9383 ( .A1(n7746), .A2(n7736), .ZN(n7697) );
  NAND2_X1 U9384 ( .A1(n7848), .A2(n7697), .ZN(n7698) );
  NOR2_X1 U9385 ( .A1(n7698), .A2(n7737), .ZN(n7850) );
  AOI21_X1 U9386 ( .B1(n7737), .B2(n7698), .A(n7850), .ZN(n7703) );
  OAI22_X1 U9387 ( .A1(n9298), .A2(n10286), .B1(n9320), .B2(n6139), .ZN(n7699)
         );
  AOI211_X1 U9388 ( .C1(n9322), .C2(n9647), .A(n7700), .B(n7699), .ZN(n7702)
         );
  NAND2_X1 U9389 ( .A1(n9305), .A2(n7781), .ZN(n7701) );
  OAI211_X1 U9390 ( .C1(n7703), .C2(n9340), .A(n7702), .B(n7701), .ZN(P1_U3225) );
  XOR2_X1 U9391 ( .A(n8621), .B(P2_REG1_REG_16__SCAN_IN), .Z(n7709) );
  OAI22_X1 U9392 ( .A1(n7707), .A2(n7706), .B1(n7705), .B2(n7704), .ZN(n7708)
         );
  NOR2_X1 U9393 ( .A1(n7708), .A2(n7709), .ZN(n8612) );
  AOI21_X1 U9394 ( .B1(n7709), .B2(n7708), .A(n8612), .ZN(n7720) );
  INV_X1 U9395 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7711) );
  MUX2_X1 U9396 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n7711), .S(n8621), .Z(n7712)
         );
  AOI21_X1 U9397 ( .B1(n7713), .B2(n7712), .A(n8637), .ZN(n7717) );
  NOR2_X1 U9398 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8480), .ZN(n7714) );
  AOI21_X1 U9399 ( .B1(n10347), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7714), .ZN(
        n7715) );
  OAI21_X1 U9400 ( .B1(n8626), .B2(n8621), .A(n7715), .ZN(n7716) );
  AOI21_X1 U9401 ( .B1(n7717), .B2(n8620), .A(n7716), .ZN(n7718) );
  OAI21_X1 U9402 ( .B1(n7720), .B2(n7719), .A(n7718), .ZN(P2_U3261) );
  OAI21_X1 U9403 ( .B1(n7721), .B2(n9471), .A(n7956), .ZN(n7887) );
  AOI21_X1 U9404 ( .B1(n8029), .B2(n8077), .A(n10320), .ZN(n7722) );
  NAND2_X1 U9405 ( .A1(n7722), .A2(n5002), .ZN(n7885) );
  OAI21_X1 U9406 ( .B1(n4479), .B2(n10285), .A(n7885), .ZN(n7726) );
  OAI211_X1 U9407 ( .C1(n5003), .C2(n6411), .A(n7723), .B(n9981), .ZN(n7725)
         );
  AOI22_X1 U9408 ( .A1(n9938), .A2(n9640), .B1(n9936), .B2(n9642), .ZN(n7724)
         );
  NAND2_X1 U9409 ( .A1(n7725), .A2(n7724), .ZN(n7882) );
  AOI211_X1 U9410 ( .C1(n10325), .C2(n7887), .A(n7726), .B(n7882), .ZN(n7729)
         );
  NAND2_X1 U9411 ( .A1(n10326), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7727) );
  OAI21_X1 U9412 ( .B1(n7729), .B2(n10326), .A(n7727), .ZN(P1_U3484) );
  NAND2_X1 U9413 ( .A1(n10341), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7728) );
  OAI21_X1 U9414 ( .B1(n7729), .B2(n10341), .A(n7728), .ZN(P1_U3533) );
  NAND2_X1 U9415 ( .A1(n9159), .A2(n10298), .ZN(n7731) );
  OR2_X1 U9416 ( .A1(n8217), .A2(n7876), .ZN(n7730) );
  NAND2_X1 U9417 ( .A1(n7731), .A2(n7730), .ZN(n7732) );
  XNOR2_X1 U9418 ( .A(n7732), .B(n9157), .ZN(n8046) );
  OR2_X1 U9419 ( .A1(n8297), .A2(n7876), .ZN(n7735) );
  NAND2_X1 U9420 ( .A1(n4378), .A2(n10298), .ZN(n7734) );
  NAND2_X1 U9421 ( .A1(n7735), .A2(n7734), .ZN(n8047) );
  XNOR2_X1 U9422 ( .A(n8046), .B(n8047), .ZN(n7755) );
  AND2_X1 U9423 ( .A1(n7736), .A2(n7737), .ZN(n7745) );
  INV_X1 U9424 ( .A(n7736), .ZN(n7739) );
  INV_X1 U9425 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U9426 ( .A1(n7739), .A2(n7738), .ZN(n7743) );
  NOR2_X1 U9427 ( .A1(n8217), .A2(n6421), .ZN(n7740) );
  AOI21_X1 U9428 ( .B1(n7733), .B2(n9645), .A(n7740), .ZN(n7748) );
  OR2_X1 U9429 ( .A1(n8217), .A2(n6139), .ZN(n7741) );
  OAI21_X1 U9430 ( .B1(n7022), .B2(n6421), .A(n7741), .ZN(n7742) );
  XNOR2_X1 U9431 ( .A(n8295), .B(n7742), .ZN(n7747) );
  NAND2_X1 U9432 ( .A1(n7748), .A2(n7747), .ZN(n7847) );
  AND2_X1 U9433 ( .A1(n7743), .A2(n7847), .ZN(n7744) );
  INV_X1 U9434 ( .A(n7747), .ZN(n7750) );
  INV_X1 U9435 ( .A(n7748), .ZN(n7749) );
  NAND2_X1 U9436 ( .A1(n7750), .A2(n7749), .ZN(n7846) );
  INV_X1 U9437 ( .A(n7751), .ZN(n7753) );
  INV_X1 U9438 ( .A(n8051), .ZN(n7754) );
  AOI21_X1 U9439 ( .B1(n7755), .B2(n7751), .A(n7754), .ZN(n7761) );
  AOI21_X1 U9440 ( .B1(n9322), .B2(n9645), .A(n7756), .ZN(n7758) );
  NAND2_X1 U9441 ( .A1(n9305), .A2(n7902), .ZN(n7757) );
  OAI211_X1 U9442 ( .C1(n8054), .C2(n9320), .A(n7758), .B(n7757), .ZN(n7759)
         );
  AOI21_X1 U9443 ( .B1(n9338), .B2(n10298), .A(n7759), .ZN(n7760) );
  OAI21_X1 U9444 ( .B1(n7761), .B2(n9340), .A(n7760), .ZN(P1_U3211) );
  INV_X1 U9445 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7764) );
  OAI22_X1 U9446 ( .A1(n7765), .A2(n7764), .B1(n7763), .B2(n7762), .ZN(n7937)
         );
  XOR2_X1 U9447 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n7941), .Z(n7936) );
  XNOR2_X1 U9448 ( .A(n7937), .B(n7936), .ZN(n7777) );
  INV_X1 U9449 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U9450 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9230) );
  OAI21_X1 U9451 ( .B1(n10244), .B2(n7766), .A(n9230), .ZN(n7767) );
  AOI21_X1 U9452 ( .B1(n7941), .B2(n9716), .A(n7767), .ZN(n7776) );
  INV_X1 U9453 ( .A(n7768), .ZN(n7770) );
  NAND2_X1 U9454 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  NAND2_X1 U9455 ( .A1(n7772), .A2(n7771), .ZN(n7774) );
  INV_X1 U9456 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9967) );
  XNOR2_X1 U9457 ( .A(n7941), .B(n9967), .ZN(n7773) );
  NAND2_X1 U9458 ( .A1(n7774), .A2(n7773), .ZN(n7943) );
  OAI211_X1 U9459 ( .C1(n7774), .C2(n7773), .A(n7943), .B(n9733), .ZN(n7775)
         );
  OAI211_X1 U9460 ( .C1(n7777), .C2(n9735), .A(n7776), .B(n7775), .ZN(P1_U3257) );
  INV_X1 U9461 ( .A(n7788), .ZN(n9587) );
  OAI222_X1 U9462 ( .A1(n10016), .A2(n6139), .B1(n10014), .B2(n7780), .C1(
        n10012), .C2(n7779), .ZN(n10288) );
  INV_X1 U9463 ( .A(n10288), .ZN(n7794) );
  INV_X1 U9464 ( .A(n7781), .ZN(n7782) );
  OAI22_X1 U9465 ( .A1(n10036), .A2(n7783), .B1(n7782), .B2(n9999), .ZN(n7785)
         );
  OAI211_X1 U9466 ( .C1(n8013), .C2(n10286), .A(n10307), .B(n7830), .ZN(n10283) );
  NOR2_X1 U9467 ( .A1(n7917), .A2(n10283), .ZN(n7784) );
  AOI211_X1 U9468 ( .C1(n10032), .C2(n7786), .A(n7785), .B(n7784), .ZN(n7793)
         );
  INV_X1 U9469 ( .A(n7787), .ZN(n7789) );
  NAND2_X1 U9470 ( .A1(n7789), .A2(n7788), .ZN(n10282) );
  AND2_X1 U9471 ( .A1(n7790), .A2(n9157), .ZN(n7791) );
  NAND2_X1 U9472 ( .A1(n7787), .A2(n9587), .ZN(n10281) );
  NAND3_X1 U9473 ( .A1(n10282), .A2(n10041), .A3(n10281), .ZN(n7792) );
  OAI211_X1 U9474 ( .C1(n7794), .C2(n10021), .A(n7793), .B(n7792), .ZN(
        P1_U3286) );
  INV_X1 U9475 ( .A(n7795), .ZN(n7800) );
  NOR2_X1 U9476 ( .A1(n7796), .A2(P1_U3084), .ZN(n9625) );
  AOI21_X1 U9477 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10176), .A(n9625), .ZN(
        n7797) );
  OAI21_X1 U9478 ( .B1(n7800), .B2(n10186), .A(n7797), .ZN(P1_U3330) );
  AOI21_X1 U9479 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9093), .A(n7798), .ZN(
        n7799) );
  OAI21_X1 U9480 ( .B1(n7800), .B2(n9101), .A(n7799), .ZN(P2_U3335) );
  NAND2_X1 U9481 ( .A1(n4523), .A2(n8604), .ZN(n7801) );
  INV_X1 U9482 ( .A(n8001), .ZN(n7803) );
  NAND2_X1 U9483 ( .A1(n7803), .A2(n7805), .ZN(n8122) );
  OAI21_X1 U9484 ( .B1(n7803), .B2(n7805), .A(n8122), .ZN(n7810) );
  INV_X1 U9485 ( .A(n7810), .ZN(n9065) );
  OAI22_X1 U9486 ( .A1(n7866), .A2(n8793), .B1(n7922), .B2(n8795), .ZN(n7809)
         );
  NAND3_X1 U9487 ( .A1(n7676), .A2(n7806), .A3(n7805), .ZN(n7807) );
  AOI21_X1 U9488 ( .B1(n8126), .B2(n7807), .A(n8868), .ZN(n7808) );
  AOI211_X1 U9489 ( .C1(n7811), .C2(n7810), .A(n7809), .B(n7808), .ZN(n9064)
         );
  MUX2_X1 U9490 ( .A(n7812), .B(n9064), .S(n8945), .Z(n7817) );
  AOI21_X1 U9491 ( .B1(n9061), .B2(n7813), .A(n8137), .ZN(n9062) );
  INV_X1 U9492 ( .A(n9061), .ZN(n7871) );
  INV_X1 U9493 ( .A(n7814), .ZN(n7865) );
  OAI22_X1 U9494 ( .A1(n8920), .A2(n7871), .B1(n8877), .B2(n7865), .ZN(n7815)
         );
  AOI21_X1 U9495 ( .B1(n9062), .B2(n8944), .A(n7815), .ZN(n7816) );
  OAI211_X1 U9496 ( .C1(n9065), .C2(n8898), .A(n7817), .B(n7816), .ZN(P2_U3287) );
  INV_X1 U9497 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7824) );
  OR2_X1 U9498 ( .A1(n7818), .A2(n9623), .ZN(n7819) );
  OAI21_X1 U9499 ( .B1(n9990), .B2(n10032), .A(n7820), .ZN(n7823) );
  INV_X1 U9500 ( .A(n9999), .ZN(n10029) );
  AOI22_X1 U9501 ( .A1(n10036), .A2(n7821), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10029), .ZN(n7822) );
  OAI211_X1 U9502 ( .C1(n7824), .C2(n10036), .A(n7823), .B(n7822), .ZN(
        P1_U3291) );
  NAND2_X1 U9503 ( .A1(n10282), .A2(n7825), .ZN(n7826) );
  XNOR2_X1 U9504 ( .A(n7826), .B(n9584), .ZN(n10292) );
  NAND2_X1 U9505 ( .A1(n9437), .A2(n9439), .ZN(n7827) );
  INV_X1 U9506 ( .A(n9584), .ZN(n9438) );
  XNOR2_X1 U9507 ( .A(n7827), .B(n9438), .ZN(n7828) );
  AOI222_X1 U9508 ( .A1(n9981), .A2(n7828), .B1(n9644), .B2(n9938), .C1(n9646), 
        .C2(n9936), .ZN(n10293) );
  MUX2_X1 U9509 ( .A(n6844), .B(n10293), .S(n10036), .Z(n7834) );
  INV_X1 U9510 ( .A(n7899), .ZN(n7829) );
  AOI21_X1 U9511 ( .B1(n7853), .B2(n7830), .A(n7829), .ZN(n10289) );
  INV_X1 U9512 ( .A(n7858), .ZN(n7831) );
  OAI22_X1 U9513 ( .A1(n10024), .A2(n6421), .B1(n7831), .B2(n9999), .ZN(n7832)
         );
  AOI21_X1 U9514 ( .B1(n10289), .B2(n9990), .A(n7832), .ZN(n7833) );
  OAI211_X1 U9515 ( .C1(n10028), .C2(n10292), .A(n7834), .B(n7833), .ZN(
        P1_U3285) );
  XOR2_X1 U9516 ( .A(n7836), .B(n7835), .Z(n7837) );
  NAND2_X1 U9517 ( .A1(n7837), .A2(n8583), .ZN(n7844) );
  OAI22_X1 U9518 ( .A1(n7839), .A2(n8565), .B1(n8564), .B2(n7838), .ZN(n7842)
         );
  OAI21_X1 U9519 ( .B1(n8537), .B2(n8132), .A(n7840), .ZN(n7841) );
  NOR2_X1 U9520 ( .A1(n7842), .A2(n7841), .ZN(n7843) );
  OAI211_X1 U9521 ( .C1(n7845), .C2(n8570), .A(n7844), .B(n7843), .ZN(P2_U3223) );
  NAND2_X1 U9522 ( .A1(n7847), .A2(n7846), .ZN(n7852) );
  INV_X1 U9523 ( .A(n7848), .ZN(n7849) );
  NOR2_X1 U9524 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  XOR2_X1 U9525 ( .A(n7852), .B(n7851), .Z(n7860) );
  NAND2_X1 U9526 ( .A1(n10299), .A2(n7853), .ZN(n10290) );
  OAI22_X1 U9527 ( .A1(n9320), .A2(n7876), .B1(n9264), .B2(n10290), .ZN(n7857)
         );
  INV_X1 U9528 ( .A(n9322), .ZN(n9332) );
  OAI21_X1 U9529 ( .B1(n9332), .B2(n7855), .A(n7854), .ZN(n7856) );
  AOI211_X1 U9530 ( .C1(n7858), .C2(n9305), .A(n7857), .B(n7856), .ZN(n7859)
         );
  OAI21_X1 U9531 ( .B1(n7860), .B2(n9340), .A(n7859), .ZN(P1_U3237) );
  OAI21_X1 U9532 ( .B1(n7863), .B2(n7862), .A(n7861), .ZN(n7864) );
  NAND2_X1 U9533 ( .A1(n7864), .A2(n8583), .ZN(n7870) );
  OAI22_X1 U9534 ( .A1(n7866), .A2(n8565), .B1(n8564), .B2(n7865), .ZN(n7867)
         );
  AOI211_X1 U9535 ( .C1(n8589), .C2(n8602), .A(n7868), .B(n7867), .ZN(n7869)
         );
  OAI211_X1 U9536 ( .C1(n7871), .C2(n8570), .A(n7870), .B(n7869), .ZN(P2_U3233) );
  OAI21_X1 U9537 ( .B1(n7872), .B2(n6155), .A(n7873), .ZN(n10312) );
  NAND2_X1 U9538 ( .A1(n7892), .A2(n9454), .ZN(n7874) );
  XOR2_X1 U9539 ( .A(n9590), .B(n7874), .Z(n7875) );
  OAI222_X1 U9540 ( .A1(n10016), .A2(n8061), .B1(n10014), .B2(n7876), .C1(
        n7875), .C2(n10012), .ZN(n10313) );
  NAND2_X1 U9541 ( .A1(n10313), .A2(n10036), .ZN(n7881) );
  AOI21_X1 U9542 ( .B1(n9177), .B2(n7900), .A(n8031), .ZN(n10308) );
  INV_X1 U9543 ( .A(n9177), .ZN(n7878) );
  AOI22_X1 U9544 ( .A1(n10021), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9184), .B2(
        n10029), .ZN(n7877) );
  OAI21_X1 U9545 ( .B1(n7878), .B2(n10024), .A(n7877), .ZN(n7879) );
  AOI21_X1 U9546 ( .B1(n10308), .B2(n9990), .A(n7879), .ZN(n7880) );
  OAI211_X1 U9547 ( .C1(n10028), .C2(n10312), .A(n7881), .B(n7880), .ZN(
        P1_U3283) );
  INV_X1 U9548 ( .A(n7882), .ZN(n7889) );
  INV_X1 U9549 ( .A(n10019), .ZN(n7917) );
  AOI22_X1 U9550 ( .A1(n10021), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8078), .B2(
        n10029), .ZN(n7884) );
  NAND2_X1 U9551 ( .A1(n10032), .A2(n8077), .ZN(n7883) );
  OAI211_X1 U9552 ( .C1(n7885), .C2(n7917), .A(n7884), .B(n7883), .ZN(n7886)
         );
  AOI21_X1 U9553 ( .B1(n7887), .B2(n10041), .A(n7886), .ZN(n7888) );
  OAI21_X1 U9554 ( .B1(n10021), .B2(n7889), .A(n7888), .ZN(P1_U3281) );
  NAND2_X1 U9555 ( .A1(n7890), .A2(n6410), .ZN(n7891) );
  NAND2_X1 U9556 ( .A1(n7892), .A2(n7891), .ZN(n7894) );
  OAI22_X1 U9557 ( .A1(n6139), .A2(n10014), .B1(n10016), .B2(n8054), .ZN(n7893) );
  AOI21_X1 U9558 ( .B1(n7894), .B2(n9981), .A(n7893), .ZN(n10305) );
  INV_X1 U9559 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U9560 ( .A1(n7897), .A2(n7896), .ZN(n7898) );
  XNOR2_X1 U9561 ( .A(n7898), .B(n6410), .ZN(n10303) );
  AOI21_X1 U9562 ( .B1(n7899), .B2(n10298), .A(n10320), .ZN(n7901) );
  NAND2_X1 U9563 ( .A1(n7901), .A2(n7900), .ZN(n10301) );
  AOI22_X1 U9564 ( .A1(n10021), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7902), .B2(
        n10029), .ZN(n7904) );
  NAND2_X1 U9565 ( .A1(n10032), .A2(n10298), .ZN(n7903) );
  OAI211_X1 U9566 ( .C1(n10301), .C2(n7917), .A(n7904), .B(n7903), .ZN(n7905)
         );
  AOI21_X1 U9567 ( .B1(n10303), .B2(n10041), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9568 ( .B1(n10305), .B2(n10021), .A(n7906), .ZN(P1_U3284) );
  INV_X1 U9569 ( .A(n7908), .ZN(n7909) );
  AOI21_X1 U9570 ( .B1(n7961), .B2(n9472), .A(n7909), .ZN(n7910) );
  XOR2_X1 U9571 ( .A(n9595), .B(n7910), .Z(n7911) );
  OAI222_X1 U9572 ( .A1(n10016), .A2(n9996), .B1(n10014), .B2(n8196), .C1(
        n10012), .C2(n7911), .ZN(n10147) );
  INV_X1 U9573 ( .A(n10147), .ZN(n7920) );
  INV_X1 U9574 ( .A(n7912), .ZN(n7913) );
  AOI21_X1 U9575 ( .B1(n9595), .B2(n7914), .A(n7913), .ZN(n10149) );
  OAI211_X1 U9576 ( .C1(n7958), .C2(n10146), .A(n10018), .B(n10307), .ZN(
        n10145) );
  AOI22_X1 U9577 ( .A1(n10021), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9207), .B2(
        n10029), .ZN(n7916) );
  NAND2_X1 U9578 ( .A1(n10032), .A2(n8206), .ZN(n7915) );
  OAI211_X1 U9579 ( .C1(n10145), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7918)
         );
  AOI21_X1 U9580 ( .B1(n10149), .B2(n10041), .A(n7918), .ZN(n7919) );
  OAI21_X1 U9581 ( .B1(n7920), .B2(n10021), .A(n7919), .ZN(P1_U3279) );
  INV_X1 U9582 ( .A(n8132), .ZN(n8603) );
  OR2_X1 U9583 ( .A1(n8603), .A2(n9061), .ZN(n8121) );
  NAND2_X1 U9584 ( .A1(n8124), .A2(n8121), .ZN(n7998) );
  INV_X1 U9585 ( .A(n7998), .ZN(n7925) );
  NAND3_X1 U9586 ( .A1(n7921), .A2(n8124), .A3(n8121), .ZN(n7924) );
  OR2_X1 U9587 ( .A1(n7922), .A2(n8142), .ZN(n7923) );
  NAND2_X1 U9588 ( .A1(n7924), .A2(n7923), .ZN(n8002) );
  AOI21_X1 U9589 ( .B1(n8001), .B2(n7925), .A(n8002), .ZN(n7926) );
  XNOR2_X1 U9590 ( .A(n7926), .B(n7999), .ZN(n9055) );
  INV_X1 U9591 ( .A(n7999), .ZN(n8003) );
  XNOR2_X1 U9592 ( .A(n8131), .B(n8003), .ZN(n7929) );
  OR2_X1 U9593 ( .A1(n8153), .A2(n8795), .ZN(n7928) );
  NAND2_X1 U9594 ( .A1(n8602), .A2(n8907), .ZN(n7927) );
  NAND2_X1 U9595 ( .A1(n7928), .A2(n7927), .ZN(n8547) );
  AOI21_X1 U9596 ( .B1(n7929), .B2(n8902), .A(n8547), .ZN(n9054) );
  MUX2_X1 U9597 ( .A(n9054), .B(n7930), .S(n8924), .Z(n7935) );
  NAND2_X1 U9598 ( .A1(n8137), .A2(n8142), .ZN(n8138) );
  INV_X1 U9599 ( .A(n5014), .ZN(n7931) );
  AOI211_X1 U9600 ( .C1(n9052), .C2(n8138), .A(n10400), .B(n7931), .ZN(n9051)
         );
  INV_X1 U9601 ( .A(n9052), .ZN(n8554) );
  INV_X1 U9602 ( .A(n8551), .ZN(n7932) );
  OAI22_X1 U9603 ( .A1(n8920), .A2(n8554), .B1(n8877), .B2(n7932), .ZN(n7933)
         );
  AOI21_X1 U9604 ( .B1(n9051), .B2(n8818), .A(n7933), .ZN(n7934) );
  OAI211_X1 U9605 ( .C1(n9055), .C2(n8860), .A(n7935), .B(n7934), .ZN(P2_U3285) );
  AOI22_X1 U9606 ( .A1(n7937), .A2(n7936), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n7941), .ZN(n8106) );
  XNOR2_X1 U9607 ( .A(n8112), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8105) );
  XNOR2_X1 U9608 ( .A(n8106), .B(n8105), .ZN(n7949) );
  NOR2_X1 U9609 ( .A1(n7938), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9251) );
  INV_X1 U9610 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7939) );
  NOR2_X1 U9611 ( .A1(n10244), .A2(n7939), .ZN(n7940) );
  AOI211_X1 U9612 ( .C1(n9716), .C2(n8112), .A(n9251), .B(n7940), .ZN(n7948)
         );
  NAND2_X1 U9613 ( .A1(n7941), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U9614 ( .A1(n7943), .A2(n7942), .ZN(n7946) );
  INV_X1 U9615 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7944) );
  XNOR2_X1 U9616 ( .A(n8112), .B(n7944), .ZN(n7945) );
  NAND2_X1 U9617 ( .A1(n7946), .A2(n7945), .ZN(n8114) );
  OAI211_X1 U9618 ( .C1(n7946), .C2(n7945), .A(n8114), .B(n9733), .ZN(n7947)
         );
  OAI211_X1 U9619 ( .C1(n7949), .C2(n9735), .A(n7948), .B(n7947), .ZN(P1_U3258) );
  INV_X1 U9620 ( .A(n7950), .ZN(n7982) );
  OAI222_X1 U9621 ( .A1(n10186), .A2(n7982), .B1(P1_U3084), .B2(n7952), .C1(
        n7951), .C2(n10182), .ZN(P1_U3329) );
  NAND2_X1 U9622 ( .A1(n7954), .A2(n7953), .ZN(n9593) );
  NAND2_X1 U9623 ( .A1(n7956), .A2(n7955), .ZN(n7957) );
  XOR2_X1 U9624 ( .A(n9593), .B(n7957), .Z(n10040) );
  AND2_X1 U9625 ( .A1(n5002), .A2(n10031), .ZN(n7959) );
  OR2_X1 U9626 ( .A1(n7959), .A2(n7958), .ZN(n10035) );
  INV_X1 U9627 ( .A(n10031), .ZN(n7960) );
  OAI22_X1 U9628 ( .A1(n10035), .A2(n10320), .B1(n7960), .B2(n10285), .ZN(
        n7963) );
  XNOR2_X1 U9629 ( .A(n7961), .B(n9593), .ZN(n7962) );
  OAI222_X1 U9630 ( .A1(n10016), .A2(n10013), .B1(n10014), .B2(n8073), .C1(
        n7962), .C2(n10012), .ZN(n10037) );
  AOI211_X1 U9631 ( .C1(n10040), .C2(n10325), .A(n7963), .B(n10037), .ZN(n7966) );
  NAND2_X1 U9632 ( .A1(n10341), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7964) );
  OAI21_X1 U9633 ( .B1(n7966), .B2(n10341), .A(n7964), .ZN(P1_U3534) );
  NAND2_X1 U9634 ( .A1(n10326), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7965) );
  OAI21_X1 U9635 ( .B1(n7966), .B2(n10326), .A(n7965), .ZN(P1_U3487) );
  XOR2_X1 U9636 ( .A(n7967), .B(n9581), .Z(n7971) );
  AOI22_X1 U9637 ( .A1(n9936), .A2(n7075), .B1(n9938), .B2(n9647), .ZN(n7970)
         );
  OAI21_X1 U9638 ( .B1(n9581), .B2(n9554), .A(n8010), .ZN(n7968) );
  NAND2_X1 U9639 ( .A1(n7968), .A2(n9981), .ZN(n7969) );
  OAI211_X1 U9640 ( .C1(n7971), .C2(n10311), .A(n7970), .B(n7969), .ZN(n10268)
         );
  INV_X1 U9641 ( .A(n10268), .ZN(n7980) );
  INV_X1 U9642 ( .A(n7971), .ZN(n10270) );
  INV_X1 U9643 ( .A(n10265), .ZN(n7974) );
  NAND2_X1 U9644 ( .A1(n7973), .A2(n7972), .ZN(n10264) );
  NAND3_X1 U9645 ( .A1(n9990), .A2(n7974), .A3(n10264), .ZN(n7976) );
  AOI22_X1 U9646 ( .A1(n10021), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10029), .B2(
        n6078), .ZN(n7975) );
  OAI211_X1 U9647 ( .C1(n10267), .C2(n10024), .A(n7976), .B(n7975), .ZN(n7977)
         );
  AOI21_X1 U9648 ( .B1(n7978), .B2(n10270), .A(n7977), .ZN(n7979) );
  OAI21_X1 U9649 ( .B1(n7980), .B2(n10021), .A(n7979), .ZN(P1_U3288) );
  OAI222_X1 U9650 ( .A1(P2_U3152), .A2(n7983), .B1(n9101), .B2(n7982), .C1(
        n7981), .C2(n9099), .ZN(P2_U3334) );
  AOI22_X1 U9651 ( .A1(n10021), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10029), .ZN(n7984) );
  OAI21_X1 U9652 ( .B1(n10034), .B2(n7985), .A(n7984), .ZN(n7986) );
  AOI21_X1 U9653 ( .B1(n10032), .B2(n7987), .A(n7986), .ZN(n7990) );
  NAND2_X1 U9654 ( .A1(n7988), .A2(n10036), .ZN(n7989) );
  OAI211_X1 U9655 ( .C1(n7991), .C2(n9987), .A(n7990), .B(n7989), .ZN(P1_U3289) );
  OAI211_X1 U9656 ( .C1(n8148), .C2(n7993), .A(n7992), .B(n8902), .ZN(n7995)
         );
  INV_X1 U9657 ( .A(n8458), .ZN(n8599) );
  INV_X1 U9658 ( .A(n8455), .ZN(n8601) );
  AOI22_X1 U9659 ( .A1(n8908), .A2(n8599), .B1(n8601), .B2(n8907), .ZN(n7994)
         );
  AND2_X1 U9660 ( .A1(n7995), .A2(n7994), .ZN(n9049) );
  AOI21_X1 U9661 ( .B1(n9046), .B2(n5014), .A(n8158), .ZN(n9047) );
  INV_X1 U9662 ( .A(n9046), .ZN(n7997) );
  INV_X1 U9663 ( .A(n8877), .ZN(n8942) );
  AOI22_X1 U9664 ( .A1(n8924), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n8456), .B2(
        n8942), .ZN(n7996) );
  OAI21_X1 U9665 ( .B1(n8920), .B2(n7997), .A(n7996), .ZN(n8007) );
  NOR2_X1 U9666 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  NAND2_X1 U9667 ( .A1(n8001), .A2(n8000), .ZN(n8005) );
  XOR2_X1 U9668 ( .A(n8149), .B(n8148), .Z(n9050) );
  NOR2_X1 U9669 ( .A1(n9050), .A2(n8860), .ZN(n8006) );
  AOI211_X1 U9670 ( .C1(n9047), .C2(n8944), .A(n8007), .B(n8006), .ZN(n8008)
         );
  OAI21_X1 U9671 ( .B1(n8924), .B2(n9049), .A(n8008), .ZN(P2_U3284) );
  XOR2_X1 U9672 ( .A(n8009), .B(n9583), .Z(n10273) );
  NAND2_X1 U9673 ( .A1(n8010), .A2(n9558), .ZN(n8011) );
  XOR2_X1 U9674 ( .A(n9583), .B(n8011), .Z(n8012) );
  AOI222_X1 U9675 ( .A1(n9981), .A2(n8012), .B1(n9646), .B2(n9938), .C1(n9648), 
        .C2(n9936), .ZN(n10276) );
  MUX2_X1 U9676 ( .A(n6836), .B(n10276), .S(n10036), .Z(n8021) );
  INV_X1 U9677 ( .A(n8013), .ZN(n8014) );
  OAI21_X1 U9678 ( .B1(n8015), .B2(n10265), .A(n8014), .ZN(n10275) );
  INV_X1 U9679 ( .A(n8016), .ZN(n8017) );
  OAI22_X1 U9680 ( .A1(n10034), .A2(n10275), .B1(n8017), .B2(n9999), .ZN(n8018) );
  AOI21_X1 U9681 ( .B1(n10032), .B2(n8019), .A(n8018), .ZN(n8020) );
  OAI211_X1 U9682 ( .C1(n10273), .C2(n10028), .A(n8021), .B(n8020), .ZN(
        P1_U3287) );
  NAND2_X1 U9683 ( .A1(n8022), .A2(n9457), .ZN(n8026) );
  INV_X1 U9684 ( .A(n8023), .ZN(n8025) );
  OR2_X1 U9685 ( .A1(n8025), .A2(n8024), .ZN(n9586) );
  XNOR2_X1 U9686 ( .A(n8026), .B(n9586), .ZN(n8027) );
  OAI222_X1 U9687 ( .A1(n10014), .A2(n8054), .B1(n10016), .B2(n8073), .C1(
        n8027), .C2(n10012), .ZN(n10322) );
  INV_X1 U9688 ( .A(n10322), .ZN(n8036) );
  XNOR2_X1 U9689 ( .A(n8028), .B(n9586), .ZN(n10324) );
  OAI21_X1 U9690 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n10321) );
  AOI22_X1 U9691 ( .A1(n10021), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8095), .B2(
        n10029), .ZN(n8033) );
  NAND2_X1 U9692 ( .A1(n10032), .A2(n8093), .ZN(n8032) );
  OAI211_X1 U9693 ( .C1(n10321), .C2(n10034), .A(n8033), .B(n8032), .ZN(n8034)
         );
  AOI21_X1 U9694 ( .B1(n10324), .B2(n10041), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9695 ( .B1(n8036), .B2(n10021), .A(n8035), .ZN(P1_U3282) );
  XOR2_X1 U9696 ( .A(n8038), .B(n8037), .Z(n8039) );
  NAND2_X1 U9697 ( .A1(n8039), .A2(n8583), .ZN(n8045) );
  INV_X1 U9698 ( .A(n8040), .ZN(n8141) );
  OAI22_X1 U9699 ( .A1(n8132), .A2(n8565), .B1(n8564), .B2(n8141), .ZN(n8043)
         );
  OAI21_X1 U9700 ( .B1(n8537), .B2(n8455), .A(n8041), .ZN(n8042) );
  NOR2_X1 U9701 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  OAI211_X1 U9702 ( .C1(n8142), .C2(n8570), .A(n8045), .B(n8044), .ZN(P2_U3219) );
  INV_X1 U9703 ( .A(n8046), .ZN(n8049) );
  INV_X1 U9704 ( .A(n8047), .ZN(n8048) );
  NAND2_X1 U9705 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  OR2_X1 U9706 ( .A1(n8297), .A2(n8054), .ZN(n8053) );
  NAND2_X1 U9707 ( .A1(n9177), .A2(n8237), .ZN(n8052) );
  NAND2_X1 U9708 ( .A1(n8053), .A2(n8052), .ZN(n8086) );
  NAND2_X1 U9709 ( .A1(n9177), .A2(n9159), .ZN(n8056) );
  OR2_X1 U9710 ( .A1(n8217), .A2(n8054), .ZN(n8055) );
  NAND2_X1 U9711 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  XNOR2_X1 U9712 ( .A(n8057), .B(n9157), .ZN(n9181) );
  NAND2_X1 U9713 ( .A1(n8093), .A2(n9159), .ZN(n8059) );
  NAND2_X1 U9714 ( .A1(n4378), .A2(n9642), .ZN(n8058) );
  NAND2_X1 U9715 ( .A1(n8059), .A2(n8058), .ZN(n8060) );
  XNOR2_X1 U9716 ( .A(n8060), .B(n9157), .ZN(n8065) );
  OR2_X1 U9717 ( .A1(n8297), .A2(n8061), .ZN(n8063) );
  NAND2_X1 U9718 ( .A1(n8093), .A2(n4378), .ZN(n8062) );
  NAND2_X1 U9719 ( .A1(n8063), .A2(n8062), .ZN(n8089) );
  AOI22_X1 U9720 ( .A1(n8086), .A2(n9181), .B1(n8065), .B2(n8089), .ZN(n8064)
         );
  OAI21_X1 U9721 ( .B1(n9181), .B2(n8086), .A(n8089), .ZN(n8068) );
  INV_X1 U9722 ( .A(n8065), .ZN(n8090) );
  INV_X1 U9723 ( .A(n9181), .ZN(n8067) );
  NOR2_X1 U9724 ( .A1(n8086), .A2(n8089), .ZN(n8066) );
  AOI22_X1 U9725 ( .A1(n8068), .A2(n8090), .B1(n8067), .B2(n8066), .ZN(n8069)
         );
  NAND2_X1 U9726 ( .A1(n8077), .A2(n9159), .ZN(n8071) );
  OR2_X1 U9727 ( .A1(n8217), .A2(n8073), .ZN(n8070) );
  NAND2_X1 U9728 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  XNOR2_X1 U9729 ( .A(n8072), .B(n8295), .ZN(n8191) );
  OR2_X1 U9730 ( .A1(n8297), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U9731 ( .A1(n8077), .A2(n8237), .ZN(n8074) );
  NAND2_X1 U9732 ( .A1(n8075), .A2(n8074), .ZN(n8189) );
  XNOR2_X1 U9733 ( .A(n8191), .B(n8189), .ZN(n8187) );
  XNOR2_X1 U9734 ( .A(n8188), .B(n8187), .ZN(n8084) );
  AOI21_X1 U9735 ( .B1(n9322), .B2(n9642), .A(n8076), .ZN(n8082) );
  NAND2_X1 U9736 ( .A1(n9338), .A2(n8077), .ZN(n8081) );
  NAND2_X1 U9737 ( .A1(n9305), .A2(n8078), .ZN(n8080) );
  NAND2_X1 U9738 ( .A1(n9334), .A2(n9640), .ZN(n8079) );
  NAND4_X1 U9739 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n8083)
         );
  AOI21_X1 U9740 ( .B1(n8084), .B2(n9311), .A(n8083), .ZN(n8085) );
  INV_X1 U9741 ( .A(n8085), .ZN(P1_U3215) );
  INV_X1 U9742 ( .A(n8086), .ZN(n8087) );
  NOR2_X1 U9743 ( .A1(n8088), .A2(n8087), .ZN(n9178) );
  NAND2_X1 U9744 ( .A1(n8088), .A2(n8087), .ZN(n9179) );
  OAI21_X1 U9745 ( .B1(n9178), .B2(n9181), .A(n9179), .ZN(n8092) );
  XNOR2_X1 U9746 ( .A(n8090), .B(n8089), .ZN(n8091) );
  XNOR2_X1 U9747 ( .A(n8092), .B(n8091), .ZN(n8101) );
  AND2_X1 U9748 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9695) );
  AOI21_X1 U9749 ( .B1(n9322), .B2(n9643), .A(n9695), .ZN(n8099) );
  AND2_X1 U9750 ( .A1(n10299), .A2(n8093), .ZN(n10318) );
  NAND2_X1 U9751 ( .A1(n8094), .A2(n10318), .ZN(n8098) );
  NAND2_X1 U9752 ( .A1(n9305), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U9753 ( .A1(n9334), .A2(n9641), .ZN(n8096) );
  NAND4_X1 U9754 ( .A1(n8099), .A2(n8098), .A3(n8097), .A4(n8096), .ZN(n8100)
         );
  AOI21_X1 U9755 ( .B1(n8101), .B2(n9311), .A(n8100), .ZN(n8102) );
  INV_X1 U9756 ( .A(n8102), .ZN(P1_U3229) );
  OAI22_X1 U9757 ( .A1(n8106), .A2(n8105), .B1(n8104), .B2(n8103), .ZN(n8110)
         );
  INV_X1 U9758 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U9759 ( .A1(n8108), .A2(n8107), .ZN(n9723) );
  OAI21_X1 U9760 ( .B1(n8108), .B2(n8107), .A(n9723), .ZN(n8109) );
  AOI21_X1 U9761 ( .B1(n8110), .B2(n8109), .A(n9725), .ZN(n8120) );
  NAND2_X1 U9762 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9319) );
  OAI21_X1 U9763 ( .B1(n10244), .B2(n10479), .A(n9319), .ZN(n8111) );
  AOI21_X1 U9764 ( .B1(n9728), .B2(n9716), .A(n8111), .ZN(n8119) );
  NAND2_X1 U9765 ( .A1(n8112), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U9766 ( .A1(n8114), .A2(n8113), .ZN(n8117) );
  INV_X1 U9767 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8115) );
  MUX2_X1 U9768 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n8115), .S(n9728), .Z(n8116)
         );
  NAND2_X1 U9769 ( .A1(n8117), .A2(n8116), .ZN(n9730) );
  OAI211_X1 U9770 ( .C1(n8117), .C2(n8116), .A(n9730), .B(n9733), .ZN(n8118)
         );
  OAI211_X1 U9771 ( .C1(n8120), .C2(n9735), .A(n8119), .B(n8118), .ZN(P1_U3259) );
  NAND2_X1 U9772 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  XOR2_X1 U9773 ( .A(n8124), .B(n8123), .Z(n9060) );
  OAI211_X1 U9774 ( .C1(n8128), .C2(n8127), .A(n8126), .B(n8125), .ZN(n8129)
         );
  OAI21_X1 U9775 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8135) );
  OAI22_X1 U9776 ( .A1(n8132), .A2(n8793), .B1(n8455), .B2(n8795), .ZN(n8134)
         );
  NOR2_X1 U9777 ( .A1(n9060), .A2(n8890), .ZN(n8133) );
  AOI211_X1 U9778 ( .C1(n8902), .C2(n8135), .A(n8134), .B(n8133), .ZN(n9059)
         );
  MUX2_X1 U9779 ( .A(n8136), .B(n9059), .S(n8945), .Z(n8145) );
  INV_X1 U9780 ( .A(n8137), .ZN(n8140) );
  INV_X1 U9781 ( .A(n8138), .ZN(n8139) );
  AOI21_X1 U9782 ( .B1(n9056), .B2(n8140), .A(n8139), .ZN(n9057) );
  OAI22_X1 U9783 ( .A1(n8920), .A2(n8142), .B1(n8877), .B2(n8141), .ZN(n8143)
         );
  AOI21_X1 U9784 ( .B1(n9057), .B2(n8944), .A(n8143), .ZN(n8144) );
  OAI211_X1 U9785 ( .C1(n9060), .C2(n8898), .A(n8145), .B(n8144), .ZN(P2_U3286) );
  OAI21_X1 U9786 ( .B1(n8150), .B2(n4470), .A(n8146), .ZN(n8157) );
  INV_X1 U9787 ( .A(n8153), .ZN(n8600) );
  NAND2_X1 U9788 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND2_X1 U9789 ( .A1(n8182), .A2(n8152), .ZN(n9045) );
  NOR2_X1 U9790 ( .A1(n9045), .A2(n8890), .ZN(n8156) );
  OR2_X1 U9791 ( .A1(n8153), .A2(n8793), .ZN(n8155) );
  OR2_X1 U9792 ( .A1(n8335), .A2(n8795), .ZN(n8154) );
  NAND2_X1 U9793 ( .A1(n8155), .A2(n8154), .ZN(n8521) );
  AOI211_X1 U9794 ( .C1(n8157), .C2(n8902), .A(n8156), .B(n8521), .ZN(n9044)
         );
  INV_X1 U9795 ( .A(n9045), .ZN(n8163) );
  INV_X1 U9796 ( .A(n8898), .ZN(n8929) );
  INV_X1 U9797 ( .A(n8180), .ZN(n9040) );
  NOR2_X1 U9798 ( .A1(n8158), .A2(n9040), .ZN(n8159) );
  OR2_X1 U9799 ( .A1(n8175), .A2(n8159), .ZN(n9041) );
  AOI22_X1 U9800 ( .A1(n8924), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8525), .B2(
        n8942), .ZN(n8161) );
  NAND2_X1 U9801 ( .A1(n8939), .A2(n8180), .ZN(n8160) );
  OAI211_X1 U9802 ( .C1(n9041), .C2(n8932), .A(n8161), .B(n8160), .ZN(n8162)
         );
  AOI21_X1 U9803 ( .B1(n8163), .B2(n8929), .A(n8162), .ZN(n8164) );
  OAI21_X1 U9804 ( .B1(n9044), .B2(n8924), .A(n8164), .ZN(P2_U3283) );
  INV_X1 U9805 ( .A(n8165), .ZN(n8169) );
  OAI222_X1 U9806 ( .A1(n10182), .A2(n8167), .B1(n10186), .B2(n8169), .C1(
        n8166), .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9807 ( .A1(n9099), .A2(n8170), .B1(n9101), .B2(n8169), .C1(n4369), 
        .C2(n8168), .ZN(P2_U3333) );
  OAI211_X1 U9808 ( .C1(n4485), .C2(n8172), .A(n8171), .B(n8902), .ZN(n8174)
         );
  INV_X1 U9809 ( .A(n8481), .ZN(n8887) );
  AOI22_X1 U9810 ( .A1(n8908), .A2(n8887), .B1(n8599), .B2(n8907), .ZN(n8173)
         );
  INV_X1 U9811 ( .A(n8175), .ZN(n8177) );
  INV_X1 U9812 ( .A(n9035), .ZN(n8179) );
  INV_X1 U9813 ( .A(n8916), .ZN(n8176) );
  AOI21_X1 U9814 ( .B1(n9035), .B2(n8177), .A(n8176), .ZN(n9036) );
  AOI22_X1 U9815 ( .A1(n8924), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8395), .B2(
        n8942), .ZN(n8178) );
  OAI21_X1 U9816 ( .B1(n8179), .B2(n8920), .A(n8178), .ZN(n8184) );
  NAND2_X1 U9817 ( .A1(n8180), .A2(n8599), .ZN(n8181) );
  XNOR2_X1 U9818 ( .A(n8332), .B(n8333), .ZN(n9039) );
  NOR2_X1 U9819 ( .A1(n9039), .A2(n8860), .ZN(n8183) );
  AOI211_X1 U9820 ( .C1(n9036), .C2(n8944), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI21_X1 U9821 ( .B1(n9038), .B2(n8924), .A(n8185), .ZN(P2_U3282) );
  INV_X1 U9822 ( .A(n9342), .ZN(n8380) );
  OAI222_X1 U9823 ( .A1(n10186), .A2(n8380), .B1(n8186), .B2(P1_U3084), .C1(
        n9343), .C2(n10182), .ZN(P1_U3324) );
  INV_X1 U9824 ( .A(n8189), .ZN(n8190) );
  NAND2_X1 U9825 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  NAND2_X1 U9826 ( .A1(n10031), .A2(n9159), .ZN(n8194) );
  NAND2_X1 U9827 ( .A1(n8237), .A2(n9640), .ZN(n8193) );
  NAND2_X1 U9828 ( .A1(n8194), .A2(n8193), .ZN(n8195) );
  XNOR2_X1 U9829 ( .A(n8195), .B(n8295), .ZN(n9300) );
  NAND2_X1 U9830 ( .A1(n10031), .A2(n8237), .ZN(n8198) );
  OR2_X1 U9831 ( .A1(n8297), .A2(n8196), .ZN(n8197) );
  AND2_X1 U9832 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  AND2_X1 U9833 ( .A1(n9300), .A2(n8199), .ZN(n8201) );
  INV_X1 U9834 ( .A(n9300), .ZN(n8200) );
  INV_X1 U9835 ( .A(n8199), .ZN(n9299) );
  NAND2_X1 U9836 ( .A1(n8206), .A2(n9159), .ZN(n8203) );
  OR2_X1 U9837 ( .A1(n8217), .A2(n10013), .ZN(n8202) );
  NAND2_X1 U9838 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  XNOR2_X1 U9839 ( .A(n8204), .B(n8295), .ZN(n8207) );
  NOR2_X1 U9840 ( .A1(n8297), .A2(n10013), .ZN(n8205) );
  AOI21_X1 U9841 ( .B1(n8206), .B2(n8237), .A(n8205), .ZN(n8208) );
  NAND2_X1 U9842 ( .A1(n8207), .A2(n8208), .ZN(n9199) );
  INV_X1 U9843 ( .A(n8207), .ZN(n8210) );
  INV_X1 U9844 ( .A(n8208), .ZN(n8209) );
  NAND2_X1 U9845 ( .A1(n8210), .A2(n8209), .ZN(n9200) );
  NAND2_X1 U9846 ( .A1(n8211), .A2(n9200), .ZN(n9279) );
  NAND2_X1 U9847 ( .A1(n10141), .A2(n9159), .ZN(n8213) );
  NAND2_X1 U9848 ( .A1(n8237), .A2(n9638), .ZN(n8212) );
  NAND2_X1 U9849 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  XNOR2_X1 U9850 ( .A(n8214), .B(n9157), .ZN(n9276) );
  NAND2_X1 U9851 ( .A1(n10141), .A2(n8237), .ZN(n8216) );
  OR2_X1 U9852 ( .A1(n8297), .A2(n9996), .ZN(n8215) );
  NAND2_X1 U9853 ( .A1(n8216), .A2(n8215), .ZN(n9277) );
  NAND2_X1 U9854 ( .A1(n10119), .A2(n9159), .ZN(n8219) );
  OR2_X1 U9855 ( .A1(n9962), .A2(n8217), .ZN(n8218) );
  NAND2_X1 U9856 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  XNOR2_X1 U9857 ( .A(n8220), .B(n9157), .ZN(n8245) );
  NOR2_X1 U9858 ( .A1(n9962), .A2(n8297), .ZN(n8221) );
  AOI21_X1 U9859 ( .B1(n10119), .B2(n8237), .A(n8221), .ZN(n8247) );
  XNOR2_X1 U9860 ( .A(n8245), .B(n8247), .ZN(n9235) );
  NAND2_X1 U9861 ( .A1(n10128), .A2(n9159), .ZN(n8223) );
  NAND2_X1 U9862 ( .A1(n4378), .A2(n9636), .ZN(n8222) );
  NAND2_X1 U9863 ( .A1(n8223), .A2(n8222), .ZN(n8224) );
  XNOR2_X1 U9864 ( .A(n8224), .B(n8295), .ZN(n9242) );
  NOR2_X1 U9865 ( .A1(n8297), .A2(n9997), .ZN(n8225) );
  AOI21_X1 U9866 ( .B1(n10128), .B2(n4378), .A(n8225), .ZN(n9237) );
  NAND2_X1 U9867 ( .A1(n10125), .A2(n9159), .ZN(n8227) );
  NAND2_X1 U9868 ( .A1(n9937), .A2(n4378), .ZN(n8226) );
  NAND2_X1 U9869 ( .A1(n8227), .A2(n8226), .ZN(n8228) );
  XNOR2_X1 U9870 ( .A(n8228), .B(n9157), .ZN(n8231) );
  NAND2_X1 U9871 ( .A1(n10125), .A2(n8237), .ZN(n8230) );
  NAND2_X1 U9872 ( .A1(n9937), .A2(n7733), .ZN(n8229) );
  NAND2_X1 U9873 ( .A1(n8230), .A2(n8229), .ZN(n8232) );
  NAND2_X1 U9874 ( .A1(n8231), .A2(n8232), .ZN(n9225) );
  OAI21_X1 U9875 ( .B1(n9242), .B2(n9237), .A(n9225), .ZN(n8235) );
  INV_X1 U9876 ( .A(n8231), .ZN(n8234) );
  INV_X1 U9877 ( .A(n8232), .ZN(n8233) );
  NAND2_X1 U9878 ( .A1(n8235), .A2(n9238), .ZN(n8236) );
  NAND2_X1 U9879 ( .A1(n10136), .A2(n9159), .ZN(n8239) );
  NAND2_X1 U9880 ( .A1(n4378), .A2(n9637), .ZN(n8238) );
  NAND2_X1 U9881 ( .A1(n8239), .A2(n8238), .ZN(n8240) );
  XNOR2_X1 U9882 ( .A(n8240), .B(n9157), .ZN(n9220) );
  NAND2_X1 U9883 ( .A1(n10136), .A2(n4378), .ZN(n8242) );
  OR2_X1 U9884 ( .A1(n8297), .A2(n10015), .ZN(n8241) );
  NAND2_X1 U9885 ( .A1(n8242), .A2(n8241), .ZN(n9224) );
  NAND2_X1 U9886 ( .A1(n4373), .A2(n4431), .ZN(n8250) );
  INV_X1 U9887 ( .A(n9220), .ZN(n8243) );
  INV_X1 U9888 ( .A(n9224), .ZN(n9219) );
  AOI22_X1 U9889 ( .A1(n9242), .A2(n9237), .B1(n8243), .B2(n9219), .ZN(n8244)
         );
  NAND2_X1 U9890 ( .A1(n9238), .A2(n8244), .ZN(n8248) );
  INV_X1 U9891 ( .A(n8245), .ZN(n8246) );
  AOI22_X1 U9892 ( .A1(n4373), .A2(n8248), .B1(n8247), .B2(n8246), .ZN(n8249)
         );
  NAND2_X1 U9893 ( .A1(n10108), .A2(n9159), .ZN(n8252) );
  NAND2_X1 U9894 ( .A1(n9925), .A2(n8237), .ZN(n8251) );
  NAND2_X1 U9895 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  XNOR2_X1 U9896 ( .A(n8253), .B(n9157), .ZN(n8262) );
  NAND2_X1 U9897 ( .A1(n10108), .A2(n8237), .ZN(n8255) );
  NAND2_X1 U9898 ( .A1(n9925), .A2(n7733), .ZN(n8254) );
  NAND2_X1 U9899 ( .A1(n8255), .A2(n8254), .ZN(n8263) );
  NAND2_X1 U9900 ( .A1(n8262), .A2(n8263), .ZN(n9147) );
  INV_X1 U9901 ( .A(n9147), .ZN(n8261) );
  NAND2_X1 U9902 ( .A1(n10113), .A2(n9159), .ZN(n8257) );
  INV_X1 U9903 ( .A(n9918), .ZN(n9939) );
  NAND2_X1 U9904 ( .A1(n9939), .A2(n8237), .ZN(n8256) );
  NAND2_X1 U9905 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  XNOR2_X1 U9906 ( .A(n8258), .B(n8295), .ZN(n9143) );
  NOR2_X1 U9907 ( .A1(n9918), .A2(n8297), .ZN(n8259) );
  AOI21_X1 U9908 ( .B1(n10113), .B2(n8237), .A(n8259), .ZN(n9317) );
  NOR2_X1 U9909 ( .A1(n9143), .A2(n9317), .ZN(n8260) );
  NAND3_X1 U9910 ( .A1(n9147), .A2(n9143), .A3(n9317), .ZN(n8266) );
  INV_X1 U9911 ( .A(n8262), .ZN(n8265) );
  INV_X1 U9912 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U9913 ( .A1(n8265), .A2(n8264), .ZN(n9146) );
  AND2_X1 U9914 ( .A1(n8266), .A2(n9146), .ZN(n8267) );
  NAND2_X1 U9915 ( .A1(n10103), .A2(n9159), .ZN(n8270) );
  OR2_X1 U9916 ( .A1(n9917), .A2(n8217), .ZN(n8269) );
  NAND2_X1 U9917 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  XNOR2_X1 U9918 ( .A(n8271), .B(n9157), .ZN(n8274) );
  NAND2_X1 U9919 ( .A1(n10103), .A2(n8237), .ZN(n8273) );
  OR2_X1 U9920 ( .A1(n9917), .A2(n8297), .ZN(n8272) );
  NAND2_X1 U9921 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  NAND2_X1 U9922 ( .A1(n8274), .A2(n8275), .ZN(n9267) );
  INV_X1 U9923 ( .A(n8274), .ZN(n8277) );
  INV_X1 U9924 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U9925 ( .A1(n8277), .A2(n8276), .ZN(n9269) );
  OAI22_X1 U9926 ( .A1(n9876), .A2(n7022), .B1(n9866), .B2(n8217), .ZN(n8278)
         );
  XNOR2_X1 U9927 ( .A(n8278), .B(n8295), .ZN(n8283) );
  OR2_X1 U9928 ( .A1(n9876), .A2(n8217), .ZN(n8280) );
  NAND2_X1 U9929 ( .A1(n4839), .A2(n7733), .ZN(n8279) );
  NAND2_X1 U9930 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  XNOR2_X1 U9931 ( .A(n8283), .B(n8281), .ZN(n9192) );
  INV_X1 U9932 ( .A(n8281), .ZN(n8282) );
  NAND2_X1 U9933 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  NAND2_X1 U9934 ( .A1(n9190), .A2(n8284), .ZN(n8289) );
  NOR2_X1 U9935 ( .A1(n9886), .A2(n8297), .ZN(n8285) );
  AOI21_X1 U9936 ( .B1(n10092), .B2(n8237), .A(n8285), .ZN(n8290) );
  NAND2_X1 U9937 ( .A1(n10092), .A2(n9159), .ZN(n8287) );
  INV_X1 U9938 ( .A(n9886), .ZN(n9634) );
  NAND2_X1 U9939 ( .A1(n9634), .A2(n8237), .ZN(n8286) );
  NAND2_X1 U9940 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  XNOR2_X1 U9941 ( .A(n8288), .B(n9157), .ZN(n9288) );
  NAND2_X1 U9942 ( .A1(n10089), .A2(n9159), .ZN(n8294) );
  NAND2_X1 U9943 ( .A1(n9825), .A2(n8237), .ZN(n8293) );
  NAND2_X1 U9944 ( .A1(n8294), .A2(n8293), .ZN(n8296) );
  XNOR2_X1 U9945 ( .A(n8296), .B(n8295), .ZN(n8298) );
  INV_X1 U9946 ( .A(n10089), .ZN(n9419) );
  OAI22_X1 U9947 ( .A1(n9419), .A2(n8217), .B1(n9867), .B2(n8297), .ZN(n9135)
         );
  NAND3_X1 U9948 ( .A1(n9287), .A2(n8298), .A3(n9289), .ZN(n9132) );
  OAI22_X1 U9949 ( .A1(n9833), .A2(n8217), .B1(n9852), .B2(n8297), .ZN(n8303)
         );
  NAND2_X1 U9950 ( .A1(n9836), .A2(n9159), .ZN(n8300) );
  NAND2_X1 U9951 ( .A1(n9633), .A2(n8237), .ZN(n8299) );
  NAND2_X1 U9952 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  XNOR2_X1 U9953 ( .A(n8301), .B(n9157), .ZN(n8302) );
  XOR2_X1 U9954 ( .A(n8303), .B(n8302), .Z(n9256) );
  INV_X1 U9955 ( .A(n8302), .ZN(n8305) );
  INV_X1 U9956 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U9957 ( .A1(n10079), .A2(n9159), .ZN(n8307) );
  NAND2_X1 U9958 ( .A1(n9824), .A2(n8237), .ZN(n8306) );
  NAND2_X1 U9959 ( .A1(n8307), .A2(n8306), .ZN(n8308) );
  XNOR2_X1 U9960 ( .A(n8308), .B(n9157), .ZN(n8310) );
  OAI22_X1 U9961 ( .A1(n9819), .A2(n8217), .B1(n9799), .B2(n8297), .ZN(n8309)
         );
  XNOR2_X1 U9962 ( .A(n8310), .B(n8309), .ZN(n9211) );
  NOR2_X1 U9963 ( .A1(n9215), .A2(n8297), .ZN(n8311) );
  AOI21_X1 U9964 ( .B1(n10072), .B2(n8237), .A(n8311), .ZN(n9104) );
  NAND2_X1 U9965 ( .A1(n10072), .A2(n9159), .ZN(n8313) );
  NAND2_X1 U9966 ( .A1(n6361), .A2(n8237), .ZN(n8312) );
  NAND2_X1 U9967 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  XNOR2_X1 U9968 ( .A(n8314), .B(n9157), .ZN(n9106) );
  XOR2_X1 U9969 ( .A(n9104), .B(n9106), .Z(n8315) );
  OAI22_X1 U9970 ( .A1(n9795), .A2(n9336), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8316), .ZN(n8317) );
  AOI21_X1 U9971 ( .B1(n9824), .B2(n9322), .A(n8317), .ZN(n8318) );
  OAI21_X1 U9972 ( .B1(n9800), .B2(n9320), .A(n8318), .ZN(n8319) );
  INV_X1 U9973 ( .A(n8319), .ZN(n8320) );
  INV_X1 U9974 ( .A(n8323), .ZN(P1_U3238) );
  XNOR2_X1 U9975 ( .A(n8324), .B(n8657), .ZN(n8325) );
  OAI21_X1 U9976 ( .B1(n9097), .B2(n8326), .A(n8908), .ZN(n8647) );
  NAND2_X1 U9977 ( .A1(n8334), .A2(n8333), .ZN(n8337) );
  INV_X1 U9978 ( .A(n8335), .ZN(n8906) );
  OR2_X1 U9979 ( .A1(n9035), .A2(n8906), .ZN(n8336) );
  NAND2_X1 U9980 ( .A1(n8337), .A2(n8336), .ZN(n8912) );
  OR2_X1 U9981 ( .A1(n9030), .A2(n8887), .ZN(n8338) );
  NAND2_X1 U9982 ( .A1(n8913), .A2(n8338), .ZN(n8884) );
  INV_X1 U9983 ( .A(n8884), .ZN(n8340) );
  INV_X1 U9984 ( .A(n4435), .ZN(n8339) );
  INV_X1 U9985 ( .A(n8487), .ZN(n8909) );
  NAND2_X1 U9986 ( .A1(n9024), .A2(n8909), .ZN(n8341) );
  NAND2_X1 U9987 ( .A1(n9014), .A2(n8598), .ZN(n8342) );
  NAND2_X1 U9988 ( .A1(n8858), .A2(n8342), .ZN(n8344) );
  OR2_X1 U9989 ( .A1(n9014), .A2(n8598), .ZN(n8343) );
  NAND2_X1 U9990 ( .A1(n8344), .A2(n8343), .ZN(n8832) );
  NAND2_X1 U9991 ( .A1(n8837), .A2(n8848), .ZN(n8345) );
  NAND2_X1 U9992 ( .A1(n8832), .A2(n8345), .ZN(n8347) );
  OR2_X1 U9993 ( .A1(n8837), .A2(n8848), .ZN(n8346) );
  NAND2_X1 U9994 ( .A1(n8347), .A2(n8346), .ZN(n8808) );
  NAND2_X1 U9995 ( .A1(n9004), .A2(n8597), .ZN(n8348) );
  INV_X1 U9996 ( .A(n8536), .ZN(n8773) );
  NAND2_X1 U9997 ( .A1(n9000), .A2(n8773), .ZN(n8349) );
  INV_X1 U9998 ( .A(n8794), .ZN(n8758) );
  OR2_X1 U9999 ( .A1(n8982), .A2(n8757), .ZN(n8351) );
  NAND2_X1 U10000 ( .A1(n8731), .A2(n8730), .ZN(n8729) );
  INV_X1 U10001 ( .A(n8502), .ZN(n8596) );
  NAND2_X1 U10002 ( .A1(n4962), .A2(n8502), .ZN(n8352) );
  INV_X1 U10003 ( .A(n8677), .ZN(n8355) );
  INV_X1 U10004 ( .A(n8669), .ZN(n8363) );
  INV_X1 U10005 ( .A(n9014), .ZN(n8857) );
  NAND2_X1 U10006 ( .A1(n8815), .A2(n5771), .ZN(n8817) );
  INV_X1 U10007 ( .A(n8992), .ZN(n8779) );
  INV_X1 U10008 ( .A(n8987), .ZN(n8764) );
  NOR2_X2 U10009 ( .A1(n4375), .A2(n8732), .ZN(n8718) );
  NAND2_X1 U10010 ( .A1(n8662), .A2(n8671), .ZN(n8358) );
  NAND3_X1 U10011 ( .A1(n8657), .A2(n8656), .A3(n8356), .ZN(n8360) );
  NAND2_X1 U10012 ( .A1(n8662), .A2(n10423), .ZN(n8359) );
  OAI211_X1 U10013 ( .C1(n10400), .C2(n8664), .A(n8360), .B(n8359), .ZN(n8361)
         );
  MUX2_X1 U10014 ( .A(n8365), .B(P2_REG0_REG_29__SCAN_IN), .S(n10431), .Z(
        P2_U3517) );
  INV_X1 U10015 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9402) );
  INV_X1 U10016 ( .A(n9401), .ZN(n8369) );
  OAI222_X1 U10017 ( .A1(n10182), .A2(n9402), .B1(n10186), .B2(n8369), .C1(
        P1_U3084), .C2(n8366), .ZN(P1_U3323) );
  INV_X1 U10018 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8368) );
  INV_X1 U10019 ( .A(n9757), .ZN(n8373) );
  NAND2_X1 U10020 ( .A1(n8370), .A2(n10019), .ZN(n8372) );
  AOI22_X1 U10021 ( .A1(n9166), .A2(n10029), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10021), .ZN(n8371) );
  OAI211_X1 U10022 ( .C1(n8373), .C2(n10024), .A(n8372), .B(n8371), .ZN(n8374)
         );
  AOI21_X1 U10023 ( .B1(n8375), .B2(n10036), .A(n8374), .ZN(n8376) );
  OAI21_X1 U10024 ( .B1(n8377), .B2(n10028), .A(n8376), .ZN(P1_U3263) );
  OAI222_X1 U10025 ( .A1(n8381), .A2(P2_U3152), .B1(n9101), .B2(n8380), .C1(
        n8379), .C2(n8378), .ZN(P2_U3329) );
  XNOR2_X1 U10026 ( .A(n8383), .B(n4929), .ZN(n8384) );
  NAND2_X1 U10027 ( .A1(n8384), .A2(n8583), .ZN(n8389) );
  OAI22_X1 U10028 ( .A1(n8698), .A2(n8565), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8385), .ZN(n8387) );
  NOR2_X1 U10029 ( .A1(n8699), .A2(n8537), .ZN(n8386) );
  AOI211_X1 U10030 ( .C1(n8464), .C2(n8690), .A(n8387), .B(n8386), .ZN(n8388)
         );
  OAI211_X1 U10031 ( .C1(n8692), .C2(n8570), .A(n8389), .B(n8388), .ZN(
        P2_U3216) );
  INV_X1 U10032 ( .A(n8518), .ZN(n8392) );
  NOR3_X1 U10033 ( .A1(n8390), .A2(n8458), .A3(n8559), .ZN(n8391) );
  AOI21_X1 U10034 ( .B1(n8392), .B2(n8583), .A(n8391), .ZN(n8403) );
  NOR2_X1 U10035 ( .A1(n8393), .A2(n8579), .ZN(n8400) );
  AND2_X1 U10036 ( .A1(n8590), .A2(n9035), .ZN(n8399) );
  OAI22_X1 U10037 ( .A1(n8537), .A2(n8481), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8394), .ZN(n8398) );
  INV_X1 U10038 ( .A(n8395), .ZN(n8396) );
  OAI22_X1 U10039 ( .A1(n8458), .A2(n8565), .B1(n8564), .B2(n8396), .ZN(n8397)
         );
  NOR4_X1 U10040 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n8401)
         );
  OAI21_X1 U10041 ( .B1(n8403), .B2(n8402), .A(n8401), .ZN(P2_U3217) );
  AOI22_X1 U10042 ( .A1(n8405), .A2(n8583), .B1(n8581), .B2(n8774), .ZN(n8411)
         );
  OAI22_X1 U10043 ( .A1(n8499), .A2(n8537), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8406), .ZN(n8409) );
  INV_X1 U10044 ( .A(n8464), .ZN(n8575) );
  INV_X1 U10045 ( .A(n8762), .ZN(n8407) );
  OAI22_X1 U10046 ( .A1(n8575), .A2(n8407), .B1(n8794), .B2(n8565), .ZN(n8408)
         );
  AOI211_X1 U10047 ( .C1(n8987), .C2(n8590), .A(n8409), .B(n8408), .ZN(n8410)
         );
  OAI21_X1 U10048 ( .B1(n8496), .B2(n8411), .A(n8410), .ZN(P2_U3218) );
  NOR3_X1 U10049 ( .A1(n8559), .A2(n8412), .A3(n5754), .ZN(n8417) );
  INV_X1 U10050 ( .A(n8413), .ZN(n8414) );
  AOI21_X1 U10051 ( .B1(n7561), .B2(n8414), .A(n8579), .ZN(n8416) );
  OAI21_X1 U10052 ( .B1(n8417), .B2(n8416), .A(n8415), .ZN(n8421) );
  AOI22_X1 U10053 ( .A1(n8590), .A2(n8927), .B1(n8510), .B2(n8418), .ZN(n8420)
         );
  MUX2_X1 U10054 ( .A(P2_STATE_REG_SCAN_IN), .B(n8564), .S(n8930), .Z(n8419)
         );
  NAND3_X1 U10055 ( .A1(n8421), .A2(n8420), .A3(n8419), .ZN(P2_U3220) );
  OR2_X1 U10056 ( .A1(n8426), .A2(n8423), .ZN(n8491) );
  NOR2_X1 U10057 ( .A1(n8422), .A2(n8491), .ZN(n8555) );
  AND2_X1 U10058 ( .A1(n8425), .A2(n8424), .ZN(n8556) );
  OAI21_X1 U10059 ( .B1(n8555), .B2(n8426), .A(n8556), .ZN(n8561) );
  NAND3_X1 U10060 ( .A1(n8427), .A2(n8581), .A3(n8598), .ZN(n8428) );
  OAI21_X1 U10061 ( .B1(n8561), .B2(n8579), .A(n8428), .ZN(n8431) );
  INV_X1 U10062 ( .A(n8429), .ZN(n8430) );
  NAND2_X1 U10063 ( .A1(n8431), .A2(n8430), .ZN(n8436) );
  AOI22_X1 U10064 ( .A1(n8597), .A2(n8908), .B1(n8598), .B2(n8907), .ZN(n8830)
         );
  OAI22_X1 U10065 ( .A1(n8830), .A2(n8573), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8432), .ZN(n8434) );
  INV_X1 U10066 ( .A(n8837), .ZN(n9011) );
  NOR2_X1 U10067 ( .A1(n9011), .A2(n8570), .ZN(n8433) );
  AOI211_X1 U10068 ( .C1(n8836), .C2(n8588), .A(n8434), .B(n8433), .ZN(n8435)
         );
  OAI211_X1 U10069 ( .C1(n8579), .C2(n8437), .A(n8436), .B(n8435), .ZN(
        P2_U3221) );
  INV_X1 U10070 ( .A(n9000), .ZN(n8449) );
  AOI21_X1 U10071 ( .B1(n8438), .B2(n4941), .A(n8579), .ZN(n8443) );
  NOR3_X1 U10072 ( .A1(n8440), .A2(n8792), .A3(n8559), .ZN(n8442) );
  OAI21_X1 U10073 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8448) );
  NOR2_X1 U10074 ( .A1(n8565), .A2(n8792), .ZN(n8446) );
  OAI22_X1 U10075 ( .A1(n8794), .A2(n8537), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8444), .ZN(n8445) );
  AOI211_X1 U10076 ( .C1(n8464), .C2(n8798), .A(n8446), .B(n8445), .ZN(n8447)
         );
  OAI211_X1 U10077 ( .C1(n8449), .C2(n8570), .A(n8448), .B(n8447), .ZN(
        P2_U3225) );
  NAND2_X1 U10078 ( .A1(n8451), .A2(n8450), .ZN(n8453) );
  XOR2_X1 U10079 ( .A(n8453), .B(n8452), .Z(n8462) );
  OAI22_X1 U10080 ( .A1(n8565), .A2(n8455), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8454), .ZN(n8460) );
  INV_X1 U10081 ( .A(n8456), .ZN(n8457) );
  OAI22_X1 U10082 ( .A1(n8458), .A2(n8537), .B1(n8564), .B2(n8457), .ZN(n8459)
         );
  AOI211_X1 U10083 ( .C1(n9046), .C2(n8590), .A(n8460), .B(n8459), .ZN(n8461)
         );
  OAI21_X1 U10084 ( .B1(n8462), .B2(n8579), .A(n8461), .ZN(P2_U3226) );
  NOR2_X1 U10085 ( .A1(n8499), .A2(n8793), .ZN(n8463) );
  AOI21_X1 U10086 ( .B1(n4532), .B2(n8908), .A(n8463), .ZN(n8727) );
  AOI22_X1 U10087 ( .A1(n8734), .A2(n8464), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        n4369), .ZN(n8465) );
  OAI21_X1 U10088 ( .B1(n8727), .B2(n8573), .A(n8465), .ZN(n8472) );
  NAND3_X1 U10089 ( .A1(n8467), .A2(n8581), .A3(n8596), .ZN(n8468) );
  OAI21_X1 U10090 ( .B1(n8469), .B2(n8579), .A(n8468), .ZN(n8471) );
  XNOR2_X1 U10091 ( .A(n8474), .B(n8473), .ZN(n8584) );
  AOI22_X1 U10092 ( .A1(n8584), .A2(n8582), .B1(n8475), .B2(n8474), .ZN(n8479)
         );
  XNOR2_X1 U10093 ( .A(n8477), .B(n8476), .ZN(n8478) );
  XNOR2_X1 U10094 ( .A(n8479), .B(n8478), .ZN(n8485) );
  OAI22_X1 U10095 ( .A1(n8565), .A2(n8481), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8480), .ZN(n8483) );
  OAI22_X1 U10096 ( .A1(n8566), .A2(n8537), .B1(n8564), .B2(n8894), .ZN(n8482)
         );
  AOI211_X1 U10097 ( .C1(n9024), .C2(n8590), .A(n8483), .B(n8482), .ZN(n8484)
         );
  OAI21_X1 U10098 ( .B1(n8485), .B2(n8579), .A(n8484), .ZN(P2_U3228) );
  INV_X1 U10099 ( .A(n8486), .ZN(n8878) );
  OAI22_X1 U10100 ( .A1(n8488), .A2(n8795), .B1(n8487), .B2(n8793), .ZN(n8871)
         );
  NAND2_X1 U10101 ( .A1(n8510), .A2(n8871), .ZN(n8490) );
  NAND2_X1 U10102 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10345)
         );
  OAI211_X1 U10103 ( .C1(n8564), .C2(n8878), .A(n8490), .B(n10345), .ZN(n8493)
         );
  AOI211_X1 U10104 ( .C1(n8422), .C2(n8491), .A(n8579), .B(n8555), .ZN(n8492)
         );
  AOI211_X1 U10105 ( .C1(n9020), .C2(n8590), .A(n8493), .B(n8492), .ZN(n8494)
         );
  INV_X1 U10106 ( .A(n8494), .ZN(P2_U3230) );
  NOR2_X1 U10107 ( .A1(n8496), .A2(n8495), .ZN(n8498) );
  XNOR2_X1 U10108 ( .A(n8498), .B(n8497), .ZN(n8501) );
  OR2_X1 U10109 ( .A1(n8502), .A2(n8795), .ZN(n8504) );
  NAND2_X1 U10110 ( .A1(n8774), .A2(n8907), .ZN(n8503) );
  NAND2_X1 U10111 ( .A1(n8504), .A2(n8503), .ZN(n8742) );
  OAI22_X1 U10112 ( .A1(n8746), .A2(n8575), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8505), .ZN(n8506) );
  AOI21_X1 U10113 ( .B1(n8742), .B2(n8510), .A(n8506), .ZN(n8507) );
  OAI211_X1 U10114 ( .C1(n8748), .C2(n8570), .A(n8508), .B(n8507), .ZN(
        P2_U3231) );
  OAI22_X1 U10115 ( .A1(n8536), .A2(n8795), .B1(n8509), .B2(n8793), .ZN(n8806)
         );
  AOI22_X1 U10116 ( .A1(n8806), .A2(n8510), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        n4369), .ZN(n8511) );
  OAI21_X1 U10117 ( .B1(n8812), .B2(n8575), .A(n8511), .ZN(n8516) );
  INV_X1 U10118 ( .A(n8438), .ZN(n8512) );
  AOI211_X1 U10119 ( .C1(n8514), .C2(n8513), .A(n8579), .B(n8512), .ZN(n8515)
         );
  AOI211_X1 U10120 ( .C1(n9004), .C2(n8590), .A(n8516), .B(n8515), .ZN(n8517)
         );
  INV_X1 U10121 ( .A(n8517), .ZN(P2_U3235) );
  OAI211_X1 U10122 ( .C1(n8520), .C2(n8519), .A(n8518), .B(n8583), .ZN(n8527)
         );
  INV_X1 U10123 ( .A(n8521), .ZN(n8523) );
  OAI22_X1 U10124 ( .A1(n8573), .A2(n8523), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8522), .ZN(n8524) );
  AOI21_X1 U10125 ( .B1(n8525), .B2(n8588), .A(n8524), .ZN(n8526) );
  OAI211_X1 U10126 ( .C1(n9040), .C2(n8570), .A(n8527), .B(n8526), .ZN(
        P2_U3236) );
  INV_X1 U10127 ( .A(n8528), .ZN(n8529) );
  NAND2_X1 U10128 ( .A1(n8441), .A2(n8529), .ZN(n8531) );
  XNOR2_X1 U10129 ( .A(n8531), .B(n8530), .ZN(n8533) );
  NAND3_X1 U10130 ( .A1(n8533), .A2(n8583), .A3(n8532), .ZN(n8543) );
  INV_X1 U10131 ( .A(n8533), .ZN(n8534) );
  NAND3_X1 U10132 ( .A1(n8534), .A2(n8581), .A3(n8758), .ZN(n8542) );
  OAI22_X1 U10133 ( .A1(n8565), .A2(n8536), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8535), .ZN(n8540) );
  OAI22_X1 U10134 ( .A1(n8538), .A2(n8537), .B1(n8780), .B2(n8575), .ZN(n8539)
         );
  AOI211_X1 U10135 ( .C1(n8992), .C2(n8590), .A(n8540), .B(n8539), .ZN(n8541)
         );
  NAND3_X1 U10136 ( .A1(n8543), .A2(n8542), .A3(n8541), .ZN(P2_U3237) );
  XOR2_X1 U10137 ( .A(n8545), .B(n8544), .Z(n8546) );
  NAND2_X1 U10138 ( .A1(n8546), .A2(n8583), .ZN(n8553) );
  INV_X1 U10139 ( .A(n8547), .ZN(n8549) );
  OAI21_X1 U10140 ( .B1(n8573), .B2(n8549), .A(n8548), .ZN(n8550) );
  AOI21_X1 U10141 ( .B1(n8551), .B2(n8588), .A(n8550), .ZN(n8552) );
  OAI211_X1 U10142 ( .C1(n8554), .C2(n8570), .A(n8553), .B(n8552), .ZN(
        P2_U3238) );
  INV_X1 U10143 ( .A(n8555), .ZN(n8558) );
  INV_X1 U10144 ( .A(n8556), .ZN(n8557) );
  AOI21_X1 U10145 ( .B1(n8558), .B2(n8557), .A(n8579), .ZN(n8563) );
  NOR3_X1 U10146 ( .A1(n8560), .A2(n8566), .A3(n8559), .ZN(n8562) );
  OAI21_X1 U10147 ( .B1(n8563), .B2(n8562), .A(n8561), .ZN(n8569) );
  OAI22_X1 U10148 ( .A1(n8566), .A2(n8565), .B1(n8564), .B2(n8854), .ZN(n8567)
         );
  AOI211_X1 U10149 ( .C1(n8589), .C2(n8848), .A(n8618), .B(n8567), .ZN(n8568)
         );
  OAI211_X1 U10150 ( .C1(n8857), .C2(n8570), .A(n8569), .B(n8568), .ZN(
        P2_U3240) );
  XNOR2_X1 U10151 ( .A(n8571), .B(n8572), .ZN(n8580) );
  AOI22_X1 U10152 ( .A1(n8595), .A2(n8908), .B1(n8907), .B2(n8596), .ZN(n8714)
         );
  NOR2_X1 U10153 ( .A1(n8714), .A2(n8573), .ZN(n8577) );
  OAI22_X1 U10154 ( .A1(n8720), .A2(n8575), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8574), .ZN(n8576) );
  AOI211_X1 U10155 ( .C1(n4375), .C2(n8590), .A(n8577), .B(n8576), .ZN(n8578)
         );
  OAI21_X1 U10156 ( .B1(n8580), .B2(n8579), .A(n8578), .ZN(P2_U3242) );
  NAND2_X1 U10157 ( .A1(n8581), .A2(n8887), .ZN(n8586) );
  NAND2_X1 U10158 ( .A1(n8583), .A2(n8582), .ZN(n8585) );
  MUX2_X1 U10159 ( .A(n8586), .B(n8585), .S(n8584), .Z(n8594) );
  AOI22_X1 U10160 ( .A1(n8587), .A2(n8906), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8593) );
  AOI22_X1 U10161 ( .A1(n8589), .A2(n8909), .B1(n8588), .B2(n8917), .ZN(n8592)
         );
  NAND2_X1 U10162 ( .A1(n9030), .A2(n8590), .ZN(n8591) );
  NAND4_X1 U10163 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(
        P2_U3243) );
  MUX2_X1 U10164 ( .A(n8329), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8610), .Z(
        P2_U3580) );
  MUX2_X1 U10165 ( .A(n8595), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8610), .Z(
        P2_U3579) );
  MUX2_X1 U10166 ( .A(n4532), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8610), .Z(
        P2_U3578) );
  MUX2_X1 U10167 ( .A(n8596), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8610), .Z(
        P2_U3577) );
  MUX2_X1 U10168 ( .A(n8757), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8610), .Z(
        P2_U3576) );
  MUX2_X1 U10169 ( .A(n8774), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8610), .Z(
        P2_U3575) );
  MUX2_X1 U10170 ( .A(n8758), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8610), .Z(
        P2_U3574) );
  MUX2_X1 U10171 ( .A(n8773), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8610), .Z(
        P2_U3573) );
  MUX2_X1 U10172 ( .A(n8597), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8610), .Z(
        P2_U3572) );
  MUX2_X1 U10173 ( .A(n8848), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8610), .Z(
        P2_U3571) );
  MUX2_X1 U10174 ( .A(n8598), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8610), .Z(
        P2_U3570) );
  MUX2_X1 U10175 ( .A(n8888), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8610), .Z(
        P2_U3569) );
  MUX2_X1 U10176 ( .A(n8909), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8610), .Z(
        P2_U3568) );
  MUX2_X1 U10177 ( .A(n8887), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8610), .Z(
        P2_U3567) );
  MUX2_X1 U10178 ( .A(n8906), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8610), .Z(
        P2_U3566) );
  MUX2_X1 U10179 ( .A(n8599), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8610), .Z(
        P2_U3565) );
  MUX2_X1 U10180 ( .A(n8600), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8610), .Z(
        P2_U3564) );
  MUX2_X1 U10181 ( .A(n8601), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8610), .Z(
        P2_U3563) );
  MUX2_X1 U10182 ( .A(n8602), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8610), .Z(
        P2_U3562) );
  MUX2_X1 U10183 ( .A(n8603), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8610), .Z(
        P2_U3561) );
  MUX2_X1 U10184 ( .A(n8604), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8610), .Z(
        P2_U3560) );
  MUX2_X1 U10185 ( .A(n8605), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8610), .Z(
        P2_U3559) );
  MUX2_X1 U10186 ( .A(n8606), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8610), .Z(
        P2_U3558) );
  MUX2_X1 U10187 ( .A(n8607), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8610), .Z(
        P2_U3557) );
  MUX2_X1 U10188 ( .A(n8608), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8610), .Z(
        P2_U3556) );
  MUX2_X1 U10189 ( .A(n8609), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8610), .Z(
        P2_U3555) );
  MUX2_X1 U10190 ( .A(n5753), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8610), .Z(
        P2_U3554) );
  MUX2_X1 U10191 ( .A(n7336), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8610), .Z(
        P2_U3553) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n4973), .S(P2_U3966), .Z(
        P2_U3552) );
  OR2_X1 U10193 ( .A1(n8627), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U10194 ( .A1(n8627), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8611) );
  AND2_X1 U10195 ( .A1(n8632), .A2(n8611), .ZN(n8615) );
  INV_X1 U10196 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8614) );
  INV_X1 U10197 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8613) );
  XNOR2_X1 U10198 ( .A(n10352), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U10199 ( .A1(n10358), .A2(n10357), .ZN(n10356) );
  OAI21_X1 U10200 ( .B1(n8615), .B2(n4413), .A(n8633), .ZN(n8619) );
  INV_X1 U10201 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8616) );
  NOR2_X1 U10202 ( .A1(n8643), .A2(n8616), .ZN(n8617) );
  AOI211_X1 U10203 ( .C1(n10355), .C2(n8619), .A(n8618), .B(n8617), .ZN(n8625)
         );
  MUX2_X1 U10204 ( .A(n8622), .B(P2_REG2_REG_17__SCAN_IN), .S(n10352), .Z(
        n10350) );
  NAND2_X1 U10205 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8623), .ZN(n8630) );
  OAI211_X1 U10206 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n8623), .A(n10349), .B(
        n8630), .ZN(n8624) );
  OAI211_X1 U10207 ( .C1(n8626), .C2(n4695), .A(n8625), .B(n8624), .ZN(
        P2_U3263) );
  NAND2_X1 U10208 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  NAND2_X1 U10209 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  XOR2_X1 U10210 ( .A(n8631), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8638) );
  NAND2_X1 U10211 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  INV_X1 U10212 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8634) );
  XNOR2_X1 U10213 ( .A(n8635), .B(n8634), .ZN(n8639) );
  INV_X1 U10214 ( .A(n8639), .ZN(n8636) );
  AOI22_X1 U10215 ( .A1(n8638), .A2(n10349), .B1(n10355), .B2(n8636), .ZN(
        n8641) );
  NAND2_X1 U10216 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8642) );
  NOR2_X1 U10217 ( .A1(n8647), .A2(n8646), .ZN(n8951) );
  INV_X1 U10218 ( .A(n8951), .ZN(n8956) );
  NOR2_X1 U10219 ( .A1(n8924), .A2(n8956), .ZN(n8653) );
  AOI21_X1 U10220 ( .B1(n8924), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8653), .ZN(
        n8649) );
  NAND2_X1 U10221 ( .A1(n8952), .A2(n8939), .ZN(n8648) );
  OAI211_X1 U10222 ( .C1(n8954), .C2(n8932), .A(n8649), .B(n8648), .ZN(
        P2_U3265) );
  INV_X1 U10223 ( .A(n8652), .ZN(n8958) );
  AOI21_X1 U10224 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(n8955) );
  NAND2_X1 U10225 ( .A1(n8955), .A2(n8944), .ZN(n8655) );
  AOI21_X1 U10226 ( .B1(n8924), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8653), .ZN(
        n8654) );
  OAI211_X1 U10227 ( .C1(n8958), .C2(n8920), .A(n8655), .B(n8654), .ZN(
        P2_U3266) );
  NOR2_X1 U10228 ( .A1(n8669), .A2(n8656), .ZN(n8658) );
  XNOR2_X1 U10229 ( .A(n8658), .B(n8657), .ZN(n8668) );
  OAI22_X1 U10230 ( .A1(n8660), .A2(n8877), .B1(n8659), .B2(n8945), .ZN(n8661)
         );
  AOI21_X1 U10231 ( .B1(n8662), .B2(n8939), .A(n8661), .ZN(n8663) );
  OAI21_X1 U10232 ( .B1(n8664), .B2(n8932), .A(n8663), .ZN(n8665) );
  AOI21_X1 U10233 ( .B1(n8666), .B2(n8945), .A(n8665), .ZN(n8667) );
  OAI21_X1 U10234 ( .B1(n8668), .B2(n8860), .A(n8667), .ZN(P2_U3267) );
  AOI21_X2 U10235 ( .B1(n8670), .B2(n8677), .A(n8669), .ZN(n8963) );
  INV_X1 U10236 ( .A(n8671), .ZN(n8672) );
  AOI21_X1 U10237 ( .B1(n8959), .B2(n8689), .A(n8672), .ZN(n8960) );
  AOI22_X1 U10238 ( .A1(n8673), .A2(n8942), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8924), .ZN(n8674) );
  OAI21_X1 U10239 ( .B1(n8675), .B2(n8920), .A(n8674), .ZN(n8682) );
  NOR2_X1 U10240 ( .A1(n8677), .A2(n8676), .ZN(n8680) );
  INV_X1 U10241 ( .A(n8730), .ZN(n8726) );
  INV_X1 U10242 ( .A(n8706), .ZN(n8710) );
  NAND3_X1 U10243 ( .A1(n8709), .A2(n8694), .A3(n8695), .ZN(n8693) );
  INV_X1 U10244 ( .A(n8678), .ZN(n8679) );
  OAI21_X1 U10245 ( .B1(n8963), .B2(n8860), .A(n8683), .ZN(P2_U3268) );
  OAI21_X1 U10246 ( .B1(n8684), .B2(n8686), .A(n8685), .ZN(n8687) );
  INV_X1 U10247 ( .A(n8687), .ZN(n8968) );
  OR2_X1 U10248 ( .A1(n8692), .A2(n8718), .ZN(n8688) );
  AND2_X1 U10249 ( .A1(n8689), .A2(n8688), .ZN(n8965) );
  AOI22_X1 U10250 ( .A1(n8690), .A2(n8942), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8924), .ZN(n8691) );
  OAI21_X1 U10251 ( .B1(n8692), .B2(n8920), .A(n8691), .ZN(n8703) );
  INV_X1 U10252 ( .A(n8693), .ZN(n8697) );
  AOI21_X1 U10253 ( .B1(n8709), .B2(n8695), .A(n8694), .ZN(n8696) );
  NOR3_X1 U10254 ( .A1(n8697), .A2(n8696), .A3(n8868), .ZN(n8701) );
  OAI22_X1 U10255 ( .A1(n8699), .A2(n8795), .B1(n8698), .B2(n8793), .ZN(n8700)
         );
  NOR2_X1 U10256 ( .A1(n8967), .A2(n8924), .ZN(n8702) );
  OAI21_X1 U10257 ( .B1(n8968), .B2(n8860), .A(n8704), .ZN(P2_U3269) );
  OAI21_X1 U10258 ( .B1(n8707), .B2(n8706), .A(n8705), .ZN(n8708) );
  INV_X1 U10259 ( .A(n8708), .ZN(n8973) );
  INV_X1 U10260 ( .A(n8709), .ZN(n8713) );
  AOI21_X1 U10261 ( .B1(n8724), .B2(n8711), .A(n8710), .ZN(n8712) );
  OAI21_X1 U10262 ( .B1(n8715), .B2(n8868), .A(n8714), .ZN(n8975) );
  NAND2_X1 U10263 ( .A1(n4375), .A2(n8732), .ZN(n8716) );
  NAND2_X1 U10264 ( .A1(n8716), .A2(n10424), .ZN(n8717) );
  NOR2_X1 U10265 ( .A1(n8718), .A2(n8717), .ZN(n8971) );
  NAND2_X1 U10266 ( .A1(n8971), .A2(n8874), .ZN(n8719) );
  OAI21_X1 U10267 ( .B1(n8877), .B2(n8720), .A(n8719), .ZN(n8721) );
  OAI21_X1 U10268 ( .B1(n8975), .B2(n8721), .A(n8945), .ZN(n8723) );
  AOI22_X1 U10269 ( .A1(n4375), .A2(n8939), .B1(n8924), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8722) );
  OAI211_X1 U10270 ( .C1(n8973), .C2(n8860), .A(n8723), .B(n8722), .ZN(
        P2_U3270) );
  OAI211_X1 U10271 ( .C1(n8726), .C2(n8725), .A(n8724), .B(n8902), .ZN(n8728)
         );
  OAI21_X1 U10272 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n8979) );
  INV_X1 U10273 ( .A(n8860), .ZN(n8940) );
  AOI21_X1 U10274 ( .B1(n8749), .B2(n4387), .A(n10400), .ZN(n8733) );
  NAND2_X1 U10275 ( .A1(n8733), .A2(n8732), .ZN(n8977) );
  AOI22_X1 U10276 ( .A1(n8734), .A2(n8942), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8924), .ZN(n8736) );
  NAND2_X1 U10277 ( .A1(n4387), .A2(n8939), .ZN(n8735) );
  OAI211_X1 U10278 ( .C1(n8977), .C2(n8840), .A(n8736), .B(n8735), .ZN(n8737)
         );
  AOI21_X1 U10279 ( .B1(n8979), .B2(n8940), .A(n8737), .ZN(n8738) );
  OAI21_X1 U10280 ( .B1(n8981), .B2(n8924), .A(n8738), .ZN(P2_U3271) );
  XNOR2_X1 U10281 ( .A(n8739), .B(n8740), .ZN(n8986) );
  AOI21_X1 U10282 ( .B1(n8741), .B2(n8740), .A(n8868), .ZN(n8744) );
  AOI21_X1 U10283 ( .B1(n8744), .B2(n8743), .A(n8742), .ZN(n8985) );
  OAI22_X1 U10284 ( .A1(n8746), .A2(n8877), .B1(n8745), .B2(n8945), .ZN(n8747)
         );
  AOI21_X1 U10285 ( .B1(n8982), .B2(n8939), .A(n8747), .ZN(n8752) );
  OR2_X1 U10286 ( .A1(n8760), .A2(n8748), .ZN(n8750) );
  AND2_X1 U10287 ( .A1(n8750), .A2(n8749), .ZN(n8983) );
  NAND2_X1 U10288 ( .A1(n8983), .A2(n8944), .ZN(n8751) );
  OAI211_X1 U10289 ( .C1(n8985), .C2(n8924), .A(n8752), .B(n8751), .ZN(n8753)
         );
  INV_X1 U10290 ( .A(n8753), .ZN(n8754) );
  OAI21_X1 U10291 ( .B1(n8860), .B2(n8986), .A(n8754), .ZN(P2_U3272) );
  OAI21_X1 U10292 ( .B1(n4826), .B2(n8756), .A(n8755), .ZN(n8759) );
  AOI222_X1 U10293 ( .A1(n8902), .A2(n8759), .B1(n8758), .B2(n8907), .C1(n8757), .C2(n8908), .ZN(n8990) );
  INV_X1 U10294 ( .A(n8777), .ZN(n8761) );
  AOI21_X1 U10295 ( .B1(n8987), .B2(n8761), .A(n8760), .ZN(n8988) );
  AOI22_X1 U10296 ( .A1(n8762), .A2(n8942), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n8924), .ZN(n8763) );
  OAI21_X1 U10297 ( .B1(n8764), .B2(n8920), .A(n8763), .ZN(n8768) );
  OAI21_X1 U10298 ( .B1(n4424), .B2(n8766), .A(n8765), .ZN(n8991) );
  NOR2_X1 U10299 ( .A1(n8991), .A2(n8860), .ZN(n8767) );
  AOI211_X1 U10300 ( .C1(n8988), .C2(n8944), .A(n8768), .B(n8767), .ZN(n8769)
         );
  OAI21_X1 U10301 ( .B1(n8990), .B2(n8924), .A(n8769), .ZN(P2_U3273) );
  OAI211_X1 U10302 ( .C1(n8772), .C2(n8771), .A(n8770), .B(n8902), .ZN(n8776)
         );
  AOI22_X1 U10303 ( .A1(n8774), .A2(n8908), .B1(n8907), .B2(n8773), .ZN(n8775)
         );
  INV_X1 U10304 ( .A(n8796), .ZN(n8778) );
  AOI21_X1 U10305 ( .B1(n8992), .B2(n8778), .A(n8777), .ZN(n8993) );
  NOR2_X1 U10306 ( .A1(n8779), .A2(n8920), .ZN(n8783) );
  OAI22_X1 U10307 ( .A1(n8781), .A2(n8945), .B1(n8780), .B2(n8877), .ZN(n8782)
         );
  AOI211_X1 U10308 ( .C1(n8993), .C2(n8944), .A(n8783), .B(n8782), .ZN(n8786)
         );
  XNOR2_X1 U10309 ( .A(n8784), .B(n4988), .ZN(n8996) );
  OR2_X1 U10310 ( .A1(n8996), .A2(n8860), .ZN(n8785) );
  OAI211_X1 U10311 ( .C1(n8995), .C2(n8924), .A(n8786), .B(n8785), .ZN(
        P2_U3274) );
  XNOR2_X1 U10312 ( .A(n8787), .B(n8790), .ZN(n9002) );
  AOI21_X1 U10313 ( .B1(n8790), .B2(n8789), .A(n8788), .ZN(n8791) );
  OAI222_X1 U10314 ( .A1(n8795), .A2(n8794), .B1(n8793), .B2(n8792), .C1(n8868), .C2(n8791), .ZN(n8998) );
  AND2_X1 U10315 ( .A1(n8817), .A2(n9000), .ZN(n8797) );
  OR2_X1 U10316 ( .A1(n8797), .A2(n8796), .ZN(n8997) );
  AOI22_X1 U10317 ( .A1(n8924), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8798), .B2(
        n8942), .ZN(n8800) );
  NAND2_X1 U10318 ( .A1(n9000), .A2(n8939), .ZN(n8799) );
  OAI211_X1 U10319 ( .C1(n8997), .C2(n8932), .A(n8800), .B(n8799), .ZN(n8801)
         );
  AOI21_X1 U10320 ( .B1(n8998), .B2(n8945), .A(n8801), .ZN(n8802) );
  OAI21_X1 U10321 ( .B1(n9002), .B2(n8860), .A(n8802), .ZN(P2_U3275) );
  AOI21_X1 U10322 ( .B1(n8803), .B2(n8804), .A(n8868), .ZN(n8807) );
  AOI21_X1 U10323 ( .B1(n8807), .B2(n8805), .A(n8806), .ZN(n9006) );
  NAND2_X1 U10324 ( .A1(n8809), .A2(n5772), .ZN(n8810) );
  NAND2_X1 U10325 ( .A1(n8811), .A2(n8810), .ZN(n9007) );
  INV_X1 U10326 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8813) );
  OAI22_X1 U10327 ( .A1(n8945), .A2(n8813), .B1(n8812), .B2(n8877), .ZN(n8814)
         );
  AOI21_X1 U10328 ( .B1(n9004), .B2(n8939), .A(n8814), .ZN(n8820) );
  AOI21_X1 U10329 ( .B1(n8834), .B2(n9004), .A(n10400), .ZN(n8816) );
  AND2_X1 U10330 ( .A1(n8817), .A2(n8816), .ZN(n9003) );
  NAND2_X1 U10331 ( .A1(n9003), .A2(n8818), .ZN(n8819) );
  OAI211_X1 U10332 ( .C1(n9007), .C2(n8860), .A(n8820), .B(n8819), .ZN(n8821)
         );
  INV_X1 U10333 ( .A(n8821), .ZN(n8822) );
  OAI21_X1 U10334 ( .B1(n9006), .B2(n8924), .A(n8822), .ZN(P2_U3276) );
  AOI21_X1 U10335 ( .B1(n8844), .B2(n8824), .A(n8823), .ZN(n8826) );
  OR2_X1 U10336 ( .A1(n8826), .A2(n4806), .ZN(n8828) );
  INV_X1 U10337 ( .A(n8833), .ZN(n8827) );
  XNOR2_X1 U10338 ( .A(n8828), .B(n8827), .ZN(n8829) );
  NAND2_X1 U10339 ( .A1(n8829), .A2(n8902), .ZN(n8831) );
  NAND2_X1 U10340 ( .A1(n8831), .A2(n8830), .ZN(n9013) );
  INV_X1 U10341 ( .A(n9013), .ZN(n8843) );
  XNOR2_X1 U10342 ( .A(n8832), .B(n8833), .ZN(n9008) );
  AOI21_X1 U10343 ( .B1(n8851), .B2(n8837), .A(n10400), .ZN(n8835) );
  NAND2_X1 U10344 ( .A1(n8835), .A2(n8834), .ZN(n9009) );
  AOI22_X1 U10345 ( .A1(n8924), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8836), .B2(
        n8942), .ZN(n8839) );
  NAND2_X1 U10346 ( .A1(n8837), .A2(n8939), .ZN(n8838) );
  OAI211_X1 U10347 ( .C1(n9009), .C2(n8840), .A(n8839), .B(n8838), .ZN(n8841)
         );
  AOI21_X1 U10348 ( .B1(n9008), .B2(n8940), .A(n8841), .ZN(n8842) );
  OAI21_X1 U10349 ( .B1(n8843), .B2(n8924), .A(n8842), .ZN(P2_U3277) );
  INV_X1 U10350 ( .A(n8844), .ZN(n8883) );
  NAND2_X1 U10351 ( .A1(n8883), .A2(n4435), .ZN(n8882) );
  NAND2_X1 U10352 ( .A1(n8882), .A2(n8845), .ZN(n8869) );
  NOR2_X1 U10353 ( .A1(n8869), .A2(n8870), .ZN(n8867) );
  NOR2_X1 U10354 ( .A1(n8867), .A2(n8846), .ZN(n8847) );
  XNOR2_X1 U10355 ( .A(n8847), .B(n8859), .ZN(n8849) );
  AOI222_X1 U10356 ( .A1(n8902), .A2(n8849), .B1(n8848), .B2(n8908), .C1(n8888), .C2(n8907), .ZN(n9017) );
  INV_X1 U10357 ( .A(n8850), .ZN(n8853) );
  INV_X1 U10358 ( .A(n8851), .ZN(n8852) );
  AOI21_X1 U10359 ( .B1(n9014), .B2(n8853), .A(n8852), .ZN(n9015) );
  INV_X1 U10360 ( .A(n8854), .ZN(n8855) );
  AOI22_X1 U10361 ( .A1(n8924), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8855), .B2(
        n8942), .ZN(n8856) );
  OAI21_X1 U10362 ( .B1(n8857), .B2(n8920), .A(n8856), .ZN(n8862) );
  XNOR2_X1 U10363 ( .A(n8858), .B(n8859), .ZN(n9018) );
  NOR2_X1 U10364 ( .A1(n9018), .A2(n8860), .ZN(n8861) );
  AOI211_X1 U10365 ( .C1(n9015), .C2(n8944), .A(n8862), .B(n8861), .ZN(n8863)
         );
  OAI21_X1 U10366 ( .B1(n9017), .B2(n8924), .A(n8863), .ZN(P2_U3278) );
  NAND2_X1 U10367 ( .A1(n4466), .A2(n8864), .ZN(n8866) );
  AND2_X1 U10368 ( .A1(n8866), .A2(n8865), .ZN(n9023) );
  AOI211_X1 U10369 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8867), .ZN(n8872)
         );
  NOR2_X1 U10370 ( .A1(n8872), .A2(n8871), .ZN(n9022) );
  INV_X1 U10371 ( .A(n8893), .ZN(n8873) );
  AOI211_X1 U10372 ( .C1(n9020), .C2(n8873), .A(n10400), .B(n8850), .ZN(n9019)
         );
  NAND2_X1 U10373 ( .A1(n9019), .A2(n8874), .ZN(n8875) );
  OAI211_X1 U10374 ( .C1(n9023), .C2(n8890), .A(n9022), .B(n8875), .ZN(n8876)
         );
  NAND2_X1 U10375 ( .A1(n8876), .A2(n8945), .ZN(n8881) );
  OAI22_X1 U10376 ( .A1(n8945), .A2(n8622), .B1(n8878), .B2(n8877), .ZN(n8879)
         );
  AOI21_X1 U10377 ( .B1(n9020), .B2(n8939), .A(n8879), .ZN(n8880) );
  OAI211_X1 U10378 ( .C1(n9023), .C2(n8898), .A(n8881), .B(n8880), .ZN(
        P2_U3279) );
  OAI21_X1 U10379 ( .B1(n4435), .B2(n8883), .A(n8882), .ZN(n8892) );
  NAND2_X1 U10380 ( .A1(n8884), .A2(n4435), .ZN(n8885) );
  NAND2_X1 U10381 ( .A1(n8886), .A2(n8885), .ZN(n9028) );
  AOI22_X1 U10382 ( .A1(n8888), .A2(n8908), .B1(n8907), .B2(n8887), .ZN(n8889)
         );
  OAI21_X1 U10383 ( .B1(n9028), .B2(n8890), .A(n8889), .ZN(n8891) );
  AOI21_X1 U10384 ( .B1(n8892), .B2(n8902), .A(n8891), .ZN(n9027) );
  AOI21_X1 U10385 ( .B1(n9024), .B2(n8915), .A(n8893), .ZN(n9025) );
  INV_X1 U10386 ( .A(n9024), .ZN(n8897) );
  INV_X1 U10387 ( .A(n8894), .ZN(n8895) );
  AOI22_X1 U10388 ( .A1(n8924), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8895), .B2(
        n8942), .ZN(n8896) );
  OAI21_X1 U10389 ( .B1(n8897), .B2(n8920), .A(n8896), .ZN(n8900) );
  NOR2_X1 U10390 ( .A1(n9028), .A2(n8898), .ZN(n8899) );
  AOI211_X1 U10391 ( .C1(n9025), .C2(n8944), .A(n8900), .B(n8899), .ZN(n8901)
         );
  OAI21_X1 U10392 ( .B1(n9027), .B2(n8924), .A(n8901), .ZN(P2_U3280) );
  OAI211_X1 U10393 ( .C1(n8905), .C2(n8904), .A(n8903), .B(n8902), .ZN(n8911)
         );
  AOI22_X1 U10394 ( .A1(n8909), .A2(n8908), .B1(n8907), .B2(n8906), .ZN(n8910)
         );
  OAI21_X1 U10395 ( .B1(n8912), .B2(n8914), .A(n8913), .ZN(n9029) );
  INV_X1 U10396 ( .A(n9030), .ZN(n8921) );
  AOI21_X1 U10397 ( .B1(n9030), .B2(n8916), .A(n4972), .ZN(n9031) );
  NAND2_X1 U10398 ( .A1(n9031), .A2(n8944), .ZN(n8919) );
  AOI22_X1 U10399 ( .A1(n8924), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8917), .B2(
        n8942), .ZN(n8918) );
  OAI211_X1 U10400 ( .C1(n8921), .C2(n8920), .A(n8919), .B(n8918), .ZN(n8922)
         );
  AOI21_X1 U10401 ( .B1(n9029), .B2(n8940), .A(n8922), .ZN(n8923) );
  OAI21_X1 U10402 ( .B1(n9033), .B2(n8924), .A(n8923), .ZN(P2_U3281) );
  MUX2_X1 U10403 ( .A(n8926), .B(n8925), .S(n8924), .Z(n8936) );
  AOI22_X1 U10404 ( .A1(n8929), .A2(n8928), .B1(n8939), .B2(n8927), .ZN(n8935)
         );
  NAND2_X1 U10405 ( .A1(n8942), .A2(n8930), .ZN(n8934) );
  OR2_X1 U10406 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NAND4_X1 U10407 ( .A1(n8936), .A2(n8935), .A3(n8934), .A4(n8933), .ZN(
        P2_U3293) );
  INV_X1 U10408 ( .A(n8937), .ZN(n8941) );
  AOI22_X1 U10409 ( .A1(n8941), .A2(n8940), .B1(n8939), .B2(n8938), .ZN(n8950)
         );
  AOI22_X1 U10410 ( .A1(n8944), .A2(n8943), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8942), .ZN(n8949) );
  MUX2_X1 U10411 ( .A(n8947), .B(n8946), .S(n8945), .Z(n8948) );
  NAND3_X1 U10412 ( .A1(n8950), .A2(n8949), .A3(n8948), .ZN(P2_U3295) );
  AOI21_X1 U10413 ( .B1(n8952), .B2(n10423), .A(n8951), .ZN(n8953) );
  OAI21_X1 U10414 ( .B1(n8954), .B2(n10400), .A(n8953), .ZN(n9066) );
  MUX2_X1 U10415 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9066), .S(n10444), .Z(
        P2_U3551) );
  NAND2_X1 U10416 ( .A1(n8955), .A2(n10424), .ZN(n8957) );
  OAI211_X1 U10417 ( .C1(n8958), .C2(n10398), .A(n8957), .B(n8956), .ZN(n9067)
         );
  MUX2_X1 U10418 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9067), .S(n10444), .Z(
        P2_U3550) );
  AOI22_X1 U10419 ( .A1(n8960), .A2(n10424), .B1(n10423), .B2(n8959), .ZN(
        n8961) );
  OAI211_X1 U10420 ( .C1(n8963), .C2(n10418), .A(n8962), .B(n8961), .ZN(n9068)
         );
  MUX2_X1 U10421 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9068), .S(n10444), .Z(
        P2_U3548) );
  AOI22_X1 U10422 ( .A1(n8965), .A2(n10424), .B1(n10423), .B2(n8964), .ZN(
        n8966) );
  OAI211_X1 U10423 ( .C1(n10418), .C2(n8968), .A(n8967), .B(n8966), .ZN(n9069)
         );
  MUX2_X1 U10424 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9069), .S(n10444), .Z(
        P2_U3547) );
  MUX2_X1 U10425 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9070), .S(n10444), .Z(
        P2_U3546) );
  OAI21_X1 U10426 ( .B1(n4962), .B2(n10398), .A(n8977), .ZN(n8978) );
  AOI21_X1 U10427 ( .B1(n8979), .B2(n8356), .A(n8978), .ZN(n8980) );
  NAND2_X1 U10428 ( .A1(n8981), .A2(n8980), .ZN(n9071) );
  MUX2_X1 U10429 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9071), .S(n10444), .Z(
        P2_U3545) );
  AOI22_X1 U10430 ( .A1(n8983), .A2(n10424), .B1(n10423), .B2(n8982), .ZN(
        n8984) );
  OAI211_X1 U10431 ( .C1(n10418), .C2(n8986), .A(n8985), .B(n8984), .ZN(n9072)
         );
  MUX2_X1 U10432 ( .A(n9072), .B(P2_REG1_REG_24__SCAN_IN), .S(n10441), .Z(
        P2_U3544) );
  AOI22_X1 U10433 ( .A1(n8988), .A2(n10424), .B1(n10423), .B2(n8987), .ZN(
        n8989) );
  OAI211_X1 U10434 ( .C1(n10418), .C2(n8991), .A(n8990), .B(n8989), .ZN(n9073)
         );
  MUX2_X1 U10435 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9073), .S(n10444), .Z(
        P2_U3543) );
  AOI22_X1 U10436 ( .A1(n8993), .A2(n10424), .B1(n10423), .B2(n8992), .ZN(
        n8994) );
  OAI211_X1 U10437 ( .C1(n10418), .C2(n8996), .A(n8995), .B(n8994), .ZN(n9074)
         );
  MUX2_X1 U10438 ( .A(n9074), .B(P2_REG1_REG_22__SCAN_IN), .S(n10441), .Z(
        P2_U3542) );
  NOR2_X1 U10439 ( .A1(n8997), .A2(n10400), .ZN(n8999) );
  AOI211_X1 U10440 ( .C1(n10423), .C2(n9000), .A(n8999), .B(n8998), .ZN(n9001)
         );
  OAI21_X1 U10441 ( .B1(n10418), .B2(n9002), .A(n9001), .ZN(n9075) );
  MUX2_X1 U10442 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9075), .S(n10444), .Z(
        P2_U3541) );
  AOI21_X1 U10443 ( .B1(n10423), .B2(n9004), .A(n9003), .ZN(n9005) );
  OAI211_X1 U10444 ( .C1(n10418), .C2(n9007), .A(n9006), .B(n9005), .ZN(n9076)
         );
  MUX2_X1 U10445 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9076), .S(n10444), .Z(
        P2_U3540) );
  NAND2_X1 U10446 ( .A1(n9008), .A2(n8356), .ZN(n9010) );
  OAI211_X1 U10447 ( .C1(n9011), .C2(n10398), .A(n9010), .B(n9009), .ZN(n9012)
         );
  MUX2_X1 U10448 ( .A(n9077), .B(P2_REG1_REG_19__SCAN_IN), .S(n10441), .Z(
        P2_U3539) );
  AOI22_X1 U10449 ( .A1(n9015), .A2(n10424), .B1(n10423), .B2(n9014), .ZN(
        n9016) );
  OAI211_X1 U10450 ( .C1(n10418), .C2(n9018), .A(n9017), .B(n9016), .ZN(n9078)
         );
  MUX2_X1 U10451 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9078), .S(n10444), .Z(
        P2_U3538) );
  AOI21_X1 U10452 ( .B1(n10423), .B2(n9020), .A(n9019), .ZN(n9021) );
  OAI211_X1 U10453 ( .C1(n10418), .C2(n9023), .A(n9022), .B(n9021), .ZN(n9079)
         );
  MUX2_X1 U10454 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9079), .S(n10444), .Z(
        P2_U3537) );
  AOI22_X1 U10455 ( .A1(n9025), .A2(n10424), .B1(n10423), .B2(n9024), .ZN(
        n9026) );
  OAI211_X1 U10456 ( .C1(n10429), .C2(n9028), .A(n9027), .B(n9026), .ZN(n9080)
         );
  MUX2_X1 U10457 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9080), .S(n10444), .Z(
        P2_U3536) );
  INV_X1 U10458 ( .A(n9029), .ZN(n9034) );
  AOI22_X1 U10459 ( .A1(n9031), .A2(n10424), .B1(n10423), .B2(n9030), .ZN(
        n9032) );
  OAI211_X1 U10460 ( .C1(n10418), .C2(n9034), .A(n9033), .B(n9032), .ZN(n9081)
         );
  MUX2_X1 U10461 ( .A(n9081), .B(P2_REG1_REG_15__SCAN_IN), .S(n10441), .Z(
        P2_U3535) );
  AOI22_X1 U10462 ( .A1(n9036), .A2(n10424), .B1(n10423), .B2(n9035), .ZN(
        n9037) );
  OAI211_X1 U10463 ( .C1(n10418), .C2(n9039), .A(n9038), .B(n9037), .ZN(n9082)
         );
  MUX2_X1 U10464 ( .A(n9082), .B(P2_REG1_REG_14__SCAN_IN), .S(n10441), .Z(
        P2_U3534) );
  OAI22_X1 U10465 ( .A1(n9041), .A2(n10400), .B1(n9040), .B2(n10398), .ZN(
        n9042) );
  INV_X1 U10466 ( .A(n9042), .ZN(n9043) );
  OAI211_X1 U10467 ( .C1(n10429), .C2(n9045), .A(n9044), .B(n9043), .ZN(n9083)
         );
  MUX2_X1 U10468 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9083), .S(n10444), .Z(
        P2_U3533) );
  AOI22_X1 U10469 ( .A1(n9047), .A2(n10424), .B1(n10423), .B2(n9046), .ZN(
        n9048) );
  OAI211_X1 U10470 ( .C1(n10418), .C2(n9050), .A(n9049), .B(n9048), .ZN(n9084)
         );
  MUX2_X1 U10471 ( .A(n9084), .B(P2_REG1_REG_12__SCAN_IN), .S(n10441), .Z(
        P2_U3532) );
  AOI21_X1 U10472 ( .B1(n10423), .B2(n9052), .A(n9051), .ZN(n9053) );
  OAI211_X1 U10473 ( .C1(n10418), .C2(n9055), .A(n9054), .B(n9053), .ZN(n9085)
         );
  MUX2_X1 U10474 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9085), .S(n10444), .Z(
        P2_U3531) );
  AOI22_X1 U10475 ( .A1(n9057), .A2(n10424), .B1(n10423), .B2(n9056), .ZN(
        n9058) );
  OAI211_X1 U10476 ( .C1(n9060), .C2(n10429), .A(n9059), .B(n9058), .ZN(n9086)
         );
  MUX2_X1 U10477 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9086), .S(n10444), .Z(
        P2_U3530) );
  AOI22_X1 U10478 ( .A1(n9062), .A2(n10424), .B1(n10423), .B2(n9061), .ZN(
        n9063) );
  OAI211_X1 U10479 ( .C1(n9065), .C2(n10429), .A(n9064), .B(n9063), .ZN(n9087)
         );
  MUX2_X1 U10480 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9087), .S(n10444), .Z(
        P2_U3529) );
  MUX2_X1 U10481 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9066), .S(n10433), .Z(
        P2_U3519) );
  MUX2_X1 U10482 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9067), .S(n10433), .Z(
        P2_U3518) );
  MUX2_X1 U10483 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9068), .S(n10433), .Z(
        P2_U3516) );
  MUX2_X1 U10484 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9069), .S(n10433), .Z(
        P2_U3515) );
  MUX2_X1 U10485 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9070), .S(n10433), .Z(
        P2_U3514) );
  MUX2_X1 U10486 ( .A(n9071), .B(P2_REG0_REG_25__SCAN_IN), .S(n10431), .Z(
        P2_U3513) );
  MUX2_X1 U10487 ( .A(n9072), .B(P2_REG0_REG_24__SCAN_IN), .S(n10431), .Z(
        P2_U3512) );
  MUX2_X1 U10488 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9073), .S(n10433), .Z(
        P2_U3511) );
  MUX2_X1 U10489 ( .A(n9074), .B(P2_REG0_REG_22__SCAN_IN), .S(n10431), .Z(
        P2_U3510) );
  MUX2_X1 U10490 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9075), .S(n10433), .Z(
        P2_U3509) );
  MUX2_X1 U10491 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9076), .S(n10433), .Z(
        P2_U3508) );
  MUX2_X1 U10492 ( .A(n9077), .B(P2_REG0_REG_19__SCAN_IN), .S(n10431), .Z(
        P2_U3507) );
  MUX2_X1 U10493 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9078), .S(n10433), .Z(
        P2_U3505) );
  MUX2_X1 U10494 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9079), .S(n10433), .Z(
        P2_U3502) );
  MUX2_X1 U10495 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9080), .S(n10433), .Z(
        P2_U3499) );
  MUX2_X1 U10496 ( .A(n9081), .B(P2_REG0_REG_15__SCAN_IN), .S(n10431), .Z(
        P2_U3496) );
  MUX2_X1 U10497 ( .A(n9082), .B(P2_REG0_REG_14__SCAN_IN), .S(n10431), .Z(
        P2_U3493) );
  MUX2_X1 U10498 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9083), .S(n10433), .Z(
        P2_U3490) );
  MUX2_X1 U10499 ( .A(n9084), .B(P2_REG0_REG_12__SCAN_IN), .S(n10431), .Z(
        P2_U3487) );
  MUX2_X1 U10500 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9085), .S(n10433), .Z(
        P2_U3484) );
  MUX2_X1 U10501 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9086), .S(n10433), .Z(
        P2_U3481) );
  MUX2_X1 U10502 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9087), .S(n10433), .Z(
        P2_U3478) );
  INV_X1 U10503 ( .A(n9408), .ZN(n10178) );
  NOR4_X1 U10504 ( .A1(n5032), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9088), .A4(
        n4369), .ZN(n9089) );
  AOI21_X1 U10505 ( .B1(n9093), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9089), .ZN(
        n9090) );
  OAI21_X1 U10506 ( .B1(n10178), .B2(n9101), .A(n9090), .ZN(P2_U3327) );
  INV_X1 U10507 ( .A(n9091), .ZN(n10181) );
  AOI21_X1 U10508 ( .B1(n9093), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9092), .ZN(
        n9094) );
  OAI21_X1 U10509 ( .B1(n10181), .B2(n9101), .A(n9094), .ZN(P2_U3330) );
  INV_X1 U10510 ( .A(n9095), .ZN(n10185) );
  OAI222_X1 U10511 ( .A1(n9097), .A2(n4369), .B1(n9101), .B2(n10185), .C1(
        n9096), .C2(n9099), .ZN(P2_U3331) );
  INV_X1 U10512 ( .A(n9098), .ZN(n10189) );
  OAI222_X1 U10513 ( .A1(n4369), .A2(n9102), .B1(n9101), .B2(n10189), .C1(
        n9100), .C2(n9099), .ZN(P2_U3332) );
  MUX2_X1 U10514 ( .A(n9103), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10515 ( .A(n9104), .ZN(n9105) );
  NAND2_X1 U10516 ( .A1(n10067), .A2(n9159), .ZN(n9109) );
  OR2_X1 U10517 ( .A1(n9800), .A2(n8217), .ZN(n9108) );
  NAND2_X1 U10518 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  XNOR2_X1 U10519 ( .A(n9110), .B(n9157), .ZN(n9116) );
  INV_X1 U10520 ( .A(n9116), .ZN(n9114) );
  NAND2_X1 U10521 ( .A1(n10067), .A2(n8237), .ZN(n9112) );
  OR2_X1 U10522 ( .A1(n9800), .A2(n7299), .ZN(n9111) );
  NAND2_X1 U10523 ( .A1(n9112), .A2(n9111), .ZN(n9115) );
  INV_X1 U10524 ( .A(n9115), .ZN(n9113) );
  NAND2_X1 U10525 ( .A1(n9114), .A2(n9113), .ZN(n9169) );
  NAND2_X1 U10526 ( .A1(n9116), .A2(n9115), .ZN(n9164) );
  NAND2_X1 U10527 ( .A1(n9169), .A2(n9164), .ZN(n9117) );
  XNOR2_X1 U10528 ( .A(n9165), .B(n9117), .ZN(n9123) );
  OAI22_X1 U10529 ( .A1(n9215), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9118), .ZN(n9119) );
  AOI21_X1 U10530 ( .B1(n9777), .B2(n9305), .A(n9119), .ZN(n9120) );
  OAI21_X1 U10531 ( .B1(n9769), .B2(n9320), .A(n9120), .ZN(n9121) );
  AOI21_X1 U10532 ( .B1(n10067), .B2(n9338), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10533 ( .B1(n9123), .B2(n9340), .A(n9122), .ZN(P1_U3212) );
  XNOR2_X1 U10534 ( .A(n9220), .B(n9219), .ZN(n9125) );
  XNOR2_X1 U10535 ( .A(n9124), .B(n9125), .ZN(n9131) );
  OAI21_X1 U10536 ( .B1(n9332), .B2(n9996), .A(n9126), .ZN(n9127) );
  AOI21_X1 U10537 ( .B1(n9334), .B2(n9636), .A(n9127), .ZN(n9128) );
  OAI21_X1 U10538 ( .B1(n9336), .B2(n10000), .A(n9128), .ZN(n9129) );
  AOI21_X1 U10539 ( .B1(n9338), .B2(n10136), .A(n9129), .ZN(n9130) );
  OAI21_X1 U10540 ( .B1(n9131), .B2(n9340), .A(n9130), .ZN(P1_U3213) );
  INV_X1 U10541 ( .A(n9132), .ZN(n9134) );
  NOR2_X1 U10542 ( .A1(n9134), .A2(n9133), .ZN(n9136) );
  XNOR2_X1 U10543 ( .A(n9136), .B(n9135), .ZN(n9142) );
  NOR2_X1 U10544 ( .A1(n9847), .A2(n9336), .ZN(n9139) );
  OAI22_X1 U10545 ( .A1(n9886), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9137), .ZN(n9138) );
  AOI211_X1 U10546 ( .C1(n9334), .C2(n9633), .A(n9139), .B(n9138), .ZN(n9141)
         );
  NAND2_X1 U10547 ( .A1(n10089), .A2(n9338), .ZN(n9140) );
  OAI211_X1 U10548 ( .C1(n9142), .C2(n9340), .A(n9141), .B(n9140), .ZN(
        P1_U3214) );
  INV_X1 U10549 ( .A(n9317), .ZN(n9145) );
  NAND2_X1 U10550 ( .A1(n9144), .A2(n9143), .ZN(n9315) );
  NOR2_X1 U10551 ( .A1(n9144), .A2(n9143), .ZN(n9314) );
  AOI21_X1 U10552 ( .B1(n9145), .B2(n9315), .A(n9314), .ZN(n9149) );
  NAND2_X1 U10553 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  XNOR2_X1 U10554 ( .A(n9149), .B(n9148), .ZN(n9154) );
  NAND2_X1 U10555 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9743) );
  OAI21_X1 U10556 ( .B1(n9917), .B2(n9320), .A(n9743), .ZN(n9150) );
  AOI21_X1 U10557 ( .B1(n9322), .B2(n9939), .A(n9150), .ZN(n9151) );
  OAI21_X1 U10558 ( .B1(n9336), .B2(n9910), .A(n9151), .ZN(n9152) );
  AOI21_X1 U10559 ( .B1(n10108), .B2(n9338), .A(n9152), .ZN(n9153) );
  OAI21_X1 U10560 ( .B1(n9154), .B2(n9340), .A(n9153), .ZN(P1_U3217) );
  NAND2_X1 U10561 ( .A1(n9757), .A2(n8237), .ZN(n9156) );
  OR2_X1 U10562 ( .A1(n9769), .A2(n8297), .ZN(n9155) );
  NAND2_X1 U10563 ( .A1(n9156), .A2(n9155), .ZN(n9158) );
  XNOR2_X1 U10564 ( .A(n9158), .B(n9157), .ZN(n9162) );
  NAND2_X1 U10565 ( .A1(n9757), .A2(n9159), .ZN(n9160) );
  OAI21_X1 U10566 ( .B1(n9769), .B2(n8217), .A(n9160), .ZN(n9161) );
  XNOR2_X1 U10567 ( .A(n9162), .B(n9161), .ZN(n9170) );
  INV_X1 U10568 ( .A(n9170), .ZN(n9163) );
  NAND2_X1 U10569 ( .A1(n9163), .A2(n9311), .ZN(n9176) );
  INV_X1 U10570 ( .A(n9800), .ZN(n9632) );
  NAND2_X1 U10571 ( .A1(n9632), .A2(n9322), .ZN(n9168) );
  AOI22_X1 U10572 ( .A1(n9166), .A2(n9305), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9167) );
  OAI211_X1 U10573 ( .C1(n10051), .C2(n9320), .A(n9168), .B(n9167), .ZN(n9172)
         );
  NOR3_X1 U10574 ( .A1(n9170), .A2(n9340), .A3(n9169), .ZN(n9171) );
  AOI211_X1 U10575 ( .C1(n9338), .C2(n9757), .A(n9172), .B(n9171), .ZN(n9173)
         );
  OAI211_X1 U10576 ( .C1(n9176), .C2(n9175), .A(n9174), .B(n9173), .ZN(
        P1_U3218) );
  NAND2_X1 U10577 ( .A1(n10299), .A2(n9177), .ZN(n10309) );
  INV_X1 U10578 ( .A(n9178), .ZN(n9180) );
  NAND2_X1 U10579 ( .A1(n9180), .A2(n9179), .ZN(n9182) );
  XNOR2_X1 U10580 ( .A(n9182), .B(n9181), .ZN(n9183) );
  NAND2_X1 U10581 ( .A1(n9183), .A2(n9311), .ZN(n9189) );
  NAND2_X1 U10582 ( .A1(n9305), .A2(n9184), .ZN(n9187) );
  NAND2_X1 U10583 ( .A1(n9334), .A2(n9642), .ZN(n9186) );
  NAND2_X1 U10584 ( .A1(n9322), .A2(n9644), .ZN(n9185) );
  NAND2_X1 U10585 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10237) );
  AND4_X1 U10586 ( .A1(n9187), .A2(n9186), .A3(n9185), .A4(n10237), .ZN(n9188)
         );
  OAI211_X1 U10587 ( .C1(n9264), .C2(n10309), .A(n9189), .B(n9188), .ZN(
        P1_U3219) );
  OAI21_X1 U10588 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9193) );
  NAND2_X1 U10589 ( .A1(n9193), .A2(n9311), .ZN(n9198) );
  NOR2_X1 U10590 ( .A1(n9336), .A2(n9877), .ZN(n9196) );
  OAI22_X1 U10591 ( .A1(n9886), .A2(n9320), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9194), .ZN(n9195) );
  AOI211_X1 U10592 ( .C1(n9322), .C2(n9635), .A(n9196), .B(n9195), .ZN(n9197)
         );
  OAI211_X1 U10593 ( .C1(n9876), .C2(n9298), .A(n9198), .B(n9197), .ZN(
        P1_U3221) );
  NAND2_X1 U10594 ( .A1(n9200), .A2(n9199), .ZN(n9202) );
  XOR2_X1 U10595 ( .A(n9202), .B(n9201), .Z(n9209) );
  NOR2_X1 U10596 ( .A1(n10146), .A2(n9298), .ZN(n9206) );
  NAND2_X1 U10597 ( .A1(n9322), .A2(n9640), .ZN(n9204) );
  OAI211_X1 U10598 ( .C1(n9996), .C2(n9320), .A(n9204), .B(n9203), .ZN(n9205)
         );
  AOI211_X1 U10599 ( .C1(n9207), .C2(n9305), .A(n9206), .B(n9205), .ZN(n9208)
         );
  OAI21_X1 U10600 ( .B1(n9209), .B2(n9340), .A(n9208), .ZN(P1_U3222) );
  XOR2_X1 U10601 ( .A(n9211), .B(n9210), .Z(n9218) );
  INV_X1 U10602 ( .A(n9212), .ZN(n9816) );
  AOI22_X1 U10603 ( .A1(n9816), .A2(n9305), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9214) );
  NAND2_X1 U10604 ( .A1(n9633), .A2(n9322), .ZN(n9213) );
  OAI211_X1 U10605 ( .C1(n9215), .C2(n9320), .A(n9214), .B(n9213), .ZN(n9216)
         );
  AOI21_X1 U10606 ( .B1(n10079), .B2(n9338), .A(n9216), .ZN(n9217) );
  OAI21_X1 U10607 ( .B1(n9218), .B2(n9340), .A(n9217), .ZN(P1_U3223) );
  NOR2_X1 U10608 ( .A1(n9124), .A2(n9220), .ZN(n9222) );
  NOR2_X1 U10609 ( .A1(n9222), .A2(n9219), .ZN(n9248) );
  INV_X1 U10610 ( .A(n9242), .ZN(n9221) );
  NOR3_X1 U10611 ( .A1(n9248), .A2(n9239), .A3(n9221), .ZN(n9328) );
  NOR2_X1 U10612 ( .A1(n9328), .A2(n9237), .ZN(n9227) );
  INV_X1 U10613 ( .A(n9222), .ZN(n9223) );
  OAI21_X1 U10614 ( .B1(n9239), .B2(n9224), .A(n9223), .ZN(n9244) );
  NOR2_X1 U10615 ( .A1(n9244), .A2(n9242), .ZN(n9327) );
  NAND2_X1 U10616 ( .A1(n9238), .A2(n9225), .ZN(n9226) );
  NOR3_X1 U10617 ( .A1(n9227), .A2(n9327), .A3(n9226), .ZN(n9236) );
  OAI21_X1 U10618 ( .B1(n9227), .B2(n9327), .A(n9226), .ZN(n9228) );
  INV_X1 U10619 ( .A(n9228), .ZN(n9229) );
  OAI21_X1 U10620 ( .B1(n9236), .B2(n9229), .A(n9311), .ZN(n9234) );
  OAI21_X1 U10621 ( .B1(n9320), .B2(n9962), .A(n9230), .ZN(n9232) );
  NOR2_X1 U10622 ( .A1(n9336), .A2(n9966), .ZN(n9231) );
  AOI211_X1 U10623 ( .C1(n9322), .C2(n9636), .A(n9232), .B(n9231), .ZN(n9233)
         );
  OAI211_X1 U10624 ( .C1(n9965), .C2(n9298), .A(n9234), .B(n9233), .ZN(
        P1_U3224) );
  INV_X1 U10625 ( .A(n9238), .ZN(n9243) );
  NOR3_X1 U10626 ( .A1(n9236), .A2(n9243), .A3(n9235), .ZN(n9250) );
  INV_X1 U10627 ( .A(n9237), .ZN(n9329) );
  NAND2_X1 U10628 ( .A1(n9238), .A2(n9329), .ZN(n9240) );
  INV_X1 U10629 ( .A(n9240), .ZN(n9247) );
  INV_X1 U10630 ( .A(n9239), .ZN(n9241) );
  OAI21_X1 U10631 ( .B1(n9241), .B2(n9240), .A(n4373), .ZN(n9246) );
  NOR3_X1 U10632 ( .A1(n9244), .A2(n9243), .A3(n9242), .ZN(n9245) );
  AOI211_X1 U10633 ( .C1(n9248), .C2(n9247), .A(n9246), .B(n9245), .ZN(n9249)
         );
  OAI21_X1 U10634 ( .B1(n9250), .B2(n9249), .A(n9311), .ZN(n9255) );
  AOI21_X1 U10635 ( .B1(n9334), .B2(n9939), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10636 ( .B1(n9332), .B2(n9974), .A(n9252), .ZN(n9253) );
  AOI21_X1 U10637 ( .B1(n9945), .B2(n9305), .A(n9253), .ZN(n9254) );
  OAI211_X1 U10638 ( .C1(n9948), .C2(n9298), .A(n9255), .B(n9254), .ZN(
        P1_U3226) );
  NAND2_X1 U10639 ( .A1(n9836), .A2(n10299), .ZN(n10084) );
  XNOR2_X1 U10640 ( .A(n9257), .B(n9256), .ZN(n9258) );
  NAND2_X1 U10641 ( .A1(n9258), .A2(n9311), .ZN(n9263) );
  OAI22_X1 U10642 ( .A1(n9867), .A2(n9332), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9259), .ZN(n9261) );
  NOR2_X1 U10643 ( .A1(n9799), .A2(n9320), .ZN(n9260) );
  AOI211_X1 U10644 ( .C1(n9829), .C2(n9305), .A(n9261), .B(n9260), .ZN(n9262)
         );
  OAI211_X1 U10645 ( .C1(n9264), .C2(n10084), .A(n9263), .B(n9262), .ZN(
        P1_U3227) );
  INV_X1 U10646 ( .A(n9265), .ZN(n9270) );
  AOI21_X1 U10647 ( .B1(n9269), .B2(n9267), .A(n9266), .ZN(n9268) );
  AOI21_X1 U10648 ( .B1(n9270), .B2(n9269), .A(n9268), .ZN(n9275) );
  AOI22_X1 U10649 ( .A1(n4839), .A2(n9334), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9272) );
  NAND2_X1 U10650 ( .A1(n9322), .A2(n9925), .ZN(n9271) );
  OAI211_X1 U10651 ( .C1(n9336), .C2(n9895), .A(n9272), .B(n9271), .ZN(n9273)
         );
  AOI21_X1 U10652 ( .B1(n10103), .B2(n9338), .A(n9273), .ZN(n9274) );
  OAI21_X1 U10653 ( .B1(n9275), .B2(n9340), .A(n9274), .ZN(P1_U3231) );
  XOR2_X1 U10654 ( .A(n9277), .B(n9276), .Z(n9278) );
  XNOR2_X1 U10655 ( .A(n9279), .B(n9278), .ZN(n9285) );
  NOR2_X1 U10656 ( .A1(n9280), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9714) );
  AOI21_X1 U10657 ( .B1(n9322), .B2(n9639), .A(n9714), .ZN(n9282) );
  NAND2_X1 U10658 ( .A1(n9305), .A2(n10020), .ZN(n9281) );
  OAI211_X1 U10659 ( .C1(n10015), .C2(n9320), .A(n9282), .B(n9281), .ZN(n9283)
         );
  AOI21_X1 U10660 ( .B1(n9338), .B2(n10141), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10661 ( .B1(n9285), .B2(n9340), .A(n9284), .ZN(P1_U3232) );
  AOI21_X1 U10662 ( .B1(n9289), .B2(n9286), .A(n9288), .ZN(n9292) );
  INV_X1 U10663 ( .A(n9287), .ZN(n9291) );
  INV_X1 U10664 ( .A(n9288), .ZN(n9290) );
  OAI22_X1 U10665 ( .A1(n9292), .A2(n9291), .B1(n9290), .B2(n9289), .ZN(n9293)
         );
  NAND2_X1 U10666 ( .A1(n9293), .A2(n9311), .ZN(n9297) );
  AOI22_X1 U10667 ( .A1(n9825), .A2(n9334), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9294) );
  OAI21_X1 U10668 ( .B1(n9866), .B2(n9332), .A(n9294), .ZN(n9295) );
  AOI21_X1 U10669 ( .B1(n9858), .B2(n9305), .A(n9295), .ZN(n9296) );
  OAI211_X1 U10670 ( .C1(n9860), .C2(n9298), .A(n9297), .B(n9296), .ZN(
        P1_U3233) );
  XNOR2_X1 U10671 ( .A(n9300), .B(n9299), .ZN(n9301) );
  XNOR2_X1 U10672 ( .A(n9302), .B(n9301), .ZN(n9312) );
  INV_X1 U10673 ( .A(n9303), .ZN(n9304) );
  AOI21_X1 U10674 ( .B1(n9334), .B2(n9639), .A(n9304), .ZN(n9309) );
  NAND2_X1 U10675 ( .A1(n9338), .A2(n10031), .ZN(n9308) );
  NAND2_X1 U10676 ( .A1(n9305), .A2(n10030), .ZN(n9307) );
  NAND2_X1 U10677 ( .A1(n9322), .A2(n9641), .ZN(n9306) );
  NAND4_X1 U10678 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n9310)
         );
  AOI21_X1 U10679 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9313) );
  INV_X1 U10680 ( .A(n9313), .ZN(P1_U3234) );
  INV_X1 U10681 ( .A(n9314), .ZN(n9316) );
  NAND2_X1 U10682 ( .A1(n9316), .A2(n9315), .ZN(n9318) );
  XNOR2_X1 U10683 ( .A(n9318), .B(n9317), .ZN(n9326) );
  OAI21_X1 U10684 ( .B1(n9320), .B2(n9508), .A(n9319), .ZN(n9321) );
  AOI21_X1 U10685 ( .B1(n9322), .B2(n6264), .A(n9321), .ZN(n9323) );
  OAI21_X1 U10686 ( .B1(n9336), .B2(n9930), .A(n9323), .ZN(n9324) );
  AOI21_X1 U10687 ( .B1(n10113), .B2(n9338), .A(n9324), .ZN(n9325) );
  OAI21_X1 U10688 ( .B1(n9326), .B2(n9340), .A(n9325), .ZN(P1_U3236) );
  NOR2_X1 U10689 ( .A1(n9328), .A2(n9327), .ZN(n9330) );
  XNOR2_X1 U10690 ( .A(n9330), .B(n9329), .ZN(n9341) );
  OAI21_X1 U10691 ( .B1(n9332), .B2(n10015), .A(n9331), .ZN(n9333) );
  AOI21_X1 U10692 ( .B1(n9334), .B2(n9937), .A(n9333), .ZN(n9335) );
  OAI21_X1 U10693 ( .B1(n9336), .B2(n9983), .A(n9335), .ZN(n9337) );
  AOI21_X1 U10694 ( .B1(n9338), .B2(n10128), .A(n9337), .ZN(n9339) );
  OAI21_X1 U10695 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(P1_U3239) );
  NAND2_X1 U10696 ( .A1(n9342), .A2(n4620), .ZN(n9345) );
  OR2_X1 U10697 ( .A1(n9409), .A2(n9343), .ZN(n9344) );
  OR2_X1 U10698 ( .A1(n10050), .A2(n10051), .ZN(n9346) );
  NAND2_X1 U10699 ( .A1(n9346), .A2(n9535), .ZN(n9398) );
  AND2_X1 U10700 ( .A1(n9527), .A2(n9524), .ZN(n9392) );
  NAND3_X1 U10701 ( .A1(n9531), .A2(n9392), .A3(n9347), .ZN(n9348) );
  NOR2_X1 U10702 ( .A1(n9398), .A2(n9348), .ZN(n9573) );
  INV_X1 U10703 ( .A(n9573), .ZN(n9406) );
  NAND2_X1 U10704 ( .A1(n9876), .A2(n4839), .ZN(n9427) );
  INV_X1 U10705 ( .A(n9514), .ZN(n9349) );
  NAND2_X1 U10706 ( .A1(n9427), .A2(n9349), .ZN(n9350) );
  AND2_X1 U10707 ( .A1(n9431), .A2(n9350), .ZN(n9353) );
  OAI211_X1 U10708 ( .C1(n9508), .C2(n10108), .A(n9427), .B(n9516), .ZN(n9352)
         );
  INV_X1 U10709 ( .A(n9864), .ZN(n9351) );
  AOI21_X1 U10710 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9357) );
  INV_X1 U10711 ( .A(n9353), .ZN(n9354) );
  OR2_X1 U10712 ( .A1(n9354), .A2(n9900), .ZN(n9552) );
  OR2_X1 U10713 ( .A1(n9552), .A2(n9355), .ZN(n9356) );
  NAND2_X1 U10714 ( .A1(n9357), .A2(n9356), .ZN(n9569) );
  NAND2_X1 U10715 ( .A1(n10136), .A2(n10015), .ZN(n9449) );
  NAND2_X1 U10716 ( .A1(n9449), .A2(n9380), .ZN(n9451) );
  INV_X1 U10717 ( .A(n9451), .ZN(n9359) );
  AND4_X1 U10718 ( .A1(n9459), .A2(n9462), .A3(n9461), .A4(n9454), .ZN(n9358)
         );
  NAND4_X1 U10719 ( .A1(n9433), .A2(n9359), .A3(n9444), .A4(n9358), .ZN(n9360)
         );
  OR3_X1 U10720 ( .A1(n9491), .A2(n4864), .A3(n9360), .ZN(n9568) );
  INV_X1 U10721 ( .A(n9361), .ZN(n9362) );
  OAI211_X1 U10722 ( .C1(n9364), .C2(n4386), .A(n6393), .B(n9362), .ZN(n9365)
         );
  INV_X1 U10723 ( .A(n9365), .ZN(n9367) );
  OAI21_X1 U10724 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9370) );
  NAND3_X1 U10725 ( .A1(n9370), .A2(n9369), .A3(n9558), .ZN(n9372) );
  AND2_X1 U10726 ( .A1(n9555), .A2(n9371), .ZN(n9553) );
  NAND2_X1 U10727 ( .A1(n9372), .A2(n9553), .ZN(n9377) );
  AND2_X1 U10728 ( .A1(n9373), .A2(n9556), .ZN(n9376) );
  AND2_X1 U10729 ( .A1(n9374), .A2(n9456), .ZN(n9563) );
  NAND2_X1 U10730 ( .A1(n9563), .A2(n9561), .ZN(n9375) );
  AOI21_X1 U10731 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9387) );
  OAI21_X1 U10732 ( .B1(n9441), .B2(n4507), .A(n9466), .ZN(n9378) );
  NAND3_X1 U10733 ( .A1(n9444), .A2(n9459), .A3(n9378), .ZN(n9379) );
  NAND2_X1 U10734 ( .A1(n9379), .A2(n9478), .ZN(n9381) );
  AND2_X1 U10735 ( .A1(n9381), .A2(n9380), .ZN(n9383) );
  NAND2_X1 U10736 ( .A1(n9450), .A2(n9382), .ZN(n9480) );
  OAI211_X1 U10737 ( .C1(n9383), .C2(n9480), .A(n9433), .B(n9449), .ZN(n9384)
         );
  NAND2_X1 U10738 ( .A1(n9435), .A2(n9384), .ZN(n9385) );
  NAND2_X1 U10739 ( .A1(n9385), .A2(n9492), .ZN(n9386) );
  OR2_X1 U10740 ( .A1(n9491), .A2(n9386), .ZN(n9566) );
  OAI21_X1 U10741 ( .B1(n9568), .B2(n9387), .A(n9566), .ZN(n9388) );
  INV_X1 U10742 ( .A(n9388), .ZN(n9389) );
  NOR2_X1 U10743 ( .A1(n9552), .A2(n9389), .ZN(n9390) );
  OAI21_X1 U10744 ( .B1(n9569), .B2(n9390), .A(n9551), .ZN(n9391) );
  NAND2_X1 U10745 ( .A1(n9391), .A2(n9572), .ZN(n9405) );
  INV_X1 U10746 ( .A(n9392), .ZN(n9394) );
  AND2_X1 U10747 ( .A1(n9523), .A2(n9393), .ZN(n9418) );
  OAI211_X1 U10748 ( .C1(n9394), .C2(n9418), .A(n9532), .B(n9528), .ZN(n9395)
         );
  NAND2_X1 U10749 ( .A1(n9395), .A2(n9531), .ZN(n9396) );
  AND2_X1 U10750 ( .A1(n9396), .A2(n9764), .ZN(n9397) );
  OR2_X1 U10751 ( .A1(n9398), .A2(n9397), .ZN(n9400) );
  NAND2_X1 U10752 ( .A1(n10050), .A2(n10051), .ZN(n9399) );
  NAND2_X1 U10753 ( .A1(n9401), .A2(n4620), .ZN(n9404) );
  OR2_X1 U10754 ( .A1(n9409), .A2(n9402), .ZN(n9403) );
  NAND2_X1 U10755 ( .A1(n9407), .A2(n9768), .ZN(n9608) );
  OAI211_X1 U10756 ( .C1(n9406), .C2(n9405), .A(n9577), .B(n9608), .ZN(n9415)
         );
  OR2_X1 U10757 ( .A1(n9407), .A2(n9768), .ZN(n9412) );
  NAND2_X1 U10758 ( .A1(n9408), .A2(n4620), .ZN(n9411) );
  OR2_X1 U10759 ( .A1(n9409), .A2(n6778), .ZN(n9410) );
  NAND2_X1 U10760 ( .A1(n10043), .A2(n9749), .ZN(n9537) );
  NAND2_X1 U10761 ( .A1(n9412), .A2(n9537), .ZN(n9609) );
  INV_X1 U10762 ( .A(n9609), .ZN(n9414) );
  INV_X1 U10763 ( .A(n9606), .ZN(n9413) );
  AOI21_X1 U10764 ( .B1(n9415), .B2(n9414), .A(n9413), .ZN(n9620) );
  INV_X1 U10765 ( .A(n9620), .ZN(n9624) );
  OAI21_X1 U10766 ( .B1(n9749), .B2(n9768), .A(n9407), .ZN(n9576) );
  INV_X1 U10767 ( .A(n9576), .ZN(n9538) );
  INV_X1 U10768 ( .A(n10050), .ZN(n10052) );
  INV_X1 U10769 ( .A(n9605), .ZN(n9534) );
  INV_X1 U10770 ( .A(n9827), .ZN(n9823) );
  MUX2_X1 U10771 ( .A(n9825), .B(n10089), .S(n9540), .Z(n9416) );
  INV_X1 U10772 ( .A(n9416), .ZN(n9417) );
  OAI21_X1 U10773 ( .B1(n9425), .B2(n9419), .A(n9418), .ZN(n9421) );
  OAI211_X1 U10774 ( .C1(n9425), .C2(n9867), .A(n9572), .B(n9524), .ZN(n9420)
         );
  INV_X1 U10775 ( .A(n9422), .ZN(n9423) );
  NAND2_X1 U10776 ( .A1(n9823), .A2(n9423), .ZN(n9424) );
  NAND2_X1 U10777 ( .A1(n9425), .A2(n9424), .ZN(n9522) );
  AND2_X1 U10778 ( .A1(n9864), .A2(n9540), .ZN(n9517) );
  INV_X1 U10779 ( .A(n9517), .ZN(n9430) );
  INV_X1 U10780 ( .A(n9540), .ZN(n9530) );
  AND2_X1 U10781 ( .A1(n9426), .A2(n9530), .ZN(n9506) );
  NAND2_X1 U10782 ( .A1(n9864), .A2(n9427), .ZN(n9428) );
  NAND2_X1 U10783 ( .A1(n9506), .A2(n9428), .ZN(n9429) );
  OAI21_X1 U10784 ( .B1(n9431), .B2(n9430), .A(n9429), .ZN(n9432) );
  INV_X1 U10785 ( .A(n9432), .ZN(n9521) );
  NOR2_X1 U10786 ( .A1(n9955), .A2(n4872), .ZN(n9434) );
  MUX2_X1 U10787 ( .A(n9435), .B(n9434), .S(n9530), .Z(n9490) );
  INV_X1 U10788 ( .A(n9439), .ZN(n9560) );
  NAND2_X1 U10789 ( .A1(n4460), .A2(n9441), .ZN(n9448) );
  INV_X1 U10790 ( .A(n9442), .ZN(n9443) );
  NOR2_X1 U10791 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  OR2_X1 U10792 ( .A1(n9451), .A2(n9445), .ZN(n9477) );
  NAND3_X1 U10793 ( .A1(n9459), .A2(n9530), .A3(n9461), .ZN(n9446) );
  NOR2_X1 U10794 ( .A1(n9477), .A2(n9446), .ZN(n9447) );
  NAND2_X1 U10795 ( .A1(n9448), .A2(n9447), .ZN(n9486) );
  INV_X1 U10796 ( .A(n9972), .ZN(n9975) );
  NAND2_X1 U10797 ( .A1(n9480), .A2(n9449), .ZN(n9453) );
  NAND2_X1 U10798 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  MUX2_X1 U10799 ( .A(n9453), .B(n9452), .S(n9540), .Z(n9485) );
  NAND3_X1 U10800 ( .A1(n9455), .A2(n9454), .A3(n9557), .ZN(n9458) );
  NAND3_X1 U10801 ( .A1(n9458), .A2(n9457), .A3(n9456), .ZN(n9465) );
  NAND2_X1 U10802 ( .A1(n9460), .A2(n9459), .ZN(n9474) );
  NAND4_X1 U10803 ( .A1(n9472), .A2(n9540), .A3(n9462), .A4(n9461), .ZN(n9463)
         );
  NOR2_X1 U10804 ( .A1(n9474), .A2(n9463), .ZN(n9464) );
  NAND2_X1 U10805 ( .A1(n9465), .A2(n9464), .ZN(n9483) );
  NOR2_X1 U10806 ( .A1(n9466), .A2(n9540), .ZN(n9467) );
  NOR2_X1 U10807 ( .A1(n9468), .A2(n9467), .ZN(n9476) );
  NAND2_X1 U10808 ( .A1(n9469), .A2(n9540), .ZN(n9470) );
  OAI22_X1 U10809 ( .A1(n9472), .A2(n9530), .B1(n9471), .B2(n9470), .ZN(n9473)
         );
  AOI21_X1 U10810 ( .B1(n9474), .B2(n9540), .A(n9473), .ZN(n9475) );
  OAI21_X1 U10811 ( .B1(n9477), .B2(n9476), .A(n9475), .ZN(n9482) );
  INV_X1 U10812 ( .A(n9478), .ZN(n9479) );
  OAI21_X1 U10813 ( .B1(n9480), .B2(n9479), .A(n9540), .ZN(n9481) );
  NAND3_X1 U10814 ( .A1(n9483), .A2(n9482), .A3(n9481), .ZN(n9484) );
  NAND4_X1 U10815 ( .A1(n9486), .A2(n9975), .A3(n9485), .A4(n9484), .ZN(n9489)
         );
  NOR2_X1 U10816 ( .A1(n9487), .A2(n9540), .ZN(n9488) );
  OR2_X1 U10817 ( .A1(n9492), .A2(n9530), .ZN(n9493) );
  NAND3_X1 U10818 ( .A1(n9496), .A2(n6264), .A3(n10119), .ZN(n9497) );
  AND2_X1 U10819 ( .A1(n9502), .A2(n9508), .ZN(n9500) );
  INV_X1 U10820 ( .A(n9510), .ZN(n9498) );
  NOR2_X1 U10821 ( .A1(n9498), .A2(n10108), .ZN(n9499) );
  MUX2_X1 U10822 ( .A(n9500), .B(n9499), .S(n9540), .Z(n9501) );
  NAND2_X1 U10823 ( .A1(n9511), .A2(n9501), .ZN(n9509) );
  NAND2_X1 U10824 ( .A1(n9509), .A2(n9909), .ZN(n9505) );
  NAND2_X1 U10825 ( .A1(n9511), .A2(n9502), .ZN(n9503) );
  NAND2_X1 U10826 ( .A1(n9503), .A2(n9925), .ZN(n9504) );
  NAND3_X1 U10827 ( .A1(n9505), .A2(n9516), .A3(n9504), .ZN(n9507) );
  NAND4_X1 U10828 ( .A1(n9507), .A2(n9506), .A3(n6414), .A4(n9514), .ZN(n9520)
         );
  NAND2_X1 U10829 ( .A1(n9509), .A2(n9508), .ZN(n9515) );
  NAND2_X1 U10830 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  NAND2_X1 U10831 ( .A1(n9512), .A2(n10108), .ZN(n9513) );
  NAND3_X1 U10832 ( .A1(n9515), .A2(n9514), .A3(n9513), .ZN(n9518) );
  NAND4_X1 U10833 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n6414), .ZN(n9519)
         );
  MUX2_X1 U10834 ( .A(n9524), .B(n9523), .S(n9540), .Z(n9525) );
  MUX2_X1 U10835 ( .A(n9528), .B(n9527), .S(n9540), .Z(n9529) );
  MUX2_X1 U10836 ( .A(n9532), .B(n9531), .S(n9530), .Z(n9533) );
  MUX2_X1 U10837 ( .A(n9764), .B(n9535), .S(n9540), .Z(n9536) );
  NAND2_X1 U10838 ( .A1(n10053), .A2(n9540), .ZN(n9542) );
  OR2_X1 U10839 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  NAND4_X1 U10840 ( .A1(n9606), .A2(n6396), .A3(n9740), .A4(n9547), .ZN(n9622)
         );
  INV_X1 U10841 ( .A(n9548), .ZN(n9549) );
  NAND2_X1 U10842 ( .A1(n9550), .A2(n9740), .ZN(n9619) );
  INV_X1 U10843 ( .A(n9551), .ZN(n9575) );
  INV_X1 U10844 ( .A(n9552), .ZN(n9571) );
  NAND3_X1 U10845 ( .A1(n9554), .A2(n9553), .A3(n9561), .ZN(n9565) );
  INV_X1 U10846 ( .A(n9555), .ZN(n9559) );
  OAI211_X1 U10847 ( .C1(n9559), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9562)
         );
  AOI21_X1 U10848 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9564) );
  AOI21_X1 U10849 ( .B1(n9565), .B2(n9564), .A(n4551), .ZN(n9567) );
  OAI21_X1 U10850 ( .B1(n9568), .B2(n9567), .A(n9566), .ZN(n9570) );
  AOI21_X1 U10851 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9574) );
  OAI211_X1 U10852 ( .C1(n9575), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9578)
         );
  NAND4_X1 U10853 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9606), .ZN(n9580)
         );
  AOI21_X1 U10854 ( .B1(n9580), .B2(n9579), .A(n9611), .ZN(n9613) );
  INV_X1 U10855 ( .A(n9807), .ZN(n9806) );
  INV_X1 U10856 ( .A(n9927), .ZN(n9598) );
  INV_X1 U10857 ( .A(n9955), .ZN(n9959) );
  NAND4_X1 U10858 ( .A1(n9582), .A2(n6074), .A3(n9581), .A4(n7081), .ZN(n9585)
         );
  NOR3_X1 U10859 ( .A1(n9585), .A2(n9584), .A3(n9583), .ZN(n9589) );
  NAND4_X1 U10860 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(n9592)
         );
  NAND2_X1 U10861 ( .A1(n6411), .A2(n9590), .ZN(n9591) );
  NOR2_X1 U10862 ( .A1(n9592), .A2(n9591), .ZN(n9594) );
  NAND4_X1 U10863 ( .A1(n6412), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9596)
         );
  NOR3_X1 U10864 ( .A1(n9972), .A2(n9993), .A3(n9596), .ZN(n9597) );
  NAND4_X1 U10865 ( .A1(n9598), .A2(n9959), .A3(n9943), .A4(n9597), .ZN(n9599)
         );
  NOR3_X1 U10866 ( .A1(n9899), .A2(n9915), .A3(n9599), .ZN(n9600) );
  NAND4_X1 U10867 ( .A1(n9849), .A2(n4417), .A3(n9600), .A4(n6414), .ZN(n9601)
         );
  NOR2_X1 U10868 ( .A1(n9601), .A2(n9827), .ZN(n9602) );
  NAND4_X1 U10869 ( .A1(n9780), .A2(n9603), .A3(n9806), .A4(n9602), .ZN(n9604)
         );
  NOR2_X1 U10870 ( .A1(n9605), .A2(n9604), .ZN(n9607) );
  NAND3_X1 U10871 ( .A1(n9608), .A2(n9607), .A3(n9606), .ZN(n9610) );
  XNOR2_X1 U10872 ( .A(n10050), .B(n10053), .ZN(n10058) );
  INV_X1 U10873 ( .A(n10058), .ZN(n10061) );
  NAND2_X1 U10874 ( .A1(n9612), .A2(n9611), .ZN(n9614) );
  OAI211_X1 U10875 ( .C1(n9613), .C2(n9740), .A(n6396), .B(n9614), .ZN(n9618)
         );
  INV_X1 U10876 ( .A(n9614), .ZN(n9616) );
  NAND3_X1 U10877 ( .A1(n9616), .A2(n6396), .A3(n9615), .ZN(n9617) );
  OAI211_X1 U10878 ( .C1(n9620), .C2(n9619), .A(n9618), .B(n9617), .ZN(n9621)
         );
  INV_X1 U10879 ( .A(n9625), .ZN(n9628) );
  NAND3_X1 U10880 ( .A1(n9626), .A2(n9662), .A3(n9652), .ZN(n9627) );
  OAI211_X1 U10881 ( .C1(n9629), .C2(n9628), .A(n9627), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9630) );
  NAND2_X1 U10882 ( .A1(n9631), .A2(n9630), .ZN(P1_U3240) );
  MUX2_X1 U10883 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10053), .S(P1_U4006), .Z(
        P1_U3584) );
  INV_X1 U10884 ( .A(n9769), .ZN(n9781) );
  MUX2_X1 U10885 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9781), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10886 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9632), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10887 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n6361), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10888 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9824), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10889 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9633), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9825), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9634), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10892 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n4839), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10893 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9635), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9925), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9939), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n6264), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10897 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9937), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10898 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9636), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10899 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9637), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10900 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9638), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10901 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9639), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10902 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9640), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10903 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9641), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10904 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9642), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10905 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9643), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10906 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9644), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10907 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9645), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10908 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9646), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10909 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9647), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10910 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9648), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7075), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6057), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND2_X1 U10913 ( .A1(n9684), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9659) );
  NAND3_X1 U10914 ( .A1(n10235), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9650), .ZN(
        n9658) );
  NAND2_X1 U10915 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9657) );
  NOR2_X1 U10916 ( .A1(n10184), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9651) );
  NOR2_X1 U10917 ( .A1(n9651), .A2(n10180), .ZN(n9665) );
  XNOR2_X1 U10918 ( .A(n9665), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9654) );
  OAI21_X1 U10919 ( .B1(n9652), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6085), .ZN(
        n9653) );
  OR3_X1 U10920 ( .A1(n9655), .A2(n9654), .A3(n9653), .ZN(n9656) );
  NAND4_X1 U10921 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(
        P1_U3241) );
  MUX2_X1 U10922 ( .A(n9661), .B(n9660), .S(n10184), .Z(n9663) );
  NAND2_X1 U10923 ( .A1(n9663), .A2(n9662), .ZN(n9664) );
  OAI211_X1 U10924 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9665), .A(n9664), .B(
        P1_U4006), .ZN(n9693) );
  XNOR2_X1 U10925 ( .A(n9667), .B(n9666), .ZN(n9669) );
  INV_X1 U10926 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9668) );
  OAI22_X1 U10927 ( .A1(n9735), .A2(n9669), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9668), .ZN(n9670) );
  AOI21_X1 U10928 ( .B1(n9684), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n9670), .ZN(
        n9677) );
  NAND2_X1 U10929 ( .A1(n9716), .A2(n9671), .ZN(n9676) );
  OAI211_X1 U10930 ( .C1(n9674), .C2(n9673), .A(n9733), .B(n9672), .ZN(n9675)
         );
  NAND4_X1 U10931 ( .A1(n9693), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(
        P1_U3243) );
  NAND2_X1 U10932 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  AOI21_X1 U10933 ( .B1(n9681), .B2(n9680), .A(n9735), .ZN(n9682) );
  AOI211_X1 U10934 ( .C1(n9684), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9683), .B(
        n9682), .ZN(n9692) );
  NAND2_X1 U10935 ( .A1(n9686), .A2(n9685), .ZN(n9687) );
  AOI21_X1 U10936 ( .B1(n9688), .B2(n9687), .A(n10228), .ZN(n9689) );
  AOI21_X1 U10937 ( .B1(n9716), .B2(n9690), .A(n9689), .ZN(n9691) );
  NAND3_X1 U10938 ( .A1(n9693), .A2(n9692), .A3(n9691), .ZN(P1_U3245) );
  INV_X1 U10939 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10483) );
  NOR2_X1 U10940 ( .A1(n10244), .A2(n10483), .ZN(n9694) );
  AOI211_X1 U10941 ( .C1(n9716), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9705)
         );
  OAI211_X1 U10942 ( .C1(n9698), .C2(n10224), .A(n9733), .B(n9697), .ZN(n9704)
         );
  OAI21_X1 U10943 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9702) );
  NAND2_X1 U10944 ( .A1(n9702), .A2(n10235), .ZN(n9703) );
  NAND3_X1 U10945 ( .A1(n9705), .A2(n9704), .A3(n9703), .ZN(P1_U3250) );
  INV_X1 U10946 ( .A(n9706), .ZN(n9711) );
  NOR3_X1 U10947 ( .A1(n9709), .A2(n9708), .A3(n9707), .ZN(n9710) );
  OAI21_X1 U10948 ( .B1(n9711), .B2(n9710), .A(n10235), .ZN(n9722) );
  NOR2_X1 U10949 ( .A1(n10244), .A2(n9712), .ZN(n9713) );
  AOI211_X1 U10950 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9721)
         );
  OAI211_X1 U10951 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9733), .ZN(n9720)
         );
  NAND3_X1 U10952 ( .A1(n9722), .A2(n9721), .A3(n9720), .ZN(P1_U3254) );
  INV_X1 U10953 ( .A(n9723), .ZN(n9724) );
  NOR2_X1 U10954 ( .A1(n9725), .A2(n9724), .ZN(n9727) );
  XNOR2_X1 U10955 ( .A(n9727), .B(n9726), .ZN(n9736) );
  NAND2_X1 U10956 ( .A1(n9728), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9729) );
  NAND2_X1 U10957 ( .A1(n9730), .A2(n9729), .ZN(n9731) );
  XNOR2_X1 U10958 ( .A(n9731), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9739) );
  INV_X1 U10959 ( .A(n9739), .ZN(n9732) );
  AOI22_X1 U10960 ( .A1(n9736), .A2(n10235), .B1(n9733), .B2(n9732), .ZN(n9742) );
  INV_X1 U10961 ( .A(n9734), .ZN(n9738) );
  OAI21_X1 U10962 ( .B1(n9736), .B2(n9735), .A(n10239), .ZN(n9737) );
  AOI21_X1 U10963 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9741) );
  NAND2_X1 U10964 ( .A1(n9759), .A2(n9753), .ZN(n9746) );
  INV_X1 U10965 ( .A(P1_B_REG_SCAN_IN), .ZN(n9747) );
  NOR2_X1 U10966 ( .A1(n10184), .A2(n9747), .ZN(n9748) );
  OR2_X1 U10967 ( .A1(n10016), .A2(n9748), .ZN(n9767) );
  NOR2_X1 U10968 ( .A1(n9767), .A2(n9749), .ZN(n10046) );
  INV_X1 U10969 ( .A(n10046), .ZN(n9750) );
  NOR2_X1 U10970 ( .A1(n9750), .A2(n10021), .ZN(n9755) );
  AOI21_X1 U10971 ( .B1(n10021), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9755), .ZN(
        n9752) );
  NAND2_X1 U10972 ( .A1(n10043), .A2(n10032), .ZN(n9751) );
  OAI211_X1 U10973 ( .C1(n10045), .C2(n10034), .A(n9752), .B(n9751), .ZN(
        P1_U3261) );
  XNOR2_X1 U10974 ( .A(n9759), .B(n9753), .ZN(n10048) );
  NOR2_X1 U10975 ( .A1(n9753), .A2(n10024), .ZN(n9754) );
  AOI211_X1 U10976 ( .C1(n10021), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9755), .B(
        n9754), .ZN(n9756) );
  OAI21_X1 U10977 ( .B1(n10048), .B2(n10034), .A(n9756), .ZN(P1_U3262) );
  NAND2_X1 U10978 ( .A1(n9757), .A2(n9781), .ZN(n10060) );
  NAND2_X1 U10979 ( .A1(n10062), .A2(n10060), .ZN(n9758) );
  XNOR2_X1 U10980 ( .A(n9758), .B(n10061), .ZN(n9774) );
  AOI211_X1 U10981 ( .C1(n10050), .C2(n9760), .A(n10320), .B(n9759), .ZN(
        n10055) );
  AOI22_X1 U10982 ( .A1(n9761), .A2(n10029), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10021), .ZN(n9762) );
  OAI21_X1 U10983 ( .B1(n10052), .B2(n10024), .A(n9762), .ZN(n9772) );
  INV_X1 U10984 ( .A(n9763), .ZN(n9765) );
  NAND2_X1 U10985 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  XNOR2_X1 U10986 ( .A(n9766), .B(n10058), .ZN(n9771) );
  OAI22_X1 U10987 ( .A1(n9769), .A2(n10014), .B1(n9768), .B2(n9767), .ZN(n9770) );
  OAI21_X1 U10988 ( .B1(n9774), .B2(n10028), .A(n9773), .ZN(P1_U3355) );
  XOR2_X1 U10989 ( .A(n9780), .B(n9775), .Z(n10071) );
  AOI21_X1 U10990 ( .B1(n10067), .B2(n9792), .A(n4922), .ZN(n10068) );
  AOI22_X1 U10991 ( .A1(n9777), .A2(n10029), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10021), .ZN(n9778) );
  OAI21_X1 U10992 ( .B1(n9779), .B2(n10024), .A(n9778), .ZN(n9786) );
  AOI211_X1 U10993 ( .C1(n10068), .C2(n9990), .A(n9786), .B(n9785), .ZN(n9787)
         );
  OAI21_X1 U10994 ( .B1(n10071), .B2(n10028), .A(n9787), .ZN(P1_U3264) );
  OAI21_X1 U10995 ( .B1(n9789), .B2(n9797), .A(n9788), .ZN(n10076) );
  INV_X1 U10996 ( .A(n9815), .ZN(n9790) );
  NAND2_X1 U10997 ( .A1(n9790), .A2(n10072), .ZN(n9791) );
  AND2_X1 U10998 ( .A1(n9792), .A2(n9791), .ZN(n10073) );
  NAND2_X1 U10999 ( .A1(n10072), .A2(n10032), .ZN(n9794) );
  NAND2_X1 U11000 ( .A1(n10021), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9793) );
  OAI211_X1 U11001 ( .C1(n9999), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9796)
         );
  AOI21_X1 U11002 ( .B1(n10073), .B2(n9990), .A(n9796), .ZN(n9804) );
  XNOR2_X1 U11003 ( .A(n9797), .B(n9798), .ZN(n9802) );
  OAI22_X1 U11004 ( .A1(n9800), .A2(n10016), .B1(n9799), .B2(n10014), .ZN(
        n9801) );
  AOI21_X1 U11005 ( .B1(n9802), .B2(n9981), .A(n9801), .ZN(n10075) );
  OR2_X1 U11006 ( .A1(n10075), .A2(n10021), .ZN(n9803) );
  OAI211_X1 U11007 ( .C1(n10076), .C2(n10028), .A(n9804), .B(n9803), .ZN(
        P1_U3265) );
  XNOR2_X1 U11008 ( .A(n9805), .B(n9806), .ZN(n10081) );
  INV_X1 U11009 ( .A(n9822), .ZN(n9809) );
  OAI21_X1 U11010 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9811) );
  NAND3_X1 U11011 ( .A1(n9811), .A2(n9981), .A3(n9810), .ZN(n9813) );
  NAND2_X1 U11012 ( .A1(n6361), .A2(n9938), .ZN(n9812) );
  OAI211_X1 U11013 ( .C1(n9852), .C2(n10014), .A(n9813), .B(n9812), .ZN(n10077) );
  INV_X1 U11014 ( .A(n9814), .ZN(n9832) );
  AOI211_X1 U11015 ( .C1(n10079), .C2(n9832), .A(n10320), .B(n9815), .ZN(
        n10078) );
  NAND2_X1 U11016 ( .A1(n10078), .A2(n10019), .ZN(n9818) );
  AOI22_X1 U11017 ( .A1(n9816), .A2(n10029), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10021), .ZN(n9817) );
  OAI211_X1 U11018 ( .C1(n9819), .C2(n10024), .A(n9818), .B(n9817), .ZN(n9820)
         );
  AOI21_X1 U11019 ( .B1(n10077), .B2(n10036), .A(n9820), .ZN(n9821) );
  OAI21_X1 U11020 ( .B1(n10081), .B2(n10028), .A(n9821), .ZN(P1_U3266) );
  OAI21_X1 U11021 ( .B1(n4428), .B2(n9823), .A(n9822), .ZN(n9826) );
  AOI222_X1 U11022 ( .A1(n9981), .A2(n9826), .B1(n9825), .B2(n9936), .C1(n9824), .C2(n9938), .ZN(n10085) );
  XOR2_X1 U11023 ( .A(n9827), .B(n9828), .Z(n10082) );
  NAND2_X1 U11024 ( .A1(n10082), .A2(n10041), .ZN(n9838) );
  INV_X1 U11025 ( .A(n9829), .ZN(n9831) );
  OAI22_X1 U11026 ( .A1(n9831), .A2(n9999), .B1(n9830), .B2(n10036), .ZN(n9835) );
  OAI211_X1 U11027 ( .C1(n9833), .C2(n9844), .A(n9832), .B(n10307), .ZN(n10083) );
  NOR2_X1 U11028 ( .A1(n10083), .A2(n7917), .ZN(n9834) );
  AOI211_X1 U11029 ( .C1(n10032), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9837)
         );
  OAI211_X1 U11030 ( .C1(n10021), .C2(n10085), .A(n9838), .B(n9837), .ZN(
        P1_U3267) );
  OAI21_X1 U11031 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n10091) );
  NAND2_X1 U11032 ( .A1(n9856), .A2(n10089), .ZN(n9842) );
  NAND2_X1 U11033 ( .A1(n9842), .A2(n10307), .ZN(n9843) );
  NOR2_X1 U11034 ( .A1(n9844), .A2(n9843), .ZN(n10088) );
  NAND2_X1 U11035 ( .A1(n10089), .A2(n10032), .ZN(n9846) );
  NAND2_X1 U11036 ( .A1(n10021), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9845) );
  OAI211_X1 U11037 ( .C1(n9999), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9848)
         );
  AOI21_X1 U11038 ( .B1(n10088), .B2(n10019), .A(n9848), .ZN(n9854) );
  XNOR2_X1 U11039 ( .A(n9850), .B(n9849), .ZN(n9851) );
  OAI222_X1 U11040 ( .A1(n10016), .A2(n9852), .B1(n10014), .B2(n9886), .C1(
        n10012), .C2(n9851), .ZN(n10087) );
  NAND2_X1 U11041 ( .A1(n10087), .A2(n10036), .ZN(n9853) );
  OAI211_X1 U11042 ( .C1(n10091), .C2(n10028), .A(n9854), .B(n9853), .ZN(
        P1_U3268) );
  XNOR2_X1 U11043 ( .A(n9855), .B(n4417), .ZN(n10096) );
  INV_X1 U11044 ( .A(n9856), .ZN(n9857) );
  AOI21_X1 U11045 ( .B1(n10092), .B2(n9874), .A(n9857), .ZN(n10093) );
  AOI22_X1 U11046 ( .A1(n9858), .A2(n10029), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10021), .ZN(n9859) );
  OAI21_X1 U11047 ( .B1(n9860), .B2(n10024), .A(n9859), .ZN(n9871) );
  INV_X1 U11048 ( .A(n9861), .ZN(n9865) );
  AOI21_X1 U11049 ( .B1(n9881), .B2(n9862), .A(n4417), .ZN(n9863) );
  AOI211_X1 U11050 ( .C1(n9865), .C2(n9864), .A(n10012), .B(n9863), .ZN(n9869)
         );
  OAI22_X1 U11051 ( .A1(n9867), .A2(n10016), .B1(n9866), .B2(n10014), .ZN(
        n9868) );
  NOR2_X1 U11052 ( .A1(n9869), .A2(n9868), .ZN(n10095) );
  NOR2_X1 U11053 ( .A1(n10095), .A2(n10021), .ZN(n9870) );
  AOI211_X1 U11054 ( .C1(n10093), .C2(n9990), .A(n9871), .B(n9870), .ZN(n9872)
         );
  OAI21_X1 U11055 ( .B1(n10096), .B2(n10028), .A(n9872), .ZN(P1_U3269) );
  XNOR2_X1 U11056 ( .A(n9873), .B(n6414), .ZN(n10100) );
  INV_X1 U11057 ( .A(n9874), .ZN(n9875) );
  AOI211_X1 U11058 ( .C1(n4377), .C2(n9891), .A(n10320), .B(n9875), .ZN(n10098) );
  NOR2_X1 U11059 ( .A1(n9876), .A2(n10024), .ZN(n9880) );
  OAI22_X1 U11060 ( .A1(n10036), .A2(n9878), .B1(n9877), .B2(n9999), .ZN(n9879) );
  AOI211_X1 U11061 ( .C1(n10098), .C2(n10019), .A(n9880), .B(n9879), .ZN(n9888) );
  INV_X1 U11062 ( .A(n9881), .ZN(n9882) );
  AOI21_X1 U11063 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9885) );
  OAI222_X1 U11064 ( .A1(n10014), .A2(n9917), .B1(n10016), .B2(n9886), .C1(
        n10012), .C2(n9885), .ZN(n10097) );
  NAND2_X1 U11065 ( .A1(n10097), .A2(n10036), .ZN(n9887) );
  OAI211_X1 U11066 ( .C1(n10100), .C2(n10028), .A(n9888), .B(n9887), .ZN(
        P1_U3270) );
  XNOR2_X1 U11067 ( .A(n9889), .B(n9899), .ZN(n10105) );
  INV_X1 U11068 ( .A(n9890), .ZN(n9893) );
  INV_X1 U11069 ( .A(n9891), .ZN(n9892) );
  AOI211_X1 U11070 ( .C1(n10103), .C2(n9893), .A(n10320), .B(n9892), .ZN(
        n10102) );
  NOR2_X1 U11071 ( .A1(n9894), .A2(n10024), .ZN(n9897) );
  OAI22_X1 U11072 ( .A1(n10036), .A2(n6692), .B1(n9895), .B2(n9999), .ZN(n9896) );
  AOI211_X1 U11073 ( .C1(n10102), .C2(n10019), .A(n9897), .B(n9896), .ZN(n9906) );
  INV_X1 U11074 ( .A(n9898), .ZN(n9913) );
  OAI21_X1 U11075 ( .B1(n9913), .B2(n9900), .A(n9899), .ZN(n9902) );
  NAND3_X1 U11076 ( .A1(n9902), .A2(n9981), .A3(n9901), .ZN(n9904) );
  AOI22_X1 U11077 ( .A1(n4839), .A2(n9938), .B1(n9936), .B2(n9925), .ZN(n9903)
         );
  NAND2_X1 U11078 ( .A1(n9904), .A2(n9903), .ZN(n10101) );
  NAND2_X1 U11079 ( .A1(n10101), .A2(n10036), .ZN(n9905) );
  OAI211_X1 U11080 ( .C1(n10105), .C2(n10028), .A(n9906), .B(n9905), .ZN(
        P1_U3271) );
  XNOR2_X1 U11081 ( .A(n9907), .B(n9915), .ZN(n10110) );
  INV_X1 U11082 ( .A(n9928), .ZN(n9908) );
  AOI211_X1 U11083 ( .C1(n10108), .C2(n9908), .A(n10320), .B(n9890), .ZN(
        n10107) );
  NOR2_X1 U11084 ( .A1(n9909), .A2(n10024), .ZN(n9912) );
  OAI22_X1 U11085 ( .A1(n10036), .A2(n6517), .B1(n9910), .B2(n9999), .ZN(n9911) );
  AOI211_X1 U11086 ( .C1(n10107), .C2(n10019), .A(n9912), .B(n9911), .ZN(n9920) );
  AOI21_X1 U11087 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  OAI222_X1 U11088 ( .A1(n10014), .A2(n9918), .B1(n10016), .B2(n9917), .C1(
        n10012), .C2(n9916), .ZN(n10106) );
  NAND2_X1 U11089 ( .A1(n10106), .A2(n10036), .ZN(n9919) );
  OAI211_X1 U11090 ( .C1(n10110), .C2(n10028), .A(n9920), .B(n9919), .ZN(
        P1_U3272) );
  INV_X1 U11091 ( .A(n9921), .ZN(n9923) );
  OAI21_X1 U11092 ( .B1(n9935), .B2(n9923), .A(n9922), .ZN(n9924) );
  XNOR2_X1 U11093 ( .A(n9924), .B(n9927), .ZN(n9926) );
  AOI222_X1 U11094 ( .A1(n9981), .A2(n9926), .B1(n6264), .B2(n9936), .C1(n9925), .C2(n9938), .ZN(n10116) );
  OR2_X1 U11095 ( .A1(n4469), .A2(n9927), .ZN(n10112) );
  NAND3_X1 U11096 ( .A1(n10112), .A2(n10111), .A3(n10041), .ZN(n9934) );
  AOI21_X1 U11097 ( .B1(n10113), .B2(n4464), .A(n9928), .ZN(n10114) );
  NOR2_X1 U11098 ( .A1(n9929), .A2(n10024), .ZN(n9932) );
  OAI22_X1 U11099 ( .A1(n10036), .A2(n8115), .B1(n9930), .B2(n9999), .ZN(n9931) );
  AOI211_X1 U11100 ( .C1(n10114), .C2(n9990), .A(n9932), .B(n9931), .ZN(n9933)
         );
  OAI211_X1 U11101 ( .C1(n10021), .C2(n10116), .A(n9934), .B(n9933), .ZN(
        P1_U3273) );
  XNOR2_X1 U11102 ( .A(n9935), .B(n9943), .ZN(n9940) );
  AOI222_X1 U11103 ( .A1(n9981), .A2(n9940), .B1(n9939), .B2(n9938), .C1(n9937), .C2(n9936), .ZN(n10121) );
  AOI21_X1 U11104 ( .B1(n9943), .B2(n9942), .A(n9941), .ZN(n10122) );
  INV_X1 U11105 ( .A(n10122), .ZN(n9950) );
  AOI21_X1 U11106 ( .B1(n9964), .B2(n10119), .A(n10320), .ZN(n9944) );
  AND2_X1 U11107 ( .A1(n9944), .A2(n4464), .ZN(n10118) );
  NAND2_X1 U11108 ( .A1(n10118), .A2(n10019), .ZN(n9947) );
  AOI22_X1 U11109 ( .A1(n10021), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9945), 
        .B2(n10029), .ZN(n9946) );
  OAI211_X1 U11110 ( .C1(n9948), .C2(n10024), .A(n9947), .B(n9946), .ZN(n9949)
         );
  AOI21_X1 U11111 ( .B1(n9950), .B2(n10041), .A(n9949), .ZN(n9951) );
  OAI21_X1 U11112 ( .B1(n10021), .B2(n10121), .A(n9951), .ZN(P1_U3274) );
  INV_X1 U11113 ( .A(n9953), .ZN(n9954) );
  NAND2_X1 U11114 ( .A1(n9977), .A2(n9954), .ZN(n9956) );
  XNOR2_X1 U11115 ( .A(n9956), .B(n9955), .ZN(n10127) );
  NAND2_X1 U11116 ( .A1(n9958), .A2(n9957), .ZN(n9960) );
  XNOR2_X1 U11117 ( .A(n9960), .B(n9959), .ZN(n9961) );
  OAI222_X1 U11118 ( .A1(n10016), .A2(n9962), .B1(n10014), .B2(n9997), .C1(
        n10012), .C2(n9961), .ZN(n10123) );
  NAND2_X1 U11119 ( .A1(n10123), .A2(n10036), .ZN(n9971) );
  OR2_X1 U11120 ( .A1(n9982), .A2(n9965), .ZN(n9963) );
  AND3_X1 U11121 ( .A1(n9964), .A2(n9963), .A3(n10307), .ZN(n10124) );
  NOR2_X1 U11122 ( .A1(n9965), .A2(n10024), .ZN(n9969) );
  OAI22_X1 U11123 ( .A1(n10036), .A2(n9967), .B1(n9966), .B2(n9999), .ZN(n9968) );
  AOI211_X1 U11124 ( .C1(n10124), .C2(n10019), .A(n9969), .B(n9968), .ZN(n9970) );
  OAI211_X1 U11125 ( .C1(n10127), .C2(n10028), .A(n9971), .B(n9970), .ZN(
        P1_U3275) );
  XNOR2_X1 U11126 ( .A(n9973), .B(n9972), .ZN(n9980) );
  OAI22_X1 U11127 ( .A1(n9974), .A2(n10016), .B1(n10015), .B2(n10014), .ZN(
        n9979) );
  NAND2_X1 U11128 ( .A1(n9952), .A2(n9975), .ZN(n9976) );
  NAND2_X1 U11129 ( .A1(n9977), .A2(n9976), .ZN(n10132) );
  NOR2_X1 U11130 ( .A1(n10132), .A2(n10311), .ZN(n9978) );
  AOI211_X1 U11131 ( .C1(n9981), .C2(n9980), .A(n9979), .B(n9978), .ZN(n10131)
         );
  AOI21_X1 U11132 ( .B1(n10128), .B2(n4912), .A(n9982), .ZN(n10129) );
  INV_X1 U11133 ( .A(n9983), .ZN(n9984) );
  AOI22_X1 U11134 ( .A1(n10021), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9984), 
        .B2(n10029), .ZN(n9985) );
  OAI21_X1 U11135 ( .B1(n9986), .B2(n10024), .A(n9985), .ZN(n9989) );
  NOR2_X1 U11136 ( .A1(n10132), .A2(n9987), .ZN(n9988) );
  AOI211_X1 U11137 ( .C1(n10129), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9991)
         );
  OAI21_X1 U11138 ( .B1(n10131), .B2(n10021), .A(n9991), .ZN(P1_U3276) );
  XNOR2_X1 U11139 ( .A(n9992), .B(n9993), .ZN(n10138) );
  XNOR2_X1 U11140 ( .A(n4496), .B(n9993), .ZN(n9995) );
  OAI222_X1 U11141 ( .A1(n10016), .A2(n9997), .B1(n10014), .B2(n9996), .C1(
        n10012), .C2(n9995), .ZN(n10134) );
  NAND2_X1 U11142 ( .A1(n10134), .A2(n10036), .ZN(n10005) );
  AOI211_X1 U11143 ( .C1(n10136), .C2(n5008), .A(n10320), .B(n9998), .ZN(
        n10135) );
  NOR2_X1 U11144 ( .A1(n4910), .A2(n10024), .ZN(n10003) );
  OAI22_X1 U11145 ( .A1(n10036), .A2(n10001), .B1(n10000), .B2(n9999), .ZN(
        n10002) );
  AOI211_X1 U11146 ( .C1(n10135), .C2(n10019), .A(n10003), .B(n10002), .ZN(
        n10004) );
  OAI211_X1 U11147 ( .C1(n10138), .C2(n10028), .A(n10005), .B(n10004), .ZN(
        P1_U3277) );
  XNOR2_X1 U11148 ( .A(n10006), .B(n10010), .ZN(n10143) );
  INV_X1 U11149 ( .A(n10007), .ZN(n10008) );
  AOI21_X1 U11150 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10011) );
  OAI222_X1 U11151 ( .A1(n10016), .A2(n10015), .B1(n10014), .B2(n10013), .C1(
        n10012), .C2(n10011), .ZN(n10139) );
  INV_X1 U11152 ( .A(n10141), .ZN(n10025) );
  INV_X1 U11153 ( .A(n5008), .ZN(n10017) );
  AOI211_X1 U11154 ( .C1(n10141), .C2(n10018), .A(n10320), .B(n10017), .ZN(
        n10140) );
  NAND2_X1 U11155 ( .A1(n10140), .A2(n10019), .ZN(n10023) );
  AOI22_X1 U11156 ( .A1(n10021), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10020), 
        .B2(n10029), .ZN(n10022) );
  OAI211_X1 U11157 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10026) );
  AOI21_X1 U11158 ( .B1(n10139), .B2(n10036), .A(n10026), .ZN(n10027) );
  OAI21_X1 U11159 ( .B1(n10028), .B2(n10143), .A(n10027), .ZN(P1_U3278) );
  AOI22_X1 U11160 ( .A1(n10032), .A2(n10031), .B1(n10030), .B2(n10029), .ZN(
        n10033) );
  OAI21_X1 U11161 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(n10039) );
  MUX2_X1 U11162 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10037), .S(n10036), .Z(
        n10038) );
  AOI211_X1 U11163 ( .C1(n10041), .C2(n10040), .A(n10039), .B(n10038), .ZN(
        n10042) );
  INV_X1 U11164 ( .A(n10042), .ZN(P1_U3280) );
  AOI21_X1 U11165 ( .B1(n10043), .B2(n10299), .A(n10046), .ZN(n10044) );
  OAI21_X1 U11166 ( .B1(n10045), .B2(n10320), .A(n10044), .ZN(n10151) );
  MUX2_X1 U11167 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10151), .S(n10344), .Z(
        P1_U3554) );
  AOI21_X1 U11168 ( .B1(n9407), .B2(n10299), .A(n10046), .ZN(n10047) );
  OAI21_X1 U11169 ( .B1(n10048), .B2(n10320), .A(n10047), .ZN(n10152) );
  MUX2_X1 U11170 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10152), .S(n10344), .Z(
        P1_U3553) );
  INV_X1 U11171 ( .A(n10060), .ZN(n10049) );
  NAND2_X1 U11172 ( .A1(n10049), .A2(n10325), .ZN(n10054) );
  OAI211_X1 U11173 ( .C1(n10054), .C2(n10051), .A(n10285), .B(n10050), .ZN(
        n10057) );
  OAI21_X1 U11174 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n10056) );
  AOI21_X1 U11175 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10066) );
  INV_X1 U11176 ( .A(n10062), .ZN(n10059) );
  NAND3_X1 U11177 ( .A1(n10059), .A2(n10058), .A3(n10325), .ZN(n10064) );
  NAND4_X1 U11178 ( .A1(n10062), .A2(n10061), .A3(n10325), .A4(n10060), .ZN(
        n10063) );
  NAND4_X1 U11179 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10153) );
  MUX2_X1 U11180 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10153), .S(n10344), .Z(
        P1_U3552) );
  AOI22_X1 U11181 ( .A1(n10068), .A2(n10307), .B1(n10299), .B2(n10067), .ZN(
        n10069) );
  OAI211_X1 U11182 ( .C1(n10071), .C2(n10144), .A(n10070), .B(n10069), .ZN(
        n10155) );
  MUX2_X1 U11183 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10155), .S(n10344), .Z(
        P1_U3550) );
  AOI22_X1 U11184 ( .A1(n10073), .A2(n10307), .B1(n10299), .B2(n10072), .ZN(
        n10074) );
  OAI211_X1 U11185 ( .C1(n10076), .C2(n10144), .A(n10075), .B(n10074), .ZN(
        n10156) );
  MUX2_X1 U11186 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10156), .S(n10344), .Z(
        P1_U3549) );
  AOI211_X1 U11187 ( .C1(n10299), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10080) );
  OAI21_X1 U11188 ( .B1(n10081), .B2(n10144), .A(n10080), .ZN(n10157) );
  MUX2_X1 U11189 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10157), .S(n10344), .Z(
        P1_U3548) );
  NAND2_X1 U11190 ( .A1(n10082), .A2(n10325), .ZN(n10086) );
  NAND4_X1 U11191 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10158) );
  MUX2_X1 U11192 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10158), .S(n10344), .Z(
        P1_U3547) );
  AOI211_X1 U11193 ( .C1(n10299), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10090) );
  OAI21_X1 U11194 ( .B1(n10091), .B2(n10144), .A(n10090), .ZN(n10159) );
  MUX2_X1 U11195 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10159), .S(n10344), .Z(
        P1_U3546) );
  AOI22_X1 U11196 ( .A1(n10093), .A2(n10307), .B1(n10299), .B2(n10092), .ZN(
        n10094) );
  OAI211_X1 U11197 ( .C1(n10096), .C2(n10144), .A(n10095), .B(n10094), .ZN(
        n10160) );
  MUX2_X1 U11198 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10160), .S(n10344), .Z(
        P1_U3545) );
  AOI211_X1 U11199 ( .C1(n10299), .C2(n4377), .A(n10098), .B(n10097), .ZN(
        n10099) );
  OAI21_X1 U11200 ( .B1(n10100), .B2(n10144), .A(n10099), .ZN(n10161) );
  MUX2_X1 U11201 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10161), .S(n10344), .Z(
        P1_U3544) );
  AOI211_X1 U11202 ( .C1(n10299), .C2(n10103), .A(n10102), .B(n10101), .ZN(
        n10104) );
  OAI21_X1 U11203 ( .B1(n10105), .B2(n10144), .A(n10104), .ZN(n10162) );
  MUX2_X1 U11204 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10162), .S(n10344), .Z(
        P1_U3543) );
  AOI211_X1 U11205 ( .C1(n10299), .C2(n10108), .A(n10107), .B(n10106), .ZN(
        n10109) );
  OAI21_X1 U11206 ( .B1(n10144), .B2(n10110), .A(n10109), .ZN(n10163) );
  MUX2_X1 U11207 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10163), .S(n10344), .Z(
        P1_U3542) );
  NAND3_X1 U11208 ( .A1(n10112), .A2(n10111), .A3(n10325), .ZN(n10117) );
  AOI22_X1 U11209 ( .A1(n10114), .A2(n10307), .B1(n10299), .B2(n10113), .ZN(
        n10115) );
  NAND3_X1 U11210 ( .A1(n10117), .A2(n10116), .A3(n10115), .ZN(n10164) );
  MUX2_X1 U11211 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10164), .S(n10344), .Z(
        P1_U3541) );
  AOI21_X1 U11212 ( .B1(n10299), .B2(n10119), .A(n10118), .ZN(n10120) );
  OAI211_X1 U11213 ( .C1(n10122), .C2(n10144), .A(n10121), .B(n10120), .ZN(
        n10165) );
  MUX2_X1 U11214 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10165), .S(n10344), .Z(
        P1_U3540) );
  AOI211_X1 U11215 ( .C1(n10299), .C2(n10125), .A(n10124), .B(n10123), .ZN(
        n10126) );
  OAI21_X1 U11216 ( .B1(n10144), .B2(n10127), .A(n10126), .ZN(n10166) );
  MUX2_X1 U11217 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10166), .S(n10344), .Z(
        P1_U3539) );
  AOI22_X1 U11218 ( .A1(n10129), .A2(n10307), .B1(n10299), .B2(n10128), .ZN(
        n10130) );
  OAI211_X1 U11219 ( .C1(n10133), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10167) );
  MUX2_X1 U11220 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10167), .S(n10344), .Z(
        P1_U3538) );
  AOI211_X1 U11221 ( .C1(n10299), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10137) );
  OAI21_X1 U11222 ( .B1(n10144), .B2(n10138), .A(n10137), .ZN(n10168) );
  MUX2_X1 U11223 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10168), .S(n10344), .Z(
        P1_U3537) );
  AOI211_X1 U11224 ( .C1(n10299), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10142) );
  OAI21_X1 U11225 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(n10169) );
  MUX2_X1 U11226 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10169), .S(n10344), .Z(
        P1_U3536) );
  OAI21_X1 U11227 ( .B1(n10146), .B2(n10285), .A(n10145), .ZN(n10148) );
  AOI211_X1 U11228 ( .C1(n10149), .C2(n10325), .A(n10148), .B(n10147), .ZN(
        n10171) );
  NAND2_X1 U11229 ( .A1(n10341), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10150) );
  OAI21_X1 U11230 ( .B1(n10171), .B2(n10341), .A(n10150), .ZN(P1_U3535) );
  MUX2_X1 U11231 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10151), .S(n10328), .Z(
        P1_U3522) );
  MUX2_X1 U11232 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10152), .S(n10328), .Z(
        P1_U3521) );
  MUX2_X1 U11233 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10153), .S(n10328), .Z(
        P1_U3520) );
  MUX2_X1 U11234 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10154), .S(n10328), .Z(
        P1_U3519) );
  MUX2_X1 U11235 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10155), .S(n10328), .Z(
        P1_U3518) );
  MUX2_X1 U11236 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10156), .S(n10328), .Z(
        P1_U3517) );
  MUX2_X1 U11237 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10157), .S(n10328), .Z(
        P1_U3516) );
  MUX2_X1 U11238 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10158), .S(n10328), .Z(
        P1_U3515) );
  MUX2_X1 U11239 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10159), .S(n10328), .Z(
        P1_U3514) );
  MUX2_X1 U11240 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10160), .S(n10328), .Z(
        P1_U3513) );
  MUX2_X1 U11241 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10161), .S(n10272), .Z(
        P1_U3512) );
  MUX2_X1 U11242 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10162), .S(n10272), .Z(
        P1_U3511) );
  MUX2_X1 U11243 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10163), .S(n10272), .Z(
        P1_U3510) );
  MUX2_X1 U11244 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10164), .S(n10272), .Z(
        P1_U3508) );
  MUX2_X1 U11245 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10165), .S(n10272), .Z(
        P1_U3505) );
  MUX2_X1 U11246 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10166), .S(n10328), .Z(
        P1_U3502) );
  MUX2_X1 U11247 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10167), .S(n10328), .Z(
        P1_U3499) );
  MUX2_X1 U11248 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10168), .S(n10328), .Z(
        P1_U3496) );
  MUX2_X1 U11249 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10169), .S(n10328), .Z(
        P1_U3493) );
  NAND2_X1 U11250 ( .A1(n10326), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10170) );
  OAI21_X1 U11251 ( .B1(n10171), .B2(n10326), .A(n10170), .ZN(P1_U3490) );
  MUX2_X1 U11252 ( .A(n10172), .B(P1_D_REG_0__SCAN_IN), .S(n10255), .Z(
        P1_U3440) );
  NOR4_X1 U11253 ( .A1(n6030), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n10173), .ZN(n10175) );
  AOI21_X1 U11254 ( .B1(n10176), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10175), 
        .ZN(n10177) );
  OAI21_X1 U11255 ( .B1(n10178), .B2(n10186), .A(n10177), .ZN(P1_U3322) );
  OAI222_X1 U11256 ( .A1(n10186), .A2(n10181), .B1(n10180), .B2(P1_U3084), 
        .C1(n10179), .C2(n10182), .ZN(P1_U3325) );
  OAI222_X1 U11257 ( .A1(n10186), .A2(n10185), .B1(n10184), .B2(P1_U3084), 
        .C1(n10183), .C2(n10182), .ZN(P1_U3326) );
  OAI222_X1 U11258 ( .A1(n10186), .A2(n10189), .B1(P1_U3084), .B2(n10188), 
        .C1(n10187), .C2(n10182), .ZN(P1_U3327) );
  MUX2_X1 U11259 ( .A(n10190), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11260 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10191) );
  AOI21_X1 U11261 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10191), .ZN(n10451) );
  NOR2_X1 U11262 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10192) );
  AOI21_X1 U11263 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10192), .ZN(n10454) );
  NOR2_X1 U11264 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10193) );
  AOI21_X1 U11265 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10193), .ZN(n10457) );
  NOR2_X1 U11266 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n10194) );
  AOI21_X1 U11267 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10194), .ZN(n10460) );
  NOR2_X1 U11268 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n10195) );
  AOI21_X1 U11269 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10195), .ZN(n10463) );
  INV_X1 U11270 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10243) );
  NOR2_X1 U11271 ( .A1(n10197), .A2(n10196), .ZN(n10487) );
  NOR2_X1 U11272 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10205) );
  XNOR2_X1 U11273 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10496) );
  AOI22_X1 U11274 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10203), .B2(n6536), .ZN(n10494) );
  NAND2_X1 U11275 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10201) );
  INV_X1 U11276 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10199) );
  AOI21_X1 U11277 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10445) );
  NAND3_X1 U11278 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10447) );
  OAI21_X1 U11279 ( .B1(n10445), .B2(n7001), .A(n10447), .ZN(n10491) );
  NAND2_X1 U11280 ( .A1(n10492), .A2(n10491), .ZN(n10200) );
  NAND2_X1 U11281 ( .A1(n10201), .A2(n10200), .ZN(n10493) );
  NAND2_X1 U11282 ( .A1(n10494), .A2(n10493), .ZN(n10202) );
  NOR2_X1 U11283 ( .A1(n10496), .A2(n10495), .ZN(n10204) );
  NOR2_X1 U11284 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  NOR2_X1 U11285 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10206), .ZN(n10475) );
  NAND2_X1 U11286 ( .A1(n10208), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10210) );
  XOR2_X1 U11287 ( .A(n10208), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10473) );
  NAND2_X1 U11288 ( .A1(n10473), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10209) );
  INV_X1 U11289 ( .A(n10488), .ZN(n10211) );
  NOR2_X1 U11290 ( .A1(n10243), .A2(n10212), .ZN(n10213) );
  INV_X1 U11291 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10486) );
  XNOR2_X1 U11292 ( .A(n10243), .B(n10212), .ZN(n10485) );
  NOR2_X1 U11293 ( .A1(n10214), .A2(n10215), .ZN(n10216) );
  XNOR2_X1 U11294 ( .A(n10215), .B(n10214), .ZN(n10482) );
  NAND2_X1 U11295 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10217) );
  OAI21_X1 U11296 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10217), .ZN(n10471) );
  NAND2_X1 U11297 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10218) );
  OAI21_X1 U11298 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10218), .ZN(n10468) );
  NOR2_X1 U11299 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10219) );
  AOI21_X1 U11300 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10219), .ZN(n10465) );
  NAND2_X1 U11301 ( .A1(n10466), .A2(n10465), .ZN(n10464) );
  NAND2_X1 U11302 ( .A1(n10463), .A2(n10462), .ZN(n10461) );
  NAND2_X1 U11303 ( .A1(n10460), .A2(n10459), .ZN(n10458) );
  NAND2_X1 U11304 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  OAI21_X1 U11305 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10455), .ZN(n10453) );
  NAND2_X1 U11306 ( .A1(n10454), .A2(n10453), .ZN(n10452) );
  OAI21_X1 U11307 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10452), .ZN(n10450) );
  NAND2_X1 U11308 ( .A1(n10451), .A2(n10450), .ZN(n10449) );
  NOR2_X1 U11309 ( .A1(n10479), .A2(n10478), .ZN(n10220) );
  NAND2_X1 U11310 ( .A1(n10479), .A2(n10478), .ZN(n10477) );
  OAI21_X1 U11311 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10220), .A(n10477), 
        .ZN(n10222) );
  XOR2_X1 U11312 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n10221) );
  XNOR2_X1 U11313 ( .A(n10222), .B(n10221), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11314 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11315 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  NAND2_X1 U11316 ( .A1(n10226), .A2(n10223), .ZN(n10230) );
  INV_X1 U11317 ( .A(n10224), .ZN(n10225) );
  OAI21_X1 U11318 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(n10229) );
  AOI21_X1 U11319 ( .B1(n10230), .B2(n10229), .A(n10228), .ZN(n10241) );
  XNOR2_X1 U11320 ( .A(n10231), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n10232) );
  XNOR2_X1 U11321 ( .A(n10233), .B(n10232), .ZN(n10234) );
  NAND2_X1 U11322 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  OAI211_X1 U11323 ( .C1(n10239), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10240) );
  NOR2_X1 U11324 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  OAI21_X1 U11325 ( .B1(n10244), .B2(n10243), .A(n10242), .ZN(P1_U3249) );
  NOR2_X1 U11326 ( .A1(n10254), .A2(n10245), .ZN(P1_U3292) );
  AND2_X1 U11327 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10255), .ZN(P1_U3293) );
  AND2_X1 U11328 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10255), .ZN(P1_U3294) );
  AND2_X1 U11329 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10255), .ZN(P1_U3295) );
  AND2_X1 U11330 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10255), .ZN(P1_U3296) );
  AND2_X1 U11331 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10255), .ZN(P1_U3297) );
  AND2_X1 U11332 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10255), .ZN(P1_U3298) );
  NOR2_X1 U11333 ( .A1(n10254), .A2(n10246), .ZN(P1_U3299) );
  AND2_X1 U11334 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10255), .ZN(P1_U3300) );
  NOR2_X1 U11335 ( .A1(n10254), .A2(n10247), .ZN(P1_U3301) );
  INV_X1 U11336 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U11337 ( .A1(n10254), .A2(n10248), .ZN(P1_U3302) );
  NOR2_X1 U11338 ( .A1(n10254), .A2(n10249), .ZN(P1_U3303) );
  AND2_X1 U11339 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10255), .ZN(P1_U3304) );
  AND2_X1 U11340 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10255), .ZN(P1_U3305) );
  AND2_X1 U11341 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10255), .ZN(P1_U3306) );
  NOR2_X1 U11342 ( .A1(n10254), .A2(n10250), .ZN(P1_U3307) );
  AND2_X1 U11343 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10255), .ZN(P1_U3308) );
  AND2_X1 U11344 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10255), .ZN(P1_U3309) );
  NOR2_X1 U11345 ( .A1(n10254), .A2(n10251), .ZN(P1_U3310) );
  AND2_X1 U11346 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10255), .ZN(P1_U3311) );
  AND2_X1 U11347 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10255), .ZN(P1_U3312) );
  AND2_X1 U11348 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10255), .ZN(P1_U3313) );
  AND2_X1 U11349 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10255), .ZN(P1_U3314) );
  NOR2_X1 U11350 ( .A1(n10254), .A2(n10252), .ZN(P1_U3315) );
  AND2_X1 U11351 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10255), .ZN(P1_U3316) );
  AND2_X1 U11352 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10255), .ZN(P1_U3317) );
  NOR2_X1 U11353 ( .A1(n10254), .A2(n10253), .ZN(P1_U3318) );
  AND2_X1 U11354 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10255), .ZN(P1_U3319) );
  AND2_X1 U11355 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10255), .ZN(P1_U3320) );
  AND2_X1 U11356 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10255), .ZN(P1_U3321) );
  AOI211_X1 U11357 ( .C1(n10258), .C2(n10316), .A(n10257), .B(n10256), .ZN(
        n10259) );
  AND2_X1 U11358 ( .A1(n10260), .A2(n10259), .ZN(n10330) );
  INV_X1 U11359 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11360 ( .A1(n10272), .A2(n10330), .B1(n10261), .B2(n10326), .ZN(
        P1_U3457) );
  INV_X1 U11361 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U11362 ( .A1(n10272), .A2(n10263), .B1(n10262), .B2(n10326), .ZN(
        P1_U3460) );
  NAND2_X1 U11363 ( .A1(n10307), .A2(n10264), .ZN(n10266) );
  OAI22_X1 U11364 ( .A1(n10267), .A2(n10285), .B1(n10266), .B2(n10265), .ZN(
        n10269) );
  AOI211_X1 U11365 ( .C1(n10316), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10331) );
  INV_X1 U11366 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U11367 ( .A1(n10272), .A2(n10331), .B1(n10271), .B2(n10326), .ZN(
        P1_U3463) );
  INV_X1 U11368 ( .A(n10273), .ZN(n10279) );
  OAI21_X1 U11369 ( .B1(n10275), .B2(n10320), .A(n10274), .ZN(n10278) );
  INV_X1 U11370 ( .A(n10276), .ZN(n10277) );
  AOI211_X1 U11371 ( .C1(n10325), .C2(n10279), .A(n10278), .B(n10277), .ZN(
        n10333) );
  AOI22_X1 U11372 ( .A1(n10328), .A2(n10333), .B1(n10280), .B2(n10326), .ZN(
        P1_U3466) );
  NAND3_X1 U11373 ( .A1(n10282), .A2(n10325), .A3(n10281), .ZN(n10284) );
  OAI211_X1 U11374 ( .C1(n10286), .C2(n10285), .A(n10284), .B(n10283), .ZN(
        n10287) );
  NOR2_X1 U11375 ( .A1(n10288), .A2(n10287), .ZN(n10334) );
  AOI22_X1 U11376 ( .A1(n10328), .A2(n10334), .B1(n6119), .B2(n10326), .ZN(
        P1_U3469) );
  INV_X1 U11377 ( .A(n10292), .ZN(n10296) );
  NAND2_X1 U11378 ( .A1(n10289), .A2(n10307), .ZN(n10291) );
  OAI211_X1 U11379 ( .C1(n10292), .C2(n10311), .A(n10291), .B(n10290), .ZN(
        n10295) );
  INV_X1 U11380 ( .A(n10293), .ZN(n10294) );
  AOI211_X1 U11381 ( .C1(n10316), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10336) );
  INV_X1 U11382 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11383 ( .A1(n10328), .A2(n10336), .B1(n10297), .B2(n10326), .ZN(
        P1_U3472) );
  NAND2_X1 U11384 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  NAND2_X1 U11385 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  AOI21_X1 U11386 ( .B1(n10303), .B2(n10325), .A(n10302), .ZN(n10304) );
  AND2_X1 U11387 ( .A1(n10305), .A2(n10304), .ZN(n10338) );
  INV_X1 U11388 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U11389 ( .A1(n10328), .A2(n10338), .B1(n10306), .B2(n10326), .ZN(
        P1_U3475) );
  INV_X1 U11390 ( .A(n10312), .ZN(n10315) );
  NAND2_X1 U11391 ( .A1(n10308), .A2(n10307), .ZN(n10310) );
  OAI211_X1 U11392 ( .C1(n10312), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10314) );
  AOI211_X1 U11393 ( .C1(n10316), .C2(n10315), .A(n10314), .B(n10313), .ZN(
        n10340) );
  INV_X1 U11394 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U11395 ( .A1(n10328), .A2(n10340), .B1(n10317), .B2(n10326), .ZN(
        P1_U3478) );
  INV_X1 U11396 ( .A(n10318), .ZN(n10319) );
  OAI21_X1 U11397 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(n10323) );
  AOI211_X1 U11398 ( .C1(n10325), .C2(n10324), .A(n10323), .B(n10322), .ZN(
        n10343) );
  INV_X1 U11399 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U11400 ( .A1(n10328), .A2(n10343), .B1(n10327), .B2(n10326), .ZN(
        P1_U3481) );
  AOI22_X1 U11401 ( .A1(n10344), .A2(n10330), .B1(n10329), .B2(n10341), .ZN(
        P1_U3524) );
  AOI22_X1 U11402 ( .A1(n10344), .A2(n10331), .B1(n6855), .B2(n10341), .ZN(
        P1_U3526) );
  INV_X1 U11403 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U11404 ( .A1(n10344), .A2(n10333), .B1(n10332), .B2(n10341), .ZN(
        P1_U3527) );
  AOI22_X1 U11405 ( .A1(n10344), .A2(n10334), .B1(n6860), .B2(n10341), .ZN(
        P1_U3528) );
  AOI22_X1 U11406 ( .A1(n10344), .A2(n10336), .B1(n10335), .B2(n10341), .ZN(
        P1_U3529) );
  AOI22_X1 U11407 ( .A1(n10344), .A2(n10338), .B1(n10337), .B2(n10341), .ZN(
        P1_U3530) );
  INV_X1 U11408 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U11409 ( .A1(n10344), .A2(n10340), .B1(n10339), .B2(n10341), .ZN(
        P1_U3531) );
  AOI22_X1 U11410 ( .A1(n10344), .A2(n10343), .B1(n10342), .B2(n10341), .ZN(
        P1_U3532) );
  INV_X1 U11411 ( .A(n10345), .ZN(n10346) );
  AOI21_X1 U11412 ( .B1(n10347), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n10346), 
        .ZN(n10362) );
  OAI211_X1 U11413 ( .C1(n10351), .C2(n10350), .A(n10349), .B(n10348), .ZN(
        n10361) );
  INV_X1 U11414 ( .A(n10352), .ZN(n10353) );
  NAND2_X1 U11415 ( .A1(n10354), .A2(n10353), .ZN(n10360) );
  OAI211_X1 U11416 ( .C1(n10358), .C2(n10357), .A(n10356), .B(n10355), .ZN(
        n10359) );
  NAND4_X1 U11417 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        P2_U3262) );
  AND2_X1 U11418 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10376), .ZN(P2_U3297) );
  AND2_X1 U11419 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10376), .ZN(P2_U3298) );
  AND2_X1 U11420 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10376), .ZN(P2_U3299) );
  NOR2_X1 U11421 ( .A1(n10373), .A2(n10365), .ZN(P2_U3300) );
  NOR2_X1 U11422 ( .A1(n10373), .A2(n10366), .ZN(P2_U3301) );
  NOR2_X1 U11423 ( .A1(n10373), .A2(n10367), .ZN(P2_U3302) );
  AND2_X1 U11424 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10376), .ZN(P2_U3303) );
  AND2_X1 U11425 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10376), .ZN(P2_U3304) );
  AND2_X1 U11426 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10376), .ZN(P2_U3305) );
  NOR2_X1 U11427 ( .A1(n10373), .A2(n10368), .ZN(P2_U3306) );
  AND2_X1 U11428 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10376), .ZN(P2_U3307) );
  NOR2_X1 U11429 ( .A1(n10373), .A2(n10369), .ZN(P2_U3308) );
  AND2_X1 U11430 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10376), .ZN(P2_U3309) );
  NOR2_X1 U11431 ( .A1(n10373), .A2(n10370), .ZN(P2_U3310) );
  AND2_X1 U11432 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10376), .ZN(P2_U3311) );
  AND2_X1 U11433 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10376), .ZN(P2_U3312) );
  AND2_X1 U11434 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10376), .ZN(P2_U3313) );
  NOR2_X1 U11435 ( .A1(n10373), .A2(n10371), .ZN(P2_U3314) );
  NOR2_X1 U11436 ( .A1(n10373), .A2(n10372), .ZN(P2_U3315) );
  AND2_X1 U11437 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10376), .ZN(P2_U3316) );
  AND2_X1 U11438 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10376), .ZN(P2_U3317) );
  AND2_X1 U11439 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10376), .ZN(P2_U3318) );
  AND2_X1 U11440 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10376), .ZN(P2_U3319) );
  AND2_X1 U11441 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10376), .ZN(P2_U3320) );
  AND2_X1 U11442 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10376), .ZN(P2_U3321) );
  AND2_X1 U11443 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10376), .ZN(P2_U3322) );
  AND2_X1 U11444 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10376), .ZN(P2_U3323) );
  AND2_X1 U11445 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10376), .ZN(P2_U3324) );
  AND2_X1 U11446 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10376), .ZN(P2_U3325) );
  AND2_X1 U11447 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10376), .ZN(P2_U3326) );
  AOI22_X1 U11448 ( .A1(n10375), .A2(n10376), .B1(n10379), .B2(n10374), .ZN(
        P2_U3437) );
  AOI22_X1 U11449 ( .A1(n10379), .A2(n10378), .B1(n10377), .B2(n10376), .ZN(
        P2_U3438) );
  OAI21_X1 U11450 ( .B1(n10380), .B2(n10382), .A(n10381), .ZN(n10384) );
  AOI21_X1 U11451 ( .B1(n10382), .B2(n10381), .A(n8356), .ZN(n10383) );
  AOI21_X1 U11452 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(n10388) );
  INV_X1 U11453 ( .A(n10386), .ZN(n10387) );
  NOR2_X1 U11454 ( .A1(n10388), .A2(n10387), .ZN(n10435) );
  INV_X1 U11455 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U11456 ( .A1(n10433), .A2(n10435), .B1(n10389), .B2(n10431), .ZN(
        P2_U3451) );
  INV_X1 U11457 ( .A(n10390), .ZN(n10394) );
  AOI22_X1 U11458 ( .A1(n10392), .A2(n10424), .B1(n10423), .B2(n10391), .ZN(
        n10393) );
  OAI211_X1 U11459 ( .C1(n10418), .C2(n10395), .A(n10394), .B(n10393), .ZN(
        n10396) );
  INV_X1 U11460 ( .A(n10396), .ZN(n10436) );
  INV_X1 U11461 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U11462 ( .A1(n10433), .A2(n10436), .B1(n10397), .B2(n10431), .ZN(
        P2_U3457) );
  OAI22_X1 U11463 ( .A1(n10401), .A2(n10400), .B1(n10399), .B2(n10398), .ZN(
        n10404) );
  INV_X1 U11464 ( .A(n10402), .ZN(n10403) );
  AOI211_X1 U11465 ( .C1(n8356), .C2(n10405), .A(n10404), .B(n10403), .ZN(
        n10437) );
  AOI22_X1 U11466 ( .A1(n10433), .A2(n10437), .B1(n10406), .B2(n10431), .ZN(
        P2_U3463) );
  AOI21_X1 U11467 ( .B1(n10423), .B2(n10408), .A(n10407), .ZN(n10409) );
  OAI211_X1 U11468 ( .C1(n10418), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        n10412) );
  INV_X1 U11469 ( .A(n10412), .ZN(n10438) );
  AOI22_X1 U11470 ( .A1(n10433), .A2(n10438), .B1(n10413), .B2(n10431), .ZN(
        P2_U3466) );
  AOI22_X1 U11471 ( .A1(n10415), .A2(n10424), .B1(n10423), .B2(n10414), .ZN(
        n10416) );
  OAI211_X1 U11472 ( .C1(n10419), .C2(n10418), .A(n10417), .B(n10416), .ZN(
        n10420) );
  INV_X1 U11473 ( .A(n10420), .ZN(n10440) );
  INV_X1 U11474 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U11475 ( .A1(n10433), .A2(n10440), .B1(n10421), .B2(n10431), .ZN(
        P2_U3469) );
  AOI22_X1 U11476 ( .A1(n10425), .A2(n10424), .B1(n10423), .B2(n4523), .ZN(
        n10426) );
  OAI211_X1 U11477 ( .C1(n10429), .C2(n10428), .A(n10427), .B(n10426), .ZN(
        n10430) );
  INV_X1 U11478 ( .A(n10430), .ZN(n10443) );
  INV_X1 U11479 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11480 ( .A1(n10433), .A2(n10443), .B1(n10432), .B2(n10431), .ZN(
        P2_U3475) );
  AOI22_X1 U11481 ( .A1(n10444), .A2(n10435), .B1(n10434), .B2(n10441), .ZN(
        P2_U3520) );
  AOI22_X1 U11482 ( .A1(n10444), .A2(n10436), .B1(n7093), .B2(n10441), .ZN(
        P2_U3522) );
  AOI22_X1 U11483 ( .A1(n10444), .A2(n10437), .B1(n7118), .B2(n10441), .ZN(
        P2_U3524) );
  AOI22_X1 U11484 ( .A1(n10444), .A2(n10438), .B1(n7121), .B2(n10441), .ZN(
        P2_U3525) );
  AOI22_X1 U11485 ( .A1(n10444), .A2(n10440), .B1(n10439), .B2(n10441), .ZN(
        P2_U3526) );
  AOI22_X1 U11486 ( .A1(n10444), .A2(n10443), .B1(n10442), .B2(n10441), .ZN(
        P2_U3528) );
  INV_X1 U11487 ( .A(n10445), .ZN(n10446) );
  NAND2_X1 U11488 ( .A1(n10447), .A2(n10446), .ZN(n10448) );
  XNOR2_X1 U11489 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10448), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11490 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11491 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(ADD_1071_U56) );
  OAI21_X1 U11492 ( .B1(n10454), .B2(n10453), .A(n10452), .ZN(ADD_1071_U57) );
  OAI21_X1 U11493 ( .B1(n10457), .B2(n10456), .A(n10455), .ZN(ADD_1071_U58) );
  OAI21_X1 U11494 ( .B1(n10460), .B2(n10459), .A(n10458), .ZN(ADD_1071_U59) );
  OAI21_X1 U11495 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(ADD_1071_U60) );
  OAI21_X1 U11496 ( .B1(n10466), .B2(n10465), .A(n10464), .ZN(ADD_1071_U61) );
  AOI21_X1 U11497 ( .B1(n10469), .B2(n10468), .A(n10467), .ZN(ADD_1071_U62) );
  AOI21_X1 U11498 ( .B1(n10472), .B2(n10471), .A(n10470), .ZN(ADD_1071_U63) );
  XOR2_X1 U11499 ( .A(n10473), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11500 ( .A1(n10475), .A2(n10474), .ZN(n10476) );
  XOR2_X1 U11501 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10476), .Z(ADD_1071_U51) );
  OAI21_X1 U11502 ( .B1(n10479), .B2(n10478), .A(n10477), .ZN(n10480) );
  XNOR2_X1 U11503 ( .A(n10480), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11504 ( .B1(n10483), .B2(n10482), .A(n10481), .ZN(ADD_1071_U47) );
  AOI21_X1 U11505 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(ADD_1071_U48) );
  NOR2_X1 U11506 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  XOR2_X1 U11507 ( .A(n10490), .B(n10489), .Z(ADD_1071_U49) );
  XOR2_X1 U11508 ( .A(n10492), .B(n10491), .Z(ADD_1071_U54) );
  XOR2_X1 U11509 ( .A(n10494), .B(n10493), .Z(ADD_1071_U53) );
  XNOR2_X1 U11510 ( .A(n10496), .B(n10495), .ZN(ADD_1071_U52) );
  INV_X1 U4880 ( .A(n8640), .ZN(n8874) );
  CLKBUF_X1 U4894 ( .A(n8969), .Z(n4374) );
  CLKBUF_X1 U4906 ( .A(n8976), .Z(n4387) );
  CLKBUF_X1 U4924 ( .A(n9363), .Z(n4386) );
endmodule

