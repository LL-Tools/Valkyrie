

module b21_C_AntiSAT_k_256_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4487, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347;

  INV_X4 U4991 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4992 ( .A(n9614), .ZN(n9396) );
  NAND2_X1 U4993 ( .A1(n5329), .A2(n5328), .ZN(n9798) );
  AND2_X4 U4995 ( .A1(n5930), .A2(n6826), .ZN(n6095) );
  INV_X1 U4996 ( .A(n6260), .ZN(n5507) );
  CLKBUF_X1 U4997 ( .A(n5257), .Z(n5259) );
  NOR2_X1 U4998 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5240) );
  OAI21_X1 U4999 ( .B1(n9752), .B2(n7903), .A(n7902), .ZN(n9733) );
  NOR2_X1 U5000 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5242) );
  OR2_X1 U5001 ( .A1(n7627), .A2(n7626), .ZN(n7796) );
  OR2_X1 U5002 ( .A1(n7422), .A2(n7421), .ZN(n7594) );
  NAND2_X2 U5004 ( .A1(n6411), .A2(n8408), .ZN(n6955) );
  NAND2_X1 U5005 ( .A1(n8326), .A2(n8327), .ZN(n9008) );
  NAND2_X1 U5006 ( .A1(n8911), .A2(n4489), .ZN(n8235) );
  NAND2_X1 U5007 ( .A1(n6603), .A2(n7279), .ZN(n7274) );
  INV_X1 U5008 ( .A(n10206), .ZN(n10249) );
  NAND2_X1 U5009 ( .A1(n9325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5014) );
  OR2_X1 U5010 ( .A1(n6063), .A2(n6062), .ZN(n9353) );
  OAI21_X1 U5011 ( .B1(n6739), .B2(n5568), .A(n4541), .ZN(n6834) );
  AND3_X1 U5012 ( .A1(n5512), .A2(n4778), .A3(n4777), .ZN(n10096) );
  INV_X2 U5013 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9872) );
  CLKBUF_X3 U5014 ( .A(n5554), .Z(n4493) );
  INV_X1 U5016 ( .A(n6907), .ZN(n4781) );
  NAND4_X4 U5017 ( .A1(n4986), .A2(n4985), .A3(n4983), .A4(n4982), .ZN(n6391)
         );
  OAI21_X2 U5018 ( .B1(n7258), .B2(n4894), .A(n4895), .ZN(n7668) );
  NAND2_X4 U5019 ( .A1(n4876), .A2(n4875), .ZN(n6554) );
  NAND2_X2 U5020 ( .A1(n4610), .A2(n4877), .ZN(n4876) );
  XNOR2_X2 U5021 ( .A(n4792), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5281) );
  OAI22_X2 U5022 ( .A1(n9998), .A2(n9997), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n9996), .ZN(n10009) );
  XNOR2_X2 U5023 ( .A(n5014), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6504) );
  XNOR2_X2 U5024 ( .A(n6335), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8357) );
  NOR2_X1 U5025 ( .A1(n5964), .A2(n6831), .ZN(n4487) );
  OAI22_X2 U5026 ( .A1(n7768), .A2(n4911), .B1(n4504), .B2(n7878), .ZN(n9756)
         );
  NAND2_X1 U5027 ( .A1(n5646), .A2(n5645), .ZN(n7535) );
  NAND2_X2 U5028 ( .A1(n5878), .A2(n5711), .ZN(n6816) );
  INV_X4 U5029 ( .A(n8116), .ZN(n8094) );
  NAND2_X1 U5030 ( .A1(n6391), .A2(n10092), .ZN(n5878) );
  INV_X1 U5031 ( .A(n6889), .ZN(n6887) );
  INV_X2 U5032 ( .A(n7191), .ZN(n4489) );
  INV_X4 U5033 ( .A(n8176), .ZN(n6602) );
  NAND2_X1 U5035 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U5036 ( .A(n4724), .B(n4723), .ZN(n9936) );
  NAND2_X1 U5037 ( .A1(n4997), .A2(n4521), .ZN(n9472) );
  AOI21_X1 U5038 ( .B1(n8412), .B2(n10194), .A(n8411), .ZN(n9223) );
  NOR2_X1 U5039 ( .A1(n5874), .A2(n9775), .ZN(n5865) );
  AOI21_X1 U5040 ( .B1(n9034), .B2(n9033), .A(n9032), .ZN(n9035) );
  OAI21_X1 U5041 ( .B1(n9024), .B2(n4901), .A(n4898), .ZN(n8163) );
  AND2_X1 U5042 ( .A1(n9553), .A2(n7894), .ZN(n9778) );
  OAI21_X1 U5043 ( .B1(n8806), .B2(n4964), .A(n4960), .ZN(n8868) );
  NAND2_X1 U5044 ( .A1(n6101), .A2(n6100), .ZN(n9460) );
  XNOR2_X1 U5045 ( .A(n8056), .B(n8039), .ZN(n8426) );
  NAND2_X1 U5046 ( .A1(n4892), .A2(n4526), .ZN(n9064) );
  NOR2_X1 U5047 ( .A1(n9624), .A2(n7915), .ZN(n9610) );
  OAI21_X1 U5048 ( .B1(n9637), .B2(n9638), .A(n7914), .ZN(n9624) );
  NAND3_X1 U5049 ( .A1(n5225), .A2(n4861), .A3(n5226), .ZN(n5230) );
  OR2_X1 U5050 ( .A1(n5277), .A2(n5274), .ZN(n5225) );
  OAI21_X1 U5051 ( .B1(n8789), .B2(n4605), .A(n4603), .ZN(n8033) );
  AOI21_X1 U5052 ( .B1(n8860), .B2(n8859), .A(n7971), .ZN(n8789) );
  NAND2_X2 U5053 ( .A1(n8078), .A2(n8077), .ZN(n9237) );
  INV_X1 U5054 ( .A(n4952), .ZN(n4605) );
  OAI21_X1 U5055 ( .B1(n8823), .B2(n8824), .A(n7958), .ZN(n8860) );
  AOI21_X1 U5056 ( .B1(n4952), .B2(n4604), .A(n4525), .ZN(n4603) );
  AOI21_X1 U5057 ( .B1(n4954), .B2(n4956), .A(n4953), .ZN(n4952) );
  AOI21_X2 U5058 ( .B1(n7695), .B2(n7694), .A(n7693), .ZN(n7768) );
  NAND2_X1 U5059 ( .A1(n5341), .A2(n5340), .ZN(n9812) );
  NAND2_X1 U5060 ( .A1(n4773), .A2(n4502), .ZN(n7406) );
  NAND2_X1 U5061 ( .A1(n8023), .A2(n8022), .ZN(n9255) );
  NAND2_X1 U5062 ( .A1(n7115), .A2(n7117), .ZN(n5001) );
  NAND2_X1 U5063 ( .A1(n6013), .A2(n6012), .ZN(n7116) );
  OAI21_X1 U5064 ( .B1(n5339), .B2(n5338), .A(n5188), .ZN(n5351) );
  OAI21_X1 U5065 ( .B1(n7212), .B2(n4973), .A(n4971), .ZN(n7588) );
  AND2_X1 U5066 ( .A1(n7517), .A2(n9920), .ZN(n7707) );
  NAND2_X1 U5067 ( .A1(n7624), .A2(n7623), .ZN(n9299) );
  AND2_X2 U5068 ( .A1(n7268), .A2(n10199), .ZN(n10210) );
  AND2_X1 U5069 ( .A1(n7062), .A2(n7061), .ZN(n10260) );
  NAND2_X1 U5070 ( .A1(n7216), .A2(n7215), .ZN(n7527) );
  INV_X1 U5071 ( .A(n10253), .ZN(n8229) );
  INV_X1 U5072 ( .A(n6980), .ZN(n6985) );
  AND3_X1 U5073 ( .A1(n4582), .A2(n5536), .A3(n5535), .ZN(n6980) );
  NAND2_X1 U5074 ( .A1(n6741), .A2(n4531), .ZN(n10206) );
  XNOR2_X1 U5075 ( .A(n5629), .B(n5628), .ZN(n6916) );
  NAND2_X2 U5076 ( .A1(n10064), .A2(n5934), .ZN(n6172) );
  NAND2_X1 U5077 ( .A1(n5545), .A2(n5544), .ZN(n5629) );
  NAND2_X2 U5078 ( .A1(n8912), .A2(n10228), .ZN(n7006) );
  NAND2_X1 U5079 ( .A1(n5530), .A2(n5529), .ZN(n5545) );
  NAND2_X1 U5080 ( .A1(n5101), .A2(n5100), .ZN(n5530) );
  AND4_X2 U5081 ( .A1(n6562), .A2(n6561), .A3(n6560), .A4(n6559), .ZN(n6995)
         );
  NAND2_X2 U5082 ( .A1(n6551), .A2(n6550), .ZN(n8116) );
  NAND4_X1 U5083 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n9493)
         );
  NAND2_X1 U5084 ( .A1(n8377), .A2(n7126), .ZN(n6978) );
  NAND4_X1 U5085 ( .A1(n5560), .A2(n5559), .A3(n5558), .A4(n5557), .ZN(n9495)
         );
  AND4_X1 U5086 ( .A1(n5952), .A2(n5953), .A3(n5954), .A4(n5951), .ZN(n10059)
         );
  NOR2_X2 U5087 ( .A1(n10052), .A2(n6828), .ZN(n10048) );
  INV_X1 U5088 ( .A(n5923), .ZN(n8377) );
  XNOR2_X1 U5089 ( .A(n5710), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5923) );
  BUF_X4 U5090 ( .A(n5552), .Z(n4492) );
  NAND2_X4 U5091 ( .A1(n6955), .A2(n6556), .ZN(n8167) );
  NAND2_X1 U5092 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5710) );
  AND2_X1 U5093 ( .A1(n5929), .A2(n7102), .ZN(n6826) );
  XNOR2_X1 U5094 ( .A(n5870), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5929) );
  INV_X1 U5095 ( .A(n9879), .ZN(n5280) );
  NAND2_X1 U5096 ( .A1(n4606), .A2(n4574), .ZN(n8408) );
  XNOR2_X1 U5097 ( .A(n5914), .B(n5913), .ZN(n7781) );
  NAND2_X1 U5098 ( .A1(n5707), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  AOI21_X1 U5099 ( .B1(n5259), .B2(n4518), .A(n4791), .ZN(n4790) );
  NAND2_X1 U5100 ( .A1(n6343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  XNOR2_X1 U5101 ( .A(n5102), .B(SI_5_), .ZN(n5529) );
  MUX2_X1 U5102 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5251), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5252) );
  AOI21_X1 U5103 ( .B1(n4495), .B2(P1_IR_REG_31__SCAN_IN), .A(n4766), .ZN(
        n4765) );
  NAND2_X2 U5104 ( .A1(n6316), .A2(P1_U3084), .ZN(n9881) );
  INV_X1 U5105 ( .A(n6252), .ZN(n6249) );
  NAND2_X2 U5106 ( .A1(n6554), .A2(P1_U3084), .ZN(n8383) );
  INV_X2 U5107 ( .A(n7385), .ZN(n4490) );
  AND2_X1 U5108 ( .A1(n4941), .A2(n8474), .ZN(n4834) );
  INV_X1 U5109 ( .A(n4944), .ZN(n4941) );
  NOR2_X1 U5110 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  NAND2_X1 U5111 ( .A1(n4609), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4875) );
  NOR2_X1 U5112 ( .A1(n4510), .A2(n5010), .ZN(n4836) );
  NAND2_X1 U5113 ( .A1(n4767), .A2(n5872), .ZN(n4766) );
  AND3_X1 U5114 ( .A1(n6307), .A2(n5036), .A3(n6231), .ZN(n4980) );
  AND2_X1 U5115 ( .A1(n5244), .A2(n5531), .ZN(n5245) );
  INV_X1 U5116 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6542) );
  INV_X1 U5117 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5410) );
  NOR2_X2 U5118 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6307) );
  INV_X4 U5119 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U5120 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5083) );
  NOR2_X1 U5121 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5036) );
  NAND2_X1 U5122 ( .A1(n5922), .A2(n5924), .ZN(n4491) );
  NOR2_X2 U5123 ( .A1(n9580), .A2(n9782), .ZN(n4789) );
  NAND2_X2 U5124 ( .A1(n7510), .A2(n7509), .ZN(n7695) );
  NOR3_X2 U5125 ( .A1(n9116), .A2(n4744), .A3(n9242), .ZN(n4746) );
  OR2_X2 U5126 ( .A1(n9140), .A2(n9260), .ZN(n9116) );
  XNOR2_X1 U5127 ( .A(n5530), .B(n5529), .ZN(n6838) );
  NAND2_X1 U5128 ( .A1(n7084), .A2(n7083), .ZN(n4917) );
  OAI21_X2 U5129 ( .B1(n7030), .B2(n7029), .A(n7028), .ZN(n7084) );
  AND2_X1 U5130 ( .A1(n5281), .A2(n5280), .ZN(n5552) );
  OAI211_X1 U5131 ( .C1(n6916), .C2(n5568), .A(n5551), .B(n5550), .ZN(n6907)
         );
  NOR3_X4 U5132 ( .A1(n9658), .A2(n4786), .A3(n9798), .ZN(n4788) );
  INV_X1 U5133 ( .A(n10052), .ZN(n10092) );
  NAND2_X1 U5134 ( .A1(n5281), .A2(n9879), .ZN(n5554) );
  NAND2_X1 U5135 ( .A1(n4616), .A2(n4615), .ZN(n4619) );
  NAND2_X1 U5136 ( .A1(n4617), .A2(n8329), .ZN(n4616) );
  NAND2_X1 U5137 ( .A1(n8325), .A2(n4519), .ZN(n4615) );
  NAND2_X1 U5138 ( .A1(n4620), .A2(n4624), .ZN(n4617) );
  NAND2_X1 U5139 ( .A1(n9150), .A2(n8392), .ZN(n5046) );
  INV_X1 U5140 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5035) );
  INV_X1 U5141 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6230) );
  AND2_X1 U5142 ( .A1(n5222), .A2(n5221), .ZN(n5226) );
  NOR2_X1 U5143 ( .A1(n4857), .A2(n4854), .ZN(n4853) );
  INV_X1 U5144 ( .A(n5125), .ZN(n4854) );
  INV_X1 U5145 ( .A(n4858), .ZN(n4857) );
  AND2_X1 U5146 ( .A1(n9217), .A2(n8172), .ZN(n8200) );
  INV_X1 U5147 ( .A(n6145), .ZN(n5000) );
  NAND2_X1 U5148 ( .A1(n5216), .A2(n5215), .ZN(n5302) );
  NAND2_X1 U5149 ( .A1(n5314), .A2(n5313), .ZN(n5216) );
  NAND2_X1 U5150 ( .A1(n5195), .A2(n5194), .ZN(n5683) );
  OAI21_X1 U5151 ( .B1(n5385), .B2(n5384), .A(n5174), .ZN(n5374) );
  OAI21_X1 U5152 ( .B1(n5475), .B2(n5474), .A(n5140), .ZN(n5458) );
  NAND2_X1 U5153 ( .A1(n4644), .A2(n4648), .ZN(n4643) );
  NAND2_X1 U5154 ( .A1(n5600), .A2(n5109), .ZN(n4838) );
  OR2_X1 U5155 ( .A1(n9267), .A2(n8790), .ZN(n8310) );
  NAND2_X1 U5156 ( .A1(n5106), .A2(n5105), .ZN(n5117) );
  NAND2_X1 U5157 ( .A1(n6549), .A2(n8220), .ZN(n6551) );
  NAND2_X1 U5158 ( .A1(n6730), .A2(n8349), .ZN(n6550) );
  OAI21_X1 U5159 ( .B1(n4618), .B2(n8336), .A(n4512), .ZN(n4612) );
  AOI21_X1 U5160 ( .B1(n4619), .B2(n4621), .A(n8328), .ZN(n4618) );
  OR2_X1 U5161 ( .A1(n9293), .A2(n7930), .ZN(n8287) );
  OR2_X1 U5162 ( .A1(n7743), .A2(n7750), .ZN(n8273) );
  OR2_X1 U5163 ( .A1(n7731), .A2(n7683), .ZN(n8265) );
  NOR2_X1 U5164 ( .A1(n5020), .A2(n4511), .ZN(n5018) );
  INV_X1 U5165 ( .A(n5021), .ZN(n5020) );
  AND2_X1 U5166 ( .A1(n5046), .A2(n4497), .ZN(n5043) );
  AND2_X1 U5167 ( .A1(n9273), .A2(n9168), .ZN(n5047) );
  AND2_X1 U5168 ( .A1(n6247), .A2(n6240), .ZN(n5064) );
  AND2_X1 U5169 ( .A1(n6307), .A2(n5036), .ZN(n4979) );
  AND2_X1 U5170 ( .A1(n6231), .A2(n6235), .ZN(n4981) );
  INV_X1 U5171 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U5172 ( .A1(n6046), .A2(n4995), .ZN(n4994) );
  OR2_X1 U5173 ( .A1(n9427), .A2(n5000), .ZN(n4999) );
  AND2_X1 U5174 ( .A1(n5791), .A2(n5273), .ZN(n5874) );
  OR2_X1 U5175 ( .A1(n9789), .A2(n6213), .ZN(n5809) );
  AND2_X1 U5176 ( .A1(n4935), .A2(n4552), .ZN(n4932) );
  INV_X1 U5177 ( .A(n4800), .ZN(n4799) );
  OR2_X1 U5178 ( .A1(n9741), .A2(n9754), .ZN(n5853) );
  NOR2_X1 U5179 ( .A1(n7301), .A2(n4928), .ZN(n4927) );
  INV_X1 U5180 ( .A(n7299), .ZN(n4928) );
  NAND2_X1 U5181 ( .A1(n4916), .A2(n7697), .ZN(n4911) );
  NAND2_X1 U5182 ( .A1(n5229), .A2(n5230), .ZN(n5266) );
  NAND2_X1 U5183 ( .A1(n5224), .A2(n5223), .ZN(n5277) );
  NAND2_X1 U5184 ( .A1(n4864), .A2(n4862), .ZN(n5314) );
  AOI21_X1 U5185 ( .B1(n4866), .B2(n4869), .A(n4863), .ZN(n4862) );
  INV_X1 U5186 ( .A(n5209), .ZN(n4863) );
  NAND2_X1 U5187 ( .A1(n5915), .A2(n5011), .ZN(n5010) );
  NAND2_X1 U5188 ( .A1(n5169), .A2(n5168), .ZN(n5385) );
  NAND2_X1 U5189 ( .A1(n5161), .A2(n5160), .ZN(n5408) );
  NAND2_X1 U5190 ( .A1(n4844), .A2(n4842), .ZN(n5161) );
  AOI21_X1 U5191 ( .B1(n4845), .B2(n4506), .A(n4843), .ZN(n4842) );
  AND2_X1 U5192 ( .A1(n5160), .A2(n5159), .ZN(n5426) );
  NAND2_X1 U5193 ( .A1(n5154), .A2(n5153), .ZN(n5660) );
  XNOR2_X1 U5194 ( .A(n5147), .B(SI_14_), .ZN(n5442) );
  NAND2_X1 U5195 ( .A1(n5458), .A2(n5082), .ZN(n5146) );
  AOI21_X1 U5196 ( .B1(n4858), .B2(n4856), .A(n4545), .ZN(n4855) );
  NAND2_X1 U5197 ( .A1(n5140), .A2(n5139), .ZN(n5474) );
  NOR2_X1 U5198 ( .A1(n6555), .A2(n6316), .ZN(n4748) );
  AOI21_X1 U5199 ( .B1(n7588), .B2(n7587), .A(n7586), .ZN(n7589) );
  INV_X1 U5200 ( .A(n7322), .ZN(n6626) );
  AOI21_X1 U5201 ( .B1(n8173), .B2(n8337), .A(n8200), .ZN(n8174) );
  OAI22_X1 U5202 ( .A1(n8163), .A2(n8199), .B1(n8349), .B2(n8982), .ZN(n8164)
         );
  OR2_X1 U5203 ( .A1(n9217), .A2(n8172), .ZN(n8341) );
  INV_X1 U5205 ( .A(n8046), .ZN(n8162) );
  AND4_X1 U5206 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n7003)
         );
  OR2_X1 U5207 ( .A1(n6470), .A2(n6469), .ZN(n4701) );
  AOI21_X1 U5208 ( .B1(n10178), .B2(n10179), .A(n8972), .ZN(n8973) );
  OR2_X1 U5209 ( .A1(n9242), .A2(n9069), .ZN(n8206) );
  OR2_X1 U5210 ( .A1(n9255), .A2(n9094), .ZN(n9089) );
  NAND2_X1 U5211 ( .A1(n5067), .A2(n5065), .ZN(n9174) );
  AND2_X1 U5212 ( .A1(n9177), .A2(n5066), .ZN(n5065) );
  INV_X1 U5213 ( .A(n8389), .ZN(n5066) );
  OR2_X1 U5214 ( .A1(n9293), .A2(n9196), .ZN(n8387) );
  OR2_X1 U5215 ( .A1(n7743), .A2(n8901), .ZN(n5062) );
  INV_X1 U5216 ( .A(n8167), .ZN(n7974) );
  INV_X1 U5217 ( .A(n6955), .ZN(n7973) );
  NAND2_X1 U5218 ( .A1(n6955), .A2(n6554), .ZN(n6957) );
  XNOR2_X1 U5219 ( .A(n6368), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U5220 ( .A1(n6367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U5221 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n4949) );
  NAND2_X1 U5222 ( .A1(n6540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U5223 ( .A1(n9472), .A2(n6162), .ZN(n6169) );
  XNOR2_X1 U5224 ( .A(n5975), .B(n5992), .ZN(n5977) );
  XNOR2_X1 U5225 ( .A(n5935), .B(n6172), .ZN(n5947) );
  NOR2_X1 U5226 ( .A1(n5807), .A2(n5898), .ZN(n7921) );
  NOR2_X1 U5227 ( .A1(n9559), .A2(n9567), .ZN(n9558) );
  AND2_X1 U5228 ( .A1(n9803), .A2(n9640), .ZN(n7892) );
  OR2_X1 U5229 ( .A1(n9823), .A2(n9388), .ZN(n7909) );
  INV_X1 U5230 ( .A(n4920), .ZN(n4919) );
  NAND2_X1 U5231 ( .A1(n9716), .A2(n9722), .ZN(n9717) );
  OR2_X1 U5232 ( .A1(n5258), .A2(n9872), .ZN(n4792) );
  XNOR2_X1 U5233 ( .A(n5292), .B(n5291), .ZN(n8075) );
  NAND2_X1 U5234 ( .A1(n4865), .A2(n4871), .ZN(n5292) );
  NAND2_X1 U5235 ( .A1(n5683), .A2(n4873), .ZN(n4865) );
  XNOR2_X1 U5236 ( .A(n5327), .B(n5326), .ZN(n8062) );
  NAND2_X1 U5237 ( .A1(n4870), .A2(n5198), .ZN(n5327) );
  INV_X1 U5238 ( .A(n6549), .ZN(n8352) );
  OAI22_X2 U5239 ( .A1(n9437), .A2(n6114), .B1(n9435), .B2(n9434), .ZN(n9384)
         );
  OAI21_X1 U5240 ( .B1(n5722), .B2(n4654), .A(n4653), .ZN(n5721) );
  OR2_X1 U5241 ( .A1(n4655), .A2(n5720), .ZN(n4654) );
  AOI21_X1 U5242 ( .B1(n4546), .B2(n7291), .A(n5792), .ZN(n4653) );
  NOR2_X1 U5243 ( .A1(n4668), .A2(n5842), .ZN(n4667) );
  INV_X1 U5244 ( .A(n5733), .ZN(n4668) );
  NAND2_X1 U5245 ( .A1(n8241), .A2(n8237), .ZN(n4633) );
  NAND2_X1 U5246 ( .A1(n4631), .A2(n4630), .ZN(n4629) );
  INV_X1 U5247 ( .A(n8247), .ZN(n4631) );
  NOR2_X1 U5248 ( .A1(n4533), .A2(n4640), .ZN(n4638) );
  INV_X1 U5249 ( .A(n4640), .ZN(n4639) );
  NAND2_X1 U5250 ( .A1(n4969), .A2(n8352), .ZN(n4968) );
  INV_X1 U5251 ( .A(n8311), .ZN(n4646) );
  NOR2_X1 U5252 ( .A1(n4647), .A2(n4530), .ZN(n4644) );
  NAND2_X1 U5253 ( .A1(n8309), .A2(n8310), .ZN(n4647) );
  NOR2_X1 U5254 ( .A1(n5865), .A2(n5863), .ZN(n4676) );
  NAND2_X1 U5255 ( .A1(n4681), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U5256 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U5257 ( .A1(n5789), .A2(n5790), .ZN(n4681) );
  NOR2_X1 U5258 ( .A1(n7896), .A2(n5792), .ZN(n4679) );
  INV_X1 U5259 ( .A(n4954), .ZN(n4604) );
  NAND2_X1 U5260 ( .A1(n8407), .A2(n4903), .ZN(n4901) );
  INV_X1 U5261 ( .A(n4901), .ZN(n4900) );
  NAND2_X1 U5262 ( .A1(n5302), .A2(n5301), .ZN(n5224) );
  NOR2_X1 U5263 ( .A1(n5135), .A2(n4859), .ZN(n4858) );
  INV_X1 U5264 ( .A(n5132), .ZN(n4859) );
  NOR2_X1 U5265 ( .A1(n8842), .A2(n4958), .ZN(n4957) );
  INV_X1 U5266 ( .A(n7991), .ZN(n4958) );
  NOR2_X1 U5267 ( .A1(n6995), .A2(n6602), .ZN(n6566) );
  AND2_X1 U5268 ( .A1(n4623), .A2(n4619), .ZN(n4614) );
  NAND2_X1 U5269 ( .A1(n9001), .A2(n8330), .ZN(n4903) );
  AND2_X1 U5270 ( .A1(n8330), .A2(n8326), .ZN(n4904) );
  OR2_X1 U5271 ( .A1(n9237), .A2(n9021), .ZN(n8322) );
  OR2_X1 U5272 ( .A1(n9247), .A2(n9093), .ZN(n8319) );
  NAND2_X1 U5273 ( .A1(n9252), .A2(n8395), .ZN(n8396) );
  NOR2_X1 U5274 ( .A1(n5031), .A2(n5027), .ZN(n5024) );
  AND2_X1 U5275 ( .A1(n8319), .A2(n8318), .ZN(n8397) );
  OR2_X1 U5276 ( .A1(n9252), .A2(n9108), .ZN(n8315) );
  NAND2_X1 U5277 ( .A1(n8388), .A2(n5068), .ZN(n5067) );
  NOR2_X1 U5278 ( .A1(n9202), .A2(n5069), .ZN(n5068) );
  INV_X1 U5279 ( .A(n8387), .ZN(n5069) );
  OR2_X1 U5280 ( .A1(n9287), .A2(n9181), .ZN(n8290) );
  OR2_X1 U5281 ( .A1(n7849), .A2(n7832), .ZN(n8282) );
  OR2_X1 U5282 ( .A1(n7663), .A2(n7433), .ZN(n8254) );
  NAND2_X1 U5283 ( .A1(n7250), .A2(n7249), .ZN(n5071) );
  NAND2_X1 U5284 ( .A1(n8240), .A2(n7009), .ZN(n4883) );
  INV_X1 U5285 ( .A(n8240), .ZN(n4884) );
  NAND2_X1 U5286 ( .A1(n7174), .A2(n8908), .ZN(n8242) );
  AND2_X1 U5287 ( .A1(n8976), .A2(n8354), .ZN(n6730) );
  NAND3_X1 U5288 ( .A1(n4979), .A2(n4543), .A3(n4981), .ZN(n4978) );
  NAND2_X1 U5289 ( .A1(n4754), .A2(n4752), .ZN(n6134) );
  AOI21_X1 U5290 ( .B1(n9448), .B2(n4762), .A(n4753), .ZN(n4752) );
  NAND2_X1 U5291 ( .A1(n9384), .A2(n4755), .ZN(n4754) );
  AND2_X1 U5292 ( .A1(n4756), .A2(n9382), .ZN(n4753) );
  NAND2_X1 U5293 ( .A1(n5930), .A2(n5934), .ZN(n5964) );
  NOR2_X1 U5294 ( .A1(n5989), .A2(n4771), .ZN(n4770) );
  INV_X1 U5295 ( .A(n5981), .ZN(n4771) );
  AND2_X1 U5296 ( .A1(n4710), .A2(n4709), .ZN(n6270) );
  NAND2_X1 U5297 ( .A1(n7342), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4709) );
  INV_X1 U5298 ( .A(n5809), .ZN(n7919) );
  OR2_X1 U5299 ( .A1(n9782), .A2(n9340), .ZN(n5805) );
  NAND2_X1 U5300 ( .A1(n9782), .A2(n9340), .ZN(n7920) );
  AOI21_X1 U5301 ( .B1(n4810), .B2(n7916), .A(n5802), .ZN(n4808) );
  AND2_X1 U5302 ( .A1(n5760), .A2(n7909), .ZN(n4801) );
  AND2_X1 U5303 ( .A1(n9828), .A2(n9440), .ZN(n5857) );
  OR2_X1 U5304 ( .A1(n9832), .A2(n9420), .ZN(n5755) );
  NOR2_X1 U5305 ( .A1(n7708), .A2(n9357), .ZN(n4783) );
  OR2_X1 U5306 ( .A1(n9357), .A2(n9753), .ZN(n7900) );
  NAND2_X1 U5307 ( .A1(n9496), .A2(n10096), .ZN(n5880) );
  INV_X1 U5308 ( .A(n6826), .ZN(n5934) );
  NAND2_X1 U5309 ( .A1(n5250), .A2(n4945), .ZN(n4944) );
  OAI21_X1 U5310 ( .B1(n5408), .B2(n5165), .A(n5164), .ZN(n5396) );
  INV_X1 U5311 ( .A(n5149), .ZN(n4847) );
  INV_X1 U5312 ( .A(n4846), .ZN(n4845) );
  OAI21_X1 U5313 ( .B1(n4849), .B2(n4506), .A(n5154), .ZN(n4846) );
  NOR2_X1 U5314 ( .A1(n5150), .A2(n4850), .ZN(n4849) );
  INV_X1 U5315 ( .A(n5145), .ZN(n4850) );
  INV_X1 U5316 ( .A(n5442), .ZN(n5150) );
  XNOR2_X1 U5317 ( .A(n5133), .B(SI_11_), .ZN(n5640) );
  AND2_X1 U5318 ( .A1(n5132), .A2(n5131), .ZN(n5077) );
  NAND2_X1 U5319 ( .A1(n5120), .A2(n5119), .ZN(n5581) );
  NOR2_X1 U5320 ( .A1(n5074), .A2(n5118), .ZN(n5119) );
  AOI21_X1 U5321 ( .B1(n5110), .B2(n5545), .A(n4837), .ZN(n5120) );
  XNOR2_X1 U5322 ( .A(n5114), .B(SI_7_), .ZN(n5632) );
  NAND2_X1 U5323 ( .A1(n6547), .A2(n5520), .ZN(n5086) );
  OR2_X1 U5324 ( .A1(n8080), .A2(n8079), .ZN(n8106) );
  INV_X1 U5325 ( .A(n6932), .ZN(n6625) );
  NAND2_X1 U5326 ( .A1(n4951), .A2(n4584), .ZN(n6928) );
  AND2_X1 U5327 ( .A1(n4950), .A2(n6850), .ZN(n4584) );
  NAND2_X1 U5328 ( .A1(n6754), .A2(n6847), .ZN(n4950) );
  XNOR2_X1 U5329 ( .A(n10206), .B(n8094), .ZN(n4593) );
  NAND2_X1 U5330 ( .A1(n6744), .A2(n4593), .ZN(n6847) );
  OR2_X1 U5331 ( .A1(n6753), .A2(n6754), .ZN(n6848) );
  OR2_X1 U5332 ( .A1(n7064), .A2(n7063), .ZN(n7226) );
  NAND2_X1 U5333 ( .A1(n7212), .A2(n4508), .ZN(n7315) );
  OR2_X1 U5334 ( .A1(n7226), .A2(n7225), .ZN(n7322) );
  OR2_X1 U5335 ( .A1(n8808), .A2(n4966), .ZN(n4965) );
  INV_X1 U5336 ( .A(n8807), .ZN(n4966) );
  INV_X1 U5337 ( .A(n8121), .ZN(n8158) );
  AND4_X1 U5338 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(n8790)
         );
  AND4_X1 U5339 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n8230)
         );
  XNOR2_X1 U5340 ( .A(n8376), .B(n4688), .ZN(n8366) );
  NOR2_X1 U5341 ( .A1(n6431), .A2(n4704), .ZN(n6444) );
  AND2_X1 U5342 ( .A1(n6413), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4704) );
  OR2_X1 U5343 ( .A1(n6444), .A2(n6443), .ZN(n4703) );
  NOR2_X1 U5344 ( .A1(n6418), .A2(n6417), .ZN(n6454) );
  AND2_X1 U5345 ( .A1(n4701), .A2(n4700), .ZN(n6460) );
  NAND2_X1 U5346 ( .A1(n6457), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4700) );
  OR2_X1 U5347 ( .A1(n6460), .A2(n6459), .ZN(n4699) );
  NOR2_X1 U5348 ( .A1(n7198), .A2(n4568), .ZN(n7200) );
  NOR2_X1 U5349 ( .A1(n7200), .A2(n7199), .ZN(n7474) );
  OR2_X1 U5350 ( .A1(n9230), .A2(n9036), .ZN(n8326) );
  NAND2_X1 U5351 ( .A1(n9237), .A2(n9021), .ZN(n9019) );
  NOR2_X2 U5352 ( .A1(n9237), .A2(n9048), .ZN(n9037) );
  NAND2_X1 U5353 ( .A1(n8322), .A2(n9019), .ZN(n9034) );
  INV_X1 U5354 ( .A(n9045), .ZN(n9055) );
  NAND2_X1 U5355 ( .A1(n9056), .A2(n9055), .ZN(n9054) );
  INV_X1 U5356 ( .A(n8027), .ZN(n6631) );
  NAND2_X1 U5357 ( .A1(n4551), .A2(n4498), .ZN(n5028) );
  NAND2_X1 U5358 ( .A1(n9089), .A2(n8311), .ZN(n9106) );
  AND2_X1 U5359 ( .A1(n9166), .A2(n8295), .ZN(n4908) );
  OR2_X1 U5360 ( .A1(n9178), .A2(n9177), .ZN(n4909) );
  AND2_X1 U5361 ( .A1(n8298), .A2(n8304), .ZN(n9166) );
  INV_X1 U5362 ( .A(n5067), .ZN(n9200) );
  OR2_X1 U5363 ( .A1(n7849), .A2(n8899), .ZN(n5059) );
  NAND2_X1 U5364 ( .A1(n5052), .A2(n5058), .ZN(n5050) );
  OR2_X1 U5365 ( .A1(n7744), .A2(n5053), .ZN(n5051) );
  AOI21_X1 U5366 ( .B1(n5057), .B2(n8190), .A(n5060), .ZN(n5056) );
  NAND2_X1 U5367 ( .A1(n6627), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7627) );
  OR2_X1 U5368 ( .A1(n7744), .A2(n8190), .ZN(n5063) );
  OAI21_X1 U5369 ( .B1(n7748), .B2(n7747), .A(n8272), .ZN(n7749) );
  NAND2_X1 U5370 ( .A1(n7577), .A2(n7576), .ZN(n7743) );
  NOR2_X2 U5371 ( .A1(n7671), .A2(n7731), .ZN(n7684) );
  AOI21_X1 U5372 ( .B1(n8250), .B2(n4897), .A(n4896), .ZN(n4895) );
  NAND2_X1 U5373 ( .A1(n8259), .A2(n8250), .ZN(n4894) );
  INV_X1 U5374 ( .A(n8262), .ZN(n4896) );
  NAND2_X1 U5375 ( .A1(n4885), .A2(n8247), .ZN(n7256) );
  NAND2_X1 U5376 ( .A1(n7346), .A2(n8182), .ZN(n4885) );
  NOR2_X1 U5377 ( .A1(n7158), .A2(n5022), .ZN(n5021) );
  INV_X1 U5378 ( .A(n7004), .ZN(n5022) );
  NAND2_X1 U5379 ( .A1(n4733), .A2(n4732), .ZN(n7351) );
  INV_X1 U5380 ( .A(n4734), .ZN(n4732) );
  NAND2_X1 U5381 ( .A1(n8909), .A2(n10249), .ZN(n8240) );
  NAND2_X1 U5382 ( .A1(n7146), .A2(n8225), .ZN(n7008) );
  OR2_X1 U5383 ( .A1(n7142), .A2(n7141), .ZN(n7268) );
  OR2_X1 U5384 ( .A1(n10258), .A2(n8220), .ZN(n6725) );
  INV_X1 U5385 ( .A(n9892), .ZN(n4729) );
  NAND2_X1 U5386 ( .A1(n8155), .A2(n8154), .ZN(n9220) );
  NAND2_X1 U5387 ( .A1(n5037), .A2(n5039), .ZN(n9265) );
  AND2_X1 U5388 ( .A1(n5040), .A2(n9133), .ZN(n5039) );
  NAND2_X1 U5389 ( .A1(n5041), .A2(n5042), .ZN(n5040) );
  NAND2_X1 U5390 ( .A1(n7794), .A2(n7793), .ZN(n9293) );
  AND2_X1 U5391 ( .A1(n7313), .A2(n8349), .ZN(n7011) );
  AND2_X1 U5392 ( .A1(n5073), .A2(n6248), .ZN(n5072) );
  NOR2_X1 U5393 ( .A1(n6341), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U5394 ( .A1(n6249), .A2(n4735), .ZN(n6343) );
  NOR2_X1 U5395 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(n6341), .ZN(n4735) );
  INV_X1 U5396 ( .A(n6343), .ZN(n4576) );
  NOR2_X1 U5397 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4575) );
  NAND2_X1 U5398 ( .A1(n6249), .A2(n4910), .ZN(n6338) );
  AND2_X1 U5399 ( .A1(n6248), .A2(n6339), .ZN(n4910) );
  NAND2_X1 U5400 ( .A1(n4566), .A2(n5033), .ZN(n6385) );
  AND2_X1 U5401 ( .A1(n6334), .A2(n6352), .ZN(n6670) );
  NAND2_X1 U5402 ( .A1(n6784), .A2(n5004), .ZN(n5003) );
  INV_X1 U5403 ( .A(n6783), .ZN(n5004) );
  AOI21_X1 U5404 ( .B1(n4496), .B2(n4993), .A(n4988), .ZN(n4987) );
  INV_X1 U5405 ( .A(n7655), .ZN(n4988) );
  INV_X1 U5406 ( .A(n6717), .ZN(n4772) );
  NAND2_X1 U5407 ( .A1(n4572), .A2(n5001), .ZN(n7128) );
  AND2_X1 U5408 ( .A1(n9381), .A2(n4757), .ZN(n4756) );
  INV_X1 U5409 ( .A(n6129), .ZN(n4757) );
  NAND2_X1 U5410 ( .A1(n4763), .A2(n6129), .ZN(n4762) );
  NAND2_X1 U5411 ( .A1(n9382), .A2(n9381), .ZN(n4763) );
  AND2_X1 U5412 ( .A1(n6120), .A2(n6121), .ZN(n9382) );
  INV_X1 U5413 ( .A(n6024), .ZN(n4775) );
  AND2_X1 U5414 ( .A1(n6023), .A2(n7369), .ZN(n4776) );
  INV_X1 U5415 ( .A(n6391), .ZN(n6817) );
  AND3_X1 U5416 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5537) );
  INV_X1 U5417 ( .A(n9471), .ZN(n6157) );
  NAND2_X1 U5418 ( .A1(n5867), .A2(n6991), .ZN(n4665) );
  OR2_X1 U5419 ( .A1(n5693), .A2(n5523), .ZN(n5526) );
  NAND2_X1 U5420 ( .A1(n4492), .A2(n6719), .ZN(n5492) );
  NAND2_X1 U5421 ( .A1(n5524), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4982) );
  XNOR2_X1 U5422 ( .A(n9936), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9941) );
  OR2_X1 U5423 ( .A1(n9952), .A2(n9951), .ZN(n4714) );
  NAND2_X1 U5424 ( .A1(n4714), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U5425 ( .A1(n9946), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4713) );
  AOI21_X1 U5426 ( .B1(n6288), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7108), .ZN(
        n7340) );
  OR2_X1 U5427 ( .A1(n7340), .A2(n7339), .ZN(n4710) );
  XNOR2_X1 U5428 ( .A(n6270), .B(n7720), .ZN(n7722) );
  NOR2_X1 U5429 ( .A1(n7722), .A2(n5453), .ZN(n7721) );
  NAND2_X1 U5430 ( .A1(n4789), .A2(n7896), .ZN(n9553) );
  NAND2_X1 U5431 ( .A1(n9610), .A2(n4810), .ZN(n4807) );
  OR2_X1 U5432 ( .A1(n9798), .A2(n5337), .ZN(n9594) );
  INV_X1 U5433 ( .A(n4936), .ZN(n4935) );
  OAI22_X1 U5434 ( .A1(n9612), .A2(n4940), .B1(n9798), .B2(n9627), .ZN(n4936)
         );
  NAND2_X1 U5435 ( .A1(n4939), .A2(n4938), .ZN(n4937) );
  INV_X1 U5436 ( .A(n7892), .ZN(n4938) );
  INV_X1 U5437 ( .A(n9612), .ZN(n4939) );
  AND2_X1 U5438 ( .A1(n9594), .A2(n5773), .ZN(n9612) );
  NAND2_X1 U5439 ( .A1(n9623), .A2(n9398), .ZN(n4940) );
  INV_X1 U5440 ( .A(n4798), .ZN(n4797) );
  OAI21_X1 U5441 ( .B1(n4801), .B2(n4799), .A(n9651), .ZN(n4798) );
  OR2_X1 U5442 ( .A1(n9678), .A2(n4799), .ZN(n4793) );
  NAND2_X1 U5443 ( .A1(n4550), .A2(n5760), .ZN(n4800) );
  NAND2_X1 U5444 ( .A1(n7910), .A2(n7909), .ZN(n4803) );
  NOR2_X1 U5445 ( .A1(n5759), .A2(n7913), .ZN(n9651) );
  NOR2_X1 U5446 ( .A1(n4926), .A2(n7883), .ZN(n4925) );
  AOI21_X1 U5447 ( .B1(n4924), .B2(n4509), .A(n4923), .ZN(n4922) );
  NOR2_X1 U5448 ( .A1(n9722), .A2(n9465), .ZN(n4923) );
  INV_X1 U5449 ( .A(n7883), .ZN(n4924) );
  AND2_X1 U5450 ( .A1(n5753), .A2(n9705), .ZN(n9723) );
  OR2_X1 U5451 ( .A1(n9842), .A2(n9408), .ZN(n5079) );
  OR2_X1 U5452 ( .A1(n9760), .A2(n9736), .ZN(n4915) );
  NAND2_X1 U5453 ( .A1(n9733), .A2(n4926), .ZN(n9732) );
  NAND2_X1 U5454 ( .A1(n4783), .A2(n9842), .ZN(n9763) );
  AND2_X1 U5455 ( .A1(n7704), .A2(n7703), .ZN(n4822) );
  INV_X1 U5456 ( .A(n7879), .ZN(n7704) );
  AND2_X1 U5457 ( .A1(n7764), .A2(n7703), .ZN(n5076) );
  AND2_X1 U5458 ( .A1(n5726), .A2(n7703), .ZN(n7767) );
  NAND2_X1 U5459 ( .A1(n7765), .A2(n7767), .ZN(n7764) );
  NAND2_X1 U5460 ( .A1(n4929), .A2(n4523), .ZN(n7510) );
  AND2_X1 U5461 ( .A1(n5823), .A2(n5827), .ZN(n6986) );
  NAND2_X1 U5462 ( .A1(n5880), .A2(n5713), .ZN(n6871) );
  OAI211_X2 U5463 ( .C1(n6555), .C2(n5568), .A(n4780), .B(n4779), .ZN(n10052)
         );
  NAND2_X1 U5464 ( .A1(n5507), .A2(n9936), .ZN(n4779) );
  NAND2_X1 U5465 ( .A1(n6482), .A2(n5933), .ZN(n10064) );
  AOI21_X1 U5466 ( .B1(n8377), .B2(n5934), .A(n10054), .ZN(n5933) );
  NAND2_X1 U5467 ( .A1(n5464), .A2(n5463), .ZN(n9848) );
  OAI21_X1 U5468 ( .B1(n5266), .B2(SI_30_), .A(n5230), .ZN(n5234) );
  NAND2_X1 U5469 ( .A1(n4851), .A2(n5179), .ZN(n5363) );
  NAND2_X1 U5470 ( .A1(n5146), .A2(n5145), .ZN(n5443) );
  XNOR2_X1 U5471 ( .A(n5641), .B(n5640), .ZN(n7418) );
  NAND2_X1 U5472 ( .A1(n4860), .A2(n5132), .ZN(n5641) );
  NAND2_X1 U5473 ( .A1(n5570), .A2(n5077), .ZN(n4860) );
  NAND2_X1 U5474 ( .A1(n5494), .A2(n4608), .ZN(n5101) );
  NAND2_X1 U5475 ( .A1(n8420), .A2(n8419), .ZN(n8418) );
  NOR2_X1 U5476 ( .A1(n8119), .A2(n4589), .ZN(n4586) );
  NAND2_X1 U5477 ( .A1(n8104), .A2(n8103), .ZN(n9226) );
  NAND2_X1 U5478 ( .A1(n8361), .A2(n8153), .ZN(n8104) );
  NAND2_X1 U5479 ( .A1(n5075), .A2(n4747), .ZN(n7278) );
  OAI21_X1 U5480 ( .B1(n4748), .B2(n4749), .A(n6955), .ZN(n4747) );
  AND2_X1 U5481 ( .A1(n6556), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4749) );
  INV_X1 U5482 ( .A(n9118), .ZN(n9260) );
  NAND2_X1 U5483 ( .A1(n8061), .A2(n8060), .ZN(n8806) );
  NAND2_X1 U5484 ( .A1(n8064), .A2(n8063), .ZN(n9242) );
  NAND2_X1 U5485 ( .A1(n8062), .A2(n8153), .ZN(n8064) );
  INV_X1 U5486 ( .A(n4972), .ZN(n4971) );
  OAI21_X1 U5487 ( .B1(n4973), .B2(n4508), .A(n7415), .ZN(n4972) );
  AND2_X1 U5488 ( .A1(n8073), .A2(n8072), .ZN(n9069) );
  NOR2_X1 U5489 ( .A1(n4573), .A2(n8360), .ZN(n4888) );
  OR2_X1 U5490 ( .A1(n8359), .A2(n8358), .ZN(n4889) );
  AOI21_X1 U5491 ( .B1(n8347), .B2(n8346), .A(n8345), .ZN(n8351) );
  INV_X1 U5492 ( .A(n7011), .ZN(n8354) );
  NOR2_X1 U5493 ( .A1(n8915), .A2(n4705), .ZN(n6669) );
  AND2_X1 U5494 ( .A1(n6956), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4705) );
  NOR2_X1 U5495 ( .A1(n6669), .A2(n6668), .ZN(n6770) );
  NAND2_X1 U5496 ( .A1(n4695), .A2(n4532), .ZN(n4692) );
  NAND2_X1 U5497 ( .A1(n8974), .A2(n10181), .ZN(n4695) );
  AND2_X1 U5498 ( .A1(n10170), .A2(n9188), .ZN(n4693) );
  OAI21_X1 U5499 ( .B1(n8974), .B2(n10171), .A(n4697), .ZN(n4696) );
  AOI21_X1 U5500 ( .B1(n8975), .B2(n10185), .A(n9188), .ZN(n4697) );
  AOI21_X1 U5501 ( .B1(n8380), .B2(n8153), .A(n8156), .ZN(n8987) );
  NAND2_X1 U5502 ( .A1(n8985), .A2(n4730), .ZN(n9892) );
  OR2_X1 U5503 ( .A1(n8986), .A2(n8987), .ZN(n4730) );
  NAND2_X1 U5504 ( .A1(n7948), .A2(n7947), .ZN(n9284) );
  NAND2_X1 U5505 ( .A1(n4890), .A2(n4520), .ZN(n7191) );
  INV_X1 U5506 ( .A(n4891), .ZN(n4890) );
  NOR2_X1 U5507 ( .A1(n4947), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U5508 ( .A1(n5316), .A2(n5315), .ZN(n9789) );
  NAND2_X1 U5509 ( .A1(n8091), .A2(n5303), .ZN(n5316) );
  INV_X1 U5510 ( .A(n9494), .ZN(n6898) );
  NAND2_X1 U5511 ( .A1(n7406), .A2(n7407), .ZN(n4996) );
  NAND2_X1 U5512 ( .A1(n5433), .A2(n5432), .ZN(n9741) );
  NAND2_X1 U5513 ( .A1(n5686), .A2(n5685), .ZN(n9803) );
  NAND2_X1 U5514 ( .A1(n5376), .A2(n5375), .ZN(n9823) );
  OR2_X1 U5515 ( .A1(n7406), .A2(n4993), .ZN(n4990) );
  NAND2_X1 U5516 ( .A1(n5294), .A2(n5293), .ZN(n9792) );
  NAND2_X1 U5517 ( .A1(n8075), .A2(n5303), .ZN(n5294) );
  OR2_X1 U5518 ( .A1(n5556), .A2(n5513), .ZN(n5515) );
  OR2_X1 U5519 ( .A1(n4493), .A2(n10077), .ZN(n5514) );
  AND2_X1 U5520 ( .A1(n4707), .A2(n4706), .ZN(n10007) );
  NAND2_X1 U5521 ( .A1(n9996), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4706) );
  NOR2_X1 U5522 ( .A1(n7110), .A2(n7109), .ZN(n7108) );
  NOR2_X1 U5523 ( .A1(n9558), .A2(n4581), .ZN(n7893) );
  AND2_X1 U5524 ( .A1(n9782), .A2(n9576), .ZN(n4581) );
  AOI21_X1 U5525 ( .B1(n4828), .B2(n10061), .A(n4825), .ZN(n9780) );
  NAND2_X1 U5526 ( .A1(n4827), .A2(n4826), .ZN(n4825) );
  XNOR2_X1 U5527 ( .A(n4829), .B(n7921), .ZN(n4828) );
  NAND2_X1 U5528 ( .A1(n8132), .A2(n9483), .ZN(n4826) );
  NAND2_X1 U5529 ( .A1(n4658), .A2(n5843), .ZN(n4656) );
  INV_X1 U5530 ( .A(n5844), .ZN(n4657) );
  INV_X1 U5531 ( .A(n7291), .ZN(n4655) );
  NAND2_X1 U5532 ( .A1(n4660), .A2(n4659), .ZN(n5722) );
  AOI211_X1 U5533 ( .C1(n4669), .C2(n4522), .A(n4667), .B(n5732), .ZN(n5751)
         );
  AOI21_X1 U5534 ( .B1(n5754), .B2(n5831), .A(n4673), .ZN(n4672) );
  NAND2_X1 U5535 ( .A1(n5756), .A2(n5755), .ZN(n4673) );
  NAND2_X1 U5536 ( .A1(n4674), .A2(n4670), .ZN(n5769) );
  OAI21_X1 U5537 ( .B1(n4672), .B2(n4671), .A(n5792), .ZN(n4670) );
  NAND2_X1 U5538 ( .A1(n5758), .A2(n6207), .ZN(n4674) );
  NAND2_X1 U5539 ( .A1(n5757), .A2(n7908), .ZN(n4671) );
  OAI21_X1 U5540 ( .B1(n4632), .B2(n4514), .A(n4628), .ZN(n8260) );
  AND2_X1 U5541 ( .A1(n8246), .A2(n4629), .ZN(n4628) );
  AOI21_X1 U5542 ( .B1(n8228), .B2(n8227), .A(n4633), .ZN(n4632) );
  INV_X1 U5543 ( .A(n5773), .ZN(n4684) );
  AND2_X1 U5544 ( .A1(n4556), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5545 ( .A1(n4638), .A2(n4494), .ZN(n4637) );
  AND2_X1 U5546 ( .A1(n4639), .A2(n8275), .ZN(n4635) );
  NAND2_X1 U5547 ( .A1(n4687), .A2(n4682), .ZN(n5780) );
  NAND2_X1 U5548 ( .A1(n4685), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5549 ( .A1(n5777), .A2(n5792), .ZN(n4687) );
  NOR2_X1 U5550 ( .A1(n4684), .A2(n5792), .ZN(n4683) );
  INV_X1 U5551 ( .A(n5797), .ZN(n4680) );
  NAND2_X1 U5552 ( .A1(n4970), .A2(n4967), .ZN(n8181) );
  INV_X1 U5553 ( .A(n7273), .ZN(n4970) );
  NOR2_X1 U5554 ( .A1(n8177), .A2(n4968), .ZN(n4967) );
  AND2_X1 U5555 ( .A1(n9018), .A2(n8323), .ZN(n4627) );
  OR2_X1 U5556 ( .A1(n8326), .A2(n8343), .ZN(n4626) );
  INV_X1 U5557 ( .A(n4627), .ZN(n4620) );
  INV_X1 U5558 ( .A(n8798), .ZN(n4953) );
  AND2_X1 U5559 ( .A1(n4643), .A2(n4645), .ZN(n4642) );
  INV_X1 U5560 ( .A(n4622), .ZN(n4621) );
  AOI21_X1 U5561 ( .B1(n8325), .B2(n4627), .A(n4625), .ZN(n4622) );
  INV_X1 U5562 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6538) );
  OR2_X1 U5563 ( .A1(n4758), .A2(n4756), .ZN(n4755) );
  NOR2_X1 U5564 ( .A1(n4760), .A2(n4759), .ZN(n4758) );
  NAND2_X1 U5565 ( .A1(n4675), .A2(n5795), .ZN(n5799) );
  NAND2_X1 U5566 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  AND2_X1 U5567 ( .A1(n9775), .A2(n9482), .ZN(n5796) );
  NAND2_X1 U5568 ( .A1(n5265), .A2(n5264), .ZN(n5791) );
  NAND2_X1 U5569 ( .A1(n4914), .A2(n7697), .ZN(n4913) );
  INV_X1 U5570 ( .A(n7696), .ZN(n4914) );
  AOI21_X1 U5571 ( .B1(n4871), .B2(n4868), .A(n4867), .ZN(n4866) );
  INV_X1 U5572 ( .A(n5291), .ZN(n4867) );
  INV_X1 U5573 ( .A(n4873), .ZN(n4868) );
  INV_X1 U5574 ( .A(n4871), .ZN(n4869) );
  INV_X1 U5575 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5239) );
  INV_X1 U5576 ( .A(n5426), .ZN(n4843) );
  INV_X1 U5577 ( .A(n5077), .ZN(n4856) );
  NAND2_X1 U5578 ( .A1(n5137), .A2(n5136), .ZN(n5140) );
  AND2_X1 U5579 ( .A1(n5544), .A2(n5111), .ZN(n5110) );
  INV_X1 U5580 ( .A(n4838), .ZN(n5111) );
  NOR2_X1 U5581 ( .A1(n4838), .A2(n5628), .ZN(n4837) );
  NAND2_X1 U5582 ( .A1(n5122), .A2(n5121), .ZN(n5125) );
  OR2_X1 U5583 ( .A1(n5116), .A2(n5115), .ZN(n5599) );
  INV_X1 U5584 ( .A(n5632), .ZN(n5115) );
  XNOR2_X1 U5585 ( .A(n7278), .B(n8116), .ZN(n6565) );
  NOR2_X1 U5586 ( .A1(n7928), .A2(n4599), .ZN(n4598) );
  INV_X1 U5587 ( .A(n7840), .ZN(n4599) );
  INV_X1 U5588 ( .A(n4601), .ZN(n4596) );
  AOI21_X1 U5589 ( .B1(n4900), .B2(n4899), .A(n4536), .ZN(n4898) );
  INV_X1 U5590 ( .A(n4904), .ZN(n4899) );
  AND2_X1 U5591 ( .A1(n8341), .A2(n8171), .ZN(n8337) );
  INV_X1 U5592 ( .A(n8083), .ZN(n5013) );
  NAND2_X1 U5593 ( .A1(n4745), .A2(n9075), .ZN(n4744) );
  NOR2_X1 U5594 ( .A1(n9252), .A2(n9255), .ZN(n4745) );
  NOR2_X1 U5595 ( .A1(n9287), .A2(n9284), .ZN(n4740) );
  NAND2_X1 U5596 ( .A1(n5056), .A2(n5054), .ZN(n5053) );
  INV_X1 U5597 ( .A(n8212), .ZN(n4897) );
  NAND2_X1 U5598 ( .A1(n8238), .A2(n4489), .ZN(n4734) );
  INV_X1 U5599 ( .A(n9120), .ZN(n8142) );
  INV_X1 U5600 ( .A(n5043), .ZN(n5041) );
  INV_X1 U5601 ( .A(n6336), .ZN(n4725) );
  NAND2_X1 U5602 ( .A1(n4607), .A2(n6239), .ZN(n6336) );
  NAND2_X1 U5603 ( .A1(n5006), .A2(n6783), .ZN(n5005) );
  INV_X1 U5604 ( .A(n6172), .ZN(n5992) );
  INV_X1 U5605 ( .A(n5796), .ZN(n5903) );
  NAND2_X1 U5606 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n4767) );
  NOR2_X1 U5607 ( .A1(n5621), .A2(n5620), .ZN(n5623) );
  NOR2_X1 U5608 ( .A1(n9777), .A2(n6220), .ZN(n5807) );
  AND2_X1 U5609 ( .A1(n9777), .A2(n6220), .ZN(n5898) );
  NAND2_X1 U5610 ( .A1(n4787), .A2(n9623), .ZN(n4786) );
  INV_X1 U5611 ( .A(n5689), .ZN(n5354) );
  NOR2_X1 U5612 ( .A1(n9807), .A2(n9812), .ZN(n4787) );
  OR2_X1 U5613 ( .A1(n9807), .A2(n9450), .ZN(n7914) );
  INV_X1 U5614 ( .A(n5355), .ZN(n5342) );
  NOR2_X1 U5615 ( .A1(n9385), .A2(n5377), .ZN(n5366) );
  NAND2_X1 U5616 ( .A1(n5282), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5377) );
  INV_X1 U5617 ( .A(n5389), .ZN(n5282) );
  AOI21_X1 U5618 ( .B1(n7882), .B2(n4816), .A(n7907), .ZN(n4814) );
  OAI21_X1 U5619 ( .B1(n4921), .B2(n4925), .A(n9709), .ZN(n4920) );
  INV_X1 U5620 ( .A(n4922), .ZN(n4921) );
  NOR2_X1 U5621 ( .A1(n7905), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5622 ( .A1(n5434), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5422) );
  NOR2_X1 U5623 ( .A1(n5670), .A2(n5435), .ZN(n5434) );
  INV_X1 U5624 ( .A(n7900), .ZN(n4819) );
  NOR2_X1 U5625 ( .A1(n5467), .A2(n5450), .ZN(n5669) );
  OR2_X1 U5626 ( .A1(n5481), .A2(n5465), .ZN(n5467) );
  OR2_X1 U5627 ( .A1(n5591), .A2(n6798), .ZN(n5649) );
  OR2_X1 U5628 ( .A1(n5614), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U5629 ( .A1(n5875), .A2(n5828), .ZN(n7031) );
  OR2_X1 U5630 ( .A1(n6870), .A2(n6871), .ZN(n6868) );
  INV_X1 U5631 ( .A(n5227), .ZN(n4861) );
  NOR2_X1 U5632 ( .A1(n5326), .A2(n4874), .ZN(n4873) );
  INV_X1 U5633 ( .A(n5198), .ZN(n4874) );
  AOI21_X1 U5634 ( .B1(n4873), .B2(n5199), .A(n4872), .ZN(n4871) );
  INV_X1 U5635 ( .A(n5204), .ZN(n4872) );
  NAND2_X1 U5636 ( .A1(n5183), .A2(n5182), .ZN(n5339) );
  NAND2_X1 U5637 ( .A1(n5374), .A2(n5373), .ZN(n4851) );
  NAND2_X1 U5638 ( .A1(n5129), .A2(n5128), .ZN(n5132) );
  NAND2_X1 U5639 ( .A1(n5117), .A2(n5108), .ZN(n5604) );
  NAND2_X1 U5640 ( .A1(n5107), .A2(SI_8_), .ZN(n5108) );
  AND2_X1 U5641 ( .A1(n5630), .A2(n5113), .ZN(n5600) );
  NAND2_X1 U5642 ( .A1(n5495), .A2(n5245), .ZN(n5409) );
  INV_X1 U5643 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5244) );
  INV_X1 U5644 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4652) );
  NOR2_X1 U5645 ( .A1(n7841), .A2(n4602), .ZN(n4601) );
  INV_X1 U5646 ( .A(n7620), .ZN(n4602) );
  NAND2_X1 U5647 ( .A1(n8851), .A2(n8034), .ZN(n8056) );
  OR2_X1 U5648 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  AOI21_X1 U5649 ( .B1(n8419), .B2(n8089), .A(n8102), .ZN(n4591) );
  INV_X1 U5650 ( .A(n4591), .ZN(n4589) );
  AOI21_X1 U5651 ( .B1(n4957), .B2(n4955), .A(n4524), .ZN(n4954) );
  INV_X1 U5652 ( .A(n8788), .ZN(n4955) );
  INV_X1 U5653 ( .A(n4957), .ZN(n4956) );
  OR2_X1 U5654 ( .A1(n6962), .A2(n6961), .ZN(n7064) );
  NAND2_X1 U5655 ( .A1(n6630), .A2(n6629), .ZN(n7995) );
  OR2_X1 U5656 ( .A1(n7995), .A2(n8844), .ZN(n8009) );
  NAND2_X1 U5657 ( .A1(n8789), .A2(n8788), .ZN(n8787) );
  XNOR2_X1 U5658 ( .A(n8033), .B(n8031), .ZN(n8853) );
  NAND2_X1 U5659 ( .A1(n8853), .A2(n8852), .ZN(n8851) );
  OR2_X1 U5660 ( .A1(n7416), .A2(n4974), .ZN(n4973) );
  INV_X1 U5661 ( .A(n7314), .ZN(n4974) );
  INV_X1 U5662 ( .A(n7223), .ZN(n4975) );
  NAND2_X1 U5663 ( .A1(n6624), .A2(n6623), .ZN(n6932) );
  INV_X1 U5664 ( .A(n6854), .ZN(n6624) );
  NAND2_X1 U5665 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  OR2_X1 U5666 ( .A1(n7796), .A2(n7795), .ZN(n7804) );
  OAI21_X1 U5667 ( .B1(n7621), .B2(n4597), .A(n4594), .ZN(n8880) );
  AOI21_X1 U5668 ( .B1(n4598), .B2(n4596), .A(n4595), .ZN(n4594) );
  INV_X1 U5669 ( .A(n4598), .ZN(n4597) );
  INV_X1 U5670 ( .A(n7927), .ZN(n4595) );
  NAND2_X1 U5671 ( .A1(n8324), .A2(n4614), .ZN(n4613) );
  INV_X1 U5672 ( .A(n4612), .ZN(n4611) );
  AND2_X1 U5673 ( .A1(n4703), .A2(n4702), .ZN(n6418) );
  NAND2_X1 U5674 ( .A1(n6424), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4702) );
  AND2_X1 U5675 ( .A1(n4699), .A2(n4698), .ZN(n8917) );
  NAND2_X1 U5676 ( .A1(n6670), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4698) );
  INV_X1 U5677 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6379) );
  NOR2_X1 U5678 ( .A1(n7474), .A2(n4569), .ZN(n7478) );
  NAND2_X1 U5679 ( .A1(n7478), .A2(n7477), .ZN(n7610) );
  NAND2_X1 U5680 ( .A1(n8950), .A2(n4691), .ZN(n8952) );
  NAND2_X1 U5681 ( .A1(n8957), .A2(n8941), .ZN(n4691) );
  NOR2_X1 U5682 ( .A1(n8952), .A2(n8951), .ZN(n8970) );
  NOR2_X1 U5683 ( .A1(n8970), .A2(n4690), .ZN(n10178) );
  AND2_X1 U5684 ( .A1(n8971), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4690) );
  OR2_X1 U5685 ( .A1(n8975), .A2(n10172), .ZN(n4694) );
  NAND2_X1 U5686 ( .A1(n4902), .A2(n4903), .ZN(n8406) );
  NOR2_X1 U5687 ( .A1(n9220), .A2(n8995), .ZN(n8986) );
  OR2_X1 U5688 ( .A1(n9011), .A2(n9226), .ZN(n8995) );
  OR2_X1 U5689 ( .A1(n9242), .A2(n8897), .ZN(n8398) );
  INV_X1 U5690 ( .A(n8067), .ZN(n8065) );
  NAND2_X1 U5691 ( .A1(n5023), .A2(n5025), .ZN(n9063) );
  INV_X1 U5692 ( .A(n5026), .ZN(n5025) );
  OAI21_X1 U5693 ( .B1(n5028), .B2(n5027), .A(n8396), .ZN(n5026) );
  INV_X1 U5694 ( .A(n8397), .ZN(n9066) );
  OR2_X1 U5695 ( .A1(n8025), .A2(n8024), .ZN(n8027) );
  AND2_X1 U5696 ( .A1(n8052), .A2(n8051), .ZN(n9093) );
  NAND2_X1 U5697 ( .A1(n9102), .A2(n8144), .ZN(n9088) );
  NAND2_X1 U5698 ( .A1(n8144), .A2(n9121), .ZN(n4893) );
  NOR2_X1 U5699 ( .A1(n9116), .A2(n4743), .ZN(n9081) );
  INV_X1 U5700 ( .A(n4745), .ZN(n4743) );
  NAND2_X1 U5701 ( .A1(n8142), .A2(n8141), .ZN(n9102) );
  NOR2_X1 U5702 ( .A1(n9116), .A2(n9255), .ZN(n9098) );
  AOI21_X1 U5703 ( .B1(n4908), .B2(n9177), .A(n4906), .ZN(n4905) );
  INV_X1 U5704 ( .A(n8304), .ZN(n4906) );
  AND2_X1 U5705 ( .A1(n9208), .A2(n4736), .ZN(n9146) );
  NOR2_X1 U5706 ( .A1(n9273), .A2(n4738), .ZN(n4736) );
  NAND2_X1 U5707 ( .A1(n9208), .A2(n4740), .ZN(n9185) );
  NAND2_X1 U5708 ( .A1(n6628), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7950) );
  INV_X1 U5709 ( .A(n7804), .ZN(n6628) );
  AND4_X1 U5710 ( .A1(n7809), .A2(n7808), .A3(n7807), .A4(n7806), .ZN(n9181)
         );
  NAND2_X1 U5711 ( .A1(n9208), .A2(n9207), .ZN(n9210) );
  AND2_X1 U5712 ( .A1(n7814), .A2(n8894), .ZN(n9208) );
  OR2_X1 U5713 ( .A1(n7757), .A2(n9299), .ZN(n7823) );
  AND4_X1 U5714 ( .A1(n7802), .A2(n7801), .A3(n7800), .A4(n7799), .ZN(n7930)
         );
  AND4_X1 U5715 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n7750)
         );
  AND4_X1 U5716 ( .A1(n7632), .A2(n7631), .A3(n7630), .A4(n7629), .ZN(n7832)
         );
  AND4_X1 U5717 ( .A1(n7599), .A2(n7598), .A3(n7597), .A4(n7596), .ZN(n7846)
         );
  OR2_X1 U5718 ( .A1(n8184), .A2(n7437), .ZN(n7664) );
  AND2_X1 U5719 ( .A1(n4554), .A2(n7252), .ZN(n5070) );
  AND4_X1 U5720 ( .A1(n7327), .A2(n7326), .A3(n7325), .A4(n7324), .ZN(n7683)
         );
  AND2_X1 U5721 ( .A1(n8254), .A2(n8211), .ZN(n8184) );
  NAND2_X1 U5722 ( .A1(n4562), .A2(n8212), .ZN(n7442) );
  AND4_X1 U5723 ( .A1(n7232), .A2(n7231), .A3(n7230), .A4(n7229), .ZN(n7433)
         );
  OR2_X1 U5724 ( .A1(n7396), .A2(n7527), .ZN(n7449) );
  NAND2_X1 U5725 ( .A1(n5071), .A2(n7252), .ZN(n7436) );
  AND4_X1 U5726 ( .A1(n7070), .A2(n7069), .A3(n7068), .A4(n7067), .ZN(n7443)
         );
  AND4_X1 U5727 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n7260)
         );
  INV_X1 U5728 ( .A(n5016), .ZN(n5015) );
  OAI21_X1 U5729 ( .B1(n7157), .B2(n4511), .A(n7160), .ZN(n5016) );
  AND2_X1 U5730 ( .A1(n8248), .A2(n8258), .ZN(n8246) );
  INV_X1 U5731 ( .A(n7241), .ZN(n7251) );
  AND2_X1 U5732 ( .A1(n7352), .A2(n7251), .ZN(n7266) );
  NOR2_X1 U5733 ( .A1(n7351), .A2(n8229), .ZN(n7352) );
  NAND2_X1 U5734 ( .A1(n4880), .A2(n4878), .ZN(n7346) );
  INV_X1 U5735 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U5736 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6854) );
  NAND2_X1 U5737 ( .A1(n10198), .A2(n10249), .ZN(n10196) );
  NOR2_X1 U5738 ( .A1(n4734), .A2(n7280), .ZN(n10198) );
  NAND2_X1 U5739 ( .A1(n4731), .A2(n4489), .ZN(n7188) );
  NAND2_X1 U5740 ( .A1(n7143), .A2(n6549), .ZN(n7254) );
  NAND2_X1 U5741 ( .A1(n8093), .A2(n8092), .ZN(n9230) );
  NAND2_X1 U5742 ( .A1(n5038), .A2(n5042), .ZN(n9134) );
  NAND2_X1 U5743 ( .A1(n5045), .A2(n5043), .ZN(n5038) );
  NAND2_X1 U5744 ( .A1(n6573), .A2(n6549), .ZN(n10258) );
  INV_X1 U5745 ( .A(n4949), .ZN(n4947) );
  NOR2_X1 U5746 ( .A1(n4978), .A2(n4977), .ZN(n6694) );
  NOR2_X1 U5747 ( .A1(n4978), .A2(n4976), .ZN(n6537) );
  INV_X1 U5748 ( .A(n5033), .ZN(n4976) );
  INV_X1 U5749 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6323) );
  INV_X1 U5750 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6314) );
  INV_X1 U5751 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8770) );
  AND2_X1 U5752 ( .A1(n6307), .A2(n6231), .ZN(n6313) );
  NAND2_X1 U5753 ( .A1(n6946), .A2(n6947), .ZN(n6945) );
  NAND2_X1 U5754 ( .A1(n6137), .A2(n6136), .ZN(n9363) );
  NAND2_X1 U5755 ( .A1(n9459), .A2(n9462), .ZN(n5009) );
  INV_X1 U5756 ( .A(n9568), .ZN(n6220) );
  AND2_X1 U5757 ( .A1(n6081), .A2(n6071), .ZN(n5007) );
  NAND2_X1 U5758 ( .A1(n5354), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U5759 ( .A1(n9426), .A2(n9427), .ZN(n9425) );
  INV_X1 U5760 ( .A(n4994), .ZN(n4993) );
  AOI21_X1 U5761 ( .B1(n4994), .B2(n4992), .A(n4539), .ZN(n4991) );
  INV_X1 U5762 ( .A(n7407), .ZN(n4992) );
  XNOR2_X1 U5763 ( .A(n5957), .B(n6172), .ZN(n5959) );
  NAND2_X1 U5764 ( .A1(n6098), .A2(n6099), .ZN(n9459) );
  NAND2_X1 U5765 ( .A1(n5537), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5621) );
  AOI21_X1 U5766 ( .B1(n4770), .B2(n6718), .A(n4544), .ZN(n4769) );
  AOI21_X1 U5767 ( .B1(n4499), .B2(n5000), .A(n4534), .ZN(n4998) );
  NOR2_X1 U5768 ( .A1(n6299), .A2(n4513), .ZN(n9965) );
  INV_X1 U5769 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5531) );
  OR2_X1 U5770 ( .A1(n9992), .A2(n9993), .ZN(n4707) );
  NOR2_X1 U5771 ( .A1(n6799), .A2(n4719), .ZN(n10017) );
  AND2_X1 U5772 ( .A1(n6803), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5773 ( .A1(n10017), .A2(n10018), .ZN(n10016) );
  NOR2_X1 U5774 ( .A1(n6271), .A2(n7721), .ZN(n9497) );
  AOI21_X1 U5775 ( .B1(n9538), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9537), .ZN(
        n10035) );
  NAND2_X1 U5776 ( .A1(n5268), .A2(n5267), .ZN(n9554) );
  NOR2_X1 U5777 ( .A1(n9553), .A2(n9554), .ZN(n9552) );
  NAND2_X1 U5778 ( .A1(n9565), .A2(n7920), .ZN(n4829) );
  NAND2_X1 U5779 ( .A1(n9576), .A2(n9735), .ZN(n4827) );
  AOI21_X1 U5780 ( .B1(n4805), .B2(n7918), .A(n7919), .ZN(n4804) );
  AND2_X1 U5781 ( .A1(n7923), .A2(n5306), .ZN(n9562) );
  AND2_X1 U5782 ( .A1(n5805), .A2(n7920), .ZN(n9567) );
  NAND2_X1 U5783 ( .A1(n4931), .A2(n4930), .ZN(n9574) );
  AOI21_X1 U5784 ( .B1(n4932), .B2(n4937), .A(n4547), .ZN(n4930) );
  NAND2_X1 U5785 ( .A1(n4795), .A2(n4794), .ZN(n9637) );
  AOI21_X1 U5786 ( .B1(n4797), .B2(n4799), .A(n7913), .ZN(n4794) );
  NOR2_X1 U5787 ( .A1(n9658), .A2(n4785), .ZN(n9632) );
  INV_X1 U5788 ( .A(n4787), .ZN(n4785) );
  NOR2_X1 U5789 ( .A1(n9658), .A2(n9812), .ZN(n9645) );
  AND2_X1 U5790 ( .A1(n5757), .A2(n7909), .ZN(n9677) );
  NAND2_X1 U5791 ( .A1(n4813), .A2(n4811), .ZN(n9691) );
  AOI21_X1 U5792 ( .B1(n4814), .B2(n4815), .A(n4812), .ZN(n4811) );
  NAND2_X1 U5793 ( .A1(n9733), .A2(n4814), .ZN(n4813) );
  INV_X1 U5794 ( .A(n4816), .ZN(n4815) );
  NOR2_X1 U5795 ( .A1(n5752), .A2(n5857), .ZN(n9692) );
  AND2_X1 U5796 ( .A1(n9732), .A2(n4816), .ZN(n9707) );
  OAI21_X1 U5797 ( .B1(n7765), .B2(n4821), .A(n4818), .ZN(n9752) );
  AOI21_X1 U5798 ( .B1(n4822), .B2(n4820), .A(n4819), .ZN(n4818) );
  INV_X1 U5799 ( .A(n4822), .ZN(n4821) );
  INV_X1 U5800 ( .A(n7767), .ZN(n4820) );
  INV_X1 U5801 ( .A(n4783), .ZN(n9761) );
  NAND2_X1 U5802 ( .A1(n4832), .A2(n4830), .ZN(n7700) );
  INV_X1 U5803 ( .A(n7501), .ZN(n4831) );
  AND2_X1 U5804 ( .A1(n7292), .A2(n7291), .ZN(n7301) );
  OR2_X1 U5805 ( .A1(n7287), .A2(n4833), .ZN(n7500) );
  NAND2_X1 U5806 ( .A1(n7079), .A2(n7078), .ZN(n7287) );
  AND2_X1 U5807 ( .A1(n7463), .A2(n7288), .ZN(n7090) );
  NAND2_X1 U5808 ( .A1(n5638), .A2(n5637), .ZN(n7045) );
  OR2_X1 U5809 ( .A1(n7039), .A2(n7045), .ZN(n7091) );
  OR2_X1 U5810 ( .A1(n7034), .A2(n7083), .ZN(n7079) );
  NAND2_X1 U5811 ( .A1(n4782), .A2(n4781), .ZN(n7039) );
  AND2_X1 U5812 ( .A1(n5875), .A2(n5826), .ZN(n7029) );
  OAI21_X1 U5813 ( .B1(n6809), .B2(n6895), .A(n5820), .ZN(n6974) );
  OAI21_X1 U5814 ( .B1(n6884), .B2(n5822), .A(n5881), .ZN(n6809) );
  INV_X1 U5815 ( .A(n6834), .ZN(n6897) );
  NAND2_X1 U5816 ( .A1(n5820), .A2(n5879), .ZN(n6895) );
  NAND2_X1 U5817 ( .A1(n6868), .A2(n5713), .ZN(n6884) );
  NAND2_X1 U5818 ( .A1(n10057), .A2(n6828), .ZN(n10055) );
  INV_X1 U5819 ( .A(n5941), .ZN(n10057) );
  NAND2_X1 U5820 ( .A1(n5305), .A2(n5304), .ZN(n9782) );
  NAND2_X1 U5821 ( .A1(n8361), .A2(n5303), .ZN(n5305) );
  OR2_X1 U5822 ( .A1(n6610), .A2(n5568), .ZN(n4777) );
  NAND2_X1 U5823 ( .A1(n5563), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4778) );
  XNOR2_X1 U5824 ( .A(n5266), .B(SI_30_), .ZN(n8380) );
  XNOR2_X1 U5825 ( .A(n5277), .B(n5276), .ZN(n9329) );
  XNOR2_X1 U5826 ( .A(n5302), .B(n5301), .ZN(n8361) );
  CLKBUF_X1 U5827 ( .A(n5924), .Z(n5925) );
  XNOR2_X1 U5828 ( .A(n5314), .B(n5313), .ZN(n8091) );
  NOR2_X1 U5829 ( .A1(n4944), .A2(n5010), .ZN(n4942) );
  NAND2_X1 U5830 ( .A1(n4841), .A2(n4845), .ZN(n5427) );
  OR2_X1 U5831 ( .A1(n5146), .A2(n4506), .ZN(n4841) );
  NAND2_X1 U5832 ( .A1(n4848), .A2(n5149), .ZN(n5661) );
  NAND2_X1 U5833 ( .A1(n5146), .A2(n4849), .ZN(n4848) );
  OR2_X1 U5834 ( .A1(n5606), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5608) );
  XNOR2_X1 U5835 ( .A(n5112), .B(SI_6_), .ZN(n5628) );
  NAND2_X1 U5837 ( .A1(n5097), .A2(n5096), .ZN(n5494) );
  OR2_X1 U5838 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5564) );
  NAND2_X1 U5839 ( .A1(n6954), .A2(n6953), .ZN(n7050) );
  AND2_X1 U5840 ( .A1(n8115), .A2(n8114), .ZN(n9022) );
  NAND2_X1 U5841 ( .A1(n4600), .A2(n7840), .ZN(n7929) );
  NAND2_X1 U5842 ( .A1(n7621), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U5843 ( .A1(n7787), .A2(n7786), .ZN(n7849) );
  NAND2_X1 U5844 ( .A1(n7315), .A2(n7314), .ZN(n7417) );
  OAI22_X1 U5845 ( .A1(n4589), .A2(n4588), .B1(n8119), .B2(n4591), .ZN(n4587)
         );
  NOR2_X1 U5846 ( .A1(n8419), .A2(n8119), .ZN(n4588) );
  INV_X1 U5847 ( .A(n8119), .ZN(n4590) );
  NAND2_X1 U5848 ( .A1(n6848), .A2(n6847), .ZN(n6849) );
  NAND2_X1 U5849 ( .A1(n8043), .A2(n8042), .ZN(n9247) );
  NAND2_X1 U5850 ( .A1(n7212), .A2(n7211), .ZN(n7224) );
  NAND2_X1 U5851 ( .A1(n8787), .A2(n7991), .ZN(n8843) );
  NAND2_X1 U5852 ( .A1(n7621), .A2(n7620), .ZN(n7842) );
  NAND2_X1 U5853 ( .A1(n7420), .A2(n7419), .ZN(n7731) );
  AND2_X1 U5854 ( .A1(n8869), .A2(n4961), .ZN(n4960) );
  NAND2_X1 U5855 ( .A1(n4963), .A2(n4962), .ZN(n4961) );
  INV_X1 U5856 ( .A(n4965), .ZN(n4962) );
  NAND2_X1 U5857 ( .A1(n4959), .A2(n4963), .ZN(n8870) );
  NAND2_X1 U5858 ( .A1(n8806), .A2(n4965), .ZN(n4959) );
  AND2_X1 U5859 ( .A1(n6640), .A2(n6639), .ZN(n9108) );
  INV_X1 U5860 ( .A(n6995), .ZN(n8912) );
  INV_X1 U5861 ( .A(n4703), .ZN(n6442) );
  INV_X1 U5862 ( .A(n4701), .ZN(n6468) );
  INV_X1 U5863 ( .A(n4699), .ZN(n6666) );
  NOR2_X1 U5864 ( .A1(n6770), .A2(n4570), .ZN(n6773) );
  NOR2_X1 U5865 ( .A1(n6773), .A2(n6772), .ZN(n7017) );
  NAND2_X1 U5866 ( .A1(n6540), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U5867 ( .A1(n8169), .A2(n8168), .ZN(n9217) );
  NAND2_X1 U5868 ( .A1(n8075), .A2(n8153), .ZN(n8078) );
  NAND2_X1 U5869 ( .A1(n9054), .A2(n8206), .ZN(n9033) );
  NAND2_X1 U5870 ( .A1(n9080), .A2(n9079), .ZN(n9078) );
  NAND2_X1 U5871 ( .A1(n5029), .A2(n5028), .ZN(n9080) );
  NAND2_X1 U5872 ( .A1(n9114), .A2(n5030), .ZN(n5029) );
  AND2_X1 U5873 ( .A1(n5032), .A2(n4516), .ZN(n9097) );
  NAND2_X1 U5874 ( .A1(n9114), .A2(n8393), .ZN(n5032) );
  AND2_X1 U5875 ( .A1(n8008), .A2(n8007), .ZN(n9118) );
  NAND2_X1 U5876 ( .A1(n7994), .A2(n7993), .ZN(n9267) );
  NAND2_X1 U5877 ( .A1(n5044), .A2(n5048), .ZN(n9145) );
  NAND2_X1 U5878 ( .A1(n5045), .A2(n4497), .ZN(n5044) );
  AND2_X1 U5879 ( .A1(n4909), .A2(n8295), .ZN(n9167) );
  NOR2_X1 U5880 ( .A1(n9200), .A2(n8389), .ZN(n9175) );
  NAND2_X1 U5881 ( .A1(n8388), .A2(n8387), .ZN(n9201) );
  NAND2_X1 U5882 ( .A1(n5055), .A2(n5056), .ZN(n7820) );
  NAND2_X1 U5883 ( .A1(n5063), .A2(n5057), .ZN(n7811) );
  NAND2_X1 U5884 ( .A1(n5063), .A2(n5062), .ZN(n7745) );
  NAND2_X1 U5885 ( .A1(n7319), .A2(n7318), .ZN(n7663) );
  NAND2_X1 U5886 ( .A1(n7005), .A2(n5021), .ZN(n5019) );
  AND3_X1 U5887 ( .A1(n4649), .A2(n6840), .A3(n4553), .ZN(n7174) );
  OR2_X1 U5888 ( .A1(n6838), .A2(n6957), .ZN(n4649) );
  NAND2_X1 U5889 ( .A1(n4882), .A2(n8240), .ZN(n7162) );
  OR2_X1 U5890 ( .A1(n10192), .A2(n7009), .ZN(n4882) );
  NAND2_X1 U5891 ( .A1(n7005), .A2(n7004), .ZN(n7159) );
  INV_X1 U5892 ( .A(n9164), .ZN(n10205) );
  INV_X1 U5893 ( .A(n7278), .ZN(n10228) );
  AND2_X1 U5894 ( .A1(n4728), .A2(n4727), .ZN(n9900) );
  NAND2_X1 U5895 ( .A1(n4729), .A2(n10197), .ZN(n4728) );
  INV_X1 U5896 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U5897 ( .A1(n6338), .A2(n4535), .ZN(n4606) );
  NOR2_X1 U5898 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5899 ( .A1(n6249), .A2(n6248), .ZN(n6342) );
  AND2_X1 U5900 ( .A1(n4948), .A2(n4949), .ZN(n6545) );
  INV_X1 U5901 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U5902 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4689) );
  INV_X1 U5903 ( .A(n6169), .ZN(n9337) );
  NAND2_X1 U5904 ( .A1(n5449), .A2(n5448), .ZN(n9357) );
  NAND2_X1 U5905 ( .A1(n7128), .A2(n6024), .ZN(n7370) );
  NAND2_X1 U5906 ( .A1(n5009), .A2(n9460), .ZN(n9375) );
  NAND2_X1 U5907 ( .A1(n5388), .A2(n5387), .ZN(n9828) );
  AND2_X1 U5908 ( .A1(n6204), .A2(n6197), .ZN(n6198) );
  AND2_X1 U5909 ( .A1(n6162), .A2(n9335), .ZN(n5012) );
  NAND2_X1 U5910 ( .A1(n5940), .A2(n6172), .ZN(n5945) );
  NAND2_X1 U5911 ( .A1(n5365), .A2(n5364), .ZN(n9818) );
  NAND2_X1 U5912 ( .A1(n5480), .A2(n5479), .ZN(n7692) );
  NAND2_X1 U5913 ( .A1(n9425), .A2(n6145), .ZN(n9393) );
  NAND2_X1 U5914 ( .A1(n8062), .A2(n5303), .ZN(n5329) );
  INV_X1 U5915 ( .A(n9492), .ZN(n7037) );
  NAND2_X1 U5916 ( .A1(n6715), .A2(n5981), .ZN(n6705) );
  NAND2_X1 U5917 ( .A1(n5418), .A2(n5417), .ZN(n9837) );
  NAND2_X1 U5918 ( .A1(n5588), .A2(n5587), .ZN(n10138) );
  OAI21_X1 U5919 ( .B1(n9384), .B2(n9382), .A(n4756), .ZN(n9446) );
  INV_X1 U5920 ( .A(n4761), .ZN(n9445) );
  AOI21_X1 U5921 ( .B1(n9384), .B2(n9381), .A(n4762), .ZN(n4761) );
  NAND2_X1 U5922 ( .A1(n7369), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U5923 ( .A1(n5401), .A2(n5400), .ZN(n9832) );
  INV_X1 U5924 ( .A(n4840), .ZN(n4839) );
  OAI21_X1 U5925 ( .B1(n5871), .B2(n5929), .A(n6977), .ZN(n4840) );
  NAND4_X1 U5926 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n9494)
         );
  NAND2_X1 U5927 ( .A1(n5647), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U5928 ( .A1(n4984), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U5929 ( .A1(n4492), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4986) );
  INV_X1 U5930 ( .A(n4714), .ZN(n9950) );
  AND2_X1 U5931 ( .A1(n4712), .A2(n4711), .ZN(n6299) );
  INV_X1 U5932 ( .A(n6300), .ZN(n4711) );
  INV_X1 U5933 ( .A(n4712), .ZN(n6301) );
  NAND2_X1 U5934 ( .A1(n9980), .A2(n9981), .ZN(n9979) );
  NAND2_X1 U5935 ( .A1(n9979), .A2(n4708), .ZN(n9992) );
  NAND2_X1 U5936 ( .A1(n6326), .A2(n8450), .ZN(n4708) );
  INV_X1 U5937 ( .A(n4707), .ZN(n9991) );
  NAND2_X1 U5938 ( .A1(n10005), .A2(n4561), .ZN(n6396) );
  NOR2_X1 U5939 ( .A1(n6685), .A2(n6684), .ZN(n6683) );
  NAND2_X1 U5940 ( .A1(n4716), .A2(n4715), .ZN(n6685) );
  NAND2_X1 U5941 ( .A1(n6350), .A2(n7094), .ZN(n4715) );
  NAND2_X1 U5942 ( .A1(n6396), .A2(n4717), .ZN(n4716) );
  INV_X1 U5943 ( .A(n6397), .ZN(n4717) );
  NAND2_X1 U5944 ( .A1(n10016), .A2(n4718), .ZN(n7110) );
  OR2_X1 U5945 ( .A1(n10026), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4718) );
  INV_X1 U5946 ( .A(n4710), .ZN(n7338) );
  XNOR2_X1 U5947 ( .A(n9497), .B(n9503), .ZN(n6273) );
  NOR2_X1 U5948 ( .A1(n6273), .A2(n5673), .ZN(n9498) );
  OAI21_X1 U5949 ( .B1(n6273), .B2(n4721), .A(n4720), .ZN(n9516) );
  NAND2_X1 U5950 ( .A1(n4722), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5951 ( .A1(n9499), .A2(n4722), .ZN(n4720) );
  INV_X1 U5952 ( .A(n9501), .ZN(n4722) );
  XNOR2_X1 U5953 ( .A(n9552), .B(n5265), .ZN(n9773) );
  AND2_X1 U5954 ( .A1(n4807), .A2(n4805), .ZN(n9578) );
  NAND2_X1 U5955 ( .A1(n4933), .A2(n4935), .ZN(n9589) );
  OR2_X1 U5956 ( .A1(n9618), .A2(n4937), .ZN(n4933) );
  OR2_X1 U5957 ( .A1(n9618), .A2(n7892), .ZN(n4934) );
  INV_X1 U5958 ( .A(n9803), .ZN(n9623) );
  NAND2_X1 U5959 ( .A1(n4796), .A2(n4800), .ZN(n9650) );
  NAND2_X1 U5960 ( .A1(n4793), .A2(n4797), .ZN(n9649) );
  NAND2_X1 U5961 ( .A1(n4802), .A2(n7909), .ZN(n9664) );
  OR2_X1 U5962 ( .A1(n9678), .A2(n7910), .ZN(n4802) );
  NAND2_X1 U5963 ( .A1(n4918), .A2(n4922), .ZN(n9699) );
  NAND2_X1 U5964 ( .A1(n9731), .A2(n4925), .ZN(n4918) );
  NAND2_X1 U5965 ( .A1(n9732), .A2(n7904), .ZN(n9724) );
  AOI21_X1 U5966 ( .B1(n9731), .B2(n7882), .A(n4509), .ZN(n9715) );
  NAND2_X1 U5967 ( .A1(n4912), .A2(n7697), .ZN(n7880) );
  NAND2_X1 U5968 ( .A1(n7768), .A2(n7696), .ZN(n4912) );
  NAND2_X1 U5969 ( .A1(n7764), .A2(n4822), .ZN(n7901) );
  AND2_X1 U5970 ( .A1(n4929), .A2(n7496), .ZN(n7498) );
  NAND2_X1 U5971 ( .A1(n5574), .A2(n5573), .ZN(n7495) );
  INV_X1 U5972 ( .A(n6986), .ZN(n4580) );
  INV_X1 U5973 ( .A(n6987), .ZN(n4579) );
  AND2_X1 U5974 ( .A1(n9767), .A2(n6827), .ZN(n9750) );
  INV_X1 U5975 ( .A(n10096), .ZN(n6878) );
  NAND2_X1 U5976 ( .A1(n7041), .A2(n7922), .ZN(n10075) );
  NAND2_X1 U5977 ( .A1(n4824), .A2(n10136), .ZN(n4823) );
  INV_X1 U5978 ( .A(n5281), .ZN(n8385) );
  NAND2_X1 U5979 ( .A1(n9873), .A2(n4790), .ZN(n9879) );
  NOR2_X1 U5980 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4791) );
  OAI21_X1 U5981 ( .B1(n5906), .B2(n4835), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5251) );
  OAI21_X1 U5982 ( .B1(n4495), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  INV_X1 U5983 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8664) );
  INV_X1 U5984 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6331) );
  XNOR2_X1 U5985 ( .A(n5494), .B(n4608), .ZN(n6739) );
  INV_X1 U5986 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5987 ( .A1(n9872), .A2(n9957), .ZN(n4724) );
  XNOR2_X1 U5988 ( .A(n5504), .B(n5503), .ZN(n6555) );
  OAI21_X1 U5989 ( .B1(n8355), .B2(n4650), .A(n4542), .ZN(P2_U3244) );
  NAND2_X1 U5990 ( .A1(n4503), .A2(n6406), .ZN(n4650) );
  NAND2_X1 U5991 ( .A1(n4696), .A2(n4692), .ZN(n8979) );
  AND2_X1 U5992 ( .A1(n4578), .A2(n4577), .ZN(n9006) );
  OR2_X1 U5993 ( .A1(n9228), .A2(n10210), .ZN(n4578) );
  AOI21_X1 U5994 ( .B1(n9900), .B2(n9320), .A(n4726), .ZN(P2_U3518) );
  NOR2_X1 U5995 ( .A1(n9320), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U5996 ( .A1(n4501), .A2(n4537), .ZN(n4494) );
  NAND2_X1 U5997 ( .A1(n4943), .A2(n4945), .ZN(n4495) );
  OR2_X1 U5998 ( .A1(n9226), .A2(n9022), .ZN(n8330) );
  AND2_X1 U5999 ( .A1(n4991), .A2(n4571), .ZN(n4496) );
  NAND2_X1 U6000 ( .A1(n8315), .A2(n9065), .ZN(n9079) );
  INV_X1 U6001 ( .A(n9079), .ZN(n5027) );
  OR2_X1 U6002 ( .A1(n9278), .A2(n9153), .ZN(n4497) );
  OR2_X1 U6003 ( .A1(n9818), .A2(n9454), .ZN(n5760) );
  OR2_X1 U6004 ( .A1(n9255), .A2(n8394), .ZN(n4498) );
  AND2_X1 U6005 ( .A1(n9394), .A2(n4999), .ZN(n4499) );
  INV_X1 U6006 ( .A(n7882), .ZN(n4926) );
  AND2_X1 U6007 ( .A1(n9832), .A2(n9726), .ZN(n4500) );
  AND2_X1 U6008 ( .A1(n8285), .A2(n8284), .ZN(n4501) );
  NAND2_X1 U6009 ( .A1(n7976), .A2(n7975), .ZN(n9273) );
  AND2_X1 U6010 ( .A1(n4774), .A2(n7368), .ZN(n4502) );
  NAND2_X1 U6011 ( .A1(n8385), .A2(n9879), .ZN(n5556) );
  INV_X1 U6012 ( .A(n5556), .ZN(n4984) );
  OR2_X1 U6013 ( .A1(n8348), .A2(n4555), .ZN(n4503) );
  AND2_X1 U6014 ( .A1(n7879), .A2(n4913), .ZN(n4504) );
  INV_X1 U6015 ( .A(n7174), .ZN(n7156) );
  INV_X1 U6016 ( .A(n5034), .ZN(n6347) );
  NAND2_X1 U6017 ( .A1(n4917), .A2(n7086), .ZN(n7087) );
  AND2_X1 U6018 ( .A1(n7300), .A2(n7299), .ZN(n4505) );
  NAND2_X1 U6019 ( .A1(n5923), .A2(n5929), .ZN(n6257) );
  NAND2_X2 U6020 ( .A1(n6504), .A2(n6503), .ZN(n6634) );
  INV_X1 U6021 ( .A(n5554), .ZN(n5524) );
  INV_X2 U6022 ( .A(n5964), .ZN(n6125) );
  NOR2_X1 U6023 ( .A1(n5257), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6024 ( .A1(n5660), .A2(n4847), .ZN(n4506) );
  AND2_X1 U6025 ( .A1(n5125), .A2(n5124), .ZN(n4507) );
  AND2_X1 U6026 ( .A1(n4975), .A2(n7211), .ZN(n4508) );
  AND2_X1 U6027 ( .A1(n9741), .A2(n9727), .ZN(n4509) );
  OR3_X1 U6028 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n4510) );
  AND2_X1 U6029 ( .A1(n8230), .A2(n10253), .ZN(n4511) );
  AND2_X1 U6030 ( .A1(n8340), .A2(n8335), .ZN(n4512) );
  AND2_X1 U6032 ( .A1(n6302), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4513) );
  AND2_X1 U6033 ( .A1(n8245), .A2(n8331), .ZN(n4514) );
  OR2_X1 U6034 ( .A1(n6955), .A2(n6743), .ZN(n4515) );
  NAND2_X1 U6035 ( .A1(n9260), .A2(n9131), .ZN(n4516) );
  INV_X2 U6036 ( .A(n5568), .ZN(n5303) );
  INV_X1 U6037 ( .A(n8419), .ZN(n4592) );
  NOR2_X1 U6038 ( .A1(n7527), .A2(n8904), .ZN(n4517) );
  NAND4_X1 U6039 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n5941)
         );
  NAND2_X1 U6040 ( .A1(n7961), .A2(n7960), .ZN(n9278) );
  INV_X1 U6041 ( .A(n9278), .ZN(n4739) );
  NAND2_X1 U6042 ( .A1(n5668), .A2(n5667), .ZN(n9760) );
  NAND2_X1 U6043 ( .A1(n5256), .A2(n6260), .ZN(n9775) );
  INV_X1 U6044 ( .A(n9775), .ZN(n5265) );
  AND2_X1 U6045 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4518) );
  NAND2_X1 U6046 ( .A1(n4997), .A2(n4998), .ZN(n9469) );
  NAND2_X1 U6047 ( .A1(n5279), .A2(n5278), .ZN(n9777) );
  AND3_X1 U6048 ( .A1(n8329), .A2(n9018), .A3(n8323), .ZN(n4519) );
  OR2_X1 U6049 ( .A1(n8167), .A2(n6611), .ZN(n4520) );
  AND2_X1 U6050 ( .A1(n4998), .A2(n6157), .ZN(n4521) );
  AND2_X1 U6051 ( .A1(n5733), .A2(n7703), .ZN(n4522) );
  INV_X1 U6052 ( .A(n7918), .ZN(n4810) );
  NAND2_X1 U6053 ( .A1(n7939), .A2(n7938), .ZN(n9287) );
  AND2_X1 U6054 ( .A1(n7497), .A2(n7496), .ZN(n4523) );
  AND2_X1 U6055 ( .A1(n8004), .A2(n8003), .ZN(n4524) );
  AND2_X1 U6056 ( .A1(n8019), .A2(n8018), .ZN(n4525) );
  AND2_X1 U6057 ( .A1(n8146), .A2(n4893), .ZN(n4526) );
  AND2_X1 U6058 ( .A1(n4807), .A2(n4808), .ZN(n4527) );
  OR2_X1 U6059 ( .A1(n6744), .A2(n4593), .ZN(n4528) );
  NAND2_X1 U6061 ( .A1(n5353), .A2(n5352), .ZN(n9807) );
  INV_X1 U6062 ( .A(n7906), .ZN(n4812) );
  AND2_X1 U6063 ( .A1(n8282), .A2(n8283), .ZN(n8280) );
  INV_X1 U6064 ( .A(n8280), .ZN(n5054) );
  AND2_X1 U6065 ( .A1(n5809), .A2(n5804), .ZN(n9575) );
  INV_X1 U6066 ( .A(n9252), .ZN(n9083) );
  NAND2_X1 U6067 ( .A1(n8038), .A2(n8037), .ZN(n9252) );
  INV_X1 U6068 ( .A(n9448), .ZN(n4760) );
  INV_X1 U6069 ( .A(n4742), .ZN(n9070) );
  NOR2_X1 U6070 ( .A1(n9116), .A2(n4744), .ZN(n4742) );
  INV_X1 U6071 ( .A(n4784), .ZN(n9619) );
  NOR2_X1 U6072 ( .A1(n9658), .A2(n4786), .ZN(n4784) );
  INV_X1 U6073 ( .A(n4789), .ZN(n9561) );
  NOR2_X1 U6074 ( .A1(n4648), .A2(n8306), .ZN(n4530) );
  AND2_X1 U6075 ( .A1(n8278), .A2(n8277), .ZN(n8274) );
  AND2_X1 U6076 ( .A1(n6742), .A2(n4515), .ZN(n4531) );
  INV_X1 U6077 ( .A(n5058), .ZN(n5057) );
  NAND2_X1 U6078 ( .A1(n5061), .A2(n5062), .ZN(n5058) );
  AND2_X1 U6079 ( .A1(n4694), .A2(n4693), .ZN(n4532) );
  AND2_X1 U6080 ( .A1(n4501), .A2(n8274), .ZN(n4533) );
  AND2_X1 U6081 ( .A1(n6152), .A2(n6151), .ZN(n4534) );
  AND2_X1 U6082 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4535) );
  NOR2_X1 U6083 ( .A1(n9220), .A2(n8332), .ZN(n4536) );
  NAND2_X1 U6084 ( .A1(n8280), .A2(n8279), .ZN(n4537) );
  XNOR2_X1 U6085 ( .A(n9220), .B(n9002), .ZN(n8407) );
  INV_X1 U6086 ( .A(n5031), .ZN(n5030) );
  NAND2_X1 U6087 ( .A1(n4498), .A2(n8393), .ZN(n5031) );
  INV_X1 U6088 ( .A(n4625), .ZN(n4624) );
  INV_X1 U6089 ( .A(n5049), .ZN(n5048) );
  NOR2_X1 U6090 ( .A1(n4739), .A2(n9183), .ZN(n5049) );
  OR2_X1 U6091 ( .A1(n4921), .A2(n4500), .ZN(n4538) );
  NOR2_X1 U6092 ( .A1(n7487), .A2(n7486), .ZN(n4539) );
  OR2_X1 U6093 ( .A1(n5906), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4540) );
  AND2_X1 U6094 ( .A1(n5498), .A2(n5497), .ZN(n4541) );
  INV_X1 U6095 ( .A(n4738), .ZN(n4737) );
  NAND2_X1 U6096 ( .A1(n4740), .A2(n4739), .ZN(n4738) );
  AND2_X1 U6097 ( .A1(n4887), .A2(n4889), .ZN(n4542) );
  AND2_X1 U6098 ( .A1(n6379), .A2(n6233), .ZN(n4543) );
  INV_X1 U6099 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6364) );
  AND2_X1 U6100 ( .A1(n8212), .A2(n8249), .ZN(n8259) );
  INV_X1 U6101 ( .A(n8238), .ZN(n10241) );
  AND3_X1 U6102 ( .A1(n6651), .A2(n6650), .A3(n6649), .ZN(n8238) );
  AND2_X1 U6103 ( .A1(n5988), .A2(n5987), .ZN(n4544) );
  AND2_X1 U6104 ( .A1(n5134), .A2(SI_11_), .ZN(n4545) );
  NAND2_X1 U6105 ( .A1(n4657), .A2(n4656), .ZN(n4546) );
  AND2_X1 U6106 ( .A1(n9812), .A2(n9386), .ZN(n7913) );
  NOR2_X1 U6107 ( .A1(n9593), .A2(n9396), .ZN(n4547) );
  NOR2_X1 U6108 ( .A1(n7812), .A2(n7846), .ZN(n5060) );
  NAND2_X1 U6109 ( .A1(n8330), .A2(n8329), .ZN(n9001) );
  AND2_X1 U6110 ( .A1(n4934), .A2(n4940), .ZN(n4548) );
  OR2_X1 U6111 ( .A1(n5047), .A2(n5049), .ZN(n4549) );
  NAND2_X1 U6112 ( .A1(n7912), .A2(n4803), .ZN(n4550) );
  NAND2_X1 U6113 ( .A1(n9106), .A2(n4516), .ZN(n4551) );
  OR2_X1 U6114 ( .A1(n9792), .A2(n9614), .ZN(n4552) );
  OR2_X1 U6115 ( .A1(n6955), .A2(n6841), .ZN(n4553) );
  NOR2_X1 U6116 ( .A1(n7435), .A2(n8184), .ZN(n4554) );
  AND2_X1 U6117 ( .A1(n8350), .A2(n8349), .ZN(n4555) );
  NAND2_X1 U6118 ( .A1(n4909), .A2(n4908), .ZN(n9165) );
  INV_X1 U6119 ( .A(n7878), .ZN(n4916) );
  AND2_X1 U6120 ( .A1(n8292), .A2(n8291), .ZN(n4556) );
  AND2_X1 U6121 ( .A1(n7052), .A2(n6953), .ZN(n4557) );
  AND2_X1 U6122 ( .A1(n8150), .A2(n8206), .ZN(n4558) );
  INV_X1 U6123 ( .A(n5720), .ZN(n4658) );
  NAND2_X1 U6124 ( .A1(n4549), .A2(n5046), .ZN(n5042) );
  INV_X1 U6125 ( .A(n8336), .ZN(n4623) );
  INV_X1 U6126 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4945) );
  AND2_X1 U6127 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4559) );
  INV_X1 U6128 ( .A(n4806), .ZN(n4805) );
  NAND2_X1 U6129 ( .A1(n4808), .A2(n9575), .ZN(n4806) );
  OR2_X1 U6130 ( .A1(n4592), .A2(n4590), .ZN(n4560) );
  XNOR2_X1 U6131 ( .A(n6543), .B(n6542), .ZN(n6549) );
  INV_X1 U6132 ( .A(n9159), .ZN(n5045) );
  INV_X1 U6133 ( .A(n4943), .ZN(n5397) );
  XNOR2_X1 U6134 ( .A(n5234), .B(n5233), .ZN(n9323) );
  AND2_X1 U6135 ( .A1(n5179), .A2(n5178), .ZN(n5373) );
  INV_X1 U6136 ( .A(n7904), .ZN(n4817) );
  OAI21_X1 U6137 ( .B1(n7256), .B2(n7255), .A(n8258), .ZN(n7258) );
  OR2_X1 U6138 ( .A1(n10004), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4561) );
  INV_X1 U6139 ( .A(n9381), .ZN(n4759) );
  NAND2_X1 U6140 ( .A1(n4996), .A2(n6041), .ZN(n7485) );
  NAND2_X1 U6141 ( .A1(n4990), .A2(n4991), .ZN(n7654) );
  OR2_X1 U6142 ( .A1(n7258), .A2(n7257), .ZN(n4562) );
  AND4_X1 U6143 ( .A1(n5036), .A2(n6314), .A3(n5035), .A4(n6230), .ZN(n4563)
         );
  NAND2_X1 U6144 ( .A1(n5008), .A2(n6071), .ZN(n9403) );
  NOR2_X1 U6145 ( .A1(n9498), .A2(n9499), .ZN(n4564) );
  NOR2_X1 U6146 ( .A1(n8088), .A2(n8087), .ZN(n8089) );
  NOR2_X1 U6147 ( .A1(n7929), .A2(n7928), .ZN(n4565) );
  NAND2_X1 U6148 ( .A1(n9208), .A2(n4737), .ZN(n4741) );
  INV_X1 U6149 ( .A(n4964), .ZN(n4963) );
  NOR2_X1 U6150 ( .A1(n8074), .A2(n8807), .ZN(n4964) );
  AND2_X1 U6151 ( .A1(n4979), .A2(n4981), .ZN(n4566) );
  AND2_X1 U6152 ( .A1(n5362), .A2(n5179), .ZN(n4567) );
  NAND2_X1 U6153 ( .A1(n4563), .A2(n6313), .ZN(n5034) );
  AND2_X1 U6154 ( .A1(n7317), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4568) );
  AND2_X1 U6155 ( .A1(n7475), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U6156 ( .A1(n5019), .A2(n7157), .ZN(n7350) );
  AND2_X1 U6157 ( .A1(n7060), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U6158 ( .A1(n4772), .A2(n5976), .ZN(n6715) );
  NAND2_X1 U6159 ( .A1(n5001), .A2(n7116), .ZN(n7127) );
  NAND2_X1 U6160 ( .A1(n4943), .A2(n4941), .ZN(n5906) );
  NAND2_X1 U6161 ( .A1(n6052), .A2(n6053), .ZN(n4571) );
  AND2_X1 U6162 ( .A1(n7116), .A2(n6023), .ZN(n4572) );
  AND2_X1 U6163 ( .A1(n6549), .A2(n7011), .ZN(n10197) );
  INV_X1 U6164 ( .A(n5947), .ZN(n6588) );
  INV_X1 U6165 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5011) );
  INV_X1 U6166 ( .A(n7280), .ZN(n4731) );
  INV_X1 U6167 ( .A(n8178), .ZN(n4969) );
  AND2_X1 U6168 ( .A1(n8176), .A2(n8175), .ZN(n4573) );
  NAND2_X1 U6169 ( .A1(n6980), .A2(n6981), .ZN(n6979) );
  INV_X1 U6170 ( .A(n6979), .ZN(n4782) );
  AND2_X1 U6171 ( .A1(n6608), .A2(n6567), .ZN(n6568) );
  XNOR2_X1 U6172 ( .A(n6545), .B(n6544), .ZN(n8976) );
  INV_X1 U6173 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4651) );
  INV_X1 U6174 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4877) );
  INV_X1 U6175 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4688) );
  INV_X1 U6176 ( .A(n8343), .ZN(n4630) );
  AOI21_X1 U6177 ( .B1(n9894), .B2(n6570), .A(n9893), .ZN(n4727) );
  AOI21_X1 U6178 ( .B1(n9225), .B2(n9172), .A(n9005), .ZN(n4577) );
  INV_X2 U6179 ( .A(n10056), .ZN(n9735) );
  INV_X2 U6180 ( .A(n9327), .ZN(n9330) );
  NAND2_X2 U6181 ( .A1(n6808), .A2(n6807), .ZN(n10061) );
  NAND2_X1 U6182 ( .A1(n4980), .A2(n5033), .ZN(n6373) );
  NAND2_X1 U6183 ( .A1(n8140), .A2(n8310), .ZN(n9120) );
  NAND2_X1 U6184 ( .A1(n8149), .A2(n8319), .ZN(n9056) );
  NAND2_X1 U6185 ( .A1(n7791), .A2(n8282), .ZN(n8136) );
  OAI21_X1 U6186 ( .B1(n7681), .B2(n7680), .A(n8265), .ZN(n7748) );
  NAND2_X1 U6187 ( .A1(n10192), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U6188 ( .A1(n4907), .A2(n4905), .ZN(n9151) );
  INV_X1 U6189 ( .A(n9781), .ZN(n4824) );
  NAND2_X1 U6190 ( .A1(n10115), .A2(n6901), .ZN(n7030) );
  NAND2_X1 U6191 ( .A1(n4580), .A2(n4579), .ZN(n10115) );
  NAND2_X2 U6192 ( .A1(n7881), .A2(n5079), .ZN(n9731) );
  OAI22_X2 U6193 ( .A1(n9731), .A2(n4538), .B1(n4919), .B2(n4500), .ZN(n9684)
         );
  NAND2_X1 U6194 ( .A1(n9493), .A2(n6980), .ZN(n5827) );
  NAND2_X1 U6195 ( .A1(n4583), .A2(n5303), .ZN(n4582) );
  INV_X1 U6196 ( .A(n6838), .ZN(n4583) );
  NAND2_X1 U6197 ( .A1(n5126), .A2(n5125), .ZN(n5570) );
  NAND2_X1 U6198 ( .A1(n5083), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U6199 ( .A1(n7853), .A2(n6068), .ZN(n5008) );
  NAND2_X1 U6200 ( .A1(n4651), .A2(n4652), .ZN(n4610) );
  INV_X1 U6201 ( .A(n6041), .ZN(n4995) );
  NAND2_X1 U6202 ( .A1(n5104), .A2(SI_6_), .ZN(n5630) );
  NAND2_X1 U6203 ( .A1(n4989), .A2(n4987), .ZN(n6063) );
  NAND2_X1 U6204 ( .A1(n6929), .A2(n6930), .ZN(n6954) );
  NAND2_X1 U6205 ( .A1(n8868), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U6206 ( .A1(n8868), .A2(n8090), .ZN(n8420) );
  OAI211_X1 U6207 ( .C1(n8868), .C2(n4560), .A(n4587), .B(n4585), .ZN(n8131)
         );
  NAND2_X1 U6208 ( .A1(n6847), .A2(n4528), .ZN(n6754) );
  NAND2_X1 U6209 ( .A1(n8880), .A2(n8881), .ZN(n8879) );
  NAND2_X1 U6210 ( .A1(n7207), .A2(n7206), .ZN(n7212) );
  NAND2_X1 U6211 ( .A1(n7058), .A2(n7057), .ZN(n7207) );
  INV_X1 U6212 ( .A(n6373), .ZN(n4607) );
  NAND3_X1 U6213 ( .A1(n4607), .A2(n6239), .A3(n5064), .ZN(n6252) );
  XNOR2_X2 U6214 ( .A(n5098), .B(SI_4_), .ZN(n4608) );
  INV_X4 U6215 ( .A(n6554), .ZN(n6316) );
  NAND2_X1 U6216 ( .A1(n4613), .A2(n4611), .ZN(n8339) );
  NAND2_X1 U6217 ( .A1(n8330), .A2(n4626), .ZN(n4625) );
  NAND2_X1 U6218 ( .A1(n4634), .A2(n4636), .ZN(n8297) );
  NAND3_X1 U6219 ( .A1(n8276), .A2(n4635), .A3(n4494), .ZN(n4634) );
  NAND2_X1 U6220 ( .A1(n8288), .A2(n9202), .ZN(n4640) );
  NAND2_X1 U6221 ( .A1(n4641), .A2(n4642), .ZN(n8312) );
  NAND2_X1 U6222 ( .A1(n8307), .A2(n4644), .ZN(n4641) );
  NOR2_X1 U6223 ( .A1(n8143), .A2(n4646), .ZN(n4645) );
  NAND2_X1 U6224 ( .A1(n8308), .A2(n9128), .ZN(n4648) );
  NAND2_X1 U6225 ( .A1(n5719), .A2(n6207), .ZN(n4659) );
  NAND2_X1 U6226 ( .A1(n5718), .A2(n5792), .ZN(n4660) );
  NAND2_X1 U6227 ( .A1(n4661), .A2(n5928), .ZN(P1_U3240) );
  NAND2_X1 U6228 ( .A1(n4662), .A2(n5081), .ZN(n4661) );
  NAND2_X1 U6229 ( .A1(n4663), .A2(n4839), .ZN(n4662) );
  NAND2_X1 U6230 ( .A1(n4664), .A2(n5929), .ZN(n4663) );
  NAND2_X1 U6231 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6232 ( .A1(n5868), .A2(n5869), .ZN(n4666) );
  NAND2_X1 U6233 ( .A1(n5725), .A2(n5734), .ZN(n4669) );
  NAND4_X1 U6234 ( .A1(n4686), .A2(n5767), .A3(n5768), .A4(n9594), .ZN(n4685)
         );
  NAND4_X1 U6235 ( .A1(n5764), .A2(n5814), .A3(n9608), .A4(n5892), .ZN(n4686)
         );
  NAND3_X1 U6236 ( .A1(n4876), .A2(n4875), .A3(n4559), .ZN(n5520) );
  XNOR2_X1 U6237 ( .A(n8462), .B(n4689), .ZN(n8376) );
  NAND2_X1 U6238 ( .A1(n4725), .A2(n6240), .ZN(n6246) );
  AND3_X1 U6239 ( .A1(n4731), .A2(n10249), .A3(n7174), .ZN(n4733) );
  INV_X1 U6240 ( .A(n4741), .ZN(n9160) );
  INV_X1 U6241 ( .A(n4746), .ZN(n9048) );
  INV_X1 U6242 ( .A(n4750), .ZN(n4751) );
  XNOR2_X1 U6243 ( .A(n5959), .B(n5960), .ZN(n4750) );
  NAND2_X1 U6244 ( .A1(n6596), .A2(n4750), .ZN(n5963) );
  XNOR2_X1 U6245 ( .A(n6596), .B(n4751), .ZN(n6601) );
  INV_X1 U6246 ( .A(n6257), .ZN(n4764) );
  NAND2_X1 U6247 ( .A1(n5909), .A2(n4764), .ZN(n6482) );
  INV_X1 U6248 ( .A(n4765), .ZN(n5707) );
  NAND2_X1 U6249 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U6250 ( .A1(n6717), .A2(n4770), .ZN(n4768) );
  NAND2_X1 U6251 ( .A1(n4768), .A2(n4769), .ZN(n6786) );
  NAND3_X1 U6252 ( .A1(n5001), .A2(n4776), .A3(n7116), .ZN(n4773) );
  AND2_X1 U6254 ( .A1(n10048), .A2(n10096), .ZN(n6888) );
  MUX2_X1 U6255 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9882), .S(n6260), .Z(n6828) );
  OR2_X1 U6256 ( .A1(n5506), .A2(n5505), .ZN(n4780) );
  NAND2_X2 U6257 ( .A1(n6260), .A2(n6556), .ZN(n5568) );
  NOR2_X2 U6258 ( .A1(n6886), .A2(n6834), .ZN(n6981) );
  NOR2_X2 U6259 ( .A1(n9763), .A2(n9741), .ZN(n9716) );
  AND2_X2 U6260 ( .A1(n5246), .A2(n5247), .ZN(n4943) );
  INV_X1 U6261 ( .A(n4788), .ZN(n9604) );
  NAND2_X1 U6262 ( .A1(n9678), .A2(n4797), .ZN(n4795) );
  NAND2_X1 U6263 ( .A1(n9678), .A2(n4801), .ZN(n4796) );
  OAI21_X1 U6264 ( .B1(n9610), .B2(n4806), .A(n4804), .ZN(n4809) );
  NOR2_X1 U6265 ( .A1(n9610), .A2(n7916), .ZN(n9596) );
  INV_X1 U6266 ( .A(n4809), .ZN(n9566) );
  NAND3_X1 U6267 ( .A1(n9779), .A2(n9780), .A3(n4823), .ZN(n9856) );
  AOI21_X1 U6268 ( .B1(n7499), .B2(n4833), .A(n4831), .ZN(n4830) );
  NAND2_X1 U6269 ( .A1(n7287), .A2(n7499), .ZN(n4832) );
  INV_X1 U6270 ( .A(n7288), .ZN(n4833) );
  INV_X1 U6271 ( .A(n4836), .ZN(n4835) );
  NAND3_X1 U6272 ( .A1(n4836), .A2(n4943), .A3(n4834), .ZN(n5257) );
  OAI21_X1 U6273 ( .B1(n7700), .B2(n7699), .A(n7698), .ZN(n7702) );
  NAND2_X1 U6274 ( .A1(n5712), .A2(n5878), .ZN(n6870) );
  NAND2_X1 U6275 ( .A1(n7032), .A2(n7031), .ZN(n7034) );
  NAND2_X2 U6276 ( .A1(n5252), .A2(n5259), .ZN(n5922) );
  INV_X1 U6277 ( .A(n5506), .ZN(n5563) );
  AND2_X4 U6278 ( .A1(n5280), .A2(n8385), .ZN(n5647) );
  NAND2_X1 U6279 ( .A1(n5146), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U6280 ( .A1(n4851), .A2(n4567), .ZN(n5183) );
  NAND2_X1 U6281 ( .A1(n5126), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U6282 ( .A1(n4852), .A2(n4855), .ZN(n5475) );
  NAND2_X1 U6283 ( .A1(n5225), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6284 ( .A1(n5683), .A2(n4866), .ZN(n4864) );
  OR2_X1 U6285 ( .A1(n5683), .A2(n5199), .ZN(n4870) );
  MUX2_X1 U6286 ( .A(n5089), .B(n6611), .S(n6554), .Z(n5090) );
  NAND2_X2 U6287 ( .A1(n8235), .A2(n8234), .ZN(n8177) );
  NAND2_X1 U6288 ( .A1(n7182), .A2(n8234), .ZN(n7146) );
  OR2_X1 U6289 ( .A1(n8177), .A2(n7181), .ZN(n7182) );
  OAI21_X1 U6290 ( .B1(n7161), .B2(n4883), .A(n8217), .ZN(n4879) );
  NOR2_X1 U6291 ( .A1(n7161), .A2(n4884), .ZN(n4881) );
  NAND2_X1 U6292 ( .A1(n4886), .A2(n4888), .ZN(n4887) );
  XNOR2_X1 U6293 ( .A(n8174), .B(n8976), .ZN(n4886) );
  OAI22_X1 U6294 ( .A1(n6957), .A2(n6610), .B1(n6955), .B2(n6612), .ZN(n4891)
         );
  NAND2_X1 U6295 ( .A1(n9120), .A2(n8144), .ZN(n4892) );
  NAND2_X1 U6296 ( .A1(n9054), .A2(n4558), .ZN(n9017) );
  NAND2_X1 U6297 ( .A1(n9024), .A2(n4904), .ZN(n4902) );
  NAND2_X1 U6298 ( .A1(n9024), .A2(n8326), .ZN(n9000) );
  NAND2_X1 U6299 ( .A1(n9178), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U6300 ( .A1(n9756), .A2(n4915), .ZN(n7881) );
  NAND3_X1 U6301 ( .A1(n4917), .A2(n7086), .A3(n7088), .ZN(n7297) );
  AOI21_X2 U6302 ( .B1(n9684), .B2(n7885), .A(n7884), .ZN(n9670) );
  NAND2_X1 U6303 ( .A1(n7300), .A2(n4927), .ZN(n4929) );
  NAND2_X1 U6304 ( .A1(n9618), .A2(n4932), .ZN(n4931) );
  NAND2_X1 U6305 ( .A1(n4943), .A2(n4942), .ZN(n5253) );
  NAND2_X1 U6306 ( .A1(n4948), .A2(n4946), .ZN(n6541) );
  NAND2_X1 U6307 ( .A1(n6753), .A2(n6847), .ZN(n4951) );
  OAI21_X1 U6308 ( .B1(n8789), .B2(n4956), .A(n4954), .ZN(n8799) );
  NAND2_X1 U6309 ( .A1(n6954), .A2(n4557), .ZN(n7058) );
  NAND2_X1 U6310 ( .A1(n6536), .A2(n5033), .ZN(n4977) );
  NAND2_X1 U6311 ( .A1(n6588), .A2(n6590), .ZN(n5949) );
  NAND2_X1 U6312 ( .A1(n7406), .A2(n4496), .ZN(n4989) );
  NAND2_X1 U6313 ( .A1(n9426), .A2(n4499), .ZN(n4997) );
  NAND2_X1 U6314 ( .A1(n6786), .A2(n5005), .ZN(n5002) );
  NAND2_X1 U6315 ( .A1(n5002), .A2(n5003), .ZN(n6946) );
  NAND2_X1 U6316 ( .A1(n6945), .A2(n6006), .ZN(n6010) );
  INV_X1 U6317 ( .A(n6784), .ZN(n5006) );
  NAND2_X1 U6318 ( .A1(n5008), .A2(n5007), .ZN(n9404) );
  NAND3_X1 U6319 ( .A1(n5009), .A2(n9460), .A3(n6106), .ZN(n9373) );
  AOI21_X1 U6320 ( .B1(n9472), .B2(n5012), .A(n9334), .ZN(n6203) );
  NAND2_X1 U6321 ( .A1(n5013), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6561) );
  NAND2_X2 U6322 ( .A1(n9332), .A2(n6504), .ZN(n8083) );
  NAND2_X1 U6323 ( .A1(n7005), .A2(n5018), .ZN(n5017) );
  NAND2_X1 U6324 ( .A1(n5017), .A2(n5015), .ZN(n7248) );
  NAND2_X1 U6325 ( .A1(n9114), .A2(n5024), .ZN(n5023) );
  AND4_X2 U6326 ( .A1(n6314), .A2(n6230), .A3(n6232), .A4(n5035), .ZN(n5033)
         );
  NAND2_X1 U6327 ( .A1(n9159), .A2(n5042), .ZN(n5037) );
  INV_X1 U6328 ( .A(n8274), .ZN(n5061) );
  NAND2_X1 U6329 ( .A1(n7744), .A2(n5057), .ZN(n5055) );
  NAND3_X1 U6330 ( .A1(n5051), .A2(n5059), .A3(n5050), .ZN(n7813) );
  INV_X1 U6331 ( .A(n5053), .ZN(n5052) );
  NAND2_X1 U6332 ( .A1(n5071), .A2(n5070), .ZN(n7667) );
  NAND2_X1 U6333 ( .A1(n6249), .A2(n5072), .ZN(n6367) );
  INV_X1 U6334 ( .A(n6367), .ZN(n6366) );
  XNOR2_X1 U6335 ( .A(n5351), .B(n5350), .ZN(n8035) );
  NAND2_X1 U6336 ( .A1(n5351), .A2(n5350), .ZN(n5195) );
  OAI21_X2 U6337 ( .B1(n7891), .B2(n7890), .A(n5080), .ZN(n9618) );
  NAND2_X1 U6338 ( .A1(n8426), .A2(n8054), .ZN(n8061) );
  OAI22_X1 U6339 ( .A1(n6645), .A2(n6644), .B1(n6643), .B2(n6642), .ZN(n6746)
         );
  INV_X1 U6340 ( .A(n6504), .ZN(n8382) );
  NOR2_X1 U6341 ( .A1(n5604), .A2(n5599), .ZN(n5074) );
  OR2_X1 U6342 ( .A1(n6955), .A2(n8376), .ZN(n5075) );
  INV_X1 U6343 ( .A(n8220), .ZN(n8349) );
  INV_X1 U6344 ( .A(n9094), .ZN(n8394) );
  OR2_X1 U6345 ( .A1(n9676), .A2(n9388), .ZN(n5078) );
  OR2_X1 U6346 ( .A1(n9636), .A2(n9450), .ZN(n5080) );
  AND2_X1 U6347 ( .A1(n5912), .A2(n5911), .ZN(n5081) );
  AND2_X1 U6348 ( .A1(n5145), .A2(n5144), .ZN(n5082) );
  INV_X1 U6349 ( .A(n9121), .ZN(n8141) );
  INV_X1 U6350 ( .A(n6195), .ZN(n5909) );
  INV_X1 U6351 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9324) );
  AOI21_X1 U6352 ( .B1(n9014), .B2(n8099), .A(n8098), .ZN(n9036) );
  INV_X1 U6353 ( .A(n9034), .ZN(n8150) );
  INV_X1 U6354 ( .A(n9482), .ZN(n5264) );
  OAI21_X1 U6355 ( .B1(n8057), .B2(n9057), .A(n8831), .ZN(n8053) );
  INV_X1 U6356 ( .A(n8200), .ZN(n8344) );
  INV_X1 U6357 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U6358 ( .A1(n5794), .A2(n5863), .ZN(n5795) );
  AND2_X1 U6359 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  INV_X1 U6360 ( .A(n8053), .ZN(n8054) );
  NAND2_X1 U6361 ( .A1(n6817), .A2(n10052), .ZN(n5711) );
  AND2_X1 U6362 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n6623) );
  INV_X1 U6363 ( .A(n7980), .ZN(n6630) );
  INV_X1 U6364 ( .A(n7594), .ZN(n6627) );
  INV_X1 U6365 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6248) );
  INV_X1 U6366 ( .A(n5978), .ZN(n5979) );
  INV_X1 U6367 ( .A(n5977), .ZN(n5980) );
  INV_X1 U6368 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5620) );
  INV_X1 U6369 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6370 ( .A1(n6626), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U6371 ( .A1(n9226), .A2(n9022), .ZN(n8329) );
  NAND2_X1 U6372 ( .A1(n8065), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U6373 ( .A1(n6631), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8044) );
  AND2_X1 U6374 ( .A1(n9287), .A2(n8898), .ZN(n8389) );
  NAND2_X1 U6375 ( .A1(n6625), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6962) );
  INV_X1 U6376 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U6377 ( .A1(n6010), .A2(n6011), .ZN(n7115) );
  INV_X1 U6378 ( .A(n9406), .ZN(n6081) );
  NAND2_X1 U6379 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  NOR2_X1 U6380 ( .A1(n5687), .A2(n9395), .ZN(n5330) );
  NOR2_X1 U6381 ( .A1(n8637), .A2(n5422), .ZN(n5402) );
  NOR2_X1 U6382 ( .A1(n5649), .A2(n5648), .ZN(n5651) );
  INV_X1 U6383 ( .A(n7090), .ZN(n7088) );
  NAND2_X1 U6384 ( .A1(n5151), .A2(n8751), .ZN(n5154) );
  INV_X1 U6385 ( .A(n5640), .ZN(n5135) );
  AND2_X1 U6386 ( .A1(n7991), .A2(n7990), .ZN(n8788) );
  OR2_X1 U6387 ( .A1(n7950), .A2(n8949), .ZN(n7980) );
  AND2_X1 U6388 ( .A1(n8106), .A2(n8081), .ZN(n9038) );
  OR2_X1 U6389 ( .A1(n8009), .A2(n8800), .ZN(n8025) );
  AND2_X1 U6390 ( .A1(n8290), .A2(n8289), .ZN(n9202) );
  INV_X1 U6391 ( .A(n8976), .ZN(n9188) );
  AND2_X1 U6392 ( .A1(n8273), .A2(n8272), .ZN(n8190) );
  INV_X1 U6393 ( .A(n9576), .ZN(n9340) );
  NAND2_X1 U6394 ( .A1(n5342), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5689) );
  AND2_X1 U6395 ( .A1(n5319), .A2(n5318), .ZN(n9583) );
  NAND2_X1 U6396 ( .A1(n5402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5389) );
  INV_X1 U6397 ( .A(n5647), .ZN(n5421) );
  NOR2_X1 U6398 ( .A1(n9807), .A2(n9652), .ZN(n7890) );
  AND2_X1 U6399 ( .A1(n9818), .A2(n9680), .ZN(n7888) );
  NOR2_X1 U6400 ( .A1(n9828), .A2(n9710), .ZN(n7884) );
  INV_X1 U6401 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6402 ( .A1(n5103), .A2(SI_5_), .ZN(n5544) );
  XNOR2_X1 U6403 ( .A(n5086), .B(n5085), .ZN(n5501) );
  AND3_X1 U6404 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(n9094) );
  AND4_X1 U6405 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n8862)
         );
  AND2_X1 U6406 ( .A1(n8306), .A2(n9128), .ZN(n9152) );
  OR2_X1 U6407 ( .A1(n6725), .A2(n10212), .ZN(n10199) );
  AND2_X1 U6408 ( .A1(n7754), .A2(n10258), .ZN(n9297) );
  AND2_X1 U6409 ( .A1(n6354), .A2(n5034), .ZN(n6956) );
  INV_X1 U6410 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8462) );
  AND2_X1 U6411 ( .A1(n6496), .A2(n10139), .ZN(n9477) );
  NAND2_X1 U6412 ( .A1(n5524), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6413 ( .A1(n5524), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5490) );
  INV_X1 U6414 ( .A(n6991), .ZN(n10054) );
  INV_X1 U6415 ( .A(n9575), .ZN(n9573) );
  NAND2_X1 U6416 ( .A1(n5760), .A2(n7912), .ZN(n9663) );
  AND2_X1 U6417 ( .A1(n10064), .A2(n10145), .ZN(n9883) );
  OR2_X1 U6418 ( .A1(n6207), .A2(n6977), .ZN(n10145) );
  INV_X1 U6419 ( .A(n9093), .ZN(n9057) );
  INV_X1 U6420 ( .A(n8230), .ZN(n8907) );
  XNOR2_X1 U6421 ( .A(n8401), .B(n8407), .ZN(n9224) );
  INV_X1 U6422 ( .A(n6503), .ZN(n9332) );
  INV_X1 U6423 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6917) );
  INV_X1 U6424 ( .A(n9807), .ZN(n9636) );
  NAND2_X1 U6425 ( .A1(n6203), .A2(n6202), .ZN(n6227) );
  INV_X1 U6426 ( .A(n10169), .ZN(n10166) );
  INV_X1 U6427 ( .A(n10150), .ZN(n10149) );
  INV_X1 U6428 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8670) );
  AND2_X1 U6429 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6430 ( .A1(n6554), .A2(n5084), .ZN(n6547) );
  INV_X1 U6431 ( .A(SI_1_), .ZN(n5085) );
  MUX2_X1 U6432 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6316), .Z(n5502) );
  NAND2_X1 U6433 ( .A1(n5501), .A2(n5502), .ZN(n5088) );
  NAND2_X1 U6434 ( .A1(n5086), .A2(SI_1_), .ZN(n5087) );
  NAND2_X1 U6435 ( .A1(n5088), .A2(n5087), .ZN(n5510) );
  INV_X1 U6436 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6611) );
  INV_X1 U6437 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U6438 ( .A(n5090), .B(SI_2_), .ZN(n5509) );
  NAND2_X1 U6439 ( .A1(n5510), .A2(n5509), .ZN(n5093) );
  INV_X1 U6440 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6441 ( .A1(n5091), .A2(SI_2_), .ZN(n5092) );
  NAND2_X1 U6442 ( .A1(n5093), .A2(n5092), .ZN(n5562) );
  MUX2_X1 U6443 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6316), .Z(n5095) );
  INV_X1 U6444 ( .A(SI_3_), .ZN(n5094) );
  XNOR2_X1 U6445 ( .A(n5095), .B(n5094), .ZN(n5561) );
  NAND2_X1 U6446 ( .A1(n5562), .A2(n5561), .ZN(n5097) );
  NAND2_X1 U6447 ( .A1(n5095), .A2(SI_3_), .ZN(n5096) );
  INV_X1 U6448 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6740) );
  INV_X1 U6449 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6317) );
  BUF_X8 U6450 ( .A(n6316), .Z(n6556) );
  MUX2_X1 U6451 ( .A(n6740), .B(n6317), .S(n6556), .Z(n5098) );
  INV_X1 U6452 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6453 ( .A1(n5099), .A2(SI_4_), .ZN(n5100) );
  INV_X1 U6454 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6839) );
  INV_X1 U6455 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6327) );
  MUX2_X1 U6456 ( .A(n6839), .B(n6327), .S(n6556), .Z(n5102) );
  INV_X1 U6457 ( .A(n5102), .ZN(n5103) );
  MUX2_X1 U6458 ( .A(n6917), .B(n6331), .S(n6556), .Z(n5112) );
  INV_X1 U6459 ( .A(n5112), .ZN(n5104) );
  MUX2_X1 U6460 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6316), .Z(n5114) );
  NAND2_X1 U6461 ( .A1(n5114), .A2(SI_7_), .ZN(n5113) );
  MUX2_X1 U6462 ( .A(n6349), .B(n8664), .S(n6316), .Z(n5106) );
  INV_X1 U6463 ( .A(SI_8_), .ZN(n5105) );
  INV_X1 U6464 ( .A(n5106), .ZN(n5107) );
  INV_X1 U6465 ( .A(n5604), .ZN(n5109) );
  INV_X1 U6466 ( .A(n5113), .ZN(n5116) );
  INV_X1 U6467 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6362) );
  INV_X1 U6468 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6359) );
  MUX2_X1 U6469 ( .A(n6362), .B(n6359), .S(n6316), .Z(n5122) );
  INV_X1 U6470 ( .A(SI_9_), .ZN(n5121) );
  INV_X1 U6471 ( .A(n5122), .ZN(n5123) );
  NAND2_X1 U6472 ( .A1(n5123), .A2(SI_9_), .ZN(n5124) );
  NAND2_X1 U6473 ( .A1(n5581), .A2(n4507), .ZN(n5126) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5127) );
  MUX2_X1 U6475 ( .A(n5127), .B(n8670), .S(n6316), .Z(n5129) );
  INV_X1 U6476 ( .A(SI_10_), .ZN(n5128) );
  INV_X1 U6477 ( .A(n5129), .ZN(n5130) );
  NAND2_X1 U6478 ( .A1(n5130), .A2(SI_10_), .ZN(n5131) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6384) );
  INV_X1 U6480 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6377) );
  MUX2_X1 U6481 ( .A(n6384), .B(n6377), .S(n6316), .Z(n5133) );
  INV_X1 U6482 ( .A(n5133), .ZN(n5134) );
  INV_X1 U6483 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8475) );
  INV_X1 U6484 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6395) );
  MUX2_X1 U6485 ( .A(n8475), .B(n6395), .S(n6316), .Z(n5137) );
  INV_X1 U6486 ( .A(SI_12_), .ZN(n5136) );
  INV_X1 U6487 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6488 ( .A1(n5138), .A2(SI_12_), .ZN(n5139) );
  INV_X1 U6489 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6491) );
  INV_X1 U6490 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U6491 ( .A(n6491), .B(n6487), .S(n6316), .Z(n5142) );
  INV_X1 U6492 ( .A(SI_13_), .ZN(n5141) );
  NAND2_X1 U6493 ( .A1(n5142), .A2(n5141), .ZN(n5145) );
  INV_X1 U6494 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6495 ( .A1(n5143), .A2(SI_13_), .ZN(n5144) );
  INV_X1 U6496 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n8436) );
  INV_X1 U6497 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6502) );
  MUX2_X1 U6498 ( .A(n8436), .B(n6502), .S(n6556), .Z(n5147) );
  INV_X1 U6499 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6500 ( .A1(n5148), .A2(SI_14_), .ZN(n5149) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6701) );
  INV_X1 U6502 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6697) );
  MUX2_X1 U6503 ( .A(n6701), .B(n6697), .S(n6556), .Z(n5151) );
  INV_X1 U6504 ( .A(SI_15_), .ZN(n8751) );
  INV_X1 U6505 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6506 ( .A1(n5152), .A2(SI_15_), .ZN(n5153) );
  INV_X1 U6507 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5155) );
  INV_X1 U6508 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6714) );
  MUX2_X1 U6509 ( .A(n5155), .B(n6714), .S(n6556), .Z(n5157) );
  INV_X1 U6510 ( .A(SI_16_), .ZN(n5156) );
  NAND2_X1 U6511 ( .A1(n5157), .A2(n5156), .ZN(n5160) );
  INV_X1 U6512 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6513 ( .A1(n5158), .A2(SI_16_), .ZN(n5159) );
  INV_X1 U6514 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8667) );
  INV_X1 U6515 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6769) );
  MUX2_X1 U6516 ( .A(n8667), .B(n6769), .S(n6556), .Z(n5162) );
  XNOR2_X1 U6517 ( .A(n5162), .B(SI_17_), .ZN(n5407) );
  INV_X1 U6518 ( .A(n5407), .ZN(n5165) );
  INV_X1 U6519 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6520 ( .A1(n5163), .A2(SI_17_), .ZN(n5164) );
  MUX2_X1 U6521 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6556), .Z(n5167) );
  XNOR2_X1 U6522 ( .A(n5167), .B(SI_18_), .ZN(n5395) );
  INV_X1 U6523 ( .A(n5395), .ZN(n5166) );
  NAND2_X1 U6524 ( .A1(n5396), .A2(n5166), .ZN(n5169) );
  NAND2_X1 U6525 ( .A1(n5167), .A2(SI_18_), .ZN(n5168) );
  INV_X1 U6526 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6990) );
  INV_X1 U6527 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6993) );
  MUX2_X1 U6528 ( .A(n6990), .B(n6993), .S(n6556), .Z(n5171) );
  INV_X1 U6529 ( .A(SI_19_), .ZN(n5170) );
  NAND2_X1 U6530 ( .A1(n5171), .A2(n5170), .ZN(n5174) );
  INV_X1 U6531 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6532 ( .A1(n5172), .A2(SI_19_), .ZN(n5173) );
  NAND2_X1 U6533 ( .A1(n5174), .A2(n5173), .ZN(n5384) );
  INV_X1 U6534 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8364) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7101) );
  MUX2_X1 U6536 ( .A(n8364), .B(n7101), .S(n6556), .Z(n5176) );
  INV_X1 U6537 ( .A(SI_20_), .ZN(n5175) );
  NAND2_X1 U6538 ( .A1(n5176), .A2(n5175), .ZN(n5179) );
  INV_X1 U6539 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6540 ( .A1(n5177), .A2(SI_20_), .ZN(n5178) );
  INV_X1 U6541 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8006) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7125) );
  MUX2_X1 U6543 ( .A(n8006), .B(n7125), .S(n6556), .Z(n5180) );
  XNOR2_X1 U6544 ( .A(n5180), .B(SI_21_), .ZN(n5362) );
  INV_X1 U6545 ( .A(n5180), .ZN(n5181) );
  NAND2_X1 U6546 ( .A1(n5181), .A2(SI_21_), .ZN(n5182) );
  INV_X1 U6547 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8021) );
  INV_X1 U6548 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8379) );
  MUX2_X1 U6549 ( .A(n8021), .B(n8379), .S(n6556), .Z(n5185) );
  INV_X1 U6550 ( .A(SI_22_), .ZN(n5184) );
  NAND2_X1 U6551 ( .A1(n5185), .A2(n5184), .ZN(n5188) );
  INV_X1 U6552 ( .A(n5185), .ZN(n5186) );
  NAND2_X1 U6553 ( .A1(n5186), .A2(SI_22_), .ZN(n5187) );
  NAND2_X1 U6554 ( .A1(n5188), .A2(n5187), .ZN(n5338) );
  INV_X1 U6555 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8036) );
  INV_X1 U6556 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6557 ( .A(n8036), .B(n5189), .S(n6556), .Z(n5191) );
  INV_X1 U6558 ( .A(SI_23_), .ZN(n5190) );
  NAND2_X1 U6559 ( .A1(n5191), .A2(n5190), .ZN(n5194) );
  INV_X1 U6560 ( .A(n5191), .ZN(n5192) );
  NAND2_X1 U6561 ( .A1(n5192), .A2(SI_23_), .ZN(n5193) );
  AND2_X1 U6562 ( .A1(n5194), .A2(n5193), .ZN(n5350) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8041) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7507) );
  MUX2_X1 U6565 ( .A(n8041), .B(n7507), .S(n6556), .Z(n5196) );
  XNOR2_X1 U6566 ( .A(n5196), .B(SI_24_), .ZN(n5682) );
  INV_X1 U6567 ( .A(n5682), .ZN(n5199) );
  INV_X1 U6568 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6569 ( .A1(n5197), .A2(SI_24_), .ZN(n5198) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8444) );
  INV_X1 U6571 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7728) );
  MUX2_X1 U6572 ( .A(n8444), .B(n7728), .S(n6556), .Z(n5201) );
  INV_X1 U6573 ( .A(SI_25_), .ZN(n5200) );
  NAND2_X1 U6574 ( .A1(n5201), .A2(n5200), .ZN(n5204) );
  INV_X1 U6575 ( .A(n5201), .ZN(n5202) );
  NAND2_X1 U6576 ( .A1(n5202), .A2(SI_25_), .ZN(n5203) );
  NAND2_X1 U6577 ( .A1(n5204), .A2(n5203), .ZN(n5326) );
  INV_X1 U6578 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8076) );
  INV_X1 U6579 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7780) );
  MUX2_X1 U6580 ( .A(n8076), .B(n7780), .S(n6556), .Z(n5206) );
  INV_X1 U6581 ( .A(SI_26_), .ZN(n5205) );
  NAND2_X1 U6582 ( .A1(n5206), .A2(n5205), .ZN(n5209) );
  INV_X1 U6583 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6584 ( .A1(n5207), .A2(SI_26_), .ZN(n5208) );
  AND2_X1 U6585 ( .A1(n5209), .A2(n5208), .ZN(n5291) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8689) );
  INV_X1 U6587 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5210) );
  MUX2_X1 U6588 ( .A(n8689), .B(n5210), .S(n6556), .Z(n5212) );
  INV_X1 U6589 ( .A(SI_27_), .ZN(n5211) );
  NAND2_X1 U6590 ( .A1(n5212), .A2(n5211), .ZN(n5215) );
  INV_X1 U6591 ( .A(n5212), .ZN(n5213) );
  NAND2_X1 U6592 ( .A1(n5213), .A2(SI_27_), .ZN(n5214) );
  AND2_X1 U6593 ( .A1(n5215), .A2(n5214), .ZN(n5313) );
  INV_X1 U6594 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8417) );
  INV_X1 U6595 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8362) );
  MUX2_X1 U6596 ( .A(n8417), .B(n8362), .S(n6316), .Z(n5218) );
  XNOR2_X1 U6597 ( .A(n5218), .B(SI_28_), .ZN(n5301) );
  INV_X1 U6598 ( .A(SI_28_), .ZN(n5217) );
  NAND2_X1 U6599 ( .A1(n5218), .A2(n5217), .ZN(n5223) );
  MUX2_X1 U6600 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6554), .Z(n5275) );
  AND2_X1 U6601 ( .A1(n5223), .A2(n5275), .ZN(n5219) );
  NAND2_X1 U6602 ( .A1(n5224), .A2(n5219), .ZN(n5222) );
  INV_X1 U6603 ( .A(n5275), .ZN(n5220) );
  INV_X1 U6604 ( .A(SI_29_), .ZN(n5274) );
  OR2_X1 U6605 ( .A1(n5220), .A2(n5274), .ZN(n5221) );
  MUX2_X1 U6606 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6554), .Z(n5227) );
  NAND2_X1 U6607 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5231) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8166) );
  MUX2_X1 U6610 ( .A(n5231), .B(n8166), .S(n6554), .Z(n5232) );
  XNOR2_X1 U6611 ( .A(n5232), .B(SI_31_), .ZN(n5233) );
  MUX2_X1 U6612 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9323), .S(n6316), .Z(n5256) );
  NOR2_X1 U6613 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5238) );
  NOR2_X2 U6614 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5237) );
  NOR2_X2 U6615 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5236) );
  INV_X1 U6616 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5235) );
  NAND4_X1 U6617 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n5411)
         );
  NAND4_X1 U6618 ( .A1(n5240), .A2(n5412), .A3(n5410), .A4(n5239), .ZN(n5241)
         );
  NOR2_X1 U6619 ( .A1(n5411), .A2(n5241), .ZN(n5247) );
  AND2_X2 U6620 ( .A1(n5243), .A2(n5242), .ZN(n5495) );
  INV_X1 U6621 ( .A(n5409), .ZN(n5246) );
  NOR2_X1 U6622 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5249) );
  NOR2_X1 U6623 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5248) );
  INV_X1 U6624 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5915) );
  INV_X1 U6625 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8474) );
  OAI21_X1 U6626 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6627 ( .A1(n5918), .A2(n5254), .ZN(n5255) );
  XNOR2_X2 U6628 ( .A(n5255), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5924) );
  NAND2_X4 U6629 ( .A1(n5922), .A2(n5924), .ZN(n6260) );
  INV_X1 U6630 ( .A(n5258), .ZN(n9873) );
  INV_X1 U6631 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U6632 ( .A1(n5647), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5262) );
  INV_X2 U6633 ( .A(n4984), .ZN(n5693) );
  INV_X1 U6634 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6635 ( .A1(n5693), .A2(n5260), .ZN(n5261) );
  OAI211_X1 U6636 ( .C1(n4493), .C2(n5263), .A(n5262), .B(n5261), .ZN(n9482)
         );
  NAND2_X1 U6637 ( .A1(n8380), .A2(n5303), .ZN(n5268) );
  NAND2_X2 U6638 ( .A1(n4491), .A2(n6554), .ZN(n5506) );
  NAND2_X1 U6639 ( .A1(n5684), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5267) );
  INV_X1 U6640 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6641 ( .A1(n5647), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5271) );
  INV_X1 U6642 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5269) );
  OR2_X1 U6643 ( .A1(n5693), .A2(n5269), .ZN(n5270) );
  OAI211_X1 U6644 ( .C1(n4493), .C2(n5272), .A(n5271), .B(n5270), .ZN(n9483)
         );
  INV_X1 U6645 ( .A(n9483), .ZN(n5702) );
  OR2_X1 U6646 ( .A1(n9554), .A2(n5702), .ZN(n5273) );
  XNOR2_X1 U6647 ( .A(n5275), .B(n5274), .ZN(n5276) );
  NAND2_X1 U6648 ( .A1(n9329), .A2(n5303), .ZN(n5279) );
  NAND2_X1 U6649 ( .A1(n5684), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6650 ( .A1(n5647), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5290) );
  INV_X1 U6651 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9385) );
  INV_X1 U6652 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U6653 ( .A1(n5623), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5614) );
  INV_X1 U6654 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5589) );
  INV_X1 U6655 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6798) );
  INV_X1 U6656 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6657 ( .A1(n5651), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5481) );
  INV_X1 U6658 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5465) );
  INV_X1 U6659 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6660 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(n5669), .ZN(n5670) );
  INV_X1 U6661 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6662 ( .A1(n5366), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5355) );
  INV_X1 U6663 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U6664 ( .A1(n5330), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5317) );
  INV_X1 U6665 ( .A(n5317), .ZN(n5283) );
  NAND2_X1 U6666 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5283), .ZN(n5318) );
  INV_X1 U6667 ( .A(n5318), .ZN(n5284) );
  NAND2_X1 U6668 ( .A1(n5284), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7923) );
  INV_X1 U6669 ( .A(n7923), .ZN(n5285) );
  NAND2_X1 U6670 ( .A1(n4492), .A2(n5285), .ZN(n5289) );
  INV_X1 U6671 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5286) );
  OR2_X1 U6672 ( .A1(n5693), .A2(n5286), .ZN(n5288) );
  INV_X1 U6673 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7895) );
  OR2_X1 U6674 ( .A1(n4493), .A2(n7895), .ZN(n5287) );
  NAND4_X1 U6675 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n9568)
         );
  INV_X1 U6676 ( .A(n7921), .ZN(n5701) );
  NAND2_X1 U6677 ( .A1(n5684), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6678 ( .A1(n5647), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5300) );
  OAI21_X1 U6679 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5330), .A(n5317), .ZN(
        n5295) );
  INV_X1 U6680 ( .A(n5295), .ZN(n9591) );
  NAND2_X1 U6681 ( .A1(n4492), .A2(n9591), .ZN(n5299) );
  INV_X1 U6682 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8662) );
  OR2_X1 U6683 ( .A1(n5693), .A2(n8662), .ZN(n5298) );
  INV_X1 U6684 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5296) );
  OR2_X1 U6685 ( .A1(n4493), .A2(n5296), .ZN(n5297) );
  NAND4_X1 U6686 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n9614)
         );
  XNOR2_X1 U6687 ( .A(n9792), .B(n9396), .ZN(n9598) );
  NAND2_X1 U6688 ( .A1(n5684), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6689 ( .A1(n5647), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5312) );
  INV_X1 U6690 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U6691 ( .A1(n5318), .A2(n6212), .ZN(n5306) );
  NAND2_X1 U6692 ( .A1(n4492), .A2(n9562), .ZN(n5311) );
  INV_X1 U6693 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5307) );
  OR2_X1 U6694 ( .A1(n4493), .A2(n5307), .ZN(n5310) );
  INV_X1 U6695 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5308) );
  OR2_X1 U6696 ( .A1(n5693), .A2(n5308), .ZN(n5309) );
  NAND4_X1 U6697 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n9576)
         );
  INV_X1 U6698 ( .A(n9567), .ZN(n5700) );
  NAND2_X1 U6699 ( .A1(n5684), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6700 ( .A1(n5647), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5325) );
  INV_X1 U6701 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U6702 ( .A1(n9338), .A2(n5317), .ZN(n5319) );
  NAND2_X1 U6703 ( .A1(n4492), .A2(n9583), .ZN(n5324) );
  INV_X1 U6704 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6705 ( .A1(n5693), .A2(n5320), .ZN(n5323) );
  INV_X1 U6706 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6707 ( .A1(n4493), .A2(n5321), .ZN(n5322) );
  NAND4_X1 U6708 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n9600)
         );
  INV_X1 U6709 ( .A(n9600), .ZN(n6213) );
  NAND2_X1 U6710 ( .A1(n9789), .A2(n6213), .ZN(n5804) );
  NAND2_X1 U6711 ( .A1(n5684), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6712 ( .A1(n5647), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5336) );
  AOI21_X1 U6713 ( .B1(n9395), .B2(n5687), .A(n5330), .ZN(n9605) );
  NAND2_X1 U6714 ( .A1(n4492), .A2(n9605), .ZN(n5335) );
  INV_X1 U6715 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5331) );
  OR2_X1 U6716 ( .A1(n5693), .A2(n5331), .ZN(n5334) );
  INV_X1 U6717 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5332) );
  OR2_X1 U6718 ( .A1(n4493), .A2(n5332), .ZN(n5333) );
  NAND4_X1 U6719 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n9627)
         );
  INV_X1 U6720 ( .A(n9627), .ZN(n5337) );
  NAND2_X1 U6721 ( .A1(n9798), .A2(n5337), .ZN(n5773) );
  XNOR2_X1 U6722 ( .A(n5339), .B(n5338), .ZN(n8020) );
  NAND2_X1 U6723 ( .A1(n8020), .A2(n5303), .ZN(n5341) );
  NAND2_X1 U6724 ( .A1(n5684), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6725 ( .A1(n5647), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5349) );
  INV_X1 U6726 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9449) );
  INV_X1 U6727 ( .A(n5366), .ZN(n5343) );
  AOI21_X1 U6728 ( .B1(n9449), .B2(n5343), .A(n5342), .ZN(n9646) );
  NAND2_X1 U6729 ( .A1(n4492), .A2(n9646), .ZN(n5348) );
  INV_X1 U6730 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6731 ( .A1(n5693), .A2(n5344), .ZN(n5347) );
  INV_X1 U6732 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6733 ( .A1(n4493), .A2(n5345), .ZN(n5346) );
  NAND4_X1 U6734 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n9665)
         );
  INV_X1 U6735 ( .A(n9665), .ZN(n9386) );
  NOR2_X1 U6736 ( .A1(n9812), .A2(n9386), .ZN(n5759) );
  INV_X1 U6737 ( .A(n9651), .ZN(n5681) );
  NAND2_X1 U6738 ( .A1(n8035), .A2(n5303), .ZN(n5353) );
  NAND2_X1 U6739 ( .A1(n5684), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6740 ( .A1(n5647), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5361) );
  INV_X1 U6741 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9367) );
  AOI21_X1 U6742 ( .B1(n9367), .B2(n5355), .A(n5354), .ZN(n9634) );
  NAND2_X1 U6743 ( .A1(n4492), .A2(n9634), .ZN(n5360) );
  INV_X1 U6744 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6745 ( .A1(n5693), .A2(n5356), .ZN(n5359) );
  INV_X1 U6746 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5357) );
  OR2_X1 U6747 ( .A1(n4493), .A2(n5357), .ZN(n5358) );
  NAND4_X1 U6748 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n9652)
         );
  INV_X1 U6749 ( .A(n9652), .ZN(n9450) );
  NAND2_X1 U6750 ( .A1(n9807), .A2(n9450), .ZN(n5892) );
  NAND2_X1 U6751 ( .A1(n7914), .A2(n5892), .ZN(n9638) );
  XNOR2_X1 U6752 ( .A(n5363), .B(n5362), .ZN(n8005) );
  NAND2_X1 U6753 ( .A1(n8005), .A2(n5303), .ZN(n5365) );
  NAND2_X1 U6754 ( .A1(n5684), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6755 ( .A1(n5647), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5372) );
  AOI21_X1 U6756 ( .B1(n9385), .B2(n5377), .A(n5366), .ZN(n9660) );
  NAND2_X1 U6757 ( .A1(n4492), .A2(n9660), .ZN(n5371) );
  INV_X1 U6758 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5367) );
  OR2_X1 U6759 ( .A1(n5693), .A2(n5367), .ZN(n5370) );
  INV_X1 U6760 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5368) );
  OR2_X1 U6761 ( .A1(n4493), .A2(n5368), .ZN(n5369) );
  NAND4_X1 U6762 ( .A1(n5372), .A2(n5371), .A3(n5370), .A4(n5369), .ZN(n9680)
         );
  INV_X1 U6763 ( .A(n9680), .ZN(n9454) );
  NAND2_X1 U6764 ( .A1(n9818), .A2(n9454), .ZN(n7912) );
  XNOR2_X1 U6765 ( .A(n5374), .B(n5373), .ZN(n7992) );
  NAND2_X1 U6766 ( .A1(n7992), .A2(n5303), .ZN(n5376) );
  NAND2_X1 U6767 ( .A1(n5684), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6768 ( .A1(n5647), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5383) );
  INV_X1 U6769 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9438) );
  INV_X1 U6770 ( .A(n5377), .ZN(n5378) );
  AOI21_X1 U6771 ( .B1(n9438), .B2(n5389), .A(n5378), .ZN(n9674) );
  NAND2_X1 U6772 ( .A1(n4492), .A2(n9674), .ZN(n5382) );
  INV_X1 U6773 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8636) );
  OR2_X1 U6774 ( .A1(n4493), .A2(n8636), .ZN(n5381) );
  INV_X1 U6775 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5379) );
  OR2_X1 U6776 ( .A1(n5693), .A2(n5379), .ZN(n5380) );
  NAND4_X1 U6777 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n9693)
         );
  INV_X1 U6778 ( .A(n9693), .ZN(n9388) );
  AND2_X1 U6779 ( .A1(n9823), .A2(n9388), .ZN(n7910) );
  INV_X1 U6780 ( .A(n7910), .ZN(n5757) );
  XNOR2_X1 U6781 ( .A(n5385), .B(n5384), .ZN(n7972) );
  NAND2_X1 U6782 ( .A1(n7972), .A2(n5303), .ZN(n5388) );
  INV_X1 U6783 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5705) );
  XNOR2_X1 U6784 ( .A(n5706), .B(n5705), .ZN(n6991) );
  OAI22_X1 U6785 ( .A1(n5506), .A2(n6993), .B1(n6991), .B2(n6260), .ZN(n5386)
         );
  INV_X1 U6786 ( .A(n5386), .ZN(n5387) );
  OR2_X1 U6787 ( .A1(n5402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6788 ( .A1(n5390), .A2(n5389), .ZN(n9686) );
  INV_X1 U6789 ( .A(n4492), .ZN(n5423) );
  INV_X1 U6790 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U6791 ( .A1(n5524), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6792 ( .A1(n4984), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U6793 ( .C1(n5421), .C2(n9535), .A(n5392), .B(n5391), .ZN(n5393)
         );
  INV_X1 U6794 ( .A(n5393), .ZN(n5394) );
  OAI21_X1 U6795 ( .B1(n9686), .B2(n5423), .A(n5394), .ZN(n9710) );
  INV_X1 U6796 ( .A(n9710), .ZN(n9440) );
  NOR2_X1 U6797 ( .A1(n9828), .A2(n9440), .ZN(n5752) );
  XNOR2_X1 U6798 ( .A(n5396), .B(n5395), .ZN(n7959) );
  NAND2_X1 U6799 ( .A1(n7959), .A2(n5303), .ZN(n5401) );
  INV_X1 U6800 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U6801 ( .A1(n5397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5398) );
  XNOR2_X1 U6802 ( .A(n5398), .B(n4945), .ZN(n9539) );
  OAI22_X1 U6803 ( .A1(n5506), .A2(n6913), .B1(n6260), .B2(n9539), .ZN(n5399)
         );
  INV_X1 U6804 ( .A(n5399), .ZN(n5400) );
  INV_X1 U6805 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8433) );
  AOI21_X1 U6806 ( .B1(n8637), .B2(n5422), .A(n5402), .ZN(n9702) );
  NAND2_X1 U6807 ( .A1(n9702), .A2(n4492), .ZN(n5406) );
  NAND2_X1 U6808 ( .A1(n5647), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6809 ( .A1(n5524), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5403) );
  AND2_X1 U6810 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  OAI211_X1 U6811 ( .C1(n5693), .C2(n8433), .A(n5406), .B(n5405), .ZN(n9726)
         );
  INV_X1 U6812 ( .A(n9726), .ZN(n9420) );
  NAND2_X1 U6813 ( .A1(n9832), .A2(n9420), .ZN(n7906) );
  NAND2_X1 U6814 ( .A1(n5755), .A2(n7906), .ZN(n9709) );
  XNOR2_X1 U6815 ( .A(n5408), .B(n5407), .ZN(n7946) );
  NAND2_X1 U6816 ( .A1(n7946), .A2(n5303), .ZN(n5418) );
  NOR2_X1 U6817 ( .A1(n5546), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6818 ( .A1(n5634), .A2(n5410), .ZN(n5606) );
  OR2_X1 U6819 ( .A1(n5606), .A2(n5411), .ZN(n5662) );
  INV_X1 U6820 ( .A(n5662), .ZN(n5413) );
  NAND2_X1 U6821 ( .A1(n5413), .A2(n5412), .ZN(n5664) );
  OR2_X1 U6822 ( .A1(n5664), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6823 ( .A1(n5429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5414) );
  MUX2_X1 U6824 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5414), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5415) );
  NAND2_X1 U6825 ( .A1(n5415), .A2(n5397), .ZN(n9524) );
  OAI22_X1 U6826 ( .A1(n5506), .A2(n6769), .B1(n6260), .B2(n9524), .ZN(n5416)
         );
  INV_X1 U6827 ( .A(n5416), .ZN(n5417) );
  INV_X1 U6828 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U6829 ( .A1(n4984), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6830 ( .A1(n5524), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5419) );
  OAI211_X1 U6831 ( .C1(n5421), .C2(n9525), .A(n5420), .B(n5419), .ZN(n5425)
         );
  OAI21_X1 U6832 ( .B1(n5434), .B2(P1_REG3_REG_17__SCAN_IN), .A(n5422), .ZN(
        n9719) );
  NOR2_X1 U6833 ( .A1(n9719), .A2(n5423), .ZN(n5424) );
  OR2_X1 U6834 ( .A1(n5425), .A2(n5424), .ZN(n9738) );
  INV_X1 U6835 ( .A(n9738), .ZN(n9465) );
  AND2_X1 U6836 ( .A1(n9837), .A2(n9465), .ZN(n7905) );
  INV_X1 U6837 ( .A(n7905), .ZN(n5753) );
  OR2_X1 U6838 ( .A1(n9837), .A2(n9465), .ZN(n9705) );
  INV_X1 U6839 ( .A(n9723), .ZN(n5747) );
  XNOR2_X1 U6840 ( .A(n5427), .B(n5426), .ZN(n7937) );
  NAND2_X1 U6841 ( .A1(n7937), .A2(n5303), .ZN(n5433) );
  NAND2_X1 U6842 ( .A1(n5664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5428) );
  MUX2_X1 U6843 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5428), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5430) );
  NAND2_X1 U6844 ( .A1(n5430), .A2(n5429), .ZN(n9515) );
  OAI22_X1 U6845 ( .A1(n5506), .A2(n6714), .B1(n6260), .B2(n9515), .ZN(n5431)
         );
  INV_X1 U6846 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U6847 ( .A1(n5647), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5441) );
  AOI21_X1 U6848 ( .B1(n5670), .B2(n5435), .A(n5434), .ZN(n9745) );
  NAND2_X1 U6849 ( .A1(n4492), .A2(n9745), .ZN(n5440) );
  INV_X1 U6850 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5436) );
  OR2_X1 U6851 ( .A1(n5693), .A2(n5436), .ZN(n5439) );
  INV_X1 U6852 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5437) );
  OR2_X1 U6853 ( .A1(n4493), .A2(n5437), .ZN(n5438) );
  NAND4_X1 U6854 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n9727)
         );
  INV_X1 U6855 ( .A(n9727), .ZN(n9754) );
  NAND2_X1 U6856 ( .A1(n9741), .A2(n9754), .ZN(n7904) );
  NAND2_X1 U6857 ( .A1(n5853), .A2(n7904), .ZN(n7882) );
  XNOR2_X1 U6858 ( .A(n5443), .B(n5442), .ZN(n7785) );
  NAND2_X1 U6859 ( .A1(n7785), .A2(n5303), .ZN(n5449) );
  NOR2_X1 U6860 ( .A1(n5608), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5583) );
  INV_X1 U6861 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5444) );
  AND2_X1 U6862 ( .A1(n5583), .A2(n5444), .ZN(n5642) );
  INV_X1 U6863 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6864 ( .A1(n5642), .A2(n5445), .ZN(n5476) );
  OR2_X1 U6865 ( .A1(n5476), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U6866 ( .A1(n5446), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  INV_X1 U6867 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6868 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U6869 ( .A1(n5461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5447) );
  XNOR2_X1 U6870 ( .A(n5447), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6289) );
  AOI22_X1 U6871 ( .A1(n5507), .A2(n6289), .B1(n5684), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6872 ( .A1(n5647), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6873 ( .A1(n5467), .A2(n5450), .ZN(n5451) );
  NOR2_X1 U6874 ( .A1(n5669), .A2(n5451), .ZN(n9345) );
  NAND2_X1 U6875 ( .A1(n4492), .A2(n9345), .ZN(n5456) );
  INV_X1 U6876 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5452) );
  OR2_X1 U6877 ( .A1(n5693), .A2(n5452), .ZN(n5455) );
  INV_X1 U6878 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5453) );
  OR2_X1 U6879 ( .A1(n4493), .A2(n5453), .ZN(n5454) );
  NAND4_X1 U6880 ( .A1(n5457), .A2(n5456), .A3(n5455), .A4(n5454), .ZN(n9484)
         );
  INV_X1 U6881 ( .A(n9484), .ZN(n9753) );
  NAND2_X1 U6882 ( .A1(n9357), .A2(n9753), .ZN(n5848) );
  NAND2_X1 U6883 ( .A1(n7900), .A2(n5848), .ZN(n7879) );
  XNOR2_X1 U6884 ( .A(n5458), .B(n5082), .ZN(n7622) );
  NAND2_X1 U6885 ( .A1(n7622), .A2(n5303), .ZN(n5464) );
  OR2_X1 U6886 ( .A1(n5460), .A2(n5459), .ZN(n5462) );
  AND2_X1 U6887 ( .A1(n5462), .A2(n5461), .ZN(n7342) );
  AOI22_X1 U6888 ( .A1(n5684), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5507), .B2(
        n7342), .ZN(n5463) );
  NAND2_X1 U6889 ( .A1(n5647), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6890 ( .A1(n5481), .A2(n5465), .ZN(n5466) );
  AND2_X1 U6891 ( .A1(n5467), .A2(n5466), .ZN(n7774) );
  NAND2_X1 U6892 ( .A1(n4492), .A2(n7774), .ZN(n5472) );
  INV_X1 U6893 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5468) );
  OR2_X1 U6894 ( .A1(n5693), .A2(n5468), .ZN(n5471) );
  INV_X1 U6895 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5469) );
  OR2_X1 U6896 ( .A1(n4493), .A2(n5469), .ZN(n5470) );
  NAND4_X1 U6897 ( .A1(n5473), .A2(n5472), .A3(n5471), .A4(n5470), .ZN(n9485)
         );
  INV_X1 U6898 ( .A(n9485), .ZN(n9348) );
  OR2_X1 U6899 ( .A1(n9848), .A2(n9348), .ZN(n5726) );
  NAND2_X1 U6900 ( .A1(n9848), .A2(n9348), .ZN(n7703) );
  XNOR2_X1 U6901 ( .A(n5475), .B(n5474), .ZN(n7575) );
  NAND2_X1 U6902 ( .A1(n7575), .A2(n5303), .ZN(n5480) );
  NAND2_X1 U6903 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U6904 ( .A(n5477), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6288) );
  INV_X1 U6905 ( .A(n6288), .ZN(n7107) );
  OAI22_X1 U6906 ( .A1(n5506), .A2(n6395), .B1(n7107), .B2(n6260), .ZN(n5478)
         );
  INV_X1 U6907 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U6908 ( .A1(n5647), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5487) );
  OR2_X1 U6909 ( .A1(n5651), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5482) );
  AND2_X1 U6910 ( .A1(n5482), .A2(n5481), .ZN(n7518) );
  NAND2_X1 U6911 ( .A1(n4492), .A2(n7518), .ZN(n5486) );
  INV_X1 U6912 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6913 ( .A1(n5693), .A2(n5483), .ZN(n5485) );
  INV_X1 U6914 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6261) );
  OR2_X1 U6915 ( .A1(n4493), .A2(n6261), .ZN(n5484) );
  NAND4_X1 U6916 ( .A1(n5487), .A2(n5486), .A3(n5485), .A4(n5484), .ZN(n9486)
         );
  INV_X1 U6917 ( .A(n9486), .ZN(n7766) );
  OR2_X1 U6918 ( .A1(n7692), .A2(n7766), .ZN(n5734) );
  NAND2_X1 U6919 ( .A1(n7692), .A2(n7766), .ZN(n7701) );
  NAND2_X1 U6920 ( .A1(n5734), .A2(n7701), .ZN(n7694) );
  NAND2_X1 U6921 ( .A1(n5647), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5493) );
  INV_X1 U6922 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5488) );
  XNOR2_X1 U6923 ( .A(n5488), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6719) );
  INV_X1 U6924 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5489) );
  OR2_X1 U6925 ( .A1(n5556), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U6926 ( .A1(n5563), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5498) );
  OR2_X1 U6927 ( .A1(n5495), .A2(n9872), .ZN(n5496) );
  XNOR2_X1 U6928 ( .A(n5496), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U6929 ( .A1(n5507), .A2(n6284), .ZN(n5497) );
  NAND2_X1 U6930 ( .A1(n6898), .A2(n6834), .ZN(n5820) );
  NAND2_X1 U6931 ( .A1(n9494), .A2(n6897), .ZN(n5879) );
  INV_X1 U6932 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5499) );
  INV_X1 U6933 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5500) );
  INV_X1 U6934 ( .A(n5501), .ZN(n5504) );
  INV_X1 U6935 ( .A(n5502), .ZN(n5503) );
  INV_X1 U6936 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6937 ( .A1(n5524), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5952) );
  NAND2_X1 U6938 ( .A1(n4492), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U6939 ( .A1(n5647), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5954) );
  INV_X1 U6940 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5508) );
  OR2_X1 U6941 ( .A1(n5556), .A2(n5508), .ZN(n5951) );
  INV_X1 U6942 ( .A(n10059), .ZN(n9496) );
  XNOR2_X1 U6943 ( .A(n5510), .B(n5509), .ZN(n6610) );
  NAND2_X1 U6944 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5564), .ZN(n5511) );
  XNOR2_X1 U6945 ( .A(n5511), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U6946 ( .A1(n5507), .A2(n9946), .ZN(n5512) );
  NAND2_X1 U6947 ( .A1(n10059), .A2(n6878), .ZN(n5713) );
  NAND2_X1 U6948 ( .A1(n4492), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U6949 ( .A1(n5647), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5516) );
  INV_X1 U6950 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5513) );
  INV_X1 U6951 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10077) );
  INV_X1 U6952 ( .A(SI_0_), .ZN(n5519) );
  INV_X1 U6953 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5518) );
  OAI21_X1 U6954 ( .B1(n6554), .B2(n5519), .A(n5518), .ZN(n5521) );
  AND2_X1 U6955 ( .A1(n5521), .A2(n5520), .ZN(n9882) );
  INV_X1 U6956 ( .A(n6828), .ZN(n10050) );
  NAND2_X1 U6957 ( .A1(n5941), .A2(n10050), .ZN(n5877) );
  NAND2_X1 U6958 ( .A1(n10055), .A2(n5877), .ZN(n6483) );
  NOR4_X1 U6959 ( .A1(n6895), .A2(n6816), .A3(n6871), .A4(n6483), .ZN(n5569)
         );
  NAND2_X1 U6960 ( .A1(n5647), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5528) );
  AOI21_X1 U6961 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U6962 ( .A1(n5522), .A2(n5537), .ZN(n6707) );
  NAND2_X1 U6963 ( .A1(n4492), .A2(n6707), .ZN(n5527) );
  INV_X1 U6964 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5523) );
  INV_X1 U6965 ( .A(n9493), .ZN(n6790) );
  NAND2_X1 U6966 ( .A1(n5684), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6967 ( .A1(n5495), .A2(n5531), .ZN(n5532) );
  NAND2_X1 U6968 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5533) );
  MUX2_X1 U6969 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5533), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5534) );
  AND2_X1 U6970 ( .A1(n5534), .A2(n5546), .ZN(n9978) );
  NAND2_X1 U6971 ( .A1(n5507), .A2(n9978), .ZN(n5535) );
  NAND2_X1 U6972 ( .A1(n6790), .A2(n6985), .ZN(n5823) );
  NAND2_X1 U6973 ( .A1(n5647), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5543) );
  OAI21_X1 U6974 ( .B1(n5537), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5621), .ZN(
        n6789) );
  INV_X1 U6975 ( .A(n6789), .ZN(n6906) );
  NAND2_X1 U6976 ( .A1(n4492), .A2(n6906), .ZN(n5542) );
  INV_X1 U6977 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5538) );
  OR2_X1 U6978 ( .A1(n4493), .A2(n5538), .ZN(n5541) );
  INV_X1 U6979 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5539) );
  OR2_X1 U6980 ( .A1(n5693), .A2(n5539), .ZN(n5540) );
  NAND4_X1 U6981 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n9492)
         );
  NAND2_X1 U6982 ( .A1(n5684), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6983 ( .A1(n5546), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5547) );
  MUX2_X1 U6984 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5547), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5549) );
  INV_X1 U6985 ( .A(n5634), .ZN(n5548) );
  NAND2_X1 U6986 ( .A1(n5549), .A2(n5548), .ZN(n6330) );
  INV_X1 U6987 ( .A(n6330), .ZN(n9996) );
  NAND2_X1 U6988 ( .A1(n5507), .A2(n9996), .ZN(n5550) );
  NAND2_X1 U6989 ( .A1(n7037), .A2(n6907), .ZN(n5875) );
  NAND2_X1 U6990 ( .A1(n9492), .A2(n4781), .ZN(n5826) );
  NAND2_X1 U6991 ( .A1(n5647), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5560) );
  INV_X1 U6992 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U6993 ( .A1(n4492), .A2(n6499), .ZN(n5559) );
  INV_X1 U6994 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5553) );
  OR2_X1 U6995 ( .A1(n4493), .A2(n5553), .ZN(n5558) );
  INV_X1 U6996 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5555) );
  OR2_X1 U6997 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  XNOR2_X1 U6998 ( .A(n5562), .B(n5561), .ZN(n6646) );
  NAND2_X1 U6999 ( .A1(n5563), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5567) );
  OAI21_X1 U7000 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(n5564), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5565) );
  XNOR2_X1 U7001 ( .A(n5565), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7002 ( .A1(n5507), .A2(n6302), .ZN(n5566) );
  OAI211_X1 U7003 ( .C1(n6646), .C2(n5568), .A(n5567), .B(n5566), .ZN(n6889)
         );
  XNOR2_X1 U7004 ( .A(n9495), .B(n6887), .ZN(n6822) );
  INV_X1 U7005 ( .A(n6822), .ZN(n6883) );
  NAND4_X1 U7006 ( .A1(n5569), .A2(n6986), .A3(n7029), .A4(n6883), .ZN(n5639)
         );
  XNOR2_X1 U7007 ( .A(n5570), .B(n5077), .ZN(n7316) );
  NAND2_X1 U7008 ( .A1(n7316), .A2(n5303), .ZN(n5574) );
  OR2_X1 U7009 ( .A1(n5583), .A2(n9872), .ZN(n5571) );
  XNOR2_X1 U7010 ( .A(n5571), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6803) );
  INV_X1 U7011 ( .A(n6803), .ZN(n6375) );
  OAI22_X1 U7012 ( .A1(n5506), .A2(n8670), .B1(n6260), .B2(n6375), .ZN(n5572)
         );
  INV_X1 U7013 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7014 ( .A1(n5591), .A2(n6798), .ZN(n5575) );
  AND2_X1 U7015 ( .A1(n5649), .A2(n5575), .ZN(n7306) );
  NAND2_X1 U7016 ( .A1(n4492), .A2(n7306), .ZN(n5580) );
  NAND2_X1 U7017 ( .A1(n5647), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5579) );
  INV_X1 U7018 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7307) );
  OR2_X1 U7019 ( .A1(n4493), .A2(n7307), .ZN(n5578) );
  INV_X1 U7020 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5576) );
  OR2_X1 U7021 ( .A1(n5693), .A2(n5576), .ZN(n5577) );
  NAND4_X1 U7022 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n9488)
         );
  INV_X1 U7023 ( .A(n9488), .ZN(n7409) );
  NAND2_X1 U7024 ( .A1(n7495), .A2(n7409), .ZN(n7291) );
  XNOR2_X1 U7025 ( .A(n5581), .B(n4507), .ZN(n7213) );
  NAND2_X1 U7026 ( .A1(n7213), .A2(n5303), .ZN(n5588) );
  NAND2_X1 U7027 ( .A1(n5608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  MUX2_X1 U7028 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5582), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5585) );
  INV_X1 U7029 ( .A(n5583), .ZN(n5584) );
  AND2_X1 U7030 ( .A1(n5585), .A2(n5584), .ZN(n6687) );
  INV_X1 U7031 ( .A(n6687), .ZN(n6360) );
  OAI22_X1 U7032 ( .A1(n5506), .A2(n6359), .B1(n6260), .B2(n6360), .ZN(n5586)
         );
  INV_X1 U7033 ( .A(n5586), .ZN(n5587) );
  NAND2_X1 U7034 ( .A1(n5647), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7035 ( .A1(n5614), .A2(n5589), .ZN(n5590) );
  AND2_X1 U7036 ( .A1(n5591), .A2(n5590), .ZN(n7460) );
  NAND2_X1 U7037 ( .A1(n4492), .A2(n7460), .ZN(n5596) );
  INV_X1 U7038 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5592) );
  OR2_X1 U7039 ( .A1(n5693), .A2(n5592), .ZN(n5595) );
  INV_X1 U7040 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5593) );
  OR2_X1 U7041 ( .A1(n4493), .A2(n5593), .ZN(n5594) );
  NAND4_X1 U7042 ( .A1(n5597), .A2(n5596), .A3(n5595), .A4(n5594), .ZN(n9489)
         );
  INV_X1 U7043 ( .A(n9489), .ZN(n7376) );
  NAND2_X1 U7044 ( .A1(n10138), .A2(n7376), .ZN(n7455) );
  NAND2_X1 U7045 ( .A1(n7291), .A2(n7455), .ZN(n5833) );
  AND2_X1 U7046 ( .A1(n5628), .A2(n5599), .ZN(n5598) );
  NAND2_X1 U7047 ( .A1(n5629), .A2(n5598), .ZN(n5603) );
  INV_X1 U7048 ( .A(n5599), .ZN(n5601) );
  OR2_X1 U7049 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  NAND2_X1 U7050 ( .A1(n5603), .A2(n5602), .ZN(n5605) );
  XNOR2_X1 U7051 ( .A(n5605), .B(n5604), .ZN(n7059) );
  NAND2_X1 U7052 ( .A1(n7059), .A2(n5303), .ZN(n5612) );
  NAND2_X1 U7053 ( .A1(n5606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5607) );
  MUX2_X1 U7054 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5607), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5609) );
  NAND2_X1 U7055 ( .A1(n5609), .A2(n5608), .ZN(n6350) );
  OAI22_X1 U7056 ( .A1(n5506), .A2(n8664), .B1(n6260), .B2(n6350), .ZN(n5610)
         );
  INV_X1 U7057 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7058 ( .A1(n5612), .A2(n5611), .ZN(n7295) );
  INV_X1 U7059 ( .A(n7295), .ZN(n10131) );
  NAND2_X1 U7060 ( .A1(n5647), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5619) );
  OR2_X1 U7061 ( .A1(n5623), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5613) );
  AND2_X1 U7062 ( .A1(n5614), .A2(n5613), .ZN(n7093) );
  NAND2_X1 U7063 ( .A1(n4492), .A2(n7093), .ZN(n5618) );
  INV_X1 U7064 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7094) );
  OR2_X1 U7065 ( .A1(n4493), .A2(n7094), .ZN(n5617) );
  INV_X1 U7066 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5615) );
  OR2_X1 U7067 ( .A1(n5693), .A2(n5615), .ZN(n5616) );
  NAND4_X1 U7068 ( .A1(n5619), .A2(n5618), .A3(n5617), .A4(n5616), .ZN(n9490)
         );
  NAND2_X1 U7069 ( .A1(n10131), .A2(n9490), .ZN(n7463) );
  INV_X1 U7070 ( .A(n9490), .ZN(n7038) );
  NAND2_X1 U7071 ( .A1(n7295), .A2(n7038), .ZN(n7288) );
  NAND2_X1 U7072 ( .A1(n5647), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5627) );
  AND2_X1 U7073 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NOR2_X1 U7074 ( .A1(n5623), .A2(n5622), .ZN(n6949) );
  NAND2_X1 U7075 ( .A1(n4492), .A2(n6949), .ZN(n5626) );
  OR2_X1 U7076 ( .A1(n5693), .A2(n10129), .ZN(n5625) );
  INV_X1 U7077 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7043) );
  OR2_X1 U7078 ( .A1(n4493), .A2(n7043), .ZN(n5624) );
  NAND4_X1 U7079 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(n9491)
         );
  INV_X1 U7080 ( .A(n9491), .ZN(n7085) );
  NAND2_X1 U7081 ( .A1(n5629), .A2(n5628), .ZN(n5631) );
  NAND2_X1 U7082 ( .A1(n5631), .A2(n5630), .ZN(n5633) );
  XNOR2_X1 U7083 ( .A(n5633), .B(n5632), .ZN(n6958) );
  NAND2_X1 U7084 ( .A1(n6958), .A2(n5303), .ZN(n5638) );
  INV_X1 U7085 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6358) );
  OR2_X1 U7086 ( .A1(n5634), .A2(n9872), .ZN(n5635) );
  XNOR2_X1 U7087 ( .A(n5635), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10004) );
  INV_X1 U7088 ( .A(n10004), .ZN(n6356) );
  OAI22_X1 U7089 ( .A1(n5506), .A2(n6358), .B1(n6260), .B2(n6356), .ZN(n5636)
         );
  INV_X1 U7090 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U7091 ( .A1(n7085), .A2(n7045), .ZN(n7078) );
  INV_X1 U7092 ( .A(n7045), .ZN(n10125) );
  NAND2_X1 U7093 ( .A1(n10125), .A2(n9491), .ZN(n5884) );
  NAND2_X1 U7094 ( .A1(n7078), .A2(n5884), .ZN(n7083) );
  OR4_X1 U7095 ( .A1(n5639), .A2(n5833), .A3(n7088), .A4(n7083), .ZN(n5658) );
  NAND2_X1 U7096 ( .A1(n7418), .A2(n5303), .ZN(n5646) );
  OR2_X1 U7097 ( .A1(n5642), .A2(n9872), .ZN(n5643) );
  XNOR2_X1 U7098 ( .A(n5643), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10026) );
  INV_X1 U7099 ( .A(n10026), .ZN(n6378) );
  OAI22_X1 U7100 ( .A1(n5506), .A2(n6377), .B1(n6260), .B2(n6378), .ZN(n5644)
         );
  INV_X1 U7101 ( .A(n5644), .ZN(n5645) );
  NAND2_X1 U7102 ( .A1(n5647), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5657) );
  AND2_X1 U7103 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  NOR2_X1 U7104 ( .A1(n5651), .A2(n5650), .ZN(n7536) );
  NAND2_X1 U7105 ( .A1(n4492), .A2(n7536), .ZN(n5656) );
  INV_X1 U7106 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5652) );
  OR2_X1 U7107 ( .A1(n5693), .A2(n5652), .ZN(n5655) );
  INV_X1 U7108 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5653) );
  OR2_X1 U7109 ( .A1(n4493), .A2(n5653), .ZN(n5654) );
  NAND4_X1 U7110 ( .A1(n5657), .A2(n5656), .A3(n5655), .A4(n5654), .ZN(n9487)
         );
  INV_X1 U7111 ( .A(n9487), .ZN(n7491) );
  OR2_X1 U7112 ( .A1(n7535), .A2(n7491), .ZN(n7512) );
  NAND2_X1 U7113 ( .A1(n7535), .A2(n7491), .ZN(n7511) );
  NAND2_X1 U7114 ( .A1(n7512), .A2(n7511), .ZN(n7497) );
  OR2_X1 U7115 ( .A1(n7495), .A2(n7409), .ZN(n7292) );
  OR2_X1 U7116 ( .A1(n10138), .A2(n7376), .ZN(n7456) );
  NAND2_X1 U7117 ( .A1(n7292), .A2(n7456), .ZN(n5844) );
  NOR4_X1 U7118 ( .A1(n7694), .A2(n5658), .A3(n7497), .A4(n5844), .ZN(n5659)
         );
  NAND4_X1 U7119 ( .A1(n4926), .A2(n7704), .A3(n7767), .A4(n5659), .ZN(n5678)
         );
  XNOR2_X1 U7120 ( .A(n5661), .B(n5660), .ZN(n7792) );
  NAND2_X1 U7121 ( .A1(n7792), .A2(n5303), .ZN(n5668) );
  NAND2_X1 U7122 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5663) );
  MUX2_X1 U7123 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5663), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5665) );
  NAND2_X1 U7124 ( .A1(n5665), .A2(n5664), .ZN(n9503) );
  OAI22_X1 U7125 ( .A1(n5506), .A2(n6697), .B1(n6260), .B2(n9503), .ZN(n5666)
         );
  INV_X1 U7126 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7127 ( .A1(n5647), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5677) );
  OR2_X1 U7128 ( .A1(n5669), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5671) );
  AND2_X1 U7129 ( .A1(n5671), .A2(n5670), .ZN(n9764) );
  NAND2_X1 U7130 ( .A1(n4492), .A2(n9764), .ZN(n5676) );
  INV_X1 U7131 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5672) );
  OR2_X1 U7132 ( .A1(n5693), .A2(n5672), .ZN(n5675) );
  INV_X1 U7133 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5673) );
  OR2_X1 U7134 ( .A1(n4493), .A2(n5673), .ZN(n5674) );
  NAND4_X1 U7135 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(n9736)
         );
  INV_X1 U7136 ( .A(n9736), .ZN(n9408) );
  XNOR2_X1 U7137 ( .A(n9760), .B(n9408), .ZN(n9755) );
  NOR4_X1 U7138 ( .A1(n9709), .A2(n5747), .A3(n5678), .A4(n9755), .ZN(n5679)
         );
  NAND3_X1 U7139 ( .A1(n9677), .A2(n9692), .A3(n5679), .ZN(n5680) );
  NOR4_X1 U7140 ( .A1(n5681), .A2(n9638), .A3(n9663), .A4(n5680), .ZN(n5698)
         );
  XNOR2_X1 U7141 ( .A(n5683), .B(n5682), .ZN(n8040) );
  NAND2_X1 U7142 ( .A1(n8040), .A2(n5303), .ZN(n5686) );
  NAND2_X1 U7143 ( .A1(n5684), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7144 ( .A1(n5647), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5697) );
  INV_X1 U7145 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5690) );
  INV_X1 U7146 ( .A(n5687), .ZN(n5688) );
  AOI21_X1 U7147 ( .B1(n5690), .B2(n5689), .A(n5688), .ZN(n9621) );
  NAND2_X1 U7148 ( .A1(n4492), .A2(n9621), .ZN(n5696) );
  INV_X1 U7149 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5691) );
  OR2_X1 U7150 ( .A1(n4493), .A2(n5691), .ZN(n5695) );
  INV_X1 U7151 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5692) );
  OR2_X1 U7152 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  NAND4_X1 U7153 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n9640)
         );
  XNOR2_X1 U7154 ( .A(n9803), .B(n9640), .ZN(n9625) );
  NAND4_X1 U7155 ( .A1(n9575), .A2(n9612), .A3(n5698), .A4(n9625), .ZN(n5699)
         );
  NOR4_X1 U7156 ( .A1(n5701), .A2(n9598), .A3(n5700), .A4(n5699), .ZN(n5703)
         );
  NAND2_X1 U7157 ( .A1(n9554), .A2(n5702), .ZN(n5901) );
  NAND4_X1 U7158 ( .A1(n5874), .A2(n5703), .A3(n5901), .A4(n5903), .ZN(n5704)
         );
  XNOR2_X1 U7159 ( .A(n5704), .B(n6991), .ZN(n5871) );
  INV_X1 U7160 ( .A(n9777), .ZN(n7896) );
  INV_X1 U7161 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5872) );
  INV_X1 U7162 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7163 ( .A1(n5870), .A2(n5708), .ZN(n5709) );
  NAND2_X1 U7164 ( .A1(n8377), .A2(n10054), .ZN(n6207) );
  MUX2_X1 U7165 ( .A(n7896), .B(n6220), .S(n6207), .Z(n5790) );
  NAND2_X1 U7166 ( .A1(n10055), .A2(n5711), .ZN(n5712) );
  NOR2_X1 U7167 ( .A1(n9495), .A2(n6887), .ZN(n5822) );
  NAND2_X1 U7168 ( .A1(n9495), .A2(n6887), .ZN(n5881) );
  INV_X1 U7169 ( .A(n5823), .ZN(n5714) );
  NOR2_X1 U7170 ( .A1(n6974), .A2(n5714), .ZN(n5876) );
  INV_X1 U7171 ( .A(n5827), .ZN(n5824) );
  OR2_X1 U7172 ( .A1(n5876), .A2(n5824), .ZN(n6903) );
  AND2_X1 U7173 ( .A1(n5884), .A2(n5826), .ZN(n5841) );
  INV_X1 U7174 ( .A(n5841), .ZN(n5716) );
  INV_X1 U7175 ( .A(n5884), .ZN(n5829) );
  AND2_X1 U7176 ( .A1(n7078), .A2(n5875), .ZN(n5715) );
  OAI22_X1 U7177 ( .A1(n6903), .A2(n5716), .B1(n5829), .B2(n5715), .ZN(n5719)
         );
  NAND2_X1 U7178 ( .A1(n6903), .A2(n7029), .ZN(n6902) );
  INV_X1 U7179 ( .A(n7078), .ZN(n5717) );
  AOI21_X1 U7180 ( .B1(n6902), .B2(n5841), .A(n5717), .ZN(n5718) );
  INV_X1 U7181 ( .A(n6207), .ZN(n5792) );
  NAND2_X1 U7182 ( .A1(n7455), .A2(n7288), .ZN(n5720) );
  INV_X1 U7183 ( .A(n7497), .ZN(n7502) );
  NAND2_X1 U7184 ( .A1(n5721), .A2(n7502), .ZN(n5735) );
  NAND2_X1 U7185 ( .A1(n7456), .A2(n7463), .ZN(n7289) );
  AOI21_X1 U7186 ( .B1(n5722), .B2(n7288), .A(n7289), .ZN(n5723) );
  OAI21_X1 U7187 ( .B1(n5723), .B2(n5833), .A(n7292), .ZN(n5724) );
  OAI211_X1 U7188 ( .C1(n5735), .C2(n5724), .A(n7701), .B(n7511), .ZN(n5725)
         );
  AND2_X1 U7189 ( .A1(n7900), .A2(n5726), .ZN(n5842) );
  NAND2_X1 U7190 ( .A1(n9760), .A2(n9408), .ZN(n7902) );
  AND2_X1 U7191 ( .A1(n7902), .A2(n5792), .ZN(n5730) );
  INV_X1 U7192 ( .A(n5730), .ZN(n5728) );
  INV_X1 U7193 ( .A(n5848), .ZN(n5727) );
  NOR2_X1 U7194 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  AND2_X1 U7195 ( .A1(n7904), .A2(n5729), .ZN(n5733) );
  NAND3_X1 U7196 ( .A1(n7904), .A2(n9755), .A3(n5730), .ZN(n5731) );
  OAI21_X1 U7197 ( .B1(n5853), .B2(n6207), .A(n5731), .ZN(n5732) );
  AND2_X1 U7198 ( .A1(n5734), .A2(n7512), .ZN(n7698) );
  NAND2_X1 U7199 ( .A1(n5735), .A2(n7698), .ZN(n5736) );
  NAND2_X1 U7200 ( .A1(n5736), .A2(n7701), .ZN(n5739) );
  NAND2_X1 U7201 ( .A1(n5755), .A2(n9705), .ZN(n7907) );
  INV_X1 U7202 ( .A(n7907), .ZN(n5813) );
  NOR2_X1 U7203 ( .A1(n9760), .A2(n9408), .ZN(n7903) );
  OR2_X1 U7204 ( .A1(n7903), .A2(n5792), .ZN(n5740) );
  NAND2_X1 U7205 ( .A1(n7900), .A2(n7767), .ZN(n5737) );
  NOR2_X1 U7206 ( .A1(n5740), .A2(n5737), .ZN(n5738) );
  NAND4_X1 U7207 ( .A1(n5739), .A2(n5813), .A3(n5738), .A4(n5853), .ZN(n5750)
         );
  INV_X1 U7208 ( .A(n5740), .ZN(n5744) );
  INV_X1 U7209 ( .A(n9755), .ZN(n5742) );
  NAND2_X1 U7210 ( .A1(n5848), .A2(n7703), .ZN(n5832) );
  NAND2_X1 U7211 ( .A1(n5832), .A2(n7900), .ZN(n5741) );
  NAND2_X1 U7212 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NAND3_X1 U7213 ( .A1(n5744), .A2(n5853), .A3(n5743), .ZN(n5745) );
  OAI211_X1 U7214 ( .C1(n5792), .C2(n7904), .A(n9723), .B(n5745), .ZN(n5746)
         );
  NAND2_X1 U7215 ( .A1(n5746), .A2(n5813), .ZN(n5749) );
  NAND2_X1 U7216 ( .A1(n5747), .A2(n5792), .ZN(n5748) );
  NAND4_X1 U7217 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n5754)
         );
  OR2_X1 U7218 ( .A1(n5857), .A2(n4812), .ZN(n5812) );
  INV_X1 U7219 ( .A(n5752), .ZN(n5756) );
  AND2_X1 U7220 ( .A1(n7909), .A2(n5756), .ZN(n5811) );
  OAI21_X1 U7221 ( .B1(n5754), .B2(n5812), .A(n5811), .ZN(n5758) );
  AND2_X1 U7222 ( .A1(n7906), .A2(n5753), .ZN(n5831) );
  INV_X1 U7223 ( .A(n5857), .ZN(n7908) );
  INV_X1 U7224 ( .A(n5760), .ZN(n7911) );
  OR2_X1 U7225 ( .A1(n5759), .A2(n7911), .ZN(n5816) );
  OR2_X1 U7226 ( .A1(n5769), .A2(n5816), .ZN(n5764) );
  INV_X1 U7227 ( .A(n9640), .ZN(n9398) );
  NAND2_X1 U7228 ( .A1(n9803), .A2(n9398), .ZN(n9608) );
  INV_X1 U7229 ( .A(n5759), .ZN(n5763) );
  NAND2_X1 U7230 ( .A1(n5760), .A2(n7910), .ZN(n5761) );
  NAND2_X1 U7231 ( .A1(n5761), .A2(n7912), .ZN(n5762) );
  OR2_X1 U7232 ( .A1(n7913), .A2(n5762), .ZN(n5858) );
  NAND2_X1 U7233 ( .A1(n5763), .A2(n5858), .ZN(n5814) );
  NOR2_X1 U7234 ( .A1(n9803), .A2(n9398), .ZN(n7915) );
  INV_X1 U7235 ( .A(n7915), .ZN(n5768) );
  OR2_X1 U7236 ( .A1(n7915), .A2(n9652), .ZN(n5766) );
  NAND2_X1 U7237 ( .A1(n9608), .A2(n9636), .ZN(n5765) );
  NAND2_X1 U7238 ( .A1(n5766), .A2(n5765), .ZN(n5774) );
  NAND2_X1 U7239 ( .A1(n5774), .A2(n9652), .ZN(n5767) );
  NAND2_X1 U7240 ( .A1(n5769), .A2(n7909), .ZN(n5770) );
  AOI21_X1 U7241 ( .B1(n5770), .B2(n7912), .A(n5816), .ZN(n5772) );
  INV_X1 U7242 ( .A(n7914), .ZN(n5771) );
  NOR2_X1 U7243 ( .A1(n7915), .A2(n5771), .ZN(n5810) );
  OAI21_X1 U7244 ( .B1(n5772), .B2(n7913), .A(n5810), .ZN(n5776) );
  NAND2_X1 U7245 ( .A1(n5773), .A2(n9608), .ZN(n7916) );
  AOI21_X1 U7246 ( .B1(n9807), .B2(n5774), .A(n7916), .ZN(n5775) );
  NAND2_X1 U7247 ( .A1(n5776), .A2(n5775), .ZN(n5777) );
  OR2_X1 U7248 ( .A1(n9792), .A2(n9396), .ZN(n5778) );
  NAND2_X1 U7249 ( .A1(n5778), .A2(n9594), .ZN(n7918) );
  NAND2_X1 U7250 ( .A1(n5778), .A2(n6207), .ZN(n5782) );
  NAND2_X1 U7251 ( .A1(n9792), .A2(n9396), .ZN(n7917) );
  INV_X1 U7252 ( .A(n7917), .ZN(n5802) );
  AOI21_X1 U7253 ( .B1(n7918), .B2(n5782), .A(n5802), .ZN(n5779) );
  NAND2_X1 U7254 ( .A1(n5780), .A2(n5779), .ZN(n5784) );
  NAND2_X1 U7255 ( .A1(n7917), .A2(n5792), .ZN(n5781) );
  NAND2_X1 U7256 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  NAND3_X1 U7257 ( .A1(n5784), .A2(n9575), .A3(n5783), .ZN(n5786) );
  MUX2_X1 U7258 ( .A(n5804), .B(n5809), .S(n5792), .Z(n5785) );
  NAND3_X1 U7259 ( .A1(n5786), .A2(n9567), .A3(n5785), .ZN(n5788) );
  MUX2_X1 U7260 ( .A(n7920), .B(n5805), .S(n6207), .Z(n5787) );
  NAND2_X1 U7261 ( .A1(n5788), .A2(n5787), .ZN(n5797) );
  NAND3_X1 U7262 ( .A1(n5797), .A2(n7896), .A3(n6220), .ZN(n5789) );
  INV_X1 U7263 ( .A(n9554), .ZN(n9904) );
  AOI21_X1 U7264 ( .B1(n9482), .B2(n9483), .A(n9904), .ZN(n5863) );
  INV_X1 U7265 ( .A(n5791), .ZN(n5793) );
  NOR2_X1 U7266 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  AOI21_X1 U7267 ( .B1(n5799), .B2(n5923), .A(n5796), .ZN(n5869) );
  NOR3_X1 U7268 ( .A1(n5863), .A2(n6220), .A3(n5797), .ZN(n5798) );
  NOR3_X1 U7269 ( .A1(n5865), .A2(n5923), .A3(n5798), .ZN(n5801) );
  INV_X1 U7270 ( .A(n5799), .ZN(n5800) );
  OAI21_X1 U7271 ( .B1(n5801), .B2(n6991), .A(n5800), .ZN(n5868) );
  NAND2_X1 U7272 ( .A1(n5809), .A2(n5802), .ZN(n5803) );
  NAND3_X1 U7273 ( .A1(n7920), .A2(n5804), .A3(n5803), .ZN(n5861) );
  NOR2_X1 U7274 ( .A1(n5861), .A2(n4810), .ZN(n5808) );
  INV_X1 U7275 ( .A(n5805), .ZN(n5806) );
  NOR3_X1 U7276 ( .A1(n5808), .A2(n5807), .A3(n5806), .ZN(n5900) );
  INV_X1 U7277 ( .A(n5810), .ZN(n5819) );
  OAI21_X1 U7278 ( .B1(n5813), .B2(n5812), .A(n5811), .ZN(n5815) );
  OAI211_X1 U7279 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5892), .ZN(n5817)
         );
  INV_X1 U7280 ( .A(n5817), .ZN(n5818) );
  NOR2_X1 U7281 ( .A1(n5819), .A2(n5818), .ZN(n5895) );
  INV_X1 U7282 ( .A(n5820), .ZN(n5821) );
  AOI21_X1 U7283 ( .B1(n5822), .B2(n5879), .A(n5821), .ZN(n5825) );
  OAI211_X1 U7284 ( .C1(n5825), .C2(n5824), .A(n5875), .B(n5823), .ZN(n5840)
         );
  NAND2_X1 U7285 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  NAND4_X1 U7286 ( .A1(n6884), .A2(n5879), .A3(n7031), .A4(n5881), .ZN(n5830)
         );
  NOR2_X1 U7287 ( .A1(n5830), .A2(n5829), .ZN(n5839) );
  INV_X1 U7288 ( .A(n5831), .ZN(n5856) );
  INV_X1 U7289 ( .A(n5832), .ZN(n5837) );
  NAND2_X1 U7290 ( .A1(n5833), .A2(n7292), .ZN(n7501) );
  AND2_X1 U7291 ( .A1(n7501), .A2(n7511), .ZN(n5834) );
  NAND2_X1 U7292 ( .A1(n7701), .A2(n5834), .ZN(n5845) );
  NAND2_X1 U7293 ( .A1(n7288), .A2(n7078), .ZN(n5835) );
  NOR2_X1 U7294 ( .A1(n5845), .A2(n5835), .ZN(n5836) );
  NAND3_X1 U7295 ( .A1(n7902), .A2(n5837), .A3(n5836), .ZN(n5838) );
  OR3_X1 U7296 ( .A1(n5856), .A2(n4817), .A3(n5838), .ZN(n5890) );
  AOI211_X1 U7297 ( .C1(n5841), .C2(n5840), .A(n5839), .B(n5890), .ZN(n5859)
         );
  INV_X1 U7298 ( .A(n7903), .ZN(n5852) );
  INV_X1 U7299 ( .A(n5842), .ZN(n5850) );
  INV_X1 U7300 ( .A(n7701), .ZN(n5846) );
  INV_X1 U7301 ( .A(n7463), .ZN(n5843) );
  NOR2_X1 U7302 ( .A1(n5844), .A2(n5843), .ZN(n7499) );
  OAI22_X1 U7303 ( .A1(n7698), .A2(n5846), .B1(n5845), .B2(n7499), .ZN(n5847)
         );
  AND2_X1 U7304 ( .A1(n5847), .A2(n7703), .ZN(n5849) );
  OAI211_X1 U7305 ( .C1(n5850), .C2(n5849), .A(n5848), .B(n7902), .ZN(n5851)
         );
  NAND3_X1 U7306 ( .A1(n5853), .A2(n5852), .A3(n5851), .ZN(n5854) );
  NAND2_X1 U7307 ( .A1(n5854), .A2(n7904), .ZN(n5855) );
  NOR2_X1 U7308 ( .A1(n5856), .A2(n5855), .ZN(n5887) );
  NOR2_X1 U7309 ( .A1(n5858), .A2(n5857), .ZN(n5893) );
  OAI211_X1 U7310 ( .C1(n5859), .C2(n5887), .A(n5893), .B(n5892), .ZN(n5860)
         );
  AOI21_X1 U7311 ( .B1(n5895), .B2(n5860), .A(n7916), .ZN(n5862) );
  INV_X1 U7312 ( .A(n5861), .ZN(n5896) );
  OAI21_X1 U7313 ( .B1(n7919), .B2(n5862), .A(n5896), .ZN(n5864) );
  AOI211_X1 U7314 ( .C1(n5900), .C2(n5864), .A(n5898), .B(n5863), .ZN(n5866)
         );
  OAI21_X1 U7315 ( .B1(n5866), .B2(n5865), .A(n5903), .ZN(n5867) );
  XNOR2_X1 U7316 ( .A(n5873), .B(n5872), .ZN(n7102) );
  INV_X1 U7317 ( .A(n7102), .ZN(n6977) );
  INV_X1 U7318 ( .A(n5874), .ZN(n5905) );
  NAND2_X1 U7319 ( .A1(n5876), .A2(n5875), .ZN(n7032) );
  NAND3_X1 U7320 ( .A1(n5879), .A2(n5878), .A3(n5877), .ZN(n5883) );
  NAND3_X1 U7321 ( .A1(n5881), .A2(n5880), .A3(n5929), .ZN(n5882) );
  NOR2_X1 U7322 ( .A1(n5883), .A2(n5882), .ZN(n5885) );
  OAI211_X1 U7323 ( .C1(n7032), .C2(n5885), .A(n5884), .B(n7031), .ZN(n5886)
         );
  INV_X1 U7324 ( .A(n5886), .ZN(n5889) );
  INV_X1 U7325 ( .A(n5887), .ZN(n5888) );
  OAI21_X1 U7326 ( .B1(n5890), .B2(n5889), .A(n5888), .ZN(n5891) );
  NAND3_X1 U7327 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n5894) );
  AOI21_X1 U7328 ( .B1(n5895), .B2(n5894), .A(n7916), .ZN(n5897) );
  OAI21_X1 U7329 ( .B1(n5897), .B2(n9573), .A(n5896), .ZN(n5899) );
  AOI21_X1 U7330 ( .B1(n5900), .B2(n5899), .A(n5898), .ZN(n5902) );
  AND2_X1 U7331 ( .A1(n5902), .A2(n5901), .ZN(n5904) );
  OAI21_X1 U7332 ( .B1(n5905), .B2(n5904), .A(n5903), .ZN(n5908) );
  AND2_X1 U7333 ( .A1(n7102), .A2(n10054), .ZN(n10069) );
  NAND2_X1 U7334 ( .A1(n5906), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5907) );
  XNOR2_X1 U7335 ( .A(n5907), .B(n5011), .ZN(n6258) );
  OR2_X1 U7336 ( .A1(n6258), .A2(P1_U3084), .ZN(n7383) );
  AOI21_X1 U7337 ( .B1(n5908), .B2(n10069), .A(n7383), .ZN(n5912) );
  INV_X1 U7338 ( .A(n5908), .ZN(n5910) );
  NAND2_X1 U7339 ( .A1(n7102), .A2(n6991), .ZN(n6195) );
  NAND2_X1 U7340 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  INV_X1 U7341 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7342 ( .A1(n5918), .A2(n5917), .ZN(n5920) );
  NAND2_X1 U7343 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5914) );
  INV_X1 U7344 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7345 ( .A1(n4540), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5916) );
  XNOR2_X1 U7346 ( .A(n5916), .B(n5915), .ZN(n7508) );
  OR2_X1 U7347 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  NAND2_X1 U7348 ( .A1(n5920), .A2(n5919), .ZN(n7727) );
  AND2_X1 U7349 ( .A1(n6258), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7350 ( .A1(n5930), .A2(n5921), .ZN(n10090) );
  NOR2_X1 U7351 ( .A1(n10090), .A2(n6195), .ZN(n6210) );
  INV_X1 U7352 ( .A(n5922), .ZN(n9929) );
  NAND2_X1 U7353 ( .A1(n9929), .A2(n4764), .ZN(n10056) );
  INV_X1 U7354 ( .A(n5925), .ZN(n5926) );
  NAND3_X1 U7355 ( .A1(n6210), .A2(n9735), .A3(n5926), .ZN(n5927) );
  OAI211_X1 U7356 ( .C1(n5923), .C2(n7383), .A(n5927), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5928) );
  NAND2_X1 U7357 ( .A1(n6391), .A2(n6095), .ZN(n5932) );
  NAND2_X1 U7358 ( .A1(n10052), .A2(n6125), .ZN(n5931) );
  NAND2_X1 U7359 ( .A1(n5932), .A2(n5931), .ZN(n5935) );
  INV_X1 U7360 ( .A(n5929), .ZN(n7126) );
  NOR2_X1 U7361 ( .A1(n6978), .A2(n6195), .ZN(n6831) );
  NOR2_X4 U7362 ( .A1(n5964), .A2(n6831), .ZN(n6059) );
  NAND2_X1 U7363 ( .A1(n6391), .A2(n6059), .ZN(n5937) );
  NAND2_X1 U7364 ( .A1(n10052), .A2(n6095), .ZN(n5936) );
  NAND2_X1 U7365 ( .A1(n5937), .A2(n5936), .ZN(n5948) );
  NAND2_X1 U7366 ( .A1(n5947), .A2(n5948), .ZN(n5946) );
  NAND2_X1 U7367 ( .A1(n5941), .A2(n6095), .ZN(n5939) );
  INV_X1 U7368 ( .A(n5930), .ZN(n5942) );
  AOI22_X1 U7369 ( .A1(n6828), .A2(n6125), .B1(n5942), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7370 ( .A1(n5939), .A2(n5938), .ZN(n6389) );
  INV_X1 U7371 ( .A(n6389), .ZN(n5940) );
  NAND2_X1 U7372 ( .A1(n5941), .A2(n4487), .ZN(n5944) );
  AOI22_X1 U7373 ( .A1(n6828), .A2(n6095), .B1(n5942), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5943) );
  AND2_X1 U7374 ( .A1(n5944), .A2(n5943), .ZN(n6390) );
  NAND2_X1 U7375 ( .A1(n6390), .A2(n6389), .ZN(n6388) );
  NAND2_X1 U7376 ( .A1(n5945), .A2(n6388), .ZN(n6589) );
  NAND2_X1 U7377 ( .A1(n5946), .A2(n6589), .ZN(n5950) );
  INV_X1 U7378 ( .A(n5948), .ZN(n6590) );
  NAND2_X1 U7379 ( .A1(n5950), .A2(n5949), .ZN(n6596) );
  NAND4_X1 U7380 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n5958)
         );
  NAND2_X1 U7381 ( .A1(n5958), .A2(n6095), .ZN(n5956) );
  NAND2_X1 U7382 ( .A1(n6878), .A2(n6125), .ZN(n5955) );
  NAND2_X1 U7383 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  AOI22_X1 U7384 ( .A1(n5958), .A2(n6059), .B1(n6095), .B2(n6878), .ZN(n5960)
         );
  INV_X1 U7385 ( .A(n5959), .ZN(n5961) );
  NAND2_X1 U7386 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7387 ( .A1(n5963), .A2(n5962), .ZN(n6492) );
  NAND2_X1 U7388 ( .A1(n9495), .A2(n6095), .ZN(n5966) );
  NAND2_X1 U7389 ( .A1(n6889), .A2(n6125), .ZN(n5965) );
  NAND2_X1 U7390 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7391 ( .A(n5967), .B(n6172), .ZN(n5968) );
  AOI22_X1 U7392 ( .A1(n9495), .A2(n6059), .B1(n6095), .B2(n6889), .ZN(n5969)
         );
  XNOR2_X1 U7393 ( .A(n5968), .B(n5969), .ZN(n6493) );
  NAND2_X1 U7394 ( .A1(n6492), .A2(n6493), .ZN(n5972) );
  INV_X1 U7395 ( .A(n5968), .ZN(n5970) );
  NAND2_X1 U7396 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  NAND2_X1 U7397 ( .A1(n5972), .A2(n5971), .ZN(n6717) );
  NAND2_X1 U7398 ( .A1(n9494), .A2(n6095), .ZN(n5974) );
  NAND2_X1 U7399 ( .A1(n6834), .A2(n6125), .ZN(n5973) );
  NAND2_X1 U7400 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  AOI22_X1 U7401 ( .A1(n9494), .A2(n6059), .B1(n6095), .B2(n6834), .ZN(n5978)
         );
  XNOR2_X1 U7402 ( .A(n5977), .B(n5978), .ZN(n6718) );
  INV_X1 U7403 ( .A(n6718), .ZN(n5976) );
  NAND2_X1 U7404 ( .A1(n9493), .A2(n6095), .ZN(n5983) );
  NAND2_X1 U7405 ( .A1(n6985), .A2(n6125), .ZN(n5982) );
  NAND2_X1 U7406 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  XNOR2_X1 U7407 ( .A(n5984), .B(n6172), .ZN(n6703) );
  NAND2_X1 U7408 ( .A1(n9493), .A2(n6059), .ZN(n5986) );
  NAND2_X1 U7409 ( .A1(n6985), .A2(n6095), .ZN(n5985) );
  NAND2_X1 U7410 ( .A1(n5986), .A2(n5985), .ZN(n6702) );
  AND2_X1 U7411 ( .A1(n6703), .A2(n6702), .ZN(n5989) );
  INV_X1 U7412 ( .A(n6703), .ZN(n5988) );
  INV_X1 U7413 ( .A(n6702), .ZN(n5987) );
  NAND2_X1 U7414 ( .A1(n9492), .A2(n6095), .ZN(n5991) );
  NAND2_X1 U7415 ( .A1(n6907), .A2(n6125), .ZN(n5990) );
  NAND2_X1 U7416 ( .A1(n5991), .A2(n5990), .ZN(n5993) );
  XNOR2_X1 U7417 ( .A(n5993), .B(n6165), .ZN(n6784) );
  NAND2_X1 U7418 ( .A1(n9492), .A2(n6059), .ZN(n5995) );
  NAND2_X1 U7419 ( .A1(n6907), .A2(n6095), .ZN(n5994) );
  NAND2_X1 U7420 ( .A1(n5995), .A2(n5994), .ZN(n6783) );
  NAND2_X1 U7421 ( .A1(n9491), .A2(n6095), .ZN(n5997) );
  NAND2_X1 U7422 ( .A1(n7045), .A2(n6125), .ZN(n5996) );
  NAND2_X1 U7423 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7424 ( .A(n5998), .B(n6165), .ZN(n6001) );
  NAND2_X1 U7425 ( .A1(n9491), .A2(n6059), .ZN(n6000) );
  NAND2_X1 U7426 ( .A1(n7045), .A2(n6095), .ZN(n5999) );
  AND2_X1 U7427 ( .A1(n6000), .A2(n5999), .ZN(n6002) );
  NAND2_X1 U7428 ( .A1(n6001), .A2(n6002), .ZN(n6006) );
  INV_X1 U7429 ( .A(n6001), .ZN(n6004) );
  INV_X1 U7430 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7431 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  AND2_X1 U7432 ( .A1(n6006), .A2(n6005), .ZN(n6947) );
  AOI22_X1 U7433 ( .A1(n7295), .A2(n6095), .B1(n6059), .B2(n9490), .ZN(n6011)
         );
  NAND2_X1 U7434 ( .A1(n7295), .A2(n6125), .ZN(n6008) );
  NAND2_X1 U7435 ( .A1(n9490), .A2(n6095), .ZN(n6007) );
  NAND2_X1 U7436 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  XNOR2_X1 U7437 ( .A(n6009), .B(n6172), .ZN(n7117) );
  INV_X1 U7438 ( .A(n6010), .ZN(n6013) );
  INV_X1 U7439 ( .A(n6011), .ZN(n6012) );
  NAND2_X1 U7440 ( .A1(n10138), .A2(n6125), .ZN(n6015) );
  NAND2_X1 U7441 ( .A1(n9489), .A2(n6095), .ZN(n6014) );
  NAND2_X1 U7442 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  XNOR2_X1 U7443 ( .A(n6016), .B(n6165), .ZN(n6018) );
  AND2_X1 U7444 ( .A1(n9489), .A2(n6059), .ZN(n6017) );
  AOI21_X1 U7445 ( .B1(n10138), .B2(n6095), .A(n6017), .ZN(n6019) );
  NAND2_X1 U7446 ( .A1(n6018), .A2(n6019), .ZN(n6024) );
  INV_X1 U7447 ( .A(n6018), .ZN(n6021) );
  INV_X1 U7448 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7449 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7450 ( .A1(n6024), .A2(n6022), .ZN(n7130) );
  INV_X1 U7451 ( .A(n7130), .ZN(n6023) );
  NAND2_X1 U7452 ( .A1(n7495), .A2(n6125), .ZN(n6026) );
  NAND2_X1 U7453 ( .A1(n9488), .A2(n6095), .ZN(n6025) );
  NAND2_X1 U7454 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  XNOR2_X1 U7455 ( .A(n6027), .B(n6172), .ZN(n6030) );
  NAND2_X1 U7456 ( .A1(n7495), .A2(n6095), .ZN(n6029) );
  NAND2_X1 U7457 ( .A1(n9488), .A2(n6059), .ZN(n6028) );
  NAND2_X1 U7458 ( .A1(n6029), .A2(n6028), .ZN(n6031) );
  NAND2_X1 U7459 ( .A1(n6030), .A2(n6031), .ZN(n7369) );
  INV_X1 U7460 ( .A(n6030), .ZN(n6033) );
  INV_X1 U7461 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7462 ( .A1(n6033), .A2(n6032), .ZN(n7368) );
  NAND2_X1 U7463 ( .A1(n7535), .A2(n6125), .ZN(n6035) );
  NAND2_X1 U7464 ( .A1(n9487), .A2(n6095), .ZN(n6034) );
  NAND2_X1 U7465 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  XNOR2_X1 U7466 ( .A(n6036), .B(n6172), .ZN(n6038) );
  AND2_X1 U7467 ( .A1(n9487), .A2(n6059), .ZN(n6037) );
  AOI21_X1 U7468 ( .B1(n7535), .B2(n6095), .A(n6037), .ZN(n6039) );
  XNOR2_X1 U7469 ( .A(n6038), .B(n6039), .ZN(n7407) );
  INV_X1 U7470 ( .A(n6038), .ZN(n6040) );
  NAND2_X1 U7471 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7472 ( .A1(n7692), .A2(n6125), .ZN(n6043) );
  NAND2_X1 U7473 ( .A1(n9486), .A2(n6095), .ZN(n6042) );
  NAND2_X1 U7474 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  XNOR2_X1 U7475 ( .A(n6044), .B(n6165), .ZN(n7487) );
  AND2_X1 U7476 ( .A1(n9486), .A2(n6059), .ZN(n6045) );
  AOI21_X1 U7477 ( .B1(n7692), .B2(n6095), .A(n6045), .ZN(n7486) );
  AND2_X1 U7478 ( .A1(n7487), .A2(n7486), .ZN(n6046) );
  NAND2_X1 U7479 ( .A1(n9848), .A2(n6125), .ZN(n6048) );
  NAND2_X1 U7480 ( .A1(n9485), .A2(n6095), .ZN(n6047) );
  NAND2_X1 U7481 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  XNOR2_X1 U7482 ( .A(n6049), .B(n6172), .ZN(n6052) );
  NAND2_X1 U7483 ( .A1(n9848), .A2(n6095), .ZN(n6051) );
  NAND2_X1 U7484 ( .A1(n9485), .A2(n6059), .ZN(n6050) );
  NAND2_X1 U7485 ( .A1(n6051), .A2(n6050), .ZN(n6053) );
  INV_X1 U7486 ( .A(n6052), .ZN(n6055) );
  INV_X1 U7487 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7488 ( .A1(n6055), .A2(n6054), .ZN(n7655) );
  NAND2_X1 U7489 ( .A1(n9357), .A2(n6125), .ZN(n6057) );
  NAND2_X1 U7490 ( .A1(n9484), .A2(n6095), .ZN(n6056) );
  NAND2_X1 U7491 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  XNOR2_X1 U7492 ( .A(n6058), .B(n6165), .ZN(n6062) );
  NAND2_X1 U7493 ( .A1(n6063), .A2(n6062), .ZN(n9351) );
  NAND2_X1 U7494 ( .A1(n9357), .A2(n6095), .ZN(n6061) );
  NAND2_X1 U7495 ( .A1(n9484), .A2(n6059), .ZN(n6060) );
  NAND2_X1 U7496 ( .A1(n6061), .A2(n6060), .ZN(n9350) );
  NAND2_X1 U7497 ( .A1(n9351), .A2(n9350), .ZN(n9349) );
  NAND2_X1 U7498 ( .A1(n9349), .A2(n9353), .ZN(n7853) );
  NAND2_X1 U7499 ( .A1(n9760), .A2(n6125), .ZN(n6065) );
  NAND2_X1 U7500 ( .A1(n9736), .A2(n6095), .ZN(n6064) );
  NAND2_X1 U7501 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  XNOR2_X1 U7502 ( .A(n6066), .B(n6165), .ZN(n7855) );
  AND2_X1 U7503 ( .A1(n9736), .A2(n6059), .ZN(n6067) );
  AOI21_X1 U7504 ( .B1(n9760), .B2(n6095), .A(n6067), .ZN(n7854) );
  NAND2_X1 U7505 ( .A1(n7855), .A2(n7854), .ZN(n6068) );
  INV_X1 U7506 ( .A(n7855), .ZN(n6070) );
  INV_X1 U7507 ( .A(n7854), .ZN(n6069) );
  NAND2_X1 U7508 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U7509 ( .A1(n9741), .A2(n6125), .ZN(n6073) );
  NAND2_X1 U7510 ( .A1(n9727), .A2(n6095), .ZN(n6072) );
  NAND2_X1 U7511 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  XNOR2_X1 U7512 ( .A(n6074), .B(n6165), .ZN(n6076) );
  AND2_X1 U7513 ( .A1(n9727), .A2(n6059), .ZN(n6075) );
  AOI21_X1 U7514 ( .B1(n9741), .B2(n6095), .A(n6075), .ZN(n6077) );
  NAND2_X1 U7515 ( .A1(n6076), .A2(n6077), .ZN(n6082) );
  INV_X1 U7516 ( .A(n6076), .ZN(n6079) );
  INV_X1 U7517 ( .A(n6077), .ZN(n6078) );
  NAND2_X1 U7518 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7519 ( .A1(n6082), .A2(n6080), .ZN(n9406) );
  NAND2_X1 U7520 ( .A1(n9404), .A2(n6082), .ZN(n9415) );
  NAND2_X1 U7521 ( .A1(n9837), .A2(n6125), .ZN(n6084) );
  NAND2_X1 U7522 ( .A1(n9738), .A2(n6095), .ZN(n6083) );
  NAND2_X1 U7523 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  XNOR2_X1 U7524 ( .A(n6085), .B(n6172), .ZN(n6088) );
  NAND2_X1 U7525 ( .A1(n9837), .A2(n6095), .ZN(n6087) );
  NAND2_X1 U7526 ( .A1(n9738), .A2(n6059), .ZN(n6086) );
  NAND2_X1 U7527 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  NAND2_X1 U7528 ( .A1(n6088), .A2(n6089), .ZN(n9416) );
  NAND2_X1 U7529 ( .A1(n9415), .A2(n9416), .ZN(n9414) );
  INV_X1 U7530 ( .A(n6088), .ZN(n6091) );
  INV_X1 U7531 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7532 ( .A1(n6091), .A2(n6090), .ZN(n9418) );
  NAND2_X1 U7533 ( .A1(n9414), .A2(n9418), .ZN(n6098) );
  NAND2_X1 U7534 ( .A1(n9832), .A2(n6125), .ZN(n6093) );
  NAND2_X1 U7535 ( .A1(n9726), .A2(n6095), .ZN(n6092) );
  NAND2_X1 U7536 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  XNOR2_X1 U7537 ( .A(n6094), .B(n6165), .ZN(n6099) );
  NAND2_X1 U7538 ( .A1(n9832), .A2(n6095), .ZN(n6097) );
  NAND2_X1 U7539 ( .A1(n9726), .A2(n6059), .ZN(n6096) );
  NAND2_X1 U7540 ( .A1(n6097), .A2(n6096), .ZN(n9462) );
  INV_X1 U7541 ( .A(n6098), .ZN(n6101) );
  INV_X1 U7542 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7543 ( .A1(n9828), .A2(n6125), .ZN(n6103) );
  NAND2_X1 U7544 ( .A1(n9710), .A2(n6095), .ZN(n6102) );
  NAND2_X1 U7545 ( .A1(n6103), .A2(n6102), .ZN(n6104) );
  XNOR2_X1 U7546 ( .A(n6104), .B(n6165), .ZN(n6108) );
  AND2_X1 U7547 ( .A1(n9710), .A2(n4487), .ZN(n6105) );
  AOI21_X1 U7548 ( .B1(n9828), .B2(n6095), .A(n6105), .ZN(n6107) );
  XNOR2_X1 U7549 ( .A(n6108), .B(n6107), .ZN(n9376) );
  INV_X1 U7550 ( .A(n9376), .ZN(n6106) );
  NAND2_X1 U7551 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  NAND2_X1 U7552 ( .A1(n9373), .A2(n6109), .ZN(n9437) );
  NAND2_X1 U7553 ( .A1(n9823), .A2(n6125), .ZN(n6111) );
  NAND2_X1 U7554 ( .A1(n9693), .A2(n6095), .ZN(n6110) );
  NAND2_X1 U7555 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  XNOR2_X1 U7556 ( .A(n6112), .B(n6165), .ZN(n9435) );
  AND2_X1 U7557 ( .A1(n9693), .A2(n4487), .ZN(n6113) );
  AOI21_X1 U7558 ( .B1(n9823), .B2(n6095), .A(n6113), .ZN(n9434) );
  AND2_X1 U7559 ( .A1(n9435), .A2(n9434), .ZN(n6114) );
  NAND2_X1 U7560 ( .A1(n9818), .A2(n6125), .ZN(n6116) );
  NAND2_X1 U7561 ( .A1(n9680), .A2(n6095), .ZN(n6115) );
  NAND2_X1 U7562 ( .A1(n6116), .A2(n6115), .ZN(n6117) );
  XNOR2_X1 U7563 ( .A(n6117), .B(n6172), .ZN(n6120) );
  NAND2_X1 U7564 ( .A1(n9818), .A2(n6095), .ZN(n6119) );
  NAND2_X1 U7565 ( .A1(n9680), .A2(n4487), .ZN(n6118) );
  NAND2_X1 U7566 ( .A1(n6119), .A2(n6118), .ZN(n6121) );
  INV_X1 U7567 ( .A(n6120), .ZN(n6123) );
  INV_X1 U7568 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7569 ( .A1(n6123), .A2(n6122), .ZN(n9381) );
  AND2_X1 U7570 ( .A1(n9665), .A2(n6059), .ZN(n6124) );
  AOI21_X1 U7571 ( .B1(n9812), .B2(n6095), .A(n6124), .ZN(n6129) );
  NAND2_X1 U7572 ( .A1(n9812), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7573 ( .A1(n9665), .A2(n6095), .ZN(n6126) );
  NAND2_X1 U7574 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  XNOR2_X1 U7575 ( .A(n6128), .B(n6172), .ZN(n9448) );
  NAND2_X1 U7576 ( .A1(n9807), .A2(n6125), .ZN(n6131) );
  NAND2_X1 U7577 ( .A1(n9652), .A2(n6095), .ZN(n6130) );
  NAND2_X1 U7578 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  XNOR2_X1 U7579 ( .A(n6132), .B(n6172), .ZN(n6135) );
  NAND2_X1 U7580 ( .A1(n6134), .A2(n6135), .ZN(n9362) );
  AND2_X1 U7581 ( .A1(n9652), .A2(n6059), .ZN(n6133) );
  AOI21_X1 U7582 ( .B1(n9807), .B2(n6095), .A(n6133), .ZN(n9361) );
  NAND2_X1 U7583 ( .A1(n9362), .A2(n9361), .ZN(n9359) );
  INV_X1 U7584 ( .A(n6134), .ZN(n6137) );
  INV_X1 U7585 ( .A(n6135), .ZN(n6136) );
  NAND2_X1 U7586 ( .A1(n9359), .A2(n9363), .ZN(n9426) );
  NAND2_X1 U7587 ( .A1(n9803), .A2(n6125), .ZN(n6139) );
  NAND2_X1 U7588 ( .A1(n9640), .A2(n6095), .ZN(n6138) );
  NAND2_X1 U7589 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  XNOR2_X1 U7590 ( .A(n6140), .B(n6172), .ZN(n6142) );
  AND2_X1 U7591 ( .A1(n9640), .A2(n6059), .ZN(n6141) );
  AOI21_X1 U7592 ( .B1(n9803), .B2(n6095), .A(n6141), .ZN(n6143) );
  XNOR2_X1 U7593 ( .A(n6142), .B(n6143), .ZN(n9427) );
  INV_X1 U7594 ( .A(n6142), .ZN(n6144) );
  NAND2_X1 U7595 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  NAND2_X1 U7596 ( .A1(n9798), .A2(n6125), .ZN(n6147) );
  NAND2_X1 U7597 ( .A1(n9627), .A2(n6095), .ZN(n6146) );
  NAND2_X1 U7598 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  XNOR2_X1 U7599 ( .A(n6148), .B(n6172), .ZN(n6150) );
  AND2_X1 U7600 ( .A1(n9627), .A2(n6059), .ZN(n6149) );
  AOI21_X1 U7601 ( .B1(n9798), .B2(n6095), .A(n6149), .ZN(n6151) );
  XNOR2_X1 U7602 ( .A(n6150), .B(n6151), .ZN(n9394) );
  INV_X1 U7603 ( .A(n6150), .ZN(n6152) );
  NAND2_X1 U7604 ( .A1(n9792), .A2(n6125), .ZN(n6154) );
  NAND2_X1 U7605 ( .A1(n9614), .A2(n6095), .ZN(n6153) );
  NAND2_X1 U7606 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  XNOR2_X1 U7607 ( .A(n6155), .B(n6165), .ZN(n6158) );
  AND2_X1 U7608 ( .A1(n9614), .A2(n4487), .ZN(n6156) );
  AOI21_X1 U7609 ( .B1(n9792), .B2(n6095), .A(n6156), .ZN(n6159) );
  XNOR2_X1 U7610 ( .A(n6158), .B(n6159), .ZN(n9471) );
  INV_X1 U7611 ( .A(n6158), .ZN(n6161) );
  INV_X1 U7612 ( .A(n6159), .ZN(n6160) );
  NAND2_X1 U7613 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  NAND2_X1 U7614 ( .A1(n9789), .A2(n6125), .ZN(n6164) );
  NAND2_X1 U7615 ( .A1(n9600), .A2(n6095), .ZN(n6163) );
  NAND2_X1 U7616 ( .A1(n6164), .A2(n6163), .ZN(n6166) );
  XNOR2_X1 U7617 ( .A(n6166), .B(n6165), .ZN(n9335) );
  AND2_X1 U7618 ( .A1(n9600), .A2(n6059), .ZN(n6167) );
  AOI21_X1 U7619 ( .B1(n9789), .B2(n6095), .A(n6167), .ZN(n9334) );
  INV_X1 U7620 ( .A(n6203), .ZN(n6199) );
  INV_X1 U7621 ( .A(n9335), .ZN(n6168) );
  NAND2_X1 U7622 ( .A1(n6169), .A2(n6168), .ZN(n6204) );
  NAND2_X1 U7623 ( .A1(n9782), .A2(n6095), .ZN(n6171) );
  NAND2_X1 U7624 ( .A1(n9576), .A2(n4487), .ZN(n6170) );
  NAND2_X1 U7625 ( .A1(n6171), .A2(n6170), .ZN(n6173) );
  XNOR2_X1 U7626 ( .A(n6173), .B(n6172), .ZN(n6176) );
  AOI22_X1 U7627 ( .A1(n9782), .A2(n6125), .B1(n6095), .B2(n9576), .ZN(n6175)
         );
  XNOR2_X1 U7628 ( .A(n6176), .B(n6175), .ZN(n6200) );
  INV_X1 U7629 ( .A(n7781), .ZN(n6179) );
  NAND2_X1 U7630 ( .A1(n7727), .A2(P1_B_REG_SCAN_IN), .ZN(n6177) );
  MUX2_X1 U7631 ( .A(P1_B_REG_SCAN_IN), .B(n6177), .S(n7508), .Z(n6178) );
  NAND2_X1 U7632 ( .A1(n6179), .A2(n6178), .ZN(n10079) );
  OR2_X1 U7633 ( .A1(n10079), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7634 ( .A1(n7781), .A2(n7508), .ZN(n6180) );
  AND2_X1 U7635 ( .A1(n6181), .A2(n6180), .ZN(n9871) );
  OR2_X1 U7636 ( .A1(n10079), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7637 ( .A1(n7781), .A2(n7727), .ZN(n6182) );
  AND2_X1 U7638 ( .A1(n6183), .A2(n6182), .ZN(n6814) );
  NOR4_X1 U7639 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6187) );
  NOR4_X1 U7640 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6186) );
  NOR4_X1 U7641 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6185) );
  NOR4_X1 U7642 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6184) );
  NAND4_X1 U7643 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n6193)
         );
  NOR2_X1 U7644 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n6191) );
  NOR4_X1 U7645 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6190) );
  NOR4_X1 U7646 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6189) );
  NOR4_X1 U7647 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6188) );
  NAND4_X1 U7648 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n6192)
         );
  NOR2_X1 U7649 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  OR2_X1 U7650 ( .A1(n10079), .A2(n6194), .ZN(n6812) );
  NAND3_X1 U7651 ( .A1(n9871), .A2(n6814), .A3(n6812), .ZN(n6215) );
  NOR2_X1 U7652 ( .A1(n6215), .A2(n10090), .ZN(n6206) );
  OR2_X1 U7653 ( .A1(n6978), .A2(n5909), .ZN(n10130) );
  AND2_X1 U7654 ( .A1(n10130), .A2(n6257), .ZN(n6196) );
  AND2_X1 U7655 ( .A1(n6206), .A2(n6196), .ZN(n9428) );
  AND2_X1 U7656 ( .A1(n6200), .A2(n9428), .ZN(n6197) );
  NAND2_X1 U7657 ( .A1(n6199), .A2(n6198), .ZN(n6228) );
  INV_X1 U7658 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7659 ( .A1(n6201), .A2(n9428), .ZN(n6205) );
  INV_X1 U7660 ( .A(n6205), .ZN(n6202) );
  NOR2_X1 U7661 ( .A1(n6205), .A2(n6204), .ZN(n6225) );
  INV_X1 U7662 ( .A(n6206), .ZN(n6209) );
  INV_X1 U7663 ( .A(n10090), .ZN(n10080) );
  OR2_X1 U7664 ( .A1(n10145), .A2(n5929), .ZN(n6480) );
  INV_X1 U7665 ( .A(n6480), .ZN(n6208) );
  NAND2_X1 U7666 ( .A1(n10080), .A2(n6208), .ZN(n7922) );
  NAND2_X1 U7667 ( .A1(n6209), .A2(n7922), .ZN(n6496) );
  INV_X1 U7668 ( .A(n10130), .ZN(n10139) );
  INV_X1 U7669 ( .A(n6215), .ZN(n6211) );
  NAND2_X1 U7670 ( .A1(n6211), .A2(n6210), .ZN(n6214) );
  OR2_X1 U7671 ( .A1(n6214), .A2(n10056), .ZN(n9464) );
  OAI22_X1 U7672 ( .A1(n9464), .A2(n6213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6212), .ZN(n6222) );
  NAND2_X1 U7673 ( .A1(n5922), .A2(n4764), .ZN(n10058) );
  OR2_X1 U7674 ( .A1(n6214), .A2(n10058), .ZN(n9451) );
  NAND2_X1 U7675 ( .A1(n6215), .A2(n6480), .ZN(n6217) );
  OR2_X1 U7676 ( .A1(n6257), .A2(n5909), .ZN(n6811) );
  AND3_X1 U7677 ( .A1(n5930), .A2(n6811), .A3(n6258), .ZN(n6216) );
  NAND2_X1 U7678 ( .A1(n6217), .A2(n6216), .ZN(n6218) );
  NAND2_X1 U7679 ( .A1(n6218), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9453) );
  INV_X1 U7680 ( .A(n9562), .ZN(n6219) );
  OAI22_X1 U7681 ( .A1(n6220), .A2(n9451), .B1(n9453), .B2(n6219), .ZN(n6221)
         );
  AOI211_X1 U7682 ( .C1(n9782), .C2(n9477), .A(n6222), .B(n6221), .ZN(n6223)
         );
  INV_X1 U7683 ( .A(n6223), .ZN(n6224) );
  NOR2_X1 U7684 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND3_X1 U7685 ( .A1(n6228), .A2(n6227), .A3(n6226), .ZN(P1_U3218) );
  INV_X1 U7686 ( .A(n6258), .ZN(n6229) );
  NOR2_X1 U7687 ( .A1(n5930), .A2(n6229), .ZN(n6274) );
  AND2_X2 U7688 ( .A1(n6274), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U7689 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6233) );
  NOR2_X1 U7690 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6535) );
  NOR2_X1 U7691 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6534) );
  NOR2_X1 U7692 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6234) );
  NAND4_X1 U7693 ( .A1(n4543), .A2(n6535), .A3(n6534), .A4(n6234), .ZN(n6238)
         );
  INV_X1 U7694 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6236) );
  INV_X1 U7695 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6235) );
  NAND4_X1 U7696 ( .A1(n6236), .A2(n6538), .A3(n6235), .A4(n6542), .ZN(n6237)
         );
  NAND2_X1 U7697 ( .A1(n6246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6335) );
  INV_X1 U7698 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7699 ( .A1(n6335), .A2(n6241), .ZN(n6242) );
  NAND2_X1 U7700 ( .A1(n6242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6256) );
  INV_X1 U7701 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7702 ( .A1(n6256), .A2(n6255), .ZN(n6243) );
  NAND2_X1 U7703 ( .A1(n6243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6245) );
  INV_X1 U7704 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6244) );
  XNOR2_X1 U7705 ( .A(n6245), .B(n6244), .ZN(n7525) );
  INV_X1 U7706 ( .A(n7525), .ZN(n6517) );
  NOR3_X1 U7707 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7708 ( .A1(n6342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6250) );
  MUX2_X1 U7709 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6250), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6251) );
  NAND2_X1 U7710 ( .A1(n6251), .A2(n6338), .ZN(n7742) );
  NAND2_X1 U7711 ( .A1(n6252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6253) );
  XNOR2_X1 U7712 ( .A(n6253), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6519) );
  INV_X1 U7713 ( .A(n6519), .ZN(n7729) );
  NOR2_X1 U7714 ( .A1(n7742), .A2(n7729), .ZN(n6254) );
  AND2_X1 U7715 ( .A1(n6517), .A2(n6254), .ZN(n6407) );
  XNOR2_X1 U7716 ( .A(n6256), .B(n6255), .ZN(n6659) );
  AND2_X1 U7717 ( .A1(n6659), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10225) );
  AND2_X1 U7718 ( .A1(n6407), .A2(n10225), .ZN(P2_U3966) );
  NAND2_X1 U7719 ( .A1(n5930), .A2(n6257), .ZN(n6259) );
  NAND2_X1 U7720 ( .A1(n6259), .A2(n6258), .ZN(n6272) );
  NAND2_X1 U7721 ( .A1(n6272), .A2(n6260), .ZN(n6290) );
  NAND2_X1 U7722 ( .A1(n6290), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  MUX2_X1 U7723 ( .A(n6261), .B(P1_REG2_REG_12__SCAN_IN), .S(n6288), .Z(n7109)
         );
  NOR2_X1 U7724 ( .A1(n10026), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6262) );
  AOI21_X1 U7725 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10026), .A(n6262), .ZN(
        n10018) );
  NAND2_X1 U7726 ( .A1(n6687), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7727 ( .B1(n6687), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6263), .ZN(
        n6684) );
  XNOR2_X1 U7728 ( .A(n6350), .B(n7094), .ZN(n6397) );
  NOR2_X1 U7729 ( .A1(n10004), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6264) );
  AOI21_X1 U7730 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n10004), .A(n6264), .ZN(
        n10006) );
  INV_X1 U7731 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n8450) );
  INV_X1 U7732 ( .A(n9978), .ZN(n6326) );
  AOI22_X1 U7733 ( .A1(n9978), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n8450), .B2(
        n6326), .ZN(n9981) );
  NAND2_X1 U7734 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9956) );
  NOR2_X1 U7735 ( .A1(n9956), .A2(n9941), .ZN(n9940) );
  AOI21_X1 U7736 ( .B1(n9936), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9940), .ZN(
        n9952) );
  NAND2_X1 U7737 ( .A1(n9946), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U7738 ( .B1(n9946), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6265), .ZN(
        n9951) );
  NAND2_X1 U7739 ( .A1(n6302), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6266) );
  OAI21_X1 U7740 ( .B1(n6302), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6266), .ZN(
        n6300) );
  INV_X1 U7741 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6267) );
  INV_X1 U7742 ( .A(n6284), .ZN(n9970) );
  AOI22_X1 U7743 ( .A1(n6284), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6267), .B2(
        n9970), .ZN(n9964) );
  NAND2_X1 U7744 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  OAI21_X1 U7745 ( .B1(n6284), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9963), .ZN(
        n9980) );
  XNOR2_X1 U7746 ( .A(n9996), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7747 ( .A1(n10006), .A2(n10007), .ZN(n10005) );
  INV_X1 U7748 ( .A(n6350), .ZN(n6402) );
  AOI21_X1 U7749 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6687), .A(n6683), .ZN(
        n6801) );
  NAND2_X1 U7750 ( .A1(n6803), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7751 ( .B1(n6803), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6268), .ZN(
        n6800) );
  NOR2_X1 U7752 ( .A1(n6801), .A2(n6800), .ZN(n6799) );
  NAND2_X1 U7753 ( .A1(n7342), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6269) );
  OAI21_X1 U7754 ( .B1(n7342), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6269), .ZN(
        n7339) );
  INV_X1 U7755 ( .A(n6289), .ZN(n7720) );
  NOR2_X1 U7756 ( .A1(n6270), .A2(n7720), .ZN(n6271) );
  NOR2_X1 U7757 ( .A1(n5925), .A2(P1_U3084), .ZN(n7783) );
  NAND2_X1 U7758 ( .A1(n6272), .A2(n7783), .ZN(n9544) );
  OR2_X1 U7759 ( .A1(n9544), .A2(n5922), .ZN(n10032) );
  AOI211_X1 U7760 ( .C1(n6273), .C2(n5673), .A(n9498), .B(n10032), .ZN(n6295)
         );
  OR2_X1 U7761 ( .A1(P1_U3083), .A2(n6274), .ZN(n10046) );
  INV_X1 U7762 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6275) );
  NOR2_X1 U7763 ( .A1(n10046), .A2(n6275), .ZN(n6294) );
  INV_X1 U7764 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8529) );
  INV_X1 U7765 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6276) );
  MUX2_X1 U7766 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6276), .S(n6289), .Z(n7717)
         );
  INV_X1 U7767 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6277) );
  INV_X1 U7768 ( .A(n7342), .ZN(n6488) );
  AOI22_X1 U7769 ( .A1(n7342), .A2(P1_REG1_REG_13__SCAN_IN), .B1(n6277), .B2(
        n6488), .ZN(n7335) );
  INV_X1 U7770 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6278) );
  MUX2_X1 U7771 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6278), .S(n6288), .Z(n7104)
         );
  INV_X1 U7772 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6279) );
  AOI22_X1 U7773 ( .A1(n10026), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n6279), .B2(
        n6378), .ZN(n10025) );
  INV_X1 U7774 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U7775 ( .A1(n6803), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n9889), .B2(
        n6375), .ZN(n6795) );
  INV_X1 U7776 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U7777 ( .A1(n6687), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10167), .B2(
        n6360), .ZN(n6690) );
  INV_X1 U7778 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6286) );
  MUX2_X1 U7779 ( .A(n6286), .B(P1_REG1_REG_8__SCAN_IN), .S(n6350), .Z(n6399)
         );
  NOR2_X1 U7780 ( .A1(n10004), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6280) );
  AOI21_X1 U7781 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10004), .A(n6280), .ZN(
        n10010) );
  XNOR2_X1 U7782 ( .A(n9996), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U7783 ( .A1(n9978), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6281) );
  OAI21_X1 U7784 ( .B1(n9978), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6281), .ZN(
        n9984) );
  INV_X1 U7785 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U7786 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10157), .S(n6284), .Z(n9969)
         );
  INV_X1 U7787 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9957) );
  INV_X1 U7788 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U7789 ( .A1(n9936), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7790 ( .B1(n9936), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6282), .ZN(
        n9938) );
  NOR3_X1 U7791 ( .A1(n9957), .A2(n9930), .A3(n9938), .ZN(n9937) );
  AOI21_X1 U7792 ( .B1(n9936), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9937), .ZN(
        n9949) );
  XNOR2_X1 U7793 ( .A(n9946), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9948) );
  NOR2_X1 U7794 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  AOI21_X1 U7795 ( .B1(n9946), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9947), .ZN(
        n6298) );
  NAND2_X1 U7796 ( .A1(n6302), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6283) );
  OAI21_X1 U7797 ( .B1(n6302), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6283), .ZN(
        n6297) );
  NOR2_X1 U7798 ( .A1(n6298), .A2(n6297), .ZN(n6296) );
  AOI21_X1 U7799 ( .B1(n6302), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6296), .ZN(
        n9968) );
  NAND2_X1 U7800 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  OAI21_X1 U7801 ( .B1(n6284), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9967), .ZN(
        n9985) );
  NOR2_X1 U7802 ( .A1(n9984), .A2(n9985), .ZN(n9983) );
  AOI21_X1 U7803 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9978), .A(n9983), .ZN(
        n6285) );
  INV_X1 U7804 ( .A(n6285), .ZN(n9997) );
  NAND2_X1 U7805 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  OAI21_X1 U7806 ( .B1(n10004), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10008), .ZN(
        n6400) );
  NAND2_X1 U7807 ( .A1(n6399), .A2(n6400), .ZN(n6398) );
  NAND2_X1 U7808 ( .A1(n6350), .A2(n6286), .ZN(n6287) );
  NAND2_X1 U7809 ( .A1(n6398), .A2(n6287), .ZN(n6689) );
  NAND2_X1 U7810 ( .A1(n6690), .A2(n6689), .ZN(n6688) );
  OAI21_X1 U7811 ( .B1(n6687), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6688), .ZN(
        n6796) );
  NAND2_X1 U7812 ( .A1(n6795), .A2(n6796), .ZN(n6794) );
  OAI21_X1 U7813 ( .B1(n6803), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6794), .ZN(
        n10024) );
  NAND2_X1 U7814 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  OAI21_X1 U7815 ( .B1(n10026), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10023), .ZN(
        n7105) );
  NAND2_X1 U7816 ( .A1(n7104), .A2(n7105), .ZN(n7103) );
  OAI21_X1 U7817 ( .B1(n6288), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7103), .ZN(
        n7336) );
  NAND2_X1 U7818 ( .A1(n7335), .A2(n7336), .ZN(n7334) );
  OAI21_X1 U7819 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7342), .A(n7334), .ZN(
        n7718) );
  NAND2_X1 U7820 ( .A1(n7717), .A2(n7718), .ZN(n7716) );
  OAI21_X1 U7821 ( .B1(n6289), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7716), .ZN(
        n9502) );
  XNOR2_X1 U7822 ( .A(n9503), .B(n9502), .ZN(n6291) );
  NOR2_X1 U7823 ( .A1(n8529), .A2(n6291), .ZN(n9504) );
  NOR2_X1 U7824 ( .A1(n6290), .A2(P1_U3084), .ZN(n9932) );
  NAND2_X1 U7825 ( .A1(n9932), .A2(n5925), .ZN(n9982) );
  AOI211_X1 U7826 ( .C1(n8529), .C2(n6291), .A(n9504), .B(n9982), .ZN(n6293)
         );
  OR2_X1 U7827 ( .A1(n9544), .A2(n9929), .ZN(n9971) );
  NAND2_X1 U7828 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7858) );
  OAI21_X1 U7829 ( .B1(n9971), .B2(n9503), .A(n7858), .ZN(n6292) );
  OR4_X1 U7830 ( .A1(n6295), .A2(n6294), .A3(n6293), .A4(n6292), .ZN(P1_U3256)
         );
  NOR2_X1 U7831 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6499), .ZN(n6494) );
  AOI211_X1 U7832 ( .C1(n6298), .C2(n6297), .A(n6296), .B(n9982), .ZN(n6305)
         );
  AOI211_X1 U7833 ( .C1(n6301), .C2(n6300), .A(n6299), .B(n10032), .ZN(n6304)
         );
  INV_X1 U7834 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7550) );
  INV_X1 U7835 ( .A(n6302), .ZN(n6328) );
  OAI22_X1 U7836 ( .A1(n10046), .A2(n7550), .B1(n6328), .B2(n9971), .ZN(n6303)
         );
  OR4_X1 U7837 ( .A1(n6494), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(P1_U3244)
         );
  NOR2_X1 U7838 ( .A1(n6554), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9327) );
  INV_X1 U7839 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6306) );
  AND2_X1 U7840 ( .A1(n6554), .A2(P2_U3152), .ZN(n7385) );
  OAI222_X1 U7841 ( .A1(n9330), .A2(n6306), .B1(n4490), .B2(n6555), .C1(
        P2_U3152), .C2(n8376), .ZN(P2_U3357) );
  NOR2_X1 U7842 ( .A1(n6307), .A2(n9324), .ZN(n6308) );
  MUX2_X1 U7843 ( .A(n9324), .B(n6308), .S(P2_IR_REG_2__SCAN_IN), .Z(n6309) );
  INV_X1 U7844 ( .A(n6309), .ZN(n6311) );
  INV_X1 U7845 ( .A(n6313), .ZN(n6310) );
  NAND2_X1 U7846 ( .A1(n6311), .A2(n6310), .ZN(n6612) );
  OAI222_X1 U7847 ( .A1(n9330), .A2(n6611), .B1(n4490), .B2(n6610), .C1(
        P2_U3152), .C2(n6612), .ZN(P2_U3356) );
  INV_X1 U7848 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6647) );
  OR2_X1 U7849 ( .A1(n6313), .A2(n9324), .ZN(n6312) );
  XNOR2_X1 U7850 ( .A(n6312), .B(n8770), .ZN(n6648) );
  OAI222_X1 U7851 ( .A1(n9330), .A2(n6647), .B1(n4490), .B2(n6646), .C1(
        P2_U3152), .C2(n6648), .ZN(P2_U3355) );
  NAND2_X1 U7852 ( .A1(n6313), .A2(n8770), .ZN(n6320) );
  NAND2_X1 U7853 ( .A1(n6320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6315) );
  XNOR2_X1 U7854 ( .A(n6315), .B(n6314), .ZN(n6743) );
  OAI222_X1 U7855 ( .A1(n9330), .A2(n6740), .B1(n4490), .B2(n6739), .C1(
        P2_U3152), .C2(n6743), .ZN(P2_U3354) );
  OAI222_X1 U7856 ( .A1(n8383), .A2(n6317), .B1(n9881), .B2(n6739), .C1(
        P1_U3084), .C2(n9970), .ZN(P1_U3349) );
  INV_X1 U7857 ( .A(n8383), .ZN(n9875) );
  AOI22_X1 U7858 ( .A1(n9875), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9946), .ZN(n6318) );
  OAI21_X1 U7859 ( .B1(n6610), .B2(n9881), .A(n6318), .ZN(P1_U3351) );
  AOI22_X1 U7860 ( .A1(n9875), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9936), .ZN(n6319) );
  OAI21_X1 U7861 ( .B1(n6555), .B2(n9881), .A(n6319), .ZN(P1_U3352) );
  NOR2_X1 U7862 ( .A1(n6320), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6324) );
  INV_X1 U7863 ( .A(n6324), .ZN(n6321) );
  NAND2_X1 U7864 ( .A1(n6321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U7865 ( .A(n6322), .B(P2_IR_REG_31__SCAN_IN), .S(n6323), .Z(n6325)
         );
  NAND2_X1 U7866 ( .A1(n6324), .A2(n6323), .ZN(n6333) );
  NAND2_X1 U7867 ( .A1(n6325), .A2(n6333), .ZN(n6841) );
  OAI222_X1 U7868 ( .A1(n9330), .A2(n6839), .B1(n4490), .B2(n6838), .C1(
        P2_U3152), .C2(n6841), .ZN(P2_U3353) );
  OAI222_X1 U7869 ( .A1(n8383), .A2(n6327), .B1(n9881), .B2(n6838), .C1(
        P1_U3084), .C2(n6326), .ZN(P1_U3348) );
  INV_X1 U7870 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6329) );
  OAI222_X1 U7871 ( .A1(n8383), .A2(n6329), .B1(n9881), .B2(n6646), .C1(
        P1_U3084), .C2(n6328), .ZN(P1_U3350) );
  OAI222_X1 U7872 ( .A1(n8383), .A2(n6331), .B1(n9881), .B2(n6916), .C1(
        P1_U3084), .C2(n6330), .ZN(P1_U3347) );
  NAND2_X1 U7873 ( .A1(n6333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6332) );
  MUX2_X1 U7874 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6332), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6334) );
  OR2_X1 U7875 ( .A1(n6333), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6352) );
  INV_X1 U7876 ( .A(n6670), .ZN(n6918) );
  OAI222_X1 U7877 ( .A1(n9330), .A2(n6917), .B1(n4490), .B2(n6916), .C1(
        P2_U3152), .C2(n6918), .ZN(P2_U3352) );
  INV_X1 U7878 ( .A(n6407), .ZN(n6660) );
  NAND2_X1 U7879 ( .A1(n6660), .A2(n10225), .ZN(n10212) );
  NAND2_X1 U7880 ( .A1(n6336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6337) );
  XNOR2_X1 U7881 ( .A(n6337), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8220) );
  AND2_X1 U7882 ( .A1(n8357), .A2(n8220), .ZN(n6575) );
  INV_X1 U7883 ( .A(n6575), .ZN(n6729) );
  INV_X1 U7884 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6340) );
  INV_X1 U7885 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7886 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  XNOR2_X2 U7887 ( .A(n6344), .B(n6364), .ZN(n6411) );
  OAI21_X1 U7888 ( .B1(n10212), .B2(n6729), .A(n6955), .ZN(n6346) );
  OR2_X1 U7889 ( .A1(n6659), .A2(P2_U3152), .ZN(n8360) );
  NAND2_X1 U7890 ( .A1(n10212), .A2(n8360), .ZN(n6345) );
  AND2_X1 U7891 ( .A1(n6346), .A2(n6345), .ZN(n10187) );
  NOR2_X1 U7892 ( .A1(n10187), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7893 ( .A(n7059), .ZN(n6351) );
  OR2_X1 U7894 ( .A1(n6347), .A2(n9324), .ZN(n6348) );
  XNOR2_X1 U7895 ( .A(n6348), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7060) );
  INV_X1 U7896 ( .A(n7060), .ZN(n6775) );
  OAI222_X1 U7897 ( .A1(n9330), .A2(n6349), .B1(n4490), .B2(n6351), .C1(
        P2_U3152), .C2(n6775), .ZN(P2_U3350) );
  OAI222_X1 U7898 ( .A1(n8383), .A2(n8664), .B1(n9881), .B2(n6351), .C1(
        P1_U3084), .C2(n6350), .ZN(P1_U3345) );
  INV_X1 U7899 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6355) );
  INV_X1 U7900 ( .A(n6958), .ZN(n6357) );
  NAND2_X1 U7901 ( .A1(n6352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6353) );
  MUX2_X1 U7902 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6353), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6354) );
  INV_X1 U7903 ( .A(n6956), .ZN(n8920) );
  OAI222_X1 U7904 ( .A1(n9330), .A2(n6355), .B1(n4490), .B2(n6357), .C1(
        P2_U3152), .C2(n8920), .ZN(P2_U3351) );
  OAI222_X1 U7905 ( .A1(n8383), .A2(n6358), .B1(n9881), .B2(n6357), .C1(
        P1_U3084), .C2(n6356), .ZN(P1_U3346) );
  INV_X1 U7906 ( .A(n7213), .ZN(n6363) );
  OAI222_X1 U7907 ( .A1(n9881), .A2(n6363), .B1(n6360), .B2(P1_U3084), .C1(
        n6359), .C2(n8383), .ZN(P1_U3344) );
  NAND2_X1 U7908 ( .A1(n6373), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6361) );
  XNOR2_X1 U7909 ( .A(n6361), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7214) );
  INV_X1 U7910 ( .A(n7214), .ZN(n7023) );
  OAI222_X1 U7911 ( .A1(P2_U3152), .A2(n7023), .B1(n4490), .B2(n6363), .C1(
        n6362), .C2(n9330), .ZN(P2_U3349) );
  NAND2_X1 U7912 ( .A1(n6366), .A2(n6365), .ZN(n9325) );
  INV_X1 U7913 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8980) );
  AND2_X2 U7914 ( .A1(n8382), .A2(n6503), .ZN(n8046) );
  NAND2_X1 U7915 ( .A1(n8046), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U7916 ( .A1(n8382), .A2(n9332), .ZN(n6615) );
  INV_X1 U7917 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7918 ( .A1(n8121), .A2(n6369), .ZN(n6370) );
  OAI211_X1 U7919 ( .C1(n8083), .C2(n8980), .A(n6371), .B(n6370), .ZN(n8982)
         );
  NAND2_X1 U7920 ( .A1(n8982), .A2(P2_U3966), .ZN(n6372) );
  OAI21_X1 U7921 ( .B1(n5231), .B2(P2_U3966), .A(n6372), .ZN(P2_U3583) );
  INV_X1 U7922 ( .A(n7316), .ZN(n6376) );
  NAND2_X1 U7923 ( .A1(n6385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6380) );
  XNOR2_X1 U7924 ( .A(n6380), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7317) );
  AOI22_X1 U7925 ( .A1(n7317), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9327), .ZN(n6374) );
  OAI21_X1 U7926 ( .B1(n6376), .B2(n4490), .A(n6374), .ZN(P2_U3348) );
  OAI222_X1 U7927 ( .A1(n9881), .A2(n6376), .B1(n6375), .B2(P1_U3084), .C1(
        n8670), .C2(n8383), .ZN(P1_U3343) );
  INV_X1 U7928 ( .A(n7418), .ZN(n6383) );
  OAI222_X1 U7929 ( .A1(n9881), .A2(n6383), .B1(n6378), .B2(P1_U3084), .C1(
        n6377), .C2(n8383), .ZN(P1_U3342) );
  NAND2_X1 U7930 ( .A1(n6380), .A2(n6379), .ZN(n6381) );
  NAND2_X1 U7931 ( .A1(n6381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U7932 ( .A(n6382), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7475) );
  INV_X1 U7933 ( .A(n7475), .ZN(n7471) );
  OAI222_X1 U7934 ( .A1(n9330), .A2(n6384), .B1(n4490), .B2(n6383), .C1(n7471), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7935 ( .A(n7575), .ZN(n6394) );
  OR2_X1 U7936 ( .A1(n6537), .A2(n9324), .ZN(n6386) );
  XNOR2_X1 U7937 ( .A(n6386), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7611) );
  AOI22_X1 U7938 ( .A1(n7611), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9327), .ZN(n6387) );
  OAI21_X1 U7939 ( .B1(n6394), .B2(n4490), .A(n6387), .ZN(P2_U3346) );
  OAI21_X1 U7940 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n9955) );
  AOI22_X1 U7941 ( .A1(n9428), .A2(n9955), .B1(n9477), .B2(n6828), .ZN(n6393)
         );
  INV_X1 U7942 ( .A(n9451), .ZN(n9476) );
  NAND2_X1 U7943 ( .A1(n6496), .A2(n6811), .ZN(n6599) );
  AOI22_X1 U7944 ( .A1(n9476), .A2(n6391), .B1(n6599), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7945 ( .A1(n6393), .A2(n6392), .ZN(P1_U3230) );
  OAI222_X1 U7946 ( .A1(n8383), .A2(n6395), .B1(n9881), .B2(n6394), .C1(
        P1_U3084), .C2(n7107), .ZN(P1_U3341) );
  XNOR2_X1 U7947 ( .A(n6397), .B(n6396), .ZN(n6405) );
  INV_X1 U7948 ( .A(n9982), .ZN(n10043) );
  OAI21_X1 U7949 ( .B1(n6400), .B2(n6399), .A(n6398), .ZN(n6401) );
  INV_X1 U7950 ( .A(n10046), .ZN(n9999) );
  AOI22_X1 U7951 ( .A1(n10043), .A2(n6401), .B1(n9999), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n6404) );
  INV_X1 U7952 ( .A(n9971), .ZN(n10038) );
  INV_X1 U7953 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8588) );
  NOR2_X1 U7954 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8588), .ZN(n7122) );
  AOI21_X1 U7955 ( .B1(n10038), .B2(n6402), .A(n7122), .ZN(n6403) );
  OAI211_X1 U7956 ( .C1(n6405), .C2(n10032), .A(n6404), .B(n6403), .ZN(
        P1_U3249) );
  OR2_X1 U7957 ( .A1(n10212), .A2(n6575), .ZN(n6409) );
  INV_X1 U7958 ( .A(n8360), .ZN(n6406) );
  AOI21_X1 U7959 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6407), .A(n6406), .ZN(n6408) );
  NAND2_X1 U7960 ( .A1(n6409), .A2(n6408), .ZN(n6416) );
  NAND2_X1 U7961 ( .A1(n6416), .A2(n6955), .ZN(n6410) );
  INV_X2 U7962 ( .A(P2_U3966), .ZN(n8913) );
  NAND2_X1 U7963 ( .A1(n6410), .A2(n8913), .ZN(n6421) );
  INV_X1 U7964 ( .A(n6411), .ZN(n6515) );
  NAND2_X1 U7965 ( .A1(n6421), .A2(n6411), .ZN(n10170) );
  INV_X1 U7966 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8665) );
  NOR2_X1 U7967 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8665), .ZN(n6760) );
  INV_X1 U7968 ( .A(n6648), .ZN(n6424) );
  INV_X1 U7969 ( .A(n6612), .ZN(n6413) );
  INV_X1 U7970 ( .A(n8376), .ZN(n6412) );
  NAND2_X1 U7971 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n8367) );
  NOR2_X1 U7972 ( .A1(n8366), .A2(n8367), .ZN(n8365) );
  AOI21_X1 U7973 ( .B1(n6412), .B2(P2_REG1_REG_1__SCAN_IN), .A(n8365), .ZN(
        n6433) );
  XOR2_X1 U7974 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6612), .Z(n6432) );
  NOR2_X1 U7975 ( .A1(n6433), .A2(n6432), .ZN(n6431) );
  INV_X1 U7976 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6414) );
  MUX2_X1 U7977 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6414), .S(n6648), .Z(n6443)
         );
  XOR2_X1 U7978 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6743), .Z(n6417) );
  AND2_X1 U7979 ( .A1(n6955), .A2(n8408), .ZN(n6415) );
  AND2_X1 U7980 ( .A1(n6416), .A2(n6415), .ZN(n10181) );
  INV_X1 U7981 ( .A(n10181), .ZN(n10171) );
  AOI211_X1 U7982 ( .C1(n6418), .C2(n6417), .A(n6454), .B(n10171), .ZN(n6419)
         );
  AOI211_X1 U7983 ( .C1(n10187), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6760), .B(
        n6419), .ZN(n6430) );
  NOR2_X1 U7984 ( .A1(n6411), .A2(n8408), .ZN(n6420) );
  NAND2_X1 U7985 ( .A1(n6421), .A2(n6420), .ZN(n10172) );
  INV_X1 U7986 ( .A(n10172), .ZN(n10185) );
  INV_X1 U7987 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7187) );
  MUX2_X1 U7988 ( .A(n7187), .B(P2_REG2_REG_2__SCAN_IN), .S(n6612), .Z(n6438)
         );
  INV_X1 U7989 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8370) );
  MUX2_X1 U7990 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8370), .S(n8376), .Z(n6423)
         );
  INV_X1 U7991 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6509) );
  INV_X1 U7992 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6422) );
  OR3_X1 U7993 ( .A1(n6423), .A2(n6509), .A3(n6422), .ZN(n8371) );
  OAI21_X1 U7994 ( .B1(n8376), .B2(n8370), .A(n8371), .ZN(n6437) );
  NAND2_X1 U7995 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  INV_X1 U7996 ( .A(n6436), .ZN(n6449) );
  NOR2_X1 U7997 ( .A1(n6612), .A2(n7187), .ZN(n6448) );
  INV_X1 U7998 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7150) );
  MUX2_X1 U7999 ( .A(n7150), .B(P2_REG2_REG_3__SCAN_IN), .S(n6648), .Z(n6447)
         );
  OAI21_X1 U8000 ( .B1(n6449), .B2(n6448), .A(n6447), .ZN(n6451) );
  NAND2_X1 U8001 ( .A1(n6424), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6426) );
  INV_X1 U8002 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6463) );
  MUX2_X1 U8003 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6463), .S(n6743), .Z(n6425)
         );
  AOI21_X1 U8004 ( .B1(n6451), .B2(n6426), .A(n6425), .ZN(n6474) );
  INV_X1 U8005 ( .A(n6474), .ZN(n6428) );
  NAND3_X1 U8006 ( .A1(n6451), .A2(n6426), .A3(n6425), .ZN(n6427) );
  NAND3_X1 U8007 ( .A1(n10185), .A2(n6428), .A3(n6427), .ZN(n6429) );
  OAI211_X1 U8008 ( .C1(n10170), .C2(n6743), .A(n6430), .B(n6429), .ZN(
        P2_U3249) );
  INV_X1 U8009 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U8010 ( .A1(n7189), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6435) );
  AOI211_X1 U8011 ( .C1(n6433), .C2(n6432), .A(n6431), .B(n10171), .ZN(n6434)
         );
  AOI211_X1 U8012 ( .C1(n10187), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n6435), .B(
        n6434), .ZN(n6440) );
  OAI211_X1 U8013 ( .C1(n6438), .C2(n6437), .A(n10185), .B(n6436), .ZN(n6439)
         );
  OAI211_X1 U8014 ( .C1(n10170), .C2(n6612), .A(n6440), .B(n6439), .ZN(
        P2_U3247) );
  INV_X1 U8015 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6441) );
  NOR2_X1 U8016 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6441), .ZN(n6446) );
  AOI211_X1 U8017 ( .C1(n6444), .C2(n6443), .A(n6442), .B(n10171), .ZN(n6445)
         );
  AOI211_X1 U8018 ( .C1(n10187), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6446), .B(
        n6445), .ZN(n6453) );
  OR3_X1 U8019 ( .A1(n6449), .A2(n6448), .A3(n6447), .ZN(n6450) );
  NAND3_X1 U8020 ( .A1(n10185), .A2(n6451), .A3(n6450), .ZN(n6452) );
  OAI211_X1 U8021 ( .C1(n10170), .C2(n6648), .A(n6453), .B(n6452), .ZN(
        P2_U3248) );
  NAND2_X1 U8022 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6939) );
  INV_X1 U8023 ( .A(n6939), .ZN(n6462) );
  INV_X1 U8024 ( .A(n6841), .ZN(n6457) );
  INV_X1 U8025 ( .A(n6743), .ZN(n6455) );
  AOI21_X1 U8026 ( .B1(n6455), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6454), .ZN(
        n6470) );
  INV_X1 U8027 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6456) );
  MUX2_X1 U8028 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6456), .S(n6841), .Z(n6469)
         );
  NAND2_X1 U8029 ( .A1(n6670), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6458) );
  OAI21_X1 U8030 ( .B1(n6670), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6458), .ZN(
        n6459) );
  AOI211_X1 U8031 ( .C1(n6460), .C2(n6459), .A(n10171), .B(n6666), .ZN(n6461)
         );
  AOI211_X1 U8032 ( .C1(n10187), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6462), .B(
        n6461), .ZN(n6467) );
  INV_X1 U8033 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U8034 ( .A1(n6743), .A2(n6463), .ZN(n6473) );
  MUX2_X1 U8035 ( .A(n6464), .B(P2_REG2_REG_5__SCAN_IN), .S(n6841), .Z(n6475)
         );
  OAI21_X1 U8036 ( .B1(n6474), .B2(n6473), .A(n6475), .ZN(n6477) );
  OAI21_X1 U8037 ( .B1(n6464), .B2(n6841), .A(n6477), .ZN(n6673) );
  INV_X1 U8038 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7354) );
  MUX2_X1 U8039 ( .A(n7354), .B(P2_REG2_REG_6__SCAN_IN), .S(n6670), .Z(n6671)
         );
  XNOR2_X1 U8040 ( .A(n6673), .B(n6671), .ZN(n6465) );
  NAND2_X1 U8041 ( .A1(n10185), .A2(n6465), .ZN(n6466) );
  OAI211_X1 U8042 ( .C1(n10170), .C2(n6918), .A(n6467), .B(n6466), .ZN(
        P2_U3251) );
  NAND2_X1 U8043 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6861) );
  INV_X1 U8044 ( .A(n6861), .ZN(n6472) );
  AOI211_X1 U8045 ( .C1(n6470), .C2(n6469), .A(n10171), .B(n6468), .ZN(n6471)
         );
  AOI211_X1 U8046 ( .C1(n10187), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6472), .B(
        n6471), .ZN(n6479) );
  OR3_X1 U8047 ( .A1(n6475), .A2(n6474), .A3(n6473), .ZN(n6476) );
  NAND3_X1 U8048 ( .A1(n10185), .A2(n6477), .A3(n6476), .ZN(n6478) );
  OAI211_X1 U8049 ( .C1(n10170), .C2(n6841), .A(n6479), .B(n6478), .ZN(
        P2_U3250) );
  NOR2_X1 U8050 ( .A1(n6814), .A2(n10090), .ZN(n10088) );
  AND3_X1 U8051 ( .A1(n6812), .A2(n6480), .A3(n6811), .ZN(n6481) );
  AND2_X1 U8052 ( .A1(n10088), .A2(n6481), .ZN(n9776) );
  INV_X1 U8053 ( .A(n9871), .ZN(n6815) );
  AND2_X2 U8054 ( .A1(n9776), .A2(n6815), .ZN(n10150) );
  INV_X1 U8055 ( .A(n10058), .ZN(n9737) );
  AND3_X1 U8056 ( .A1(n6483), .A2(n6978), .A3(n6482), .ZN(n6484) );
  AOI21_X1 U8057 ( .B1(n9737), .B2(n6391), .A(n6484), .ZN(n10071) );
  INV_X1 U8058 ( .A(n6978), .ZN(n6485) );
  NAND2_X1 U8059 ( .A1(n6828), .A2(n6485), .ZN(n10070) );
  NAND2_X1 U8060 ( .A1(n10071), .A2(n10070), .ZN(n9854) );
  NAND2_X1 U8061 ( .A1(n9854), .A2(n10150), .ZN(n6486) );
  OAI21_X1 U8062 ( .B1(n10150), .B2(n5513), .A(n6486), .ZN(P1_U3454) );
  INV_X1 U8063 ( .A(n7622), .ZN(n6490) );
  OAI222_X1 U8064 ( .A1(n9881), .A2(n6490), .B1(n6488), .B2(P1_U3084), .C1(
        n6487), .C2(n8383), .ZN(P1_U3340) );
  INV_X1 U8065 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U8066 ( .A1(n6537), .A2(n8481), .ZN(n6489) );
  NAND2_X1 U8067 ( .A1(n6489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6583) );
  XNOR2_X1 U8068 ( .A(n6583), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7644) );
  INV_X1 U8069 ( .A(n7644), .ZN(n7640) );
  OAI222_X1 U8070 ( .A1(n9330), .A2(n6491), .B1(n4490), .B2(n6490), .C1(n7640), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  XOR2_X1 U8071 ( .A(n6493), .B(n6492), .Z(n6501) );
  INV_X1 U8072 ( .A(n9428), .ZN(n9470) );
  INV_X1 U8073 ( .A(n9453), .ZN(n9475) );
  INV_X1 U8074 ( .A(n6494), .ZN(n6495) );
  OAI21_X1 U8075 ( .B1(n9451), .B2(n6898), .A(n6495), .ZN(n6498) );
  INV_X1 U8076 ( .A(n6496), .ZN(n7381) );
  NAND2_X1 U8077 ( .A1(n6889), .A2(n10139), .ZN(n10103) );
  OAI22_X1 U8078 ( .A1(n7381), .A2(n10103), .B1(n9464), .B2(n10059), .ZN(n6497) );
  AOI211_X1 U8079 ( .C1(n9475), .C2(n6499), .A(n6498), .B(n6497), .ZN(n6500)
         );
  OAI21_X1 U8080 ( .B1(n6501), .B2(n9470), .A(n6500), .ZN(P1_U3216) );
  INV_X1 U8081 ( .A(n7785), .ZN(n6587) );
  OAI222_X1 U8082 ( .A1(n9881), .A2(n6587), .B1(n7720), .B2(P1_U3084), .C1(
        n6502), .C2(n8383), .ZN(P1_U3339) );
  NAND2_X1 U8083 ( .A1(n8046), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6508) );
  OR2_X1 U8084 ( .A1(n8083), .A2(n7187), .ZN(n6507) );
  OR2_X1 U8085 ( .A1(n6634), .A2(n7189), .ZN(n6506) );
  OR2_X1 U8086 ( .A1(n6615), .A2(n10238), .ZN(n6505) );
  AND4_X2 U8087 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n6998)
         );
  NAND2_X1 U8088 ( .A1(n6411), .A2(n6575), .ZN(n9184) );
  NAND2_X1 U8089 ( .A1(n8046), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6514) );
  OR2_X1 U8090 ( .A1(n8083), .A2(n6509), .ZN(n6513) );
  INV_X1 U8091 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7362) );
  OR2_X1 U8092 ( .A1(n6634), .A2(n7362), .ZN(n6512) );
  INV_X1 U8093 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6510) );
  OR2_X1 U8094 ( .A1(n6615), .A2(n6510), .ZN(n6511) );
  NAND4_X2 U8095 ( .A1(n6513), .A2(n6514), .A3(n6512), .A4(n6511), .ZN(n8914)
         );
  AND2_X1 U8096 ( .A1(n6515), .A2(n6575), .ZN(n9195) );
  NAND2_X1 U8097 ( .A1(n8914), .A2(n9195), .ZN(n6516) );
  OAI21_X1 U8098 ( .B1(n6998), .B2(n9184), .A(n6516), .ZN(n7275) );
  INV_X1 U8099 ( .A(n7275), .ZN(n6581) );
  INV_X1 U8100 ( .A(P2_B_REG_SCAN_IN), .ZN(n8453) );
  AOI22_X1 U8101 ( .A1(P2_B_REG_SCAN_IN), .A2(n7525), .B1(n6517), .B2(n8453), 
        .ZN(n6518) );
  NOR2_X1 U8102 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NOR2_X1 U8103 ( .A1(n6520), .A2(n7742), .ZN(n10211) );
  INV_X1 U8104 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10220) );
  AND2_X1 U8105 ( .A1(n7742), .A2(n7525), .ZN(n10221) );
  AOI21_X1 U8106 ( .B1(n10211), .B2(n10220), .A(n10221), .ZN(n7140) );
  NOR4_X1 U8107 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6529) );
  NOR4_X1 U8108 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6528) );
  INV_X1 U8109 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10218) );
  INV_X1 U8110 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10215) );
  INV_X1 U8111 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10216) );
  INV_X1 U8112 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U8113 ( .A1(n10218), .A2(n10215), .A3(n10216), .A4(n10214), .ZN(
        n6526) );
  NOR4_X1 U8114 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6524) );
  NOR4_X1 U8115 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6523) );
  NOR4_X1 U8116 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6522) );
  NOR4_X1 U8117 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6521) );
  NAND4_X1 U8118 ( .A1(n6524), .A2(n6523), .A3(n6522), .A4(n6521), .ZN(n6525)
         );
  NOR4_X1 U8119 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6526), .A4(n6525), .ZN(n6527) );
  AND3_X1 U8120 ( .A1(n6529), .A2(n6528), .A3(n6527), .ZN(n6531) );
  INV_X1 U8121 ( .A(n10211), .ZN(n6530) );
  NOR2_X1 U8122 ( .A1(n6531), .A2(n6530), .ZN(n6728) );
  INV_X1 U8123 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8124 ( .A1(n10211), .A2(n6532), .ZN(n6533) );
  NAND2_X1 U8125 ( .A1(n7742), .A2(n7729), .ZN(n10222) );
  NAND2_X1 U8126 ( .A1(n6533), .A2(n10222), .ZN(n6724) );
  NOR2_X1 U8127 ( .A1(n6728), .A2(n6724), .ZN(n7138) );
  NAND2_X1 U8128 ( .A1(n7140), .A2(n7138), .ZN(n6577) );
  OR2_X1 U8129 ( .A1(n6577), .A2(n10212), .ZN(n6574) );
  AND2_X1 U8130 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND2_X1 U8131 ( .A1(n6694), .A2(n6538), .ZN(n6766) );
  INV_X1 U8132 ( .A(n6766), .ZN(n6539) );
  NAND2_X1 U8133 ( .A1(n6539), .A2(n6236), .ZN(n6540) );
  INV_X1 U8134 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U8135 ( .A1(n6541), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6543) );
  NOR2_X1 U8136 ( .A1(n6574), .A2(n8356), .ZN(n6763) );
  INV_X1 U8137 ( .A(n6763), .ZN(n6969) );
  NAND2_X1 U8138 ( .A1(n6554), .A2(SI_0_), .ZN(n6546) );
  INV_X1 U8139 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8480) );
  NAND2_X1 U8140 ( .A1(n6546), .A2(n8480), .ZN(n6548) );
  AND2_X1 U8141 ( .A1(n6548), .A2(n6547), .ZN(n9333) );
  MUX2_X1 U8142 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9333), .S(n6955), .Z(n7279) );
  NAND2_X1 U8143 ( .A1(n8914), .A2(n7279), .ZN(n7277) );
  INV_X1 U8144 ( .A(n7277), .ZN(n6553) );
  INV_X1 U8145 ( .A(n8357), .ZN(n7313) );
  OR2_X2 U8146 ( .A1(n8356), .A2(n8354), .ZN(n8176) );
  NOR2_X1 U8147 ( .A1(n7279), .A2(n8116), .ZN(n6552) );
  AOI21_X1 U8148 ( .B1(n6553), .B2(n8176), .A(n6552), .ZN(n6569) );
  INV_X1 U8149 ( .A(n6565), .ZN(n6564) );
  NAND2_X1 U8150 ( .A1(n8046), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6562) );
  INV_X1 U8151 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6557) );
  OR2_X1 U8152 ( .A1(n6634), .A2(n6557), .ZN(n6560) );
  INV_X1 U8153 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6558) );
  OR2_X1 U8154 ( .A1(n6615), .A2(n6558), .ZN(n6559) );
  INV_X1 U8155 ( .A(n6566), .ZN(n6563) );
  NAND2_X1 U8156 ( .A1(n6564), .A2(n6563), .ZN(n6608) );
  NAND2_X1 U8157 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  NAND2_X1 U8158 ( .A1(n6568), .A2(n6569), .ZN(n6609) );
  OAI21_X1 U8159 ( .B1(n6569), .B2(n6568), .A(n6609), .ZN(n6572) );
  INV_X1 U8160 ( .A(n6574), .ZN(n6571) );
  AND2_X1 U8161 ( .A1(n8356), .A2(n7011), .ZN(n6570) );
  INV_X1 U8162 ( .A(n6570), .ZN(n10275) );
  NAND3_X1 U8163 ( .A1(n6571), .A2(n10275), .A3(n6729), .ZN(n8866) );
  INV_X1 U8164 ( .A(n8866), .ZN(n8882) );
  NAND2_X1 U8165 ( .A1(n6572), .A2(n8882), .ZN(n6580) );
  OR2_X1 U8166 ( .A1(n6549), .A2(n8354), .ZN(n7151) );
  AND2_X1 U8167 ( .A1(n9188), .A2(n7313), .ZN(n6573) );
  OAI21_X2 U8168 ( .B1(n6574), .B2(n7151), .A(n10199), .ZN(n8848) );
  INV_X1 U8169 ( .A(n10212), .ZN(n6576) );
  NAND2_X1 U8170 ( .A1(n8356), .A2(n6575), .ZN(n6658) );
  NAND2_X1 U8171 ( .A1(n6576), .A2(n6658), .ZN(n7142) );
  INV_X1 U8172 ( .A(n7142), .ZN(n6578) );
  NAND2_X1 U8173 ( .A1(n6725), .A2(n6577), .ZN(n6661) );
  NAND2_X1 U8174 ( .A1(n6578), .A2(n6661), .ZN(n6613) );
  AOI22_X1 U8175 ( .A1(n8848), .A2(n7278), .B1(n6613), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6579) );
  OAI211_X1 U8176 ( .C1(n6581), .C2(n6969), .A(n6580), .B(n6579), .ZN(P2_U3224) );
  INV_X1 U8177 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U8178 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  NAND2_X1 U8179 ( .A1(n6584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6585) );
  INV_X1 U8180 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U8181 ( .A1(n6585), .A2(n8592), .ZN(n6698) );
  OR2_X1 U8182 ( .A1(n6585), .A2(n8592), .ZN(n6586) );
  AND2_X1 U8183 ( .A1(n6698), .A2(n6586), .ZN(n7870) );
  INV_X1 U8184 ( .A(n7870), .ZN(n7865) );
  OAI222_X1 U8185 ( .A1(n9330), .A2(n8436), .B1(n4490), .B2(n6587), .C1(n7865), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  XNOR2_X1 U8186 ( .A(n6590), .B(n6589), .ZN(n6591) );
  XNOR2_X1 U8187 ( .A(n6588), .B(n6591), .ZN(n6595) );
  OAI22_X1 U8188 ( .A1(n10057), .A2(n9464), .B1(n9451), .B2(n10059), .ZN(n6593) );
  INV_X1 U8189 ( .A(n9477), .ZN(n9372) );
  NOR2_X1 U8190 ( .A1(n9372), .A2(n10092), .ZN(n6592) );
  AOI211_X1 U8191 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6599), .A(n6593), .B(
        n6592), .ZN(n6594) );
  OAI21_X1 U8192 ( .B1(n9470), .B2(n6595), .A(n6594), .ZN(P1_U3220) );
  INV_X1 U8193 ( .A(n9495), .ZN(n6823) );
  OAI22_X1 U8194 ( .A1(n6817), .A2(n9464), .B1(n9451), .B2(n6823), .ZN(n6598)
         );
  NOR2_X1 U8195 ( .A1(n9372), .A2(n10096), .ZN(n6597) );
  AOI211_X1 U8196 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n6599), .A(n6598), .B(
        n6597), .ZN(n6600) );
  OAI21_X1 U8197 ( .B1(n9470), .B2(n6601), .A(n6600), .ZN(P1_U3235) );
  INV_X1 U8198 ( .A(n8848), .ZN(n8893) );
  INV_X1 U8199 ( .A(n7279), .ZN(n7363) );
  NAND2_X1 U8200 ( .A1(n8914), .A2(n7363), .ZN(n8231) );
  MUX2_X1 U8201 ( .A(n8231), .B(n7363), .S(n6602), .Z(n6604) );
  INV_X1 U8202 ( .A(n8914), .ZN(n6603) );
  AOI21_X1 U8203 ( .B1(n6604), .B2(n7274), .A(n8866), .ZN(n6605) );
  INV_X1 U8204 ( .A(n6605), .ZN(n6607) );
  INV_X1 U8205 ( .A(n9184), .ZN(n9197) );
  AND2_X1 U8206 ( .A1(n6763), .A2(n9197), .ZN(n8875) );
  AOI22_X1 U8207 ( .A1(n8912), .A2(n8875), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n6613), .ZN(n6606) );
  OAI211_X1 U8208 ( .C1(n8893), .C2(n7363), .A(n6607), .B(n6606), .ZN(P2_U3234) );
  NAND2_X1 U8209 ( .A1(n6609), .A2(n6608), .ZN(n6645) );
  OR2_X1 U8210 ( .A1(n6998), .A2(n6602), .ZN(n6642) );
  XNOR2_X1 U8211 ( .A(n8094), .B(n7191), .ZN(n6643) );
  XNOR2_X1 U8212 ( .A(n6642), .B(n6643), .ZN(n6644) );
  XNOR2_X1 U8213 ( .A(n6645), .B(n6644), .ZN(n6622) );
  AOI22_X1 U8214 ( .A1(n8848), .A2(n7191), .B1(n6613), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U8215 ( .A1(n8046), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6619) );
  OR2_X1 U8216 ( .A1(n8083), .A2(n7150), .ZN(n6618) );
  OR2_X1 U8217 ( .A1(n6634), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6617) );
  INV_X1 U8218 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6614) );
  OR2_X1 U8219 ( .A1(n6615), .A2(n6614), .ZN(n6616) );
  NAND4_X1 U8220 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n8910)
         );
  INV_X1 U8221 ( .A(n8910), .ZN(n7007) );
  INV_X1 U8222 ( .A(n9195), .ZN(n9182) );
  OAI22_X1 U8223 ( .A1(n7007), .A2(n9184), .B1(n6995), .B2(n9182), .ZN(n7185)
         );
  NAND2_X1 U8224 ( .A1(n7185), .A2(n6763), .ZN(n6620) );
  OAI211_X1 U8225 ( .C1(n6622), .C2(n8866), .A(n6621), .B(n6620), .ZN(P2_U3239) );
  INV_X1 U8226 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6961) );
  INV_X1 U8227 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7063) );
  INV_X1 U8228 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7225) );
  INV_X1 U8229 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7421) );
  INV_X1 U8230 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7626) );
  INV_X1 U8231 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7795) );
  INV_X1 U8232 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8949) );
  AND2_X1 U8233 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n6629) );
  INV_X1 U8234 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8844) );
  INV_X1 U8235 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8800) );
  INV_X1 U8236 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8024) );
  INV_X1 U8237 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U8238 ( .A1(n8027), .A2(n6632), .ZN(n6633) );
  NAND2_X1 U8239 ( .A1(n8044), .A2(n6633), .ZN(n9085) );
  OR2_X1 U8240 ( .A1(n9085), .A2(n6634), .ZN(n6640) );
  INV_X1 U8241 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U8242 ( .A1(n8158), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6636) );
  INV_X1 U8243 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9084) );
  OR2_X1 U8244 ( .A1(n8083), .A2(n9084), .ZN(n6635) );
  OAI211_X1 U8245 ( .C1(n8162), .C2(n6637), .A(n6636), .B(n6635), .ZN(n6638)
         );
  INV_X1 U8246 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U8247 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8913), .ZN(n6641) );
  OAI21_X1 U8248 ( .B1(n9108), .B2(n8913), .A(n6641), .ZN(P2_U3575) );
  OR2_X1 U8249 ( .A1(n6957), .A2(n6646), .ZN(n6651) );
  OR2_X1 U8250 ( .A1(n8167), .A2(n6647), .ZN(n6650) );
  OR2_X1 U8251 ( .A1(n6955), .A2(n6648), .ZN(n6649) );
  XNOR2_X1 U8252 ( .A(n8238), .B(n8094), .ZN(n6748) );
  NAND2_X1 U8253 ( .A1(n8910), .A2(n8176), .ZN(n6747) );
  XNOR2_X1 U8254 ( .A(n6748), .B(n6747), .ZN(n6745) );
  XNOR2_X1 U8255 ( .A(n6746), .B(n6745), .ZN(n6665) );
  INV_X1 U8256 ( .A(n6998), .ZN(n8911) );
  NAND2_X1 U8257 ( .A1(n8046), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6656) );
  OR2_X1 U8258 ( .A1(n8083), .A2(n6463), .ZN(n6655) );
  OAI21_X1 U8259 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n6854), .ZN(n10200) );
  OR2_X1 U8260 ( .A1(n6634), .A2(n10200), .ZN(n6654) );
  INV_X1 U8261 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6652) );
  OR2_X1 U8262 ( .A1(n6615), .A2(n6652), .ZN(n6653) );
  INV_X1 U8263 ( .A(n7003), .ZN(n8909) );
  AOI22_X1 U8264 ( .A1(n9195), .A2(n8911), .B1(n8909), .B2(n9197), .ZN(n7147)
         );
  INV_X1 U8265 ( .A(n7147), .ZN(n6657) );
  AOI22_X1 U8266 ( .A1(n6657), .A2(n6763), .B1(n10241), .B2(n8848), .ZN(n6664)
         );
  NAND4_X1 U8267 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n6662)
         );
  AND2_X1 U8268 ( .A1(n6662), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8871) );
  INV_X1 U8269 ( .A(n8871), .ZN(n8885) );
  MUX2_X1 U8270 ( .A(n8885), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6663) );
  OAI211_X1 U8271 ( .C1(n6665), .C2(n8866), .A(n6664), .B(n6663), .ZN(P2_U3220) );
  XNOR2_X1 U8272 ( .A(n6956), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n8916) );
  NOR2_X1 U8273 ( .A1(n8917), .A2(n8916), .ZN(n8915) );
  INV_X1 U8274 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6667) );
  MUX2_X1 U8275 ( .A(n6667), .B(P2_REG1_REG_8__SCAN_IN), .S(n7060), .Z(n6668)
         );
  AOI211_X1 U8276 ( .C1(n6669), .C2(n6668), .A(n10171), .B(n6770), .ZN(n6682)
         );
  INV_X1 U8277 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U8278 ( .A1(n6670), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6675) );
  INV_X1 U8279 ( .A(n6671), .ZN(n6672) );
  NAND2_X1 U8280 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U8281 ( .A1(n6675), .A2(n6674), .ZN(n8925) );
  MUX2_X1 U8282 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7166), .S(n6956), .Z(n8924)
         );
  NAND2_X1 U8283 ( .A1(n8925), .A2(n8924), .ZN(n8923) );
  OAI21_X1 U8284 ( .B1(n7166), .B2(n8920), .A(n8923), .ZN(n6677) );
  INV_X1 U8285 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7265) );
  MUX2_X1 U8286 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7265), .S(n7060), .Z(n6676)
         );
  NAND2_X1 U8287 ( .A1(n6676), .A2(n6677), .ZN(n6774) );
  OAI211_X1 U8288 ( .C1(n6677), .C2(n6676), .A(n10185), .B(n6774), .ZN(n6680)
         );
  NAND2_X1 U8289 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7071) );
  INV_X1 U8290 ( .A(n7071), .ZN(n6678) );
  AOI21_X1 U8291 ( .B1(n10187), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6678), .ZN(
        n6679) );
  OAI211_X1 U8292 ( .C1(n10170), .C2(n6775), .A(n6680), .B(n6679), .ZN(n6681)
         );
  OR2_X1 U8293 ( .A1(n6682), .A2(n6681), .ZN(P2_U3253) );
  AND2_X1 U8294 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7133) );
  AOI211_X1 U8295 ( .C1(n6685), .C2(n6684), .A(n6683), .B(n10032), .ZN(n6686)
         );
  AOI211_X1 U8296 ( .C1(n10038), .C2(n6687), .A(n7133), .B(n6686), .ZN(n6693)
         );
  OAI21_X1 U8297 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(n6691) );
  AOI22_X1 U8298 ( .A1(n10043), .A2(n6691), .B1(n9999), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8299 ( .A1(n6693), .A2(n6692), .ZN(P1_U3250) );
  INV_X1 U8300 ( .A(n7937), .ZN(n6713) );
  OR2_X1 U8301 ( .A1(n6694), .A2(n9324), .ZN(n6695) );
  XNOR2_X1 U8302 ( .A(n6695), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8955) );
  AOI22_X1 U8303 ( .A1(n8955), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9327), .ZN(n6696) );
  OAI21_X1 U8304 ( .B1(n6713), .B2(n4490), .A(n6696), .ZN(P2_U3342) );
  INV_X1 U8305 ( .A(n7792), .ZN(n6700) );
  OAI222_X1 U8306 ( .A1(n8383), .A2(n6697), .B1(n9881), .B2(n6700), .C1(
        P1_U3084), .C2(n9503), .ZN(P1_U3338) );
  NAND2_X1 U8307 ( .A1(n6698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6699) );
  XNOR2_X1 U8308 ( .A(n6699), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8930) );
  INV_X1 U8309 ( .A(n8930), .ZN(n8938) );
  OAI222_X1 U8310 ( .A1(n9330), .A2(n6701), .B1(n4490), .B2(n6700), .C1(
        P2_U3152), .C2(n8938), .ZN(P2_U3343) );
  NAND2_X1 U8311 ( .A1(n6985), .A2(n10139), .ZN(n10118) );
  XNOR2_X1 U8312 ( .A(n6703), .B(n6702), .ZN(n6704) );
  XNOR2_X1 U8313 ( .A(n6705), .B(n6704), .ZN(n6706) );
  NAND2_X1 U8314 ( .A1(n6706), .A2(n9428), .ZN(n6712) );
  INV_X1 U8315 ( .A(n6707), .ZN(n6976) );
  OAI22_X1 U8316 ( .A1(n6898), .A2(n9464), .B1(n9453), .B2(n6976), .ZN(n6710)
         );
  AND2_X1 U8317 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9987) );
  INV_X1 U8318 ( .A(n9987), .ZN(n6708) );
  OAI21_X1 U8319 ( .B1(n9451), .B2(n7037), .A(n6708), .ZN(n6709) );
  NOR2_X1 U8320 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  OAI211_X1 U8321 ( .C1(n7381), .C2(n10118), .A(n6712), .B(n6711), .ZN(
        P1_U3225) );
  OAI222_X1 U8322 ( .A1(n8383), .A2(n6714), .B1(n9515), .B2(P1_U3084), .C1(
        n9881), .C2(n6713), .ZN(P1_U3337) );
  INV_X1 U8323 ( .A(n6715), .ZN(n6716) );
  AOI211_X1 U8324 ( .C1(n6718), .C2(n6717), .A(n9470), .B(n6716), .ZN(n6723)
         );
  NAND2_X1 U8325 ( .A1(n6834), .A2(n10139), .ZN(n10109) );
  OAI22_X1 U8326 ( .A1(n7381), .A2(n10109), .B1(n9464), .B2(n6823), .ZN(n6722)
         );
  INV_X1 U8327 ( .A(n6719), .ZN(n6832) );
  AND2_X1 U8328 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9973) );
  AOI21_X1 U8329 ( .B1(n9476), .B2(n9493), .A(n9973), .ZN(n6720) );
  OAI21_X1 U8330 ( .B1(n6832), .B2(n9453), .A(n6720), .ZN(n6721) );
  OR3_X1 U8331 ( .A1(n6723), .A2(n6722), .A3(n6721), .ZN(P1_U3228) );
  NAND2_X1 U8332 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  OR2_X1 U8333 ( .A1(n6726), .A2(n7142), .ZN(n6727) );
  NOR2_X1 U8334 ( .A1(n6728), .A2(n6727), .ZN(n6736) );
  NAND2_X1 U8335 ( .A1(n6736), .A2(n7140), .ZN(n10293) );
  INV_X2 U8336 ( .A(n10293), .ZN(n10295) );
  INV_X1 U8337 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8338 ( .A1(n7274), .A2(n8231), .ZN(n8178) );
  NAND2_X1 U8339 ( .A1(n8352), .A2(n8220), .ZN(n8175) );
  NAND2_X1 U8340 ( .A1(n9188), .A2(n8357), .ZN(n8353) );
  NAND2_X1 U8341 ( .A1(n8175), .A2(n8353), .ZN(n10194) );
  AOI22_X1 U8342 ( .A1(n8178), .A2(n10194), .B1(n9197), .B2(n8912), .ZN(n7361)
         );
  MUX2_X1 U8343 ( .A(n6729), .B(n8357), .S(n8352), .Z(n6731) );
  NAND2_X1 U8344 ( .A1(n6731), .A2(n6730), .ZN(n7754) );
  INV_X1 U8345 ( .A(n9297), .ZN(n10279) );
  AOI22_X1 U8346 ( .A1(n8178), .A2(n10279), .B1(n7011), .B2(n7279), .ZN(n6732)
         );
  NAND2_X1 U8347 ( .A1(n7361), .A2(n6732), .ZN(n6737) );
  NAND2_X1 U8348 ( .A1(n6737), .A2(n10295), .ZN(n6733) );
  OAI21_X1 U8349 ( .B1(n10295), .B2(n6734), .A(n6733), .ZN(P2_U3520) );
  INV_X1 U8350 ( .A(n7140), .ZN(n6735) );
  NAND2_X1 U8351 ( .A1(n6736), .A2(n6735), .ZN(n10281) );
  INV_X2 U8352 ( .A(n10281), .ZN(n9320) );
  NAND2_X1 U8353 ( .A1(n6737), .A2(n9320), .ZN(n6738) );
  OAI21_X1 U8354 ( .B1(n9320), .B2(n6510), .A(n6738), .ZN(P2_U3451) );
  OR2_X1 U8355 ( .A1(n7003), .A2(n6602), .ZN(n6744) );
  OR2_X1 U8356 ( .A1(n6957), .A2(n6739), .ZN(n6742) );
  OR2_X1 U8357 ( .A1(n8167), .A2(n6740), .ZN(n6741) );
  NAND2_X1 U8358 ( .A1(n6746), .A2(n6745), .ZN(n6751) );
  INV_X1 U8359 ( .A(n6747), .ZN(n6749) );
  NAND2_X1 U8360 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  NAND2_X1 U8361 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  INV_X1 U8362 ( .A(n6848), .ZN(n6752) );
  AOI21_X1 U8363 ( .B1(n6754), .B2(n6753), .A(n6752), .ZN(n6765) );
  NAND2_X1 U8364 ( .A1(n8046), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6759) );
  OR2_X1 U8365 ( .A1(n8083), .A2(n6464), .ZN(n6758) );
  INV_X1 U8366 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6853) );
  XNOR2_X1 U8367 ( .A(n6854), .B(n6853), .ZN(n7173) );
  OR2_X1 U8368 ( .A1(n6634), .A2(n7173), .ZN(n6757) );
  INV_X1 U8369 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6755) );
  OR2_X1 U8370 ( .A1(n6615), .A2(n6755), .ZN(n6756) );
  NAND4_X1 U8371 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n8908)
         );
  INV_X1 U8372 ( .A(n8908), .ZN(n6994) );
  OAI22_X1 U8373 ( .A1(n7007), .A2(n9182), .B1(n6994), .B2(n9184), .ZN(n10193)
         );
  AOI21_X1 U8374 ( .B1(n8848), .B2(n10206), .A(n6760), .ZN(n6761) );
  OAI21_X1 U8375 ( .B1(n8885), .B2(n10200), .A(n6761), .ZN(n6762) );
  AOI21_X1 U8376 ( .B1(n10193), .B2(n6763), .A(n6762), .ZN(n6764) );
  OAI21_X1 U8377 ( .B1(n6765), .B2(n8866), .A(n6764), .ZN(P2_U3232) );
  INV_X1 U8378 ( .A(n7946), .ZN(n6768) );
  NAND2_X1 U8379 ( .A1(n6766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6767) );
  XNOR2_X1 U8380 ( .A(n6767), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8971) );
  INV_X1 U8381 ( .A(n8971), .ZN(n8962) );
  OAI222_X1 U8382 ( .A1(n9330), .A2(n8667), .B1(n4490), .B2(n6768), .C1(n8962), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI222_X1 U8383 ( .A1(n8383), .A2(n6769), .B1(n9524), .B2(P1_U3084), .C1(
        n9881), .C2(n6768), .ZN(P1_U3336) );
  INV_X1 U8384 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6771) );
  MUX2_X1 U8385 ( .A(n6771), .B(P2_REG1_REG_9__SCAN_IN), .S(n7214), .Z(n6772)
         );
  AOI211_X1 U8386 ( .C1(n6773), .C2(n6772), .A(n7017), .B(n10171), .ZN(n6782)
         );
  OAI21_X1 U8387 ( .B1(n6775), .B2(n7265), .A(n6774), .ZN(n6777) );
  INV_X1 U8388 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7400) );
  MUX2_X1 U8389 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7400), .S(n7214), .Z(n6776)
         );
  NAND2_X1 U8390 ( .A1(n6776), .A2(n6777), .ZN(n7022) );
  OAI211_X1 U8391 ( .C1(n6777), .C2(n6776), .A(n10185), .B(n7022), .ZN(n6780)
         );
  NAND2_X1 U8392 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7233) );
  INV_X1 U8393 ( .A(n7233), .ZN(n6778) );
  AOI21_X1 U8394 ( .B1(n10187), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6778), .ZN(
        n6779) );
  OAI211_X1 U8395 ( .C1(n10170), .C2(n7023), .A(n6780), .B(n6779), .ZN(n6781)
         );
  OR2_X1 U8396 ( .A1(n6782), .A2(n6781), .ZN(P2_U3254) );
  XNOR2_X1 U8397 ( .A(n6784), .B(n6783), .ZN(n6785) );
  XNOR2_X1 U8398 ( .A(n6786), .B(n6785), .ZN(n6787) );
  NAND2_X1 U8399 ( .A1(n6787), .A2(n9428), .ZN(n6793) );
  INV_X1 U8400 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U8401 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6788), .ZN(n9995) );
  OAI22_X1 U8402 ( .A1(n6790), .A2(n9464), .B1(n9453), .B2(n6789), .ZN(n6791)
         );
  AOI211_X1 U8403 ( .C1(n9476), .C2(n9491), .A(n9995), .B(n6791), .ZN(n6792)
         );
  OAI211_X1 U8404 ( .C1(n4781), .C2(n9372), .A(n6793), .B(n6792), .ZN(P1_U3237) );
  INV_X1 U8405 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6806) );
  OAI21_X1 U8406 ( .B1(n6796), .B2(n6795), .A(n6794), .ZN(n6797) );
  NAND2_X1 U8407 ( .A1(n6797), .A2(n10043), .ZN(n6805) );
  NOR2_X1 U8408 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6798), .ZN(n7374) );
  AOI211_X1 U8409 ( .C1(n6801), .C2(n6800), .A(n6799), .B(n10032), .ZN(n6802)
         );
  AOI211_X1 U8410 ( .C1(n10038), .C2(n6803), .A(n7374), .B(n6802), .ZN(n6804)
         );
  OAI211_X1 U8411 ( .C1(n10046), .C2(n6806), .A(n6805), .B(n6804), .ZN(
        P1_U3251) );
  NAND2_X1 U8412 ( .A1(n5923), .A2(n10054), .ZN(n6808) );
  NAND2_X1 U8413 ( .A1(n5929), .A2(n6977), .ZN(n6807) );
  XNOR2_X1 U8414 ( .A(n6809), .B(n6895), .ZN(n6810) );
  AOI222_X1 U8415 ( .A1(n10061), .A2(n6810), .B1(n9493), .B2(n9737), .C1(n9495), .C2(n9735), .ZN(n10110) );
  AND3_X1 U8416 ( .A1(n10080), .A2(n6812), .A3(n6811), .ZN(n6813) );
  NAND3_X1 U8417 ( .A1(n6815), .A2(n6814), .A3(n6813), .ZN(n7041) );
  INV_X2 U8418 ( .A(n10075), .ZN(n10078) );
  NAND2_X1 U8419 ( .A1(n5941), .A2(n6828), .ZN(n10047) );
  NAND2_X1 U8420 ( .A1(n6816), .A2(n10047), .ZN(n6819) );
  NAND2_X1 U8421 ( .A1(n6817), .A2(n10092), .ZN(n6818) );
  NAND2_X1 U8422 ( .A1(n6819), .A2(n6818), .ZN(n6867) );
  NAND2_X1 U8423 ( .A1(n6867), .A2(n6871), .ZN(n6821) );
  NAND2_X1 U8424 ( .A1(n10059), .A2(n10096), .ZN(n6820) );
  NAND2_X1 U8425 ( .A1(n6821), .A2(n6820), .ZN(n6882) );
  NAND2_X1 U8426 ( .A1(n6882), .A2(n6822), .ZN(n6825) );
  NAND2_X1 U8427 ( .A1(n6823), .A2(n6887), .ZN(n6824) );
  NAND2_X1 U8428 ( .A1(n6825), .A2(n6824), .ZN(n6896) );
  XNOR2_X1 U8429 ( .A(n6896), .B(n6895), .ZN(n10113) );
  AND2_X1 U8430 ( .A1(n6826), .A2(n10054), .ZN(n10067) );
  NAND2_X1 U8431 ( .A1(n10075), .A2(n10067), .ZN(n9767) );
  INV_X1 U8432 ( .A(n10064), .ZN(n10148) );
  NAND2_X1 U8433 ( .A1(n10075), .A2(n10148), .ZN(n6827) );
  INV_X1 U8434 ( .A(n9750), .ZN(n7311) );
  NAND2_X1 U8435 ( .A1(n6888), .A2(n6887), .ZN(n6886) );
  INV_X1 U8436 ( .A(n6886), .ZN(n6830) );
  INV_X1 U8437 ( .A(n6981), .ZN(n6829) );
  OAI21_X1 U8438 ( .B1(n6897), .B2(n6830), .A(n6829), .ZN(n10111) );
  AND2_X1 U8439 ( .A1(n10075), .A2(n6831), .ZN(n9770) );
  INV_X1 U8440 ( .A(n9770), .ZN(n7097) );
  NOR2_X1 U8441 ( .A1(n6978), .A2(n7102), .ZN(n10051) );
  NAND2_X1 U8442 ( .A1(n10075), .A2(n10051), .ZN(n9766) );
  INV_X1 U8443 ( .A(n9766), .ZN(n7711) );
  OAI22_X1 U8444 ( .A1(n10075), .A2(n6267), .B1(n6832), .B2(n7922), .ZN(n6833)
         );
  AOI21_X1 U8445 ( .B1(n7711), .B2(n6834), .A(n6833), .ZN(n6835) );
  OAI21_X1 U8446 ( .B1(n10111), .B2(n7097), .A(n6835), .ZN(n6836) );
  AOI21_X1 U8447 ( .B1(n10113), .B2(n7311), .A(n6836), .ZN(n6837) );
  OAI21_X1 U8448 ( .B1(n10110), .B2(n10078), .A(n6837), .ZN(P1_U3287) );
  OR2_X1 U8449 ( .A1(n8167), .A2(n6839), .ZN(n6840) );
  AND2_X1 U8450 ( .A1(n8908), .A2(n8176), .ZN(n6842) );
  XNOR2_X1 U8451 ( .A(n7156), .B(n8116), .ZN(n6843) );
  NAND2_X1 U8452 ( .A1(n6842), .A2(n6843), .ZN(n6846) );
  INV_X1 U8453 ( .A(n6842), .ZN(n6845) );
  INV_X1 U8454 ( .A(n6843), .ZN(n6844) );
  NAND2_X1 U8455 ( .A1(n6845), .A2(n6844), .ZN(n6927) );
  AND2_X1 U8456 ( .A1(n6846), .A2(n6927), .ZN(n6850) );
  OAI21_X1 U8457 ( .B1(n6850), .B2(n6849), .A(n6928), .ZN(n6851) );
  NAND2_X1 U8458 ( .A1(n6851), .A2(n8882), .ZN(n6866) );
  INV_X1 U8459 ( .A(n7173), .ZN(n6864) );
  OR2_X1 U8460 ( .A1(n6969), .A2(n9182), .ZN(n8873) );
  NAND2_X1 U8461 ( .A1(n8046), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6860) );
  OR2_X1 U8462 ( .A1(n8083), .A2(n7354), .ZN(n6859) );
  INV_X1 U8463 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6852) );
  OAI21_X1 U8464 ( .B1(n6854), .B2(n6853), .A(n6852), .ZN(n6855) );
  NAND2_X1 U8465 ( .A1(n6855), .A2(n6932), .ZN(n7355) );
  OR2_X1 U8466 ( .A1(n6634), .A2(n7355), .ZN(n6858) );
  INV_X1 U8467 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6856) );
  OR2_X1 U8468 ( .A1(n8121), .A2(n6856), .ZN(n6857) );
  NAND2_X1 U8469 ( .A1(n8907), .A2(n8875), .ZN(n6862) );
  OAI211_X1 U8470 ( .C1(n7003), .C2(n8873), .A(n6862), .B(n6861), .ZN(n6863)
         );
  AOI21_X1 U8471 ( .B1(n6864), .B2(n8871), .A(n6863), .ZN(n6865) );
  OAI211_X1 U8472 ( .C1(n7174), .C2(n8893), .A(n6866), .B(n6865), .ZN(P2_U3229) );
  XNOR2_X1 U8473 ( .A(n6871), .B(n6867), .ZN(n10100) );
  INV_X1 U8474 ( .A(n10100), .ZN(n6881) );
  INV_X1 U8475 ( .A(n6868), .ZN(n6869) );
  AOI21_X1 U8476 ( .B1(n6871), .B2(n6870), .A(n6869), .ZN(n6874) );
  INV_X1 U8477 ( .A(n10061), .ZN(n7036) );
  AOI22_X1 U8478 ( .A1(n9735), .A2(n6391), .B1(n9495), .B2(n9737), .ZN(n6873)
         );
  NAND2_X1 U8479 ( .A1(n10100), .A2(n10148), .ZN(n6872) );
  OAI211_X1 U8480 ( .C1(n6874), .C2(n7036), .A(n6873), .B(n6872), .ZN(n10098)
         );
  NAND2_X1 U8481 ( .A1(n10098), .A2(n10075), .ZN(n6880) );
  INV_X1 U8482 ( .A(n6888), .ZN(n6875) );
  OAI21_X1 U8483 ( .B1(n10096), .B2(n10048), .A(n6875), .ZN(n10097) );
  INV_X1 U8484 ( .A(n7922), .ZN(n10074) );
  AOI22_X1 U8485 ( .A1(n10078), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10074), .ZN(n6876) );
  OAI21_X1 U8486 ( .B1(n7097), .B2(n10097), .A(n6876), .ZN(n6877) );
  AOI21_X1 U8487 ( .B1(n7711), .B2(n6878), .A(n6877), .ZN(n6879) );
  OAI211_X1 U8488 ( .C1(n6881), .C2(n9767), .A(n6880), .B(n6879), .ZN(P1_U3289) );
  XNOR2_X1 U8489 ( .A(n6882), .B(n6883), .ZN(n10102) );
  XNOR2_X1 U8490 ( .A(n6884), .B(n6883), .ZN(n6885) );
  AOI222_X1 U8491 ( .A1(n10061), .A2(n6885), .B1(n9494), .B2(n9737), .C1(n9496), .C2(n9735), .ZN(n10104) );
  INV_X1 U8492 ( .A(n10104), .ZN(n6893) );
  OAI21_X1 U8493 ( .B1(n6888), .B2(n6887), .A(n6886), .ZN(n10105) );
  AOI22_X1 U8494 ( .A1(n10078), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10074), .B2(
        n6499), .ZN(n6891) );
  NAND2_X1 U8495 ( .A1(n7711), .A2(n6889), .ZN(n6890) );
  OAI211_X1 U8496 ( .C1(n7097), .C2(n10105), .A(n6891), .B(n6890), .ZN(n6892)
         );
  AOI21_X1 U8497 ( .B1(n6893), .B2(n10075), .A(n6892), .ZN(n6894) );
  OAI21_X1 U8498 ( .B1(n9750), .B2(n10102), .A(n6894), .ZN(P1_U3288) );
  NAND2_X1 U8499 ( .A1(n6896), .A2(n6895), .ZN(n6900) );
  NAND2_X1 U8500 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  NAND2_X1 U8501 ( .A1(n6900), .A2(n6899), .ZN(n6987) );
  NAND2_X1 U8502 ( .A1(n9493), .A2(n6985), .ZN(n6901) );
  XNOR2_X1 U8503 ( .A(n7030), .B(n7029), .ZN(n10123) );
  INV_X1 U8504 ( .A(n10123), .ZN(n6912) );
  OAI211_X1 U8505 ( .C1(n6903), .C2(n7029), .A(n6902), .B(n10061), .ZN(n6905)
         );
  AOI22_X1 U8506 ( .A1(n9735), .A2(n9493), .B1(n9491), .B2(n9737), .ZN(n6904)
         );
  NAND2_X1 U8507 ( .A1(n6905), .A2(n6904), .ZN(n10121) );
  OAI21_X1 U8508 ( .B1(n4782), .B2(n4781), .A(n7039), .ZN(n10120) );
  AOI22_X1 U8509 ( .A1(n10078), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6906), .B2(
        n10074), .ZN(n6909) );
  NAND2_X1 U8510 ( .A1(n7711), .A2(n6907), .ZN(n6908) );
  OAI211_X1 U8511 ( .C1(n10120), .C2(n7097), .A(n6909), .B(n6908), .ZN(n6910)
         );
  AOI21_X1 U8512 ( .B1(n10121), .B2(n10075), .A(n6910), .ZN(n6911) );
  OAI21_X1 U8513 ( .B1(n9750), .B2(n6912), .A(n6911), .ZN(P1_U3285) );
  INV_X1 U8514 ( .A(n7959), .ZN(n6915) );
  OAI222_X1 U8515 ( .A1(n8383), .A2(n6913), .B1(n9881), .B2(n6915), .C1(
        P1_U3084), .C2(n9539), .ZN(P1_U3335) );
  INV_X1 U8516 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8712) );
  XNOR2_X1 U8517 ( .A(n6914), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10182) );
  INV_X1 U8518 ( .A(n10182), .ZN(n8965) );
  OAI222_X1 U8519 ( .A1(n9330), .A2(n8712), .B1(n4490), .B2(n6915), .C1(
        P2_U3152), .C2(n8965), .ZN(P2_U3340) );
  OR2_X1 U8520 ( .A1(n6957), .A2(n6916), .ZN(n6921) );
  OR2_X1 U8521 ( .A1(n8167), .A2(n6917), .ZN(n6920) );
  OR2_X1 U8522 ( .A1(n6955), .A2(n6918), .ZN(n6919) );
  AND3_X2 U8523 ( .A1(n6921), .A2(n6920), .A3(n6919), .ZN(n10253) );
  NOR2_X1 U8524 ( .A1(n8230), .A2(n6602), .ZN(n6922) );
  XNOR2_X1 U8525 ( .A(n10253), .B(n8094), .ZN(n6923) );
  NAND2_X1 U8526 ( .A1(n6922), .A2(n6923), .ZN(n6926) );
  INV_X1 U8527 ( .A(n6922), .ZN(n6925) );
  INV_X1 U8528 ( .A(n6923), .ZN(n6924) );
  NAND2_X1 U8529 ( .A1(n6925), .A2(n6924), .ZN(n6953) );
  AND2_X1 U8530 ( .A1(n6926), .A2(n6953), .ZN(n6930) );
  OAI21_X1 U8531 ( .B1(n6930), .B2(n6929), .A(n6954), .ZN(n6931) );
  NAND2_X1 U8532 ( .A1(n6931), .A2(n8882), .ZN(n6944) );
  INV_X1 U8533 ( .A(n7355), .ZN(n6942) );
  NAND2_X1 U8534 ( .A1(n8046), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6938) );
  OR2_X1 U8535 ( .A1(n8083), .A2(n7166), .ZN(n6937) );
  INV_X1 U8536 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U8537 ( .A1(n6932), .A2(n8919), .ZN(n6933) );
  NAND2_X1 U8538 ( .A1(n6962), .A2(n6933), .ZN(n7168) );
  OR2_X1 U8539 ( .A1(n6634), .A2(n7168), .ZN(n6936) );
  INV_X1 U8540 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6934) );
  OR2_X1 U8541 ( .A1(n8121), .A2(n6934), .ZN(n6935) );
  INV_X1 U8542 ( .A(n7260), .ZN(n8906) );
  NAND2_X1 U8543 ( .A1(n8906), .A2(n8875), .ZN(n6940) );
  OAI211_X1 U8544 ( .C1(n6994), .C2(n8873), .A(n6940), .B(n6939), .ZN(n6941)
         );
  AOI21_X1 U8545 ( .B1(n6942), .B2(n8871), .A(n6941), .ZN(n6943) );
  OAI211_X1 U8546 ( .C1(n10253), .C2(n8893), .A(n6944), .B(n6943), .ZN(
        P2_U3241) );
  OAI21_X1 U8547 ( .B1(n6947), .B2(n6946), .A(n6945), .ZN(n6948) );
  NAND2_X1 U8548 ( .A1(n6948), .A2(n9428), .ZN(n6952) );
  AND2_X1 U8549 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10003) );
  INV_X1 U8550 ( .A(n6949), .ZN(n7042) );
  OAI22_X1 U8551 ( .A1(n7037), .A2(n9464), .B1(n9453), .B2(n7042), .ZN(n6950)
         );
  AOI211_X1 U8552 ( .C1(n9476), .C2(n9490), .A(n10003), .B(n6950), .ZN(n6951)
         );
  OAI211_X1 U8553 ( .C1(n10125), .C2(n9372), .A(n6952), .B(n6951), .ZN(
        P1_U3211) );
  OR2_X1 U8554 ( .A1(n7260), .A2(n6602), .ZN(n7053) );
  AOI22_X1 U8555 ( .A1(n7974), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7973), .B2(
        n6956), .ZN(n6960) );
  INV_X2 U8556 ( .A(n6957), .ZN(n8153) );
  NAND2_X1 U8557 ( .A1(n6958), .A2(n8153), .ZN(n6959) );
  NAND2_X1 U8558 ( .A1(n6960), .A2(n6959), .ZN(n7241) );
  XNOR2_X1 U8559 ( .A(n7241), .B(n8094), .ZN(n7054) );
  XNOR2_X1 U8560 ( .A(n7053), .B(n7054), .ZN(n7051) );
  XNOR2_X1 U8561 ( .A(n7050), .B(n7051), .ZN(n6973) );
  OAI22_X1 U8562 ( .A1(n8885), .A2(n7168), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8919), .ZN(n6971) );
  NAND2_X1 U8563 ( .A1(n8046), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6968) );
  OR2_X1 U8564 ( .A1(n8083), .A2(n7265), .ZN(n6967) );
  NAND2_X1 U8565 ( .A1(n6962), .A2(n6961), .ZN(n6963) );
  NAND2_X1 U8566 ( .A1(n7064), .A2(n6963), .ZN(n7264) );
  OR2_X1 U8567 ( .A1(n6634), .A2(n7264), .ZN(n6966) );
  INV_X1 U8568 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6964) );
  OR2_X1 U8569 ( .A1(n8121), .A2(n6964), .ZN(n6965) );
  NAND4_X1 U8570 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n8905)
         );
  AOI22_X1 U8571 ( .A1(n8907), .A2(n9195), .B1(n9197), .B2(n8905), .ZN(n7163)
         );
  NOR2_X1 U8572 ( .A1(n7163), .A2(n6969), .ZN(n6970) );
  AOI211_X1 U8573 ( .C1(n7241), .C2(n8848), .A(n6971), .B(n6970), .ZN(n6972)
         );
  OAI21_X1 U8574 ( .B1(n6973), .B2(n8866), .A(n6972), .ZN(P2_U3215) );
  XNOR2_X1 U8575 ( .A(n6974), .B(n6986), .ZN(n6975) );
  AOI222_X1 U8576 ( .A1(n9494), .A2(n9735), .B1(n9492), .B2(n9737), .C1(n10061), .C2(n6975), .ZN(n10119) );
  OAI22_X1 U8577 ( .A1(n10075), .A2(n8450), .B1(n6976), .B2(n7922), .ZN(n6984)
         );
  OR2_X1 U8578 ( .A1(n6978), .A2(n6977), .ZN(n10132) );
  INV_X1 U8579 ( .A(n10132), .ZN(n10140) );
  OAI211_X1 U8580 ( .C1(n6981), .C2(n6980), .A(n6979), .B(n10140), .ZN(n10117)
         );
  NOR2_X1 U8581 ( .A1(n10078), .A2(n10054), .ZN(n9697) );
  INV_X1 U8582 ( .A(n9697), .ZN(n6982) );
  NOR2_X1 U8583 ( .A1(n10117), .A2(n6982), .ZN(n6983) );
  AOI211_X1 U8584 ( .C1(n7711), .C2(n6985), .A(n6984), .B(n6983), .ZN(n6989)
         );
  NAND2_X1 U8585 ( .A1(n6987), .A2(n6986), .ZN(n10114) );
  NAND3_X1 U8586 ( .A1(n10115), .A2(n10114), .A3(n7311), .ZN(n6988) );
  OAI211_X1 U8587 ( .C1(n10119), .C2(n10078), .A(n6989), .B(n6988), .ZN(
        P1_U3286) );
  INV_X1 U8588 ( .A(n7972), .ZN(n6992) );
  OAI222_X1 U8589 ( .A1(n9330), .A2(n6990), .B1(n4490), .B2(n6992), .C1(
        P2_U3152), .C2(n8976), .ZN(P2_U3339) );
  OAI222_X1 U8590 ( .A1(n8383), .A2(n6993), .B1(n9881), .B2(n6992), .C1(
        P1_U3084), .C2(n6991), .ZN(P1_U3334) );
  NAND2_X1 U8591 ( .A1(n6994), .A2(n7156), .ZN(n8217) );
  NAND2_X1 U8592 ( .A1(n8217), .A2(n8242), .ZN(n8179) );
  NAND2_X1 U8593 ( .A1(n6995), .A2(n7278), .ZN(n8233) );
  NAND2_X1 U8594 ( .A1(n7006), .A2(n8233), .ZN(n7273) );
  NAND2_X1 U8595 ( .A1(n7273), .A2(n7277), .ZN(n6997) );
  NAND2_X1 U8596 ( .A1(n6995), .A2(n10228), .ZN(n6996) );
  NAND2_X1 U8597 ( .A1(n6997), .A2(n6996), .ZN(n7180) );
  NAND2_X1 U8598 ( .A1(n6998), .A2(n7191), .ZN(n8234) );
  NAND2_X1 U8599 ( .A1(n7180), .A2(n8177), .ZN(n7000) );
  NAND2_X1 U8600 ( .A1(n6998), .A2(n4489), .ZN(n6999) );
  NAND2_X1 U8601 ( .A1(n7000), .A2(n6999), .ZN(n7145) );
  XNOR2_X1 U8602 ( .A(n8910), .B(n8238), .ZN(n8180) );
  NAND2_X1 U8603 ( .A1(n7145), .A2(n8180), .ZN(n7002) );
  NAND2_X1 U8604 ( .A1(n7007), .A2(n8238), .ZN(n7001) );
  NAND2_X1 U8605 ( .A1(n7002), .A2(n7001), .ZN(n10203) );
  NAND2_X1 U8606 ( .A1(n7003), .A2(n10206), .ZN(n8216) );
  NAND2_X1 U8607 ( .A1(n8216), .A2(n8240), .ZN(n10204) );
  NAND2_X1 U8608 ( .A1(n10203), .A2(n10204), .ZN(n7005) );
  NAND2_X1 U8609 ( .A1(n7003), .A2(n10249), .ZN(n7004) );
  XOR2_X1 U8610 ( .A(n8179), .B(n7159), .Z(n7179) );
  NAND2_X1 U8611 ( .A1(n7274), .A2(n8233), .ZN(n8222) );
  NAND2_X1 U8612 ( .A1(n8222), .A2(n7006), .ZN(n7181) );
  INV_X1 U8613 ( .A(n8180), .ZN(n8225) );
  NAND2_X1 U8614 ( .A1(n7007), .A2(n10241), .ZN(n8215) );
  NAND2_X1 U8615 ( .A1(n7008), .A2(n8215), .ZN(n10192) );
  INV_X1 U8616 ( .A(n8216), .ZN(n7009) );
  XNOR2_X1 U8617 ( .A(n7162), .B(n8179), .ZN(n7010) );
  AOI222_X1 U8618 ( .A1(n10194), .A2(n7010), .B1(n8907), .B2(n9197), .C1(n8909), .C2(n9195), .ZN(n7172) );
  NAND2_X1 U8619 ( .A1(n10228), .A2(n7363), .ZN(n7280) );
  INV_X1 U8620 ( .A(n10197), .ZN(n10261) );
  INV_X1 U8621 ( .A(n7351), .ZN(n7012) );
  AOI211_X1 U8622 ( .C1(n7156), .C2(n10196), .A(n10261), .B(n7012), .ZN(n7176)
         );
  AOI21_X1 U8623 ( .B1(n6570), .B2(n7156), .A(n7176), .ZN(n7013) );
  OAI211_X1 U8624 ( .C1(n9297), .C2(n7179), .A(n7172), .B(n7013), .ZN(n7015)
         );
  NAND2_X1 U8625 ( .A1(n7015), .A2(n10295), .ZN(n7014) );
  OAI21_X1 U8626 ( .B1(n10295), .B2(n6456), .A(n7014), .ZN(P2_U3525) );
  NAND2_X1 U8627 ( .A1(n7015), .A2(n9320), .ZN(n7016) );
  OAI21_X1 U8628 ( .B1(n9320), .B2(n6755), .A(n7016), .ZN(P2_U3466) );
  INV_X1 U8629 ( .A(n7317), .ZN(n7195) );
  NAND2_X1 U8630 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7328) );
  INV_X1 U8631 ( .A(n7328), .ZN(n7021) );
  AOI21_X1 U8632 ( .B1(n7214), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7017), .ZN(
        n7019) );
  INV_X1 U8633 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7228) );
  MUX2_X1 U8634 ( .A(n7228), .B(P2_REG1_REG_10__SCAN_IN), .S(n7317), .Z(n7018)
         );
  NOR2_X1 U8635 ( .A1(n7019), .A2(n7018), .ZN(n7198) );
  AOI211_X1 U8636 ( .C1(n7019), .C2(n7018), .A(n7198), .B(n10171), .ZN(n7020)
         );
  AOI211_X1 U8637 ( .C1(n10187), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7021), .B(
        n7020), .ZN(n7027) );
  OAI21_X1 U8638 ( .B1(n7023), .B2(n7400), .A(n7022), .ZN(n7025) );
  INV_X1 U8639 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7448) );
  MUX2_X1 U8640 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7448), .S(n7317), .Z(n7024)
         );
  NAND2_X1 U8641 ( .A1(n7024), .A2(n7025), .ZN(n7194) );
  OAI211_X1 U8642 ( .C1(n7025), .C2(n7024), .A(n10185), .B(n7194), .ZN(n7026)
         );
  OAI211_X1 U8643 ( .C1(n10170), .C2(n7195), .A(n7027), .B(n7026), .ZN(
        P2_U3255) );
  NAND2_X1 U8644 ( .A1(n7037), .A2(n4781), .ZN(n7028) );
  XNOR2_X1 U8645 ( .A(n7084), .B(n7083), .ZN(n10128) );
  INV_X1 U8646 ( .A(n10128), .ZN(n7049) );
  INV_X1 U8647 ( .A(n7079), .ZN(n7033) );
  AOI21_X1 U8648 ( .B1(n7083), .B2(n7034), .A(n7033), .ZN(n7035) );
  OAI222_X1 U8649 ( .A1(n10058), .A2(n7038), .B1(n10056), .B2(n7037), .C1(
        n7036), .C2(n7035), .ZN(n10126) );
  AOI21_X1 U8650 ( .B1(n7039), .B2(n7045), .A(n10132), .ZN(n7040) );
  NAND2_X1 U8651 ( .A1(n7040), .A2(n7091), .ZN(n10124) );
  OR2_X1 U8652 ( .A1(n7041), .A2(n10054), .ZN(n9744) );
  OAI22_X1 U8653 ( .A1(n10075), .A2(n7043), .B1(n7042), .B2(n7922), .ZN(n7044)
         );
  AOI21_X1 U8654 ( .B1(n7711), .B2(n7045), .A(n7044), .ZN(n7046) );
  OAI21_X1 U8655 ( .B1(n10124), .B2(n9744), .A(n7046), .ZN(n7047) );
  AOI21_X1 U8656 ( .B1(n10126), .B2(n10075), .A(n7047), .ZN(n7048) );
  OAI21_X1 U8657 ( .B1(n9750), .B2(n7049), .A(n7048), .ZN(P1_U3284) );
  INV_X1 U8658 ( .A(n7051), .ZN(n7052) );
  INV_X1 U8659 ( .A(n7053), .ZN(n7056) );
  INV_X1 U8660 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U8661 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U8662 ( .A1(n7059), .A2(n8153), .ZN(n7062) );
  AOI22_X1 U8663 ( .A1(n7974), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7973), .B2(
        n7060), .ZN(n7061) );
  XNOR2_X1 U8664 ( .A(n10260), .B(n8094), .ZN(n7210) );
  NAND2_X1 U8665 ( .A1(n8905), .A2(n8176), .ZN(n7208) );
  XNOR2_X1 U8666 ( .A(n7210), .B(n7208), .ZN(n7206) );
  XNOR2_X1 U8667 ( .A(n7207), .B(n7206), .ZN(n7077) );
  INV_X1 U8668 ( .A(n7264), .ZN(n7075) );
  NOR2_X1 U8669 ( .A1(n8893), .A2(n10260), .ZN(n7074) );
  NAND2_X1 U8670 ( .A1(n8046), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7070) );
  OR2_X1 U8671 ( .A1(n8083), .A2(n7400), .ZN(n7069) );
  NAND2_X1 U8672 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8673 ( .A1(n7226), .A2(n7065), .ZN(n7399) );
  OR2_X1 U8674 ( .A1(n6634), .A2(n7399), .ZN(n7068) );
  INV_X1 U8675 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7066) );
  OR2_X1 U8676 ( .A1(n8121), .A2(n7066), .ZN(n7067) );
  INV_X1 U8677 ( .A(n7443), .ZN(n8904) );
  NAND2_X1 U8678 ( .A1(n8904), .A2(n8875), .ZN(n7072) );
  OAI211_X1 U8679 ( .C1(n7260), .C2(n8873), .A(n7072), .B(n7071), .ZN(n7073)
         );
  AOI211_X1 U8680 ( .C1(n8871), .C2(n7075), .A(n7074), .B(n7073), .ZN(n7076)
         );
  OAI21_X1 U8681 ( .B1(n7077), .B2(n8866), .A(n7076), .ZN(P2_U3223) );
  XNOR2_X1 U8682 ( .A(n7287), .B(n7090), .ZN(n7080) );
  NAND2_X1 U8683 ( .A1(n7080), .A2(n10061), .ZN(n7082) );
  AOI22_X1 U8684 ( .A1(n9735), .A2(n9491), .B1(n9489), .B2(n9737), .ZN(n7081)
         );
  NAND2_X1 U8685 ( .A1(n7082), .A2(n7081), .ZN(n10134) );
  INV_X1 U8686 ( .A(n10134), .ZN(n7100) );
  NAND2_X1 U8687 ( .A1(n7085), .A2(n10125), .ZN(n7086) );
  INV_X1 U8688 ( .A(n7297), .ZN(n7089) );
  AOI21_X1 U8689 ( .B1(n7090), .B2(n7087), .A(n7089), .ZN(n10137) );
  INV_X1 U8690 ( .A(n7091), .ZN(n7092) );
  NOR2_X1 U8691 ( .A1(n7091), .A2(n7295), .ZN(n7303) );
  INV_X1 U8692 ( .A(n7303), .ZN(n7459) );
  OAI21_X1 U8693 ( .B1(n10131), .B2(n7092), .A(n7459), .ZN(n10133) );
  INV_X1 U8694 ( .A(n7093), .ZN(n7120) );
  OAI22_X1 U8695 ( .A1(n10075), .A2(n7094), .B1(n7120), .B2(n7922), .ZN(n7095)
         );
  AOI21_X1 U8696 ( .B1(n7711), .B2(n7295), .A(n7095), .ZN(n7096) );
  OAI21_X1 U8697 ( .B1(n10133), .B2(n7097), .A(n7096), .ZN(n7098) );
  AOI21_X1 U8698 ( .B1(n10137), .B2(n7311), .A(n7098), .ZN(n7099) );
  OAI21_X1 U8699 ( .B1(n10078), .B2(n7100), .A(n7099), .ZN(P1_U3283) );
  INV_X1 U8700 ( .A(n7992), .ZN(n8363) );
  OAI222_X1 U8701 ( .A1(n9881), .A2(n8363), .B1(n7102), .B2(P1_U3084), .C1(
        n7101), .C2(n8383), .ZN(P1_U3333) );
  OAI21_X1 U8702 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(n7113) );
  NAND2_X1 U8703 ( .A1(n9999), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U8704 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7489) );
  OAI211_X1 U8705 ( .C1(n7107), .C2(n9971), .A(n7106), .B(n7489), .ZN(n7112)
         );
  AOI211_X1 U8706 ( .C1(n7110), .C2(n7109), .A(n7108), .B(n10032), .ZN(n7111)
         );
  AOI211_X1 U8707 ( .C1(n10043), .C2(n7113), .A(n7112), .B(n7111), .ZN(n7114)
         );
  INV_X1 U8708 ( .A(n7114), .ZN(P1_U3253) );
  NAND2_X1 U8709 ( .A1(n7116), .A2(n7115), .ZN(n7118) );
  XNOR2_X1 U8710 ( .A(n7118), .B(n7117), .ZN(n7119) );
  NAND2_X1 U8711 ( .A1(n7119), .A2(n9428), .ZN(n7124) );
  INV_X1 U8712 ( .A(n9464), .ZN(n9474) );
  OAI22_X1 U8713 ( .A1(n7376), .A2(n9451), .B1(n9453), .B2(n7120), .ZN(n7121)
         );
  AOI211_X1 U8714 ( .C1(n9474), .C2(n9491), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OAI211_X1 U8715 ( .C1(n10131), .C2(n9372), .A(n7124), .B(n7123), .ZN(
        P1_U3219) );
  INV_X1 U8716 ( .A(n8005), .ZN(n7137) );
  OAI222_X1 U8717 ( .A1(n9881), .A2(n7137), .B1(n7126), .B2(P1_U3084), .C1(
        n7125), .C2(n8383), .ZN(P1_U3332) );
  INV_X1 U8718 ( .A(n7128), .ZN(n7129) );
  AOI21_X1 U8719 ( .B1(n7130), .B2(n7127), .A(n7129), .ZN(n7136) );
  INV_X1 U8720 ( .A(n7460), .ZN(n7131) );
  OAI22_X1 U8721 ( .A1(n7409), .A2(n9451), .B1(n9453), .B2(n7131), .ZN(n7132)
         );
  AOI211_X1 U8722 ( .C1(n9474), .C2(n9490), .A(n7133), .B(n7132), .ZN(n7135)
         );
  NAND2_X1 U8723 ( .A1(n9477), .A2(n10138), .ZN(n7134) );
  OAI211_X1 U8724 ( .C1(n7136), .C2(n9470), .A(n7135), .B(n7134), .ZN(P1_U3229) );
  OAI222_X1 U8725 ( .A1(n9330), .A2(n8006), .B1(n4490), .B2(n7137), .C1(n8349), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8726 ( .A(n7138), .ZN(n7139) );
  OR2_X1 U8727 ( .A1(n7140), .A2(n7139), .ZN(n7141) );
  OR2_X1 U8728 ( .A1(n8976), .A2(n8349), .ZN(n8203) );
  INV_X1 U8729 ( .A(n8203), .ZN(n7143) );
  NAND2_X1 U8730 ( .A1(n7754), .A2(n7254), .ZN(n7144) );
  NAND2_X1 U8731 ( .A1(n9190), .A2(n7144), .ZN(n9214) );
  XNOR2_X1 U8732 ( .A(n7145), .B(n8225), .ZN(n10243) );
  XNOR2_X1 U8733 ( .A(n7146), .B(n8180), .ZN(n7148) );
  INV_X1 U8734 ( .A(n10194), .ZN(n9180) );
  OAI21_X1 U8735 ( .B1(n7148), .B2(n9180), .A(n7147), .ZN(n10239) );
  INV_X1 U8736 ( .A(n10239), .ZN(n7149) );
  INV_X2 U8737 ( .A(n10210), .ZN(n9190) );
  MUX2_X1 U8738 ( .A(n7150), .B(n7149), .S(n9190), .Z(n7155) );
  AOI211_X1 U8739 ( .C1(n10241), .C2(n7188), .A(n10261), .B(n10198), .ZN(
        n10240) );
  NOR2_X1 U8740 ( .A1(n7268), .A2(n9188), .ZN(n9172) );
  INV_X1 U8741 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U8742 ( .A1(n9190), .A2(n7152), .ZN(n9164) );
  OAI22_X1 U8743 ( .A1(n9164), .A2(n8238), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10199), .ZN(n7153) );
  AOI21_X1 U8744 ( .B1(n10240), .B2(n9172), .A(n7153), .ZN(n7154) );
  OAI211_X1 U8745 ( .C1(n9214), .C2(n10243), .A(n7155), .B(n7154), .ZN(
        P2_U3293) );
  NOR2_X1 U8746 ( .A1(n8908), .A2(n7156), .ZN(n7158) );
  OR2_X1 U8747 ( .A1(n8179), .A2(n7174), .ZN(n7157) );
  NAND2_X1 U8748 ( .A1(n8907), .A2(n8229), .ZN(n7160) );
  NAND2_X1 U8749 ( .A1(n7260), .A2(n7241), .ZN(n8248) );
  NAND2_X1 U8750 ( .A1(n8906), .A2(n7251), .ZN(n8258) );
  XOR2_X1 U8751 ( .A(n7248), .B(n8246), .Z(n7243) );
  INV_X1 U8752 ( .A(n8242), .ZN(n7161) );
  XNOR2_X1 U8753 ( .A(n8907), .B(n8229), .ZN(n8182) );
  NAND2_X1 U8754 ( .A1(n8230), .A2(n8229), .ZN(n8247) );
  XOR2_X1 U8755 ( .A(n7256), .B(n8246), .Z(n7164) );
  OAI21_X1 U8756 ( .B1(n7164), .B2(n9180), .A(n7163), .ZN(n7239) );
  INV_X1 U8757 ( .A(n7239), .ZN(n7165) );
  MUX2_X1 U8758 ( .A(n7166), .B(n7165), .S(n9190), .Z(n7171) );
  INV_X1 U8759 ( .A(n7352), .ZN(n7167) );
  AOI211_X1 U8760 ( .C1(n7241), .C2(n7167), .A(n10261), .B(n7266), .ZN(n7240)
         );
  OAI22_X1 U8761 ( .A1(n9164), .A2(n7251), .B1(n10199), .B2(n7168), .ZN(n7169)
         );
  AOI21_X1 U8762 ( .B1(n7240), .B2(n9172), .A(n7169), .ZN(n7170) );
  OAI211_X1 U8763 ( .C1(n9214), .C2(n7243), .A(n7171), .B(n7170), .ZN(P2_U3289) );
  MUX2_X1 U8764 ( .A(n6464), .B(n7172), .S(n9190), .Z(n7178) );
  OAI22_X1 U8765 ( .A1(n9164), .A2(n7174), .B1(n7173), .B2(n10199), .ZN(n7175)
         );
  AOI21_X1 U8766 ( .B1(n7176), .B2(n9172), .A(n7175), .ZN(n7177) );
  OAI211_X1 U8767 ( .C1(n7179), .C2(n9214), .A(n7178), .B(n7177), .ZN(P2_U3291) );
  XOR2_X1 U8768 ( .A(n7180), .B(n8177), .Z(n10233) );
  INV_X1 U8769 ( .A(n7181), .ZN(n7184) );
  INV_X1 U8770 ( .A(n8177), .ZN(n7183) );
  OAI21_X1 U8771 ( .B1(n7184), .B2(n7183), .A(n7182), .ZN(n7186) );
  AOI21_X1 U8772 ( .B1(n7186), .B2(n10194), .A(n7185), .ZN(n10235) );
  MUX2_X1 U8773 ( .A(n10235), .B(n7187), .S(n10210), .Z(n7193) );
  OAI211_X1 U8774 ( .C1(n4731), .C2(n4489), .A(n10197), .B(n7188), .ZN(n10234)
         );
  INV_X1 U8775 ( .A(n9172), .ZN(n10201) );
  OAI22_X1 U8776 ( .A1(n10234), .A2(n10201), .B1(n7189), .B2(n10199), .ZN(
        n7190) );
  AOI21_X1 U8777 ( .B1(n10205), .B2(n7191), .A(n7190), .ZN(n7192) );
  OAI211_X1 U8778 ( .C1(n10233), .C2(n9214), .A(n7193), .B(n7192), .ZN(
        P2_U3294) );
  INV_X1 U8779 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7321) );
  MUX2_X1 U8780 ( .A(n7321), .B(P2_REG2_REG_11__SCAN_IN), .S(n7475), .Z(n7197)
         );
  OAI21_X1 U8781 ( .B1(n7195), .B2(n7448), .A(n7194), .ZN(n7196) );
  NOR2_X1 U8782 ( .A1(n7196), .A2(n7197), .ZN(n7470) );
  AOI21_X1 U8783 ( .B1(n7197), .B2(n7196), .A(n7470), .ZN(n7205) );
  INV_X1 U8784 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8581) );
  NOR2_X1 U8785 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8581), .ZN(n7202) );
  INV_X1 U8786 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7320) );
  MUX2_X1 U8787 ( .A(n7320), .B(P2_REG1_REG_11__SCAN_IN), .S(n7475), .Z(n7199)
         );
  AOI211_X1 U8788 ( .C1(n7200), .C2(n7199), .A(n7474), .B(n10171), .ZN(n7201)
         );
  AOI211_X1 U8789 ( .C1(n10187), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7202), .B(
        n7201), .ZN(n7204) );
  INV_X1 U8790 ( .A(n10170), .ZN(n10183) );
  NAND2_X1 U8791 ( .A1(n10183), .A2(n7475), .ZN(n7203) );
  OAI211_X1 U8792 ( .C1(n7205), .C2(n10172), .A(n7204), .B(n7203), .ZN(
        P2_U3256) );
  INV_X1 U8793 ( .A(n7208), .ZN(n7209) );
  NAND2_X1 U8794 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  NAND2_X1 U8795 ( .A1(n7213), .A2(n8153), .ZN(n7216) );
  AOI22_X1 U8796 ( .A1(n7974), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7973), .B2(
        n7214), .ZN(n7215) );
  XNOR2_X1 U8797 ( .A(n7527), .B(n8094), .ZN(n7217) );
  OR2_X1 U8798 ( .A1(n7443), .A2(n6602), .ZN(n7218) );
  NAND2_X1 U8799 ( .A1(n7217), .A2(n7218), .ZN(n7314) );
  INV_X1 U8800 ( .A(n7217), .ZN(n7220) );
  INV_X1 U8801 ( .A(n7218), .ZN(n7219) );
  NAND2_X1 U8802 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  NAND2_X1 U8803 ( .A1(n7314), .A2(n7221), .ZN(n7223) );
  INV_X1 U8804 ( .A(n7315), .ZN(n7222) );
  AOI21_X1 U8805 ( .B1(n7224), .B2(n7223), .A(n7222), .ZN(n7238) );
  NOR2_X1 U8806 ( .A1(n8885), .A2(n7399), .ZN(n7236) );
  INV_X1 U8807 ( .A(n8905), .ZN(n7392) );
  NAND2_X1 U8808 ( .A1(n8158), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7232) );
  OR2_X1 U8809 ( .A1(n8083), .A2(n7448), .ZN(n7231) );
  NAND2_X1 U8810 ( .A1(n7226), .A2(n7225), .ZN(n7227) );
  NAND2_X1 U8811 ( .A1(n7322), .A2(n7227), .ZN(n7447) );
  OR2_X1 U8812 ( .A1(n6634), .A2(n7447), .ZN(n7230) );
  OR2_X1 U8813 ( .A1(n8162), .A2(n7228), .ZN(n7229) );
  INV_X1 U8814 ( .A(n7433), .ZN(n8903) );
  NAND2_X1 U8815 ( .A1(n8903), .A2(n8875), .ZN(n7234) );
  OAI211_X1 U8816 ( .C1(n7392), .C2(n8873), .A(n7234), .B(n7233), .ZN(n7235)
         );
  AOI211_X1 U8817 ( .C1(n7527), .C2(n8848), .A(n7236), .B(n7235), .ZN(n7237)
         );
  OAI21_X1 U8818 ( .B1(n7238), .B2(n8866), .A(n7237), .ZN(P2_U3233) );
  INV_X1 U8819 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7245) );
  AOI211_X1 U8820 ( .C1(n6570), .C2(n7241), .A(n7240), .B(n7239), .ZN(n7242)
         );
  OAI21_X1 U8821 ( .B1(n9297), .B2(n7243), .A(n7242), .ZN(n7246) );
  NAND2_X1 U8822 ( .A1(n7246), .A2(n10295), .ZN(n7244) );
  OAI21_X1 U8823 ( .B1(n10295), .B2(n7245), .A(n7244), .ZN(P2_U3527) );
  NAND2_X1 U8824 ( .A1(n7246), .A2(n9320), .ZN(n7247) );
  OAI21_X1 U8825 ( .B1(n9320), .B2(n6934), .A(n7247), .ZN(P2_U3472) );
  INV_X1 U8826 ( .A(n7248), .ZN(n7250) );
  INV_X1 U8827 ( .A(n8246), .ZN(n7249) );
  NAND2_X1 U8828 ( .A1(n7260), .A2(n7251), .ZN(n7252) );
  INV_X1 U8829 ( .A(n10260), .ZN(n7387) );
  NAND2_X1 U8830 ( .A1(n7392), .A2(n7387), .ZN(n8212) );
  NAND2_X1 U8831 ( .A1(n10260), .A2(n8905), .ZN(n8249) );
  OR2_X1 U8832 ( .A1(n7436), .A2(n8259), .ZN(n7389) );
  NAND2_X1 U8833 ( .A1(n7436), .A2(n8259), .ZN(n7253) );
  NAND2_X1 U8834 ( .A1(n7389), .A2(n7253), .ZN(n10259) );
  OR2_X1 U8835 ( .A1(n10210), .A2(n7254), .ZN(n7763) );
  INV_X1 U8836 ( .A(n8248), .ZN(n7255) );
  INV_X1 U8837 ( .A(n7258), .ZN(n7259) );
  INV_X1 U8838 ( .A(n8259), .ZN(n7257) );
  OAI21_X1 U8839 ( .B1(n7259), .B2(n8259), .A(n4562), .ZN(n7262) );
  OAI22_X1 U8840 ( .A1(n7260), .A2(n9182), .B1(n7443), .B2(n9184), .ZN(n7261)
         );
  AOI21_X1 U8841 ( .B1(n7262), .B2(n10194), .A(n7261), .ZN(n7263) );
  OAI21_X1 U8842 ( .B1(n7754), .B2(n10259), .A(n7263), .ZN(n10263) );
  NAND2_X1 U8843 ( .A1(n10263), .A2(n9190), .ZN(n7272) );
  OAI22_X1 U8844 ( .A1(n9190), .A2(n7265), .B1(n7264), .B2(n10199), .ZN(n7270)
         );
  NAND2_X1 U8845 ( .A1(n7266), .A2(n10260), .ZN(n7396) );
  OR2_X1 U8846 ( .A1(n7266), .A2(n10260), .ZN(n7267) );
  NAND2_X1 U8847 ( .A1(n7396), .A2(n7267), .ZN(n10262) );
  NOR2_X1 U8848 ( .A1(n7268), .A2(n8176), .ZN(n9211) );
  INV_X1 U8849 ( .A(n9211), .ZN(n8991) );
  NOR2_X1 U8850 ( .A1(n10262), .A2(n8991), .ZN(n7269) );
  AOI211_X1 U8851 ( .C1(n10205), .C2(n7387), .A(n7270), .B(n7269), .ZN(n7271)
         );
  OAI211_X1 U8852 ( .C1(n10259), .C2(n7763), .A(n7272), .B(n7271), .ZN(
        P2_U3288) );
  XNOR2_X1 U8853 ( .A(n7273), .B(n7274), .ZN(n7276) );
  AOI21_X1 U8854 ( .B1(n7276), .B2(n10194), .A(n7275), .ZN(n10229) );
  INV_X1 U8855 ( .A(n9214), .ZN(n10207) );
  XNOR2_X1 U8856 ( .A(n7273), .B(n7277), .ZN(n10232) );
  AOI21_X1 U8857 ( .B1(n7279), .B2(n7278), .A(n10261), .ZN(n7281) );
  AND2_X1 U8858 ( .A1(n7281), .A2(n7280), .ZN(n10226) );
  NOR2_X1 U8859 ( .A1(n10199), .A2(n6557), .ZN(n7283) );
  NOR2_X1 U8860 ( .A1(n9190), .A2(n8370), .ZN(n7282) );
  AOI211_X1 U8861 ( .C1(n10226), .C2(n9172), .A(n7283), .B(n7282), .ZN(n7284)
         );
  OAI21_X1 U8862 ( .B1(n10228), .B2(n9164), .A(n7284), .ZN(n7285) );
  AOI21_X1 U8863 ( .B1(n10207), .B2(n10232), .A(n7285), .ZN(n7286) );
  OAI21_X1 U8864 ( .B1(n10210), .B2(n10229), .A(n7286), .ZN(P2_U3295) );
  INV_X1 U8865 ( .A(n7500), .ZN(n7290) );
  OAI21_X1 U8866 ( .B1(n7290), .B2(n7289), .A(n7455), .ZN(n7293) );
  XNOR2_X1 U8867 ( .A(n7293), .B(n7301), .ZN(n7294) );
  AOI222_X1 U8868 ( .A1(n9489), .A2(n9735), .B1(n9487), .B2(n9737), .C1(n10061), .C2(n7294), .ZN(n9886) );
  NAND2_X1 U8869 ( .A1(n7295), .A2(n9490), .ZN(n7296) );
  NAND2_X1 U8870 ( .A1(n7297), .A2(n7296), .ZN(n7457) );
  OR2_X1 U8871 ( .A1(n10138), .A2(n9489), .ZN(n7298) );
  NAND2_X1 U8872 ( .A1(n7457), .A2(n7298), .ZN(n7300) );
  NAND2_X1 U8873 ( .A1(n10138), .A2(n9489), .ZN(n7299) );
  INV_X1 U8874 ( .A(n7301), .ZN(n7302) );
  OAI21_X1 U8875 ( .B1(n4505), .B2(n7302), .A(n4929), .ZN(n9888) );
  INV_X1 U8876 ( .A(n10138), .ZN(n7462) );
  NAND2_X1 U8877 ( .A1(n7303), .A2(n7462), .ZN(n7304) );
  INV_X1 U8878 ( .A(n7304), .ZN(n7458) );
  INV_X1 U8879 ( .A(n7495), .ZN(n7305) );
  OR2_X2 U8880 ( .A1(n7304), .A2(n7495), .ZN(n7504) );
  OAI211_X1 U8881 ( .C1(n7458), .C2(n7305), .A(n10140), .B(n7504), .ZN(n9884)
         );
  INV_X1 U8882 ( .A(n7306), .ZN(n7373) );
  OAI22_X1 U8883 ( .A1(n10075), .A2(n7307), .B1(n7373), .B2(n7922), .ZN(n7308)
         );
  AOI21_X1 U8884 ( .B1(n7495), .B2(n7711), .A(n7308), .ZN(n7309) );
  OAI21_X1 U8885 ( .B1(n9884), .B2(n9744), .A(n7309), .ZN(n7310) );
  AOI21_X1 U8886 ( .B1(n9888), .B2(n7311), .A(n7310), .ZN(n7312) );
  OAI21_X1 U8887 ( .B1(n9886), .B2(n10078), .A(n7312), .ZN(P1_U3281) );
  INV_X1 U8888 ( .A(n8020), .ZN(n8378) );
  OAI222_X1 U8889 ( .A1(n9330), .A2(n8021), .B1(n4490), .B2(n8378), .C1(
        P2_U3152), .C2(n7313), .ZN(P2_U3336) );
  NAND2_X1 U8890 ( .A1(n7316), .A2(n8153), .ZN(n7319) );
  AOI22_X1 U8891 ( .A1(n7974), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7973), .B2(
        n7317), .ZN(n7318) );
  XNOR2_X1 U8892 ( .A(n7663), .B(n8116), .ZN(n7414) );
  NOR2_X1 U8893 ( .A1(n7433), .A2(n6602), .ZN(n7413) );
  XNOR2_X1 U8894 ( .A(n7414), .B(n7413), .ZN(n7416) );
  XNOR2_X1 U8895 ( .A(n7417), .B(n7416), .ZN(n7333) );
  INV_X1 U8896 ( .A(n8873), .ZN(n8890) );
  INV_X1 U8897 ( .A(n8875), .ZN(n8887) );
  NAND2_X1 U8898 ( .A1(n8158), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7327) );
  OR2_X1 U8899 ( .A1(n8162), .A2(n7320), .ZN(n7326) );
  OR2_X1 U8900 ( .A1(n8083), .A2(n7321), .ZN(n7325) );
  NAND2_X1 U8901 ( .A1(n7322), .A2(n8581), .ZN(n7323) );
  NAND2_X1 U8902 ( .A1(n7422), .A2(n7323), .ZN(n7732) );
  OR2_X1 U8903 ( .A1(n6634), .A2(n7732), .ZN(n7324) );
  OAI21_X1 U8904 ( .B1(n8887), .B2(n7683), .A(n7328), .ZN(n7329) );
  AOI21_X1 U8905 ( .B1(n8890), .B2(n8904), .A(n7329), .ZN(n7330) );
  OAI21_X1 U8906 ( .B1(n7447), .B2(n8885), .A(n7330), .ZN(n7331) );
  AOI21_X1 U8907 ( .B1(n7663), .B2(n8848), .A(n7331), .ZN(n7332) );
  OAI21_X1 U8908 ( .B1(n7333), .B2(n8866), .A(n7332), .ZN(P2_U3219) );
  INV_X1 U8909 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7345) );
  OAI21_X1 U8910 ( .B1(n7336), .B2(n7335), .A(n7334), .ZN(n7337) );
  NAND2_X1 U8911 ( .A1(n7337), .A2(n10043), .ZN(n7344) );
  AND2_X1 U8912 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7660) );
  AOI211_X1 U8913 ( .C1(n7340), .C2(n7339), .A(n7338), .B(n10032), .ZN(n7341)
         );
  AOI211_X1 U8914 ( .C1(n7342), .C2(n10038), .A(n7660), .B(n7341), .ZN(n7343)
         );
  OAI211_X1 U8915 ( .C1(n10046), .C2(n7345), .A(n7344), .B(n7343), .ZN(
        P1_U3254) );
  XNOR2_X1 U8916 ( .A(n7346), .B(n8182), .ZN(n7347) );
  NAND2_X1 U8917 ( .A1(n7347), .A2(n10194), .ZN(n7349) );
  AOI22_X1 U8918 ( .A1(n8906), .A2(n9197), .B1(n9195), .B2(n8908), .ZN(n7348)
         );
  NAND2_X1 U8919 ( .A1(n7349), .A2(n7348), .ZN(n10257) );
  INV_X1 U8920 ( .A(n10257), .ZN(n7360) );
  XNOR2_X1 U8921 ( .A(n7350), .B(n8182), .ZN(n10252) );
  AND2_X1 U8922 ( .A1(n7351), .A2(n8229), .ZN(n7353) );
  OR2_X1 U8923 ( .A1(n7353), .A2(n7352), .ZN(n10254) );
  OAI22_X1 U8924 ( .A1(n7355), .A2(n10199), .B1(n7354), .B2(n9190), .ZN(n7356)
         );
  AOI21_X1 U8925 ( .B1(n10205), .B2(n8229), .A(n7356), .ZN(n7357) );
  OAI21_X1 U8926 ( .B1(n10254), .B2(n8991), .A(n7357), .ZN(n7358) );
  AOI21_X1 U8927 ( .B1(n10252), .B2(n10207), .A(n7358), .ZN(n7359) );
  OAI21_X1 U8928 ( .B1(n7360), .B2(n10210), .A(n7359), .ZN(P2_U3290) );
  OAI21_X1 U8929 ( .B1(n7362), .B2(n10199), .A(n7361), .ZN(n7366) );
  AOI21_X1 U8930 ( .B1(n8991), .B2(n9164), .A(n7363), .ZN(n7365) );
  OAI22_X1 U8931 ( .A1(n4969), .A2(n9214), .B1(n6509), .B2(n9190), .ZN(n7364)
         );
  AOI211_X1 U8932 ( .C1(n9190), .C2(n7366), .A(n7365), .B(n7364), .ZN(n7367)
         );
  INV_X1 U8933 ( .A(n7367), .ZN(P2_U3296) );
  NAND2_X1 U8934 ( .A1(n7495), .A2(n10139), .ZN(n9885) );
  NAND2_X1 U8935 ( .A1(n7369), .A2(n7368), .ZN(n7371) );
  XOR2_X1 U8936 ( .A(n7371), .B(n7370), .Z(n7372) );
  NAND2_X1 U8937 ( .A1(n7372), .A2(n9428), .ZN(n7380) );
  OAI22_X1 U8938 ( .A1(n7491), .A2(n9451), .B1(n9453), .B2(n7373), .ZN(n7378)
         );
  INV_X1 U8939 ( .A(n7374), .ZN(n7375) );
  OAI21_X1 U8940 ( .B1(n9464), .B2(n7376), .A(n7375), .ZN(n7377) );
  NOR2_X1 U8941 ( .A1(n7378), .A2(n7377), .ZN(n7379) );
  OAI211_X1 U8942 ( .C1(n7381), .C2(n9885), .A(n7380), .B(n7379), .ZN(P1_U3215) );
  INV_X1 U8943 ( .A(n8035), .ZN(n7384) );
  NAND2_X1 U8944 ( .A1(n9875), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7382) );
  OAI211_X1 U8945 ( .C1(n7384), .C2(n9881), .A(n7383), .B(n7382), .ZN(P1_U3330) );
  NAND2_X1 U8946 ( .A1(n8035), .A2(n7385), .ZN(n7386) );
  OAI211_X1 U8947 ( .C1(n8036), .C2(n9330), .A(n7386), .B(n8360), .ZN(P2_U3335) );
  INV_X1 U8948 ( .A(n7754), .ZN(n10246) );
  NAND2_X1 U8949 ( .A1(n7387), .A2(n8905), .ZN(n7388) );
  AND2_X1 U8950 ( .A1(n7389), .A2(n7388), .ZN(n7391) );
  OR2_X1 U8951 ( .A1(n7527), .A2(n7443), .ZN(n8250) );
  NAND2_X1 U8952 ( .A1(n7527), .A2(n7443), .ZN(n8262) );
  NAND2_X1 U8953 ( .A1(n8250), .A2(n8262), .ZN(n8185) );
  AND2_X1 U8954 ( .A1(n8185), .A2(n7388), .ZN(n7434) );
  NAND2_X1 U8955 ( .A1(n7389), .A2(n7434), .ZN(n7390) );
  OAI21_X1 U8956 ( .B1(n7391), .B2(n8185), .A(n7390), .ZN(n7526) );
  OAI22_X1 U8957 ( .A1(n7392), .A2(n9182), .B1(n7433), .B2(n9184), .ZN(n7395)
         );
  XNOR2_X1 U8958 ( .A(n7442), .B(n8185), .ZN(n7393) );
  NOR2_X1 U8959 ( .A1(n7393), .A2(n9180), .ZN(n7394) );
  AOI211_X1 U8960 ( .C1(n10246), .C2(n7526), .A(n7395), .B(n7394), .ZN(n7530)
         );
  NAND2_X1 U8961 ( .A1(n7396), .A2(n7527), .ZN(n7397) );
  AND2_X1 U8962 ( .A1(n7449), .A2(n7397), .ZN(n7528) );
  INV_X1 U8963 ( .A(n7527), .ZN(n7398) );
  NOR2_X1 U8964 ( .A1(n7398), .A2(n9164), .ZN(n7402) );
  OAI22_X1 U8965 ( .A1(n9190), .A2(n7400), .B1(n7399), .B2(n10199), .ZN(n7401)
         );
  AOI211_X1 U8966 ( .C1(n7528), .C2(n9211), .A(n7402), .B(n7401), .ZN(n7405)
         );
  INV_X1 U8967 ( .A(n7763), .ZN(n7403) );
  NAND2_X1 U8968 ( .A1(n7526), .A2(n7403), .ZN(n7404) );
  OAI211_X1 U8969 ( .C1(n7530), .C2(n10210), .A(n7405), .B(n7404), .ZN(
        P2_U3287) );
  XOR2_X1 U8970 ( .A(n7406), .B(n7407), .Z(n7412) );
  AOI22_X1 U8971 ( .A1(n9476), .A2(n9486), .B1(n9475), .B2(n7536), .ZN(n7408)
         );
  NAND2_X1 U8972 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n10019) );
  OAI211_X1 U8973 ( .C1(n7409), .C2(n9464), .A(n7408), .B(n10019), .ZN(n7410)
         );
  AOI21_X1 U8974 ( .B1(n9477), .B2(n7535), .A(n7410), .ZN(n7411) );
  OAI21_X1 U8975 ( .B1(n7412), .B2(n9470), .A(n7411), .ZN(P1_U3234) );
  NAND2_X1 U8976 ( .A1(n7414), .A2(n7413), .ZN(n7415) );
  NAND2_X1 U8977 ( .A1(n7418), .A2(n8153), .ZN(n7420) );
  AOI22_X1 U8978 ( .A1(n7974), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7973), .B2(
        n7475), .ZN(n7419) );
  XNOR2_X1 U8979 ( .A(n7731), .B(n8094), .ZN(n7583) );
  NOR2_X1 U8980 ( .A1(n7683), .A2(n6602), .ZN(n7584) );
  XNOR2_X1 U8981 ( .A(n7583), .B(n7584), .ZN(n7587) );
  XNOR2_X1 U8982 ( .A(n7588), .B(n7587), .ZN(n7432) );
  NAND2_X1 U8983 ( .A1(n8158), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7427) );
  INV_X1 U8984 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7686) );
  OR2_X1 U8985 ( .A1(n8083), .A2(n7686), .ZN(n7426) );
  INV_X1 U8986 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7476) );
  OR2_X1 U8987 ( .A1(n8162), .A2(n7476), .ZN(n7425) );
  NAND2_X1 U8988 ( .A1(n7422), .A2(n7421), .ZN(n7423) );
  NAND2_X1 U8989 ( .A1(n7594), .A2(n7423), .ZN(n7685) );
  OR2_X1 U8990 ( .A1(n6634), .A2(n7685), .ZN(n7424) );
  OAI22_X1 U8991 ( .A1(n8887), .A2(n7750), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8581), .ZN(n7428) );
  AOI21_X1 U8992 ( .B1(n8890), .B2(n8903), .A(n7428), .ZN(n7429) );
  OAI21_X1 U8993 ( .B1(n7732), .B2(n8885), .A(n7429), .ZN(n7430) );
  AOI21_X1 U8994 ( .B1(n7731), .B2(n8848), .A(n7430), .ZN(n7431) );
  OAI21_X1 U8995 ( .B1(n7432), .B2(n8866), .A(n7431), .ZN(P2_U3238) );
  OR2_X1 U8996 ( .A1(n8259), .A2(n4517), .ZN(n7435) );
  NAND2_X1 U8997 ( .A1(n7663), .A2(n7433), .ZN(n8211) );
  OR2_X1 U8998 ( .A1(n4517), .A2(n7434), .ZN(n7437) );
  AND2_X1 U8999 ( .A1(n7667), .A2(n7664), .ZN(n7441) );
  OR2_X1 U9000 ( .A1(n7436), .A2(n7435), .ZN(n7438) );
  AND2_X1 U9001 ( .A1(n7438), .A2(n7437), .ZN(n7439) );
  NAND2_X1 U9002 ( .A1(n7439), .A2(n8184), .ZN(n7440) );
  NAND2_X1 U9003 ( .A1(n7441), .A2(n7440), .ZN(n10266) );
  XNOR2_X1 U9004 ( .A(n7668), .B(n8184), .ZN(n7445) );
  OAI22_X1 U9005 ( .A1(n7443), .A2(n9182), .B1(n7683), .B2(n9184), .ZN(n7444)
         );
  AOI21_X1 U9006 ( .B1(n7445), .B2(n10194), .A(n7444), .ZN(n7446) );
  OAI21_X1 U9007 ( .B1(n10266), .B2(n7754), .A(n7446), .ZN(n10269) );
  NAND2_X1 U9008 ( .A1(n10269), .A2(n9190), .ZN(n7454) );
  OAI22_X1 U9009 ( .A1(n9190), .A2(n7448), .B1(n7447), .B2(n10199), .ZN(n7452)
         );
  INV_X1 U9010 ( .A(n7449), .ZN(n7450) );
  INV_X1 U9011 ( .A(n7663), .ZN(n10268) );
  OR2_X2 U9012 ( .A1(n7449), .A2(n7663), .ZN(n7671) );
  OAI211_X1 U9013 ( .C1(n7450), .C2(n10268), .A(n10197), .B(n7671), .ZN(n10267) );
  NOR2_X1 U9014 ( .A1(n10267), .A2(n10201), .ZN(n7451) );
  AOI211_X1 U9015 ( .C1(n10205), .C2(n7663), .A(n7452), .B(n7451), .ZN(n7453)
         );
  OAI211_X1 U9016 ( .C1(n10266), .C2(n7763), .A(n7454), .B(n7453), .ZN(
        P2_U3286) );
  NAND2_X1 U9017 ( .A1(n7456), .A2(n7455), .ZN(n7464) );
  XNOR2_X1 U9018 ( .A(n7457), .B(n7464), .ZN(n10144) );
  AOI21_X1 U9019 ( .B1(n10138), .B2(n7459), .A(n7458), .ZN(n10141) );
  AOI22_X1 U9020 ( .A1(n10078), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7460), .B2(
        n10074), .ZN(n7461) );
  OAI21_X1 U9021 ( .B1(n7462), .B2(n9766), .A(n7461), .ZN(n7468) );
  NAND2_X1 U9022 ( .A1(n7500), .A2(n7463), .ZN(n7465) );
  XNOR2_X1 U9023 ( .A(n7465), .B(n7464), .ZN(n7466) );
  AOI222_X1 U9024 ( .A1(n10061), .A2(n7466), .B1(n9488), .B2(n9737), .C1(n9490), .C2(n9735), .ZN(n10143) );
  NOR2_X1 U9025 ( .A1(n10143), .A2(n10078), .ZN(n7467) );
  AOI211_X1 U9026 ( .C1(n10141), .C2(n9770), .A(n7468), .B(n7467), .ZN(n7469)
         );
  OAI21_X1 U9027 ( .B1(n9750), .B2(n10144), .A(n7469), .ZN(P1_U3282) );
  AOI21_X1 U9028 ( .B1(n7471), .B2(n7321), .A(n7470), .ZN(n7473) );
  MUX2_X1 U9029 ( .A(n7686), .B(P2_REG2_REG_12__SCAN_IN), .S(n7611), .Z(n7472)
         );
  NOR2_X1 U9030 ( .A1(n7472), .A2(n7473), .ZN(n7606) );
  AOI21_X1 U9031 ( .B1(n7473), .B2(n7472), .A(n7606), .ZN(n7484) );
  INV_X1 U9032 ( .A(n10187), .ZN(n7648) );
  INV_X1 U9033 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U9034 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7600) );
  MUX2_X1 U9035 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7476), .S(n7611), .Z(n7477)
         );
  OAI21_X1 U9036 ( .B1(n7478), .B2(n7477), .A(n7610), .ZN(n7479) );
  NAND2_X1 U9037 ( .A1(n10181), .A2(n7479), .ZN(n7480) );
  OAI211_X1 U9038 ( .C1(n7648), .C2(n7481), .A(n7600), .B(n7480), .ZN(n7482)
         );
  AOI21_X1 U9039 ( .B1(n7611), .B2(n10183), .A(n7482), .ZN(n7483) );
  OAI21_X1 U9040 ( .B1(n7484), .B2(n10172), .A(n7483), .ZN(P2_U3257) );
  XNOR2_X1 U9041 ( .A(n7487), .B(n7486), .ZN(n7488) );
  XNOR2_X1 U9042 ( .A(n7485), .B(n7488), .ZN(n7494) );
  AOI22_X1 U9043 ( .A1(n9476), .A2(n9485), .B1(n9475), .B2(n7518), .ZN(n7490)
         );
  OAI211_X1 U9044 ( .C1(n7491), .C2(n9464), .A(n7490), .B(n7489), .ZN(n7492)
         );
  AOI21_X1 U9045 ( .B1(n7692), .B2(n9477), .A(n7492), .ZN(n7493) );
  OAI21_X1 U9046 ( .B1(n7494), .B2(n9470), .A(n7493), .ZN(P1_U3222) );
  OR2_X1 U9047 ( .A1(n7495), .A2(n9488), .ZN(n7496) );
  OAI21_X1 U9048 ( .B1(n7498), .B2(n7497), .A(n7510), .ZN(n7544) );
  XNOR2_X1 U9049 ( .A(n7700), .B(n7502), .ZN(n7503) );
  AOI222_X1 U9050 ( .A1(n9488), .A2(n9735), .B1(n9486), .B2(n9737), .C1(n10061), .C2(n7503), .ZN(n7539) );
  NOR2_X2 U9051 ( .A1(n7504), .A2(n7535), .ZN(n7517) );
  AOI21_X1 U9052 ( .B1(n7535), .B2(n7504), .A(n7517), .ZN(n7542) );
  AOI22_X1 U9053 ( .A1(n7542), .A2(n10140), .B1(n10139), .B2(n7535), .ZN(n7505) );
  OAI211_X1 U9054 ( .C1(n9883), .C2(n7544), .A(n7539), .B(n7505), .ZN(n9853)
         );
  NAND2_X1 U9055 ( .A1(n9853), .A2(n10150), .ZN(n7506) );
  OAI21_X1 U9056 ( .B1(n10150), .B2(n5652), .A(n7506), .ZN(P1_U3487) );
  INV_X1 U9057 ( .A(n8040), .ZN(n7524) );
  OAI222_X1 U9058 ( .A1(n9881), .A2(n7524), .B1(P1_U3084), .B2(n7508), .C1(
        n7507), .C2(n8383), .ZN(P1_U3329) );
  NAND2_X1 U9059 ( .A1(n7535), .A2(n9487), .ZN(n7509) );
  XOR2_X1 U9060 ( .A(n7695), .B(n7694), .Z(n9923) );
  INV_X1 U9061 ( .A(n9923), .ZN(n7523) );
  INV_X1 U9062 ( .A(n7511), .ZN(n7699) );
  AOI21_X1 U9063 ( .B1(n7700), .B2(n7512), .A(n7699), .ZN(n7513) );
  XNOR2_X1 U9064 ( .A(n7513), .B(n7694), .ZN(n7514) );
  NAND2_X1 U9065 ( .A1(n7514), .A2(n10061), .ZN(n7516) );
  AOI22_X1 U9066 ( .A1(n9735), .A2(n9487), .B1(n9485), .B2(n9737), .ZN(n7515)
         );
  NAND2_X1 U9067 ( .A1(n7516), .A2(n7515), .ZN(n9922) );
  INV_X1 U9068 ( .A(n7692), .ZN(n9920) );
  INV_X1 U9069 ( .A(n7707), .ZN(n7773) );
  OAI211_X1 U9070 ( .C1(n9920), .C2(n7517), .A(n7773), .B(n10140), .ZN(n9919)
         );
  AOI22_X1 U9071 ( .A1(n10078), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7518), .B2(
        n10074), .ZN(n7520) );
  NAND2_X1 U9072 ( .A1(n7692), .A2(n7711), .ZN(n7519) );
  OAI211_X1 U9073 ( .C1(n9919), .C2(n9744), .A(n7520), .B(n7519), .ZN(n7521)
         );
  AOI21_X1 U9074 ( .B1(n9922), .B2(n10075), .A(n7521), .ZN(n7522) );
  OAI21_X1 U9075 ( .B1(n7523), .B2(n9750), .A(n7522), .ZN(P1_U3279) );
  OAI222_X1 U9076 ( .A1(P2_U3152), .A2(n7525), .B1(n4490), .B2(n7524), .C1(
        n8041), .C2(n9330), .ZN(P2_U3334) );
  INV_X1 U9077 ( .A(n7526), .ZN(n7531) );
  AOI22_X1 U9078 ( .A1(n7528), .A2(n10197), .B1(n6570), .B2(n7527), .ZN(n7529)
         );
  OAI211_X1 U9079 ( .C1(n7531), .C2(n10258), .A(n7530), .B(n7529), .ZN(n7533)
         );
  NAND2_X1 U9080 ( .A1(n7533), .A2(n10295), .ZN(n7532) );
  OAI21_X1 U9081 ( .B1(n10295), .B2(n6771), .A(n7532), .ZN(P2_U3529) );
  NAND2_X1 U9082 ( .A1(n7533), .A2(n9320), .ZN(n7534) );
  OAI21_X1 U9083 ( .B1(n9320), .B2(n7066), .A(n7534), .ZN(P2_U3478) );
  INV_X1 U9084 ( .A(n7535), .ZN(n7538) );
  AOI22_X1 U9085 ( .A1(n10078), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7536), .B2(
        n10074), .ZN(n7537) );
  OAI21_X1 U9086 ( .B1(n7538), .B2(n9766), .A(n7537), .ZN(n7541) );
  NOR2_X1 U9087 ( .A1(n7539), .A2(n10078), .ZN(n7540) );
  AOI211_X1 U9088 ( .C1(n7542), .C2(n9770), .A(n7541), .B(n7540), .ZN(n7543)
         );
  OAI21_X1 U9089 ( .B1(n9750), .B2(n7544), .A(n7543), .ZN(P1_U3280) );
  INV_X1 U9090 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10336) );
  NOR2_X1 U9091 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7545) );
  AOI21_X1 U9092 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7545), .ZN(n10305) );
  NOR2_X1 U9093 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7546) );
  AOI21_X1 U9094 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7546), .ZN(n10308) );
  NOR2_X1 U9095 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7547) );
  AOI21_X1 U9096 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7547), .ZN(n10311) );
  NOR2_X1 U9097 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7548) );
  AOI21_X1 U9098 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7548), .ZN(n10314) );
  NOR2_X1 U9099 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7549) );
  AOI21_X1 U9100 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7549), .ZN(n10317) );
  NOR2_X1 U9101 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7556) );
  XNOR2_X1 U9102 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10347) );
  NAND2_X1 U9103 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7554) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8691) );
  AOI22_X1 U9105 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n7550), .B2(n8691), .ZN(n10345) );
  NAND2_X1 U9106 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7552) );
  XOR2_X1 U9107 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10343) );
  AOI21_X1 U9108 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10296) );
  INV_X1 U9109 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10300) );
  NAND3_X1 U9110 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10298) );
  OAI21_X1 U9111 ( .B1(n10296), .B2(n10300), .A(n10298), .ZN(n10342) );
  NAND2_X1 U9112 ( .A1(n10343), .A2(n10342), .ZN(n7551) );
  NAND2_X1 U9113 ( .A1(n7552), .A2(n7551), .ZN(n10344) );
  NAND2_X1 U9114 ( .A1(n10345), .A2(n10344), .ZN(n7553) );
  NAND2_X1 U9115 ( .A1(n7554), .A2(n7553), .ZN(n10346) );
  NOR2_X1 U9116 ( .A1(n10347), .A2(n10346), .ZN(n7555) );
  NOR2_X1 U9117 ( .A1(n7556), .A2(n7555), .ZN(n7557) );
  NOR2_X1 U9118 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7557), .ZN(n10332) );
  AND2_X1 U9119 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7557), .ZN(n10331) );
  NOR2_X1 U9120 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10331), .ZN(n7558) );
  NOR2_X1 U9121 ( .A1(n10332), .A2(n7558), .ZN(n7559) );
  NAND2_X1 U9122 ( .A1(n7559), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7561) );
  XOR2_X1 U9123 ( .A(n7559), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10330) );
  NAND2_X1 U9124 ( .A1(n10330), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9125 ( .A1(n7561), .A2(n7560), .ZN(n7562) );
  NAND2_X1 U9126 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7562), .ZN(n7564) );
  INV_X1 U9127 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10015) );
  XNOR2_X1 U9128 ( .A(n10015), .B(n7562), .ZN(n10341) );
  NAND2_X1 U9129 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10341), .ZN(n7563) );
  NAND2_X1 U9130 ( .A1(n7564), .A2(n7563), .ZN(n7565) );
  AND2_X1 U9131 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7565), .ZN(n7566) );
  INV_X1 U9132 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10329) );
  XNOR2_X1 U9133 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7565), .ZN(n10328) );
  NOR2_X1 U9134 ( .A1(n10329), .A2(n10328), .ZN(n10327) );
  NOR2_X1 U9135 ( .A1(n7566), .A2(n10327), .ZN(n7568) );
  INV_X1 U9136 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U9137 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  INV_X1 U9138 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10340) );
  XOR2_X1 U9139 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7568), .Z(n10339) );
  NOR2_X1 U9140 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  NOR2_X1 U9141 ( .A1(n7569), .A2(n10338), .ZN(n10326) );
  INV_X1 U9142 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8764) );
  AOI22_X1 U9143 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n8764), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(n6806), .ZN(n10325) );
  NOR2_X1 U9144 ( .A1(n10326), .A2(n10325), .ZN(n10324) );
  AOI21_X1 U9145 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10324), .ZN(n10323) );
  NAND2_X1 U9146 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7570) );
  OAI21_X1 U9147 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7570), .ZN(n10322) );
  NOR2_X1 U9148 ( .A1(n10323), .A2(n10322), .ZN(n10321) );
  AOI21_X1 U9149 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10321), .ZN(n10320) );
  NOR2_X1 U9150 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7571) );
  AOI21_X1 U9151 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7571), .ZN(n10319) );
  NAND2_X1 U9152 ( .A1(n10320), .A2(n10319), .ZN(n10318) );
  OAI21_X1 U9153 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10318), .ZN(n10316) );
  NAND2_X1 U9154 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  OAI21_X1 U9155 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10315), .ZN(n10313) );
  NAND2_X1 U9156 ( .A1(n10314), .A2(n10313), .ZN(n10312) );
  OAI21_X1 U9157 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10312), .ZN(n10310) );
  NAND2_X1 U9158 ( .A1(n10311), .A2(n10310), .ZN(n10309) );
  OAI21_X1 U9159 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10309), .ZN(n10307) );
  NAND2_X1 U9160 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  OAI21_X1 U9161 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10306), .ZN(n10304) );
  NAND2_X1 U9162 ( .A1(n10305), .A2(n10304), .ZN(n10303) );
  OAI21_X1 U9163 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10303), .ZN(n10335) );
  NOR2_X1 U9164 ( .A1(n10336), .A2(n10335), .ZN(n7572) );
  NAND2_X1 U9165 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  OAI21_X1 U9166 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7572), .A(n10334), .ZN(
        n7574) );
  XNOR2_X1 U9167 ( .A(n4651), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7573) );
  XNOR2_X1 U9168 ( .A(n7574), .B(n7573), .ZN(ADD_1071_U4) );
  NAND2_X1 U9169 ( .A1(n7575), .A2(n8153), .ZN(n7577) );
  AOI22_X1 U9170 ( .A1(n7974), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7973), .B2(
        n7611), .ZN(n7576) );
  INV_X1 U9171 ( .A(n7743), .ZN(n10276) );
  XNOR2_X1 U9172 ( .A(n7743), .B(n8094), .ZN(n7578) );
  OR2_X1 U9173 ( .A1(n7750), .A2(n6602), .ZN(n7579) );
  NAND2_X1 U9174 ( .A1(n7578), .A2(n7579), .ZN(n7620) );
  INV_X1 U9175 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9176 ( .A(n7579), .ZN(n7580) );
  NAND2_X1 U9177 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  AND2_X1 U9178 ( .A1(n7620), .A2(n7582), .ZN(n7590) );
  INV_X1 U9179 ( .A(n7583), .ZN(n7585) );
  AND2_X1 U9180 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  NAND2_X1 U9181 ( .A1(n7589), .A2(n7590), .ZN(n7621) );
  OAI21_X1 U9182 ( .B1(n7590), .B2(n7589), .A(n7621), .ZN(n7591) );
  NAND2_X1 U9183 ( .A1(n7591), .A2(n8882), .ZN(n7605) );
  INV_X1 U9184 ( .A(n7685), .ZN(n7603) );
  NAND2_X1 U9185 ( .A1(n8158), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7599) );
  INV_X1 U9186 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7592) );
  OR2_X1 U9187 ( .A1(n8162), .A2(n7592), .ZN(n7598) );
  INV_X1 U9188 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7756) );
  OR2_X1 U9189 ( .A1(n8083), .A2(n7756), .ZN(n7597) );
  INV_X1 U9190 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9191 ( .A1(n7594), .A2(n7593), .ZN(n7595) );
  NAND2_X1 U9192 ( .A1(n7627), .A2(n7595), .ZN(n7755) );
  OR2_X1 U9193 ( .A1(n6634), .A2(n7755), .ZN(n7596) );
  INV_X1 U9194 ( .A(n7846), .ZN(n8900) );
  NAND2_X1 U9195 ( .A1(n8900), .A2(n8875), .ZN(n7601) );
  OAI211_X1 U9196 ( .C1(n7683), .C2(n8873), .A(n7601), .B(n7600), .ZN(n7602)
         );
  AOI21_X1 U9197 ( .B1(n7603), .B2(n8871), .A(n7602), .ZN(n7604) );
  OAI211_X1 U9198 ( .C1(n10276), .C2(n8893), .A(n7605), .B(n7604), .ZN(
        P2_U3226) );
  INV_X1 U9199 ( .A(n7611), .ZN(n7607) );
  AOI21_X1 U9200 ( .B1(n7686), .B2(n7607), .A(n7606), .ZN(n7609) );
  AOI22_X1 U9201 ( .A1(n7644), .A2(n7756), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7640), .ZN(n7608) );
  NOR2_X1 U9202 ( .A1(n7609), .A2(n7608), .ZN(n7639) );
  AOI21_X1 U9203 ( .B1(n7609), .B2(n7608), .A(n7639), .ZN(n7619) );
  INV_X1 U9204 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7616) );
  OAI21_X1 U9205 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7611), .A(n7610), .ZN(
        n7613) );
  AOI22_X1 U9206 ( .A1(n7644), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7592), .B2(
        n7640), .ZN(n7612) );
  NAND2_X1 U9207 ( .A1(n7612), .A2(n7613), .ZN(n7643) );
  OAI21_X1 U9208 ( .B1(n7613), .B2(n7612), .A(n7643), .ZN(n7614) );
  NAND2_X1 U9209 ( .A1(n10181), .A2(n7614), .ZN(n7615) );
  NAND2_X1 U9210 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7633) );
  OAI211_X1 U9211 ( .C1(n7648), .C2(n7616), .A(n7615), .B(n7633), .ZN(n7617)
         );
  AOI21_X1 U9212 ( .B1(n7644), .B2(n10183), .A(n7617), .ZN(n7618) );
  OAI21_X1 U9213 ( .B1(n7619), .B2(n10172), .A(n7618), .ZN(P2_U3258) );
  NAND2_X1 U9214 ( .A1(n7622), .A2(n8153), .ZN(n7624) );
  AOI22_X1 U9215 ( .A1(n7974), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7973), .B2(
        n7644), .ZN(n7623) );
  XNOR2_X1 U9216 ( .A(n9299), .B(n8116), .ZN(n7839) );
  NOR2_X1 U9217 ( .A1(n7846), .A2(n6602), .ZN(n7838) );
  XNOR2_X1 U9218 ( .A(n7839), .B(n7838), .ZN(n7841) );
  XNOR2_X1 U9219 ( .A(n7842), .B(n7841), .ZN(n7638) );
  INV_X1 U9220 ( .A(n7750), .ZN(n8901) );
  NAND2_X1 U9221 ( .A1(n8158), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7632) );
  INV_X1 U9222 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7826) );
  OR2_X1 U9223 ( .A1(n8083), .A2(n7826), .ZN(n7631) );
  INV_X1 U9224 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7625) );
  OR2_X1 U9225 ( .A1(n8162), .A2(n7625), .ZN(n7630) );
  NAND2_X1 U9226 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  NAND2_X1 U9227 ( .A1(n7796), .A2(n7628), .ZN(n7843) );
  OR2_X1 U9228 ( .A1(n6634), .A2(n7843), .ZN(n7629) );
  OAI21_X1 U9229 ( .B1(n8887), .B2(n7832), .A(n7633), .ZN(n7634) );
  AOI21_X1 U9230 ( .B1(n8890), .B2(n8901), .A(n7634), .ZN(n7635) );
  OAI21_X1 U9231 ( .B1(n7755), .B2(n8885), .A(n7635), .ZN(n7636) );
  AOI21_X1 U9232 ( .B1(n9299), .B2(n8848), .A(n7636), .ZN(n7637) );
  OAI21_X1 U9233 ( .B1(n7638), .B2(n8866), .A(n7637), .ZN(P2_U3236) );
  AOI21_X1 U9234 ( .B1(n7640), .B2(n7756), .A(n7639), .ZN(n7642) );
  AOI22_X1 U9235 ( .A1(n7870), .A2(n7826), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7865), .ZN(n7641) );
  NOR2_X1 U9236 ( .A1(n7642), .A2(n7641), .ZN(n7864) );
  AOI21_X1 U9237 ( .B1(n7642), .B2(n7641), .A(n7864), .ZN(n7653) );
  AOI22_X1 U9238 ( .A1(n7870), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7625), .B2(
        n7865), .ZN(n7646) );
  OAI21_X1 U9239 ( .B1(n7644), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7643), .ZN(
        n7645) );
  NAND2_X1 U9240 ( .A1(n7646), .A2(n7645), .ZN(n7869) );
  OAI21_X1 U9241 ( .B1(n7646), .B2(n7645), .A(n7869), .ZN(n7651) );
  INV_X1 U9242 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9243 ( .A1(n10183), .A2(n7870), .ZN(n7647) );
  NAND2_X1 U9244 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7844) );
  OAI211_X1 U9245 ( .C1(n7649), .C2(n7648), .A(n7647), .B(n7844), .ZN(n7650)
         );
  AOI21_X1 U9246 ( .B1(n7651), .B2(n10181), .A(n7650), .ZN(n7652) );
  OAI21_X1 U9247 ( .B1(n7653), .B2(n10172), .A(n7652), .ZN(P2_U3259) );
  INV_X1 U9248 ( .A(n9848), .ZN(n7776) );
  NAND2_X1 U9249 ( .A1(n4571), .A2(n7655), .ZN(n7656) );
  XNOR2_X1 U9250 ( .A(n7654), .B(n7656), .ZN(n7657) );
  NAND2_X1 U9251 ( .A1(n7657), .A2(n9428), .ZN(n7662) );
  INV_X1 U9252 ( .A(n7774), .ZN(n7658) );
  OAI22_X1 U9253 ( .A1(n9753), .A2(n9451), .B1(n9453), .B2(n7658), .ZN(n7659)
         );
  AOI211_X1 U9254 ( .C1(n9474), .C2(n9486), .A(n7660), .B(n7659), .ZN(n7661)
         );
  OAI211_X1 U9255 ( .C1(n7776), .C2(n9372), .A(n7662), .B(n7661), .ZN(P1_U3232) );
  NAND2_X1 U9256 ( .A1(n7663), .A2(n8903), .ZN(n7665) );
  AND2_X1 U9257 ( .A1(n7665), .A2(n7664), .ZN(n7666) );
  NAND2_X1 U9258 ( .A1(n7667), .A2(n7666), .ZN(n7677) );
  NAND2_X1 U9259 ( .A1(n7731), .A2(n7683), .ZN(n8264) );
  NAND2_X1 U9260 ( .A1(n8265), .A2(n8264), .ZN(n8188) );
  XNOR2_X1 U9261 ( .A(n7677), .B(n8188), .ZN(n7741) );
  NAND2_X1 U9262 ( .A1(n7668), .A2(n8254), .ZN(n7669) );
  NAND2_X1 U9263 ( .A1(n7669), .A2(n8211), .ZN(n7681) );
  XOR2_X1 U9264 ( .A(n7681), .B(n8188), .Z(n7670) );
  AOI222_X1 U9265 ( .A1(n10194), .A2(n7670), .B1(n8901), .B2(n9197), .C1(n8903), .C2(n9195), .ZN(n7736) );
  AOI21_X1 U9266 ( .B1(n7731), .B2(n7671), .A(n7684), .ZN(n7739) );
  AOI22_X1 U9267 ( .A1(n7739), .A2(n10197), .B1(n6570), .B2(n7731), .ZN(n7672)
         );
  OAI211_X1 U9268 ( .C1(n9297), .C2(n7741), .A(n7736), .B(n7672), .ZN(n7674)
         );
  NAND2_X1 U9269 ( .A1(n7674), .A2(n10295), .ZN(n7673) );
  OAI21_X1 U9270 ( .B1(n10295), .B2(n7320), .A(n7673), .ZN(P2_U3531) );
  INV_X1 U9271 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U9272 ( .A1(n7674), .A2(n9320), .ZN(n7675) );
  OAI21_X1 U9273 ( .B1(n9320), .B2(n7676), .A(n7675), .ZN(P2_U3484) );
  NAND2_X1 U9274 ( .A1(n7677), .A2(n8188), .ZN(n7679) );
  INV_X1 U9275 ( .A(n7683), .ZN(n8902) );
  NAND2_X1 U9276 ( .A1(n7731), .A2(n8902), .ZN(n7678) );
  NAND2_X1 U9277 ( .A1(n7679), .A2(n7678), .ZN(n7744) );
  NAND2_X1 U9278 ( .A1(n7743), .A2(n7750), .ZN(n8272) );
  XNOR2_X1 U9279 ( .A(n7744), .B(n8190), .ZN(n10280) );
  INV_X1 U9280 ( .A(n10280), .ZN(n7691) );
  INV_X1 U9281 ( .A(n8264), .ZN(n7680) );
  XNOR2_X1 U9282 ( .A(n7748), .B(n8190), .ZN(n7682) );
  OAI222_X1 U9283 ( .A1(n9184), .A2(n7846), .B1(n9182), .B2(n7683), .C1(n9180), 
        .C2(n7682), .ZN(n10277) );
  NAND2_X1 U9284 ( .A1(n7684), .A2(n10276), .ZN(n7757) );
  OAI211_X1 U9285 ( .C1(n7684), .C2(n10276), .A(n10197), .B(n7757), .ZN(n10274) );
  OAI22_X1 U9286 ( .A1(n9190), .A2(n7686), .B1(n7685), .B2(n10199), .ZN(n7687)
         );
  AOI21_X1 U9287 ( .B1(n7743), .B2(n10205), .A(n7687), .ZN(n7688) );
  OAI21_X1 U9288 ( .B1(n10274), .B2(n10201), .A(n7688), .ZN(n7689) );
  AOI21_X1 U9289 ( .B1(n10277), .B2(n9190), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9290 ( .B1(n9214), .B2(n7691), .A(n7690), .ZN(P2_U3284) );
  AND2_X1 U9291 ( .A1(n7692), .A2(n9486), .ZN(n7693) );
  NAND2_X1 U9292 ( .A1(n9848), .A2(n9485), .ZN(n7696) );
  OR2_X1 U9293 ( .A1(n9848), .A2(n9485), .ZN(n7697) );
  XNOR2_X1 U9294 ( .A(n7880), .B(n7879), .ZN(n9918) );
  INV_X1 U9295 ( .A(n9918), .ZN(n7715) );
  NAND2_X1 U9296 ( .A1(n7702), .A2(n7701), .ZN(n7765) );
  OAI211_X1 U9297 ( .C1(n5076), .C2(n7704), .A(n7901), .B(n10061), .ZN(n7706)
         );
  AOI22_X1 U9298 ( .A1(n9735), .A2(n9485), .B1(n9736), .B2(n9737), .ZN(n7705)
         );
  NAND2_X1 U9299 ( .A1(n7706), .A2(n7705), .ZN(n9917) );
  NAND2_X1 U9300 ( .A1(n7707), .A2(n7776), .ZN(n7708) );
  INV_X1 U9301 ( .A(n7708), .ZN(n7772) );
  INV_X1 U9302 ( .A(n9357), .ZN(n9915) );
  OAI211_X1 U9303 ( .C1(n7772), .C2(n9915), .A(n10140), .B(n9761), .ZN(n9914)
         );
  INV_X1 U9304 ( .A(n9345), .ZN(n7709) );
  OAI22_X1 U9305 ( .A1(n10075), .A2(n5453), .B1(n7709), .B2(n7922), .ZN(n7710)
         );
  AOI21_X1 U9306 ( .B1(n9357), .B2(n7711), .A(n7710), .ZN(n7712) );
  OAI21_X1 U9307 ( .B1(n9914), .B2(n9744), .A(n7712), .ZN(n7713) );
  AOI21_X1 U9308 ( .B1(n9917), .B2(n10075), .A(n7713), .ZN(n7714) );
  OAI21_X1 U9309 ( .B1(n7715), .B2(n9750), .A(n7714), .ZN(P1_U3277) );
  OAI21_X1 U9310 ( .B1(n7718), .B2(n7717), .A(n7716), .ZN(n7719) );
  INV_X1 U9311 ( .A(n7719), .ZN(n7726) );
  NAND2_X1 U9312 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n9346) );
  OAI21_X1 U9313 ( .B1(n9971), .B2(n7720), .A(n9346), .ZN(n7724) );
  AOI211_X1 U9314 ( .C1(n5453), .C2(n7722), .A(n7721), .B(n10032), .ZN(n7723)
         );
  AOI211_X1 U9315 ( .C1(n9999), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7724), .B(
        n7723), .ZN(n7725) );
  OAI21_X1 U9316 ( .B1(n7726), .B2(n9982), .A(n7725), .ZN(P1_U3255) );
  INV_X1 U9317 ( .A(n8062), .ZN(n7730) );
  OAI222_X1 U9318 ( .A1(n8383), .A2(n7728), .B1(n9881), .B2(n7730), .C1(n7727), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9319 ( .A1(n9330), .A2(n8444), .B1(n4490), .B2(n7730), .C1(
        P2_U3152), .C2(n7729), .ZN(P2_U3333) );
  INV_X1 U9320 ( .A(n7731), .ZN(n7735) );
  INV_X1 U9321 ( .A(n7732), .ZN(n7733) );
  INV_X1 U9322 ( .A(n10199), .ZN(n9161) );
  AOI22_X1 U9323 ( .A1(n10210), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7733), .B2(
        n9161), .ZN(n7734) );
  OAI21_X1 U9324 ( .B1(n7735), .B2(n9164), .A(n7734), .ZN(n7738) );
  NOR2_X1 U9325 ( .A1(n7736), .A2(n10210), .ZN(n7737) );
  AOI211_X1 U9326 ( .C1(n7739), .C2(n9211), .A(n7738), .B(n7737), .ZN(n7740)
         );
  OAI21_X1 U9327 ( .B1(n9214), .B2(n7741), .A(n7740), .ZN(P2_U3285) );
  INV_X1 U9328 ( .A(n8075), .ZN(n7782) );
  OAI222_X1 U9329 ( .A1(P2_U3152), .A2(n7742), .B1(n4490), .B2(n7782), .C1(
        n8076), .C2(n9330), .ZN(P2_U3332) );
  OR2_X1 U9330 ( .A1(n9299), .A2(n7846), .ZN(n8278) );
  NAND2_X1 U9331 ( .A1(n9299), .A2(n7846), .ZN(n8277) );
  NAND2_X1 U9332 ( .A1(n7745), .A2(n8274), .ZN(n7746) );
  NAND2_X1 U9333 ( .A1(n7811), .A2(n7746), .ZN(n9302) );
  INV_X1 U9334 ( .A(n8273), .ZN(n7747) );
  NAND2_X1 U9335 ( .A1(n7749), .A2(n8274), .ZN(n7790) );
  OAI21_X1 U9336 ( .B1(n8274), .B2(n7749), .A(n7790), .ZN(n7752) );
  OAI22_X1 U9337 ( .A1(n7750), .A2(n9182), .B1(n7832), .B2(n9184), .ZN(n7751)
         );
  AOI21_X1 U9338 ( .B1(n7752), .B2(n10194), .A(n7751), .ZN(n7753) );
  OAI21_X1 U9339 ( .B1(n9302), .B2(n7754), .A(n7753), .ZN(n9304) );
  NAND2_X1 U9340 ( .A1(n9304), .A2(n9190), .ZN(n7762) );
  OAI22_X1 U9341 ( .A1(n9190), .A2(n7756), .B1(n7755), .B2(n10199), .ZN(n7760)
         );
  AOI21_X1 U9342 ( .B1(n7757), .B2(n9299), .A(n10261), .ZN(n7758) );
  NAND2_X1 U9343 ( .A1(n7758), .A2(n7823), .ZN(n9300) );
  NOR2_X1 U9344 ( .A1(n9300), .A2(n10201), .ZN(n7759) );
  AOI211_X1 U9345 ( .C1(n10205), .C2(n9299), .A(n7760), .B(n7759), .ZN(n7761)
         );
  OAI211_X1 U9346 ( .C1(n9302), .C2(n7763), .A(n7762), .B(n7761), .ZN(P2_U3283) );
  OAI21_X1 U9347 ( .B1(n7767), .B2(n7765), .A(n7764), .ZN(n7771) );
  OAI22_X1 U9348 ( .A1(n9753), .A2(n10058), .B1(n7766), .B2(n10056), .ZN(n7770) );
  XNOR2_X1 U9349 ( .A(n7768), .B(n7767), .ZN(n9852) );
  NOR2_X1 U9350 ( .A1(n9852), .A2(n10064), .ZN(n7769) );
  AOI211_X1 U9351 ( .C1(n10061), .C2(n7771), .A(n7770), .B(n7769), .ZN(n9851)
         );
  AOI21_X1 U9352 ( .B1(n9848), .B2(n7773), .A(n7772), .ZN(n9849) );
  AOI22_X1 U9353 ( .A1(n10078), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7774), .B2(
        n10074), .ZN(n7775) );
  OAI21_X1 U9354 ( .B1(n7776), .B2(n9766), .A(n7775), .ZN(n7778) );
  NOR2_X1 U9355 ( .A1(n9852), .A2(n9767), .ZN(n7777) );
  AOI211_X1 U9356 ( .C1(n9849), .C2(n9770), .A(n7778), .B(n7777), .ZN(n7779)
         );
  OAI21_X1 U9357 ( .B1(n9851), .B2(n10078), .A(n7779), .ZN(P1_U3278) );
  OAI222_X1 U9358 ( .A1(n9881), .A2(n7782), .B1(P1_U3084), .B2(n7781), .C1(
        n7780), .C2(n8383), .ZN(P1_U3327) );
  INV_X1 U9359 ( .A(n8091), .ZN(n7852) );
  AOI21_X1 U9360 ( .B1(n9875), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7783), .ZN(
        n7784) );
  OAI21_X1 U9361 ( .B1(n7852), .B2(n9881), .A(n7784), .ZN(P1_U3326) );
  NAND2_X1 U9362 ( .A1(n7785), .A2(n8153), .ZN(n7787) );
  AOI22_X1 U9363 ( .A1(n7974), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7973), .B2(
        n7870), .ZN(n7786) );
  NAND2_X1 U9364 ( .A1(n7849), .A2(n7832), .ZN(n8283) );
  INV_X1 U9365 ( .A(n8277), .ZN(n7788) );
  NOR2_X1 U9366 ( .A1(n5054), .A2(n7788), .ZN(n7789) );
  NAND2_X1 U9367 ( .A1(n7790), .A2(n7789), .ZN(n7791) );
  NAND2_X1 U9368 ( .A1(n7792), .A2(n8153), .ZN(n7794) );
  AOI22_X1 U9369 ( .A1(n7974), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7973), .B2(
        n8930), .ZN(n7793) );
  INV_X1 U9370 ( .A(n8083), .ZN(n8157) );
  NAND2_X1 U9371 ( .A1(n8157), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7802) );
  INV_X1 U9372 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7872) );
  OR2_X1 U9373 ( .A1(n8162), .A2(n7872), .ZN(n7801) );
  NAND2_X1 U9374 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND2_X1 U9375 ( .A1(n7804), .A2(n7797), .ZN(n8884) );
  OR2_X1 U9376 ( .A1(n6634), .A2(n8884), .ZN(n7800) );
  INV_X1 U9377 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7798) );
  OR2_X1 U9378 ( .A1(n8121), .A2(n7798), .ZN(n7799) );
  NAND2_X1 U9379 ( .A1(n9293), .A2(n7930), .ZN(n8286) );
  NAND2_X1 U9380 ( .A1(n8287), .A2(n8286), .ZN(n8281) );
  XNOR2_X1 U9381 ( .A(n8136), .B(n8281), .ZN(n7810) );
  NAND2_X1 U9382 ( .A1(n8158), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7809) );
  INV_X1 U9383 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8941) );
  OR2_X1 U9384 ( .A1(n8162), .A2(n8941), .ZN(n7808) );
  INV_X1 U9385 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9205) );
  OR2_X1 U9386 ( .A1(n8083), .A2(n9205), .ZN(n7807) );
  INV_X1 U9387 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U9388 ( .A1(n7804), .A2(n7803), .ZN(n7805) );
  NAND2_X1 U9389 ( .A1(n7950), .A2(n7805), .ZN(n9204) );
  OR2_X1 U9390 ( .A1(n6634), .A2(n9204), .ZN(n7806) );
  INV_X1 U9391 ( .A(n9181), .ZN(n8898) );
  INV_X1 U9392 ( .A(n7832), .ZN(n8899) );
  AOI222_X1 U9393 ( .A1(n10194), .A2(n7810), .B1(n8898), .B2(n9197), .C1(n8899), .C2(n9195), .ZN(n9296) );
  INV_X1 U9394 ( .A(n9299), .ZN(n7812) );
  NAND2_X1 U9395 ( .A1(n7813), .A2(n8281), .ZN(n8388) );
  OAI21_X1 U9396 ( .B1(n7813), .B2(n8281), .A(n8388), .ZN(n9292) );
  INV_X1 U9397 ( .A(n9293), .ZN(n8894) );
  NOR2_X2 U9398 ( .A1(n7823), .A2(n7849), .ZN(n7814) );
  INV_X1 U9399 ( .A(n7814), .ZN(n7824) );
  AOI21_X1 U9400 ( .B1(n9293), .B2(n7824), .A(n9208), .ZN(n9294) );
  NAND2_X1 U9401 ( .A1(n9294), .A2(n9211), .ZN(n7817) );
  INV_X1 U9402 ( .A(n8884), .ZN(n7815) );
  AOI22_X1 U9403 ( .A1(n10210), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7815), .B2(
        n9161), .ZN(n7816) );
  OAI211_X1 U9404 ( .C1(n8894), .C2(n9164), .A(n7817), .B(n7816), .ZN(n7818)
         );
  AOI21_X1 U9405 ( .B1(n9292), .B2(n10207), .A(n7818), .ZN(n7819) );
  OAI21_X1 U9406 ( .B1(n9296), .B2(n10210), .A(n7819), .ZN(P2_U3281) );
  XNOR2_X1 U9407 ( .A(n7820), .B(n8280), .ZN(n9899) );
  INV_X1 U9408 ( .A(n9899), .ZN(n7831) );
  NAND2_X1 U9409 ( .A1(n7790), .A2(n8277), .ZN(n7821) );
  XNOR2_X1 U9410 ( .A(n7821), .B(n5054), .ZN(n7822) );
  OAI222_X1 U9411 ( .A1(n9184), .A2(n7930), .B1(n9182), .B2(n7846), .C1(n7822), 
        .C2(n9180), .ZN(n9897) );
  INV_X1 U9412 ( .A(n7849), .ZN(n9895) );
  INV_X1 U9413 ( .A(n7823), .ZN(n7825) );
  OAI21_X1 U9414 ( .B1(n9895), .B2(n7825), .A(n7824), .ZN(n9896) );
  OAI22_X1 U9415 ( .A1(n9190), .A2(n7826), .B1(n7843), .B2(n10199), .ZN(n7827)
         );
  AOI21_X1 U9416 ( .B1(n7849), .B2(n10205), .A(n7827), .ZN(n7828) );
  OAI21_X1 U9417 ( .B1(n9896), .B2(n8991), .A(n7828), .ZN(n7829) );
  AOI21_X1 U9418 ( .B1(n9897), .B2(n9190), .A(n7829), .ZN(n7830) );
  OAI21_X1 U9419 ( .B1(n9214), .B2(n7831), .A(n7830), .ZN(P2_U3282) );
  XNOR2_X1 U9420 ( .A(n7849), .B(n8094), .ZN(n7833) );
  OR2_X1 U9421 ( .A1(n7832), .A2(n6602), .ZN(n7834) );
  NAND2_X1 U9422 ( .A1(n7833), .A2(n7834), .ZN(n7927) );
  INV_X1 U9423 ( .A(n7833), .ZN(n7836) );
  INV_X1 U9424 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U9425 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  NAND2_X1 U9426 ( .A1(n7927), .A2(n7837), .ZN(n7928) );
  NAND2_X1 U9427 ( .A1(n7839), .A2(n7838), .ZN(n7840) );
  AOI21_X1 U9428 ( .B1(n7928), .B2(n7929), .A(n4565), .ZN(n7851) );
  NOR2_X1 U9429 ( .A1(n8885), .A2(n7843), .ZN(n7848) );
  INV_X1 U9430 ( .A(n7930), .ZN(n9196) );
  NAND2_X1 U9431 ( .A1(n9196), .A2(n8875), .ZN(n7845) );
  OAI211_X1 U9432 ( .C1(n7846), .C2(n8873), .A(n7845), .B(n7844), .ZN(n7847)
         );
  AOI211_X1 U9433 ( .C1(n7849), .C2(n8848), .A(n7848), .B(n7847), .ZN(n7850)
         );
  OAI21_X1 U9434 ( .B1(n7851), .B2(n8866), .A(n7850), .ZN(P2_U3217) );
  OAI222_X1 U9435 ( .A1(n9330), .A2(n8689), .B1(n4490), .B2(n7852), .C1(n8408), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9436 ( .A(n9760), .ZN(n9842) );
  XNOR2_X1 U9437 ( .A(n7855), .B(n7854), .ZN(n7856) );
  XNOR2_X1 U9438 ( .A(n7853), .B(n7856), .ZN(n7857) );
  NAND2_X1 U9439 ( .A1(n7857), .A2(n9428), .ZN(n7863) );
  INV_X1 U9440 ( .A(n7858), .ZN(n7861) );
  INV_X1 U9441 ( .A(n9764), .ZN(n7859) );
  OAI22_X1 U9442 ( .A1(n9753), .A2(n9464), .B1(n9453), .B2(n7859), .ZN(n7860)
         );
  AOI211_X1 U9443 ( .C1(n9476), .C2(n9727), .A(n7861), .B(n7860), .ZN(n7862)
         );
  OAI211_X1 U9444 ( .C1(n9842), .C2(n9372), .A(n7863), .B(n7862), .ZN(P1_U3239) );
  AOI21_X1 U9445 ( .B1(n7865), .B2(n7826), .A(n7864), .ZN(n8929) );
  XNOR2_X1 U9446 ( .A(n8929), .B(n8930), .ZN(n7866) );
  NOR2_X1 U9447 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7866), .ZN(n8931) );
  AOI21_X1 U9448 ( .B1(n7866), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8931), .ZN(
        n7877) );
  NAND2_X1 U9449 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8886) );
  INV_X1 U9450 ( .A(n8886), .ZN(n7868) );
  NOR2_X1 U9451 ( .A1(n10170), .A2(n8938), .ZN(n7867) );
  AOI211_X1 U9452 ( .C1(n10187), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7868), .B(
        n7867), .ZN(n7876) );
  OAI21_X1 U9453 ( .B1(n7870), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7869), .ZN(
        n8937) );
  XNOR2_X1 U9454 ( .A(n8937), .B(n8938), .ZN(n7871) );
  INV_X1 U9455 ( .A(n7871), .ZN(n7874) );
  NOR2_X1 U9456 ( .A1(n7872), .A2(n7871), .ZN(n8939) );
  INV_X1 U9457 ( .A(n8939), .ZN(n7873) );
  OAI211_X1 U9458 ( .C1(n7874), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10181), .B(
        n7873), .ZN(n7875) );
  OAI211_X1 U9459 ( .C1(n7877), .C2(n10172), .A(n7876), .B(n7875), .ZN(
        P2_U3260) );
  NOR2_X1 U9460 ( .A1(n9357), .A2(n9484), .ZN(n7878) );
  NOR2_X1 U9461 ( .A1(n9837), .A2(n9738), .ZN(n7883) );
  INV_X1 U9462 ( .A(n9837), .ZN(n9722) );
  NAND2_X1 U9463 ( .A1(n9828), .A2(n9710), .ZN(n7885) );
  INV_X1 U9464 ( .A(n9828), .ZN(n9689) );
  OR2_X1 U9465 ( .A1(n9823), .A2(n9693), .ZN(n7886) );
  NAND2_X1 U9466 ( .A1(n9670), .A2(n7886), .ZN(n7887) );
  INV_X1 U9467 ( .A(n9823), .ZN(n9676) );
  NAND2_X1 U9468 ( .A1(n7887), .A2(n5078), .ZN(n9657) );
  AOI21_X2 U9469 ( .B1(n9657), .B2(n9663), .A(n7888), .ZN(n9644) );
  NAND2_X1 U9470 ( .A1(n9812), .A2(n9665), .ZN(n7889) );
  INV_X1 U9471 ( .A(n9812), .ZN(n9648) );
  AOI22_X1 U9472 ( .A1(n9644), .A2(n7889), .B1(n9386), .B2(n9648), .ZN(n9631)
         );
  INV_X1 U9473 ( .A(n9631), .ZN(n7891) );
  INV_X1 U9474 ( .A(n9792), .ZN(n9593) );
  OAI22_X1 U9475 ( .A1(n9574), .A2(n9575), .B1(n9600), .B2(n9789), .ZN(n9559)
         );
  XNOR2_X1 U9476 ( .A(n7893), .B(n7921), .ZN(n9781) );
  INV_X1 U9477 ( .A(n9789), .ZN(n9586) );
  OR2_X2 U9478 ( .A1(n9717), .A2(n9832), .ZN(n9700) );
  NOR2_X2 U9479 ( .A1(n9700), .A2(n9828), .ZN(n9685) );
  NAND2_X1 U9480 ( .A1(n9685), .A2(n9676), .ZN(n9671) );
  OR2_X2 U9481 ( .A1(n9671), .A2(n9818), .ZN(n9658) );
  NOR2_X2 U9482 ( .A1(n9792), .A2(n9604), .ZN(n9590) );
  NAND2_X1 U9483 ( .A1(n9586), .A2(n9590), .ZN(n9580) );
  NAND2_X1 U9484 ( .A1(n9777), .A2(n9561), .ZN(n7894) );
  OAI22_X1 U9485 ( .A1(n7896), .A2(n9766), .B1(n7895), .B2(n10075), .ZN(n7897)
         );
  AOI21_X1 U9486 ( .B1(n9778), .B2(n9770), .A(n7897), .ZN(n7926) );
  INV_X1 U9487 ( .A(P1_B_REG_SCAN_IN), .ZN(n7898) );
  NOR2_X1 U9488 ( .A1(n5925), .A2(n7898), .ZN(n7899) );
  NOR2_X1 U9489 ( .A1(n10058), .A2(n7899), .ZN(n8132) );
  NAND2_X1 U9490 ( .A1(n9691), .A2(n9692), .ZN(n9690) );
  NAND2_X1 U9491 ( .A1(n9690), .A2(n7908), .ZN(n9678) );
  NAND2_X1 U9492 ( .A1(n9566), .A2(n9567), .ZN(n9565) );
  OAI21_X1 U9493 ( .B1(n7923), .B2(n7922), .A(n9780), .ZN(n7924) );
  NAND2_X1 U9494 ( .A1(n7924), .A2(n10075), .ZN(n7925) );
  OAI211_X1 U9495 ( .C1(n9781), .C2(n9750), .A(n7926), .B(n7925), .ZN(P1_U3355) );
  XNOR2_X1 U9496 ( .A(n9293), .B(n8094), .ZN(n7931) );
  OR2_X1 U9497 ( .A1(n7930), .A2(n6602), .ZN(n7932) );
  NAND2_X1 U9498 ( .A1(n7931), .A2(n7932), .ZN(n7936) );
  INV_X1 U9499 ( .A(n7931), .ZN(n7934) );
  INV_X1 U9500 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U9501 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  AND2_X1 U9502 ( .A1(n7936), .A2(n7935), .ZN(n8881) );
  NAND2_X1 U9503 ( .A1(n8879), .A2(n7936), .ZN(n8816) );
  NAND2_X1 U9504 ( .A1(n7937), .A2(n8153), .ZN(n7939) );
  AOI22_X1 U9505 ( .A1(n7974), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7973), .B2(
        n8955), .ZN(n7938) );
  XNOR2_X1 U9506 ( .A(n9287), .B(n8094), .ZN(n7940) );
  OR2_X1 U9507 ( .A1(n9181), .A2(n6602), .ZN(n7941) );
  NAND2_X1 U9508 ( .A1(n7940), .A2(n7941), .ZN(n7945) );
  INV_X1 U9509 ( .A(n7940), .ZN(n7943) );
  INV_X1 U9510 ( .A(n7941), .ZN(n7942) );
  NAND2_X1 U9511 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  AND2_X1 U9512 ( .A1(n7945), .A2(n7944), .ZN(n8817) );
  NAND2_X1 U9513 ( .A1(n8816), .A2(n8817), .ZN(n8815) );
  NAND2_X1 U9514 ( .A1(n8815), .A2(n7945), .ZN(n8823) );
  NAND2_X1 U9515 ( .A1(n7946), .A2(n8153), .ZN(n7948) );
  AOI22_X1 U9516 ( .A1(n7974), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7973), .B2(
        n8971), .ZN(n7947) );
  XNOR2_X1 U9517 ( .A(n9284), .B(n8116), .ZN(n7957) );
  NAND2_X1 U9518 ( .A1(n8158), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7955) );
  INV_X1 U9519 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7949) );
  OR2_X1 U9520 ( .A1(n8162), .A2(n7949), .ZN(n7954) );
  INV_X1 U9521 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8572) );
  OR2_X1 U9522 ( .A1(n8083), .A2(n8572), .ZN(n7953) );
  NAND2_X1 U9523 ( .A1(n7950), .A2(n8949), .ZN(n7951) );
  NAND2_X1 U9524 ( .A1(n7980), .A2(n7951), .ZN(n9187) );
  OR2_X1 U9525 ( .A1(n6634), .A2(n9187), .ZN(n7952) );
  NOR2_X1 U9526 ( .A1(n8862), .A2(n6602), .ZN(n7956) );
  XNOR2_X1 U9527 ( .A(n7957), .B(n7956), .ZN(n8824) );
  NAND2_X1 U9528 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U9529 ( .A1(n7959), .A2(n8153), .ZN(n7961) );
  AOI22_X1 U9530 ( .A1(n7974), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7973), .B2(
        n10182), .ZN(n7960) );
  XNOR2_X1 U9531 ( .A(n9278), .B(n8116), .ZN(n7970) );
  INV_X1 U9532 ( .A(n6634), .ZN(n8099) );
  XNOR2_X1 U9533 ( .A(n7980), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U9534 ( .A1(n8099), .A2(n9162), .ZN(n7967) );
  INV_X1 U9535 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8969) );
  OR2_X1 U9536 ( .A1(n8162), .A2(n8969), .ZN(n7966) );
  INV_X1 U9537 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7962) );
  OR2_X1 U9538 ( .A1(n8083), .A2(n7962), .ZN(n7965) );
  INV_X1 U9539 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n7963) );
  OR2_X1 U9540 ( .A1(n8121), .A2(n7963), .ZN(n7964) );
  NAND4_X1 U9541 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n9153)
         );
  NAND2_X1 U9542 ( .A1(n9153), .A2(n8176), .ZN(n7968) );
  XNOR2_X1 U9543 ( .A(n7970), .B(n7968), .ZN(n8859) );
  INV_X1 U9544 ( .A(n7968), .ZN(n7969) );
  AND2_X1 U9545 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  NAND2_X1 U9546 ( .A1(n7972), .A2(n8153), .ZN(n7976) );
  AOI22_X1 U9547 ( .A1(n7974), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9188), .B2(
        n7973), .ZN(n7975) );
  XNOR2_X1 U9548 ( .A(n9273), .B(n8094), .ZN(n7986) );
  NAND2_X1 U9549 ( .A1(n8046), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7985) );
  INV_X1 U9550 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n7977) );
  OR2_X1 U9551 ( .A1(n8083), .A2(n7977), .ZN(n7984) );
  INV_X1 U9552 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7979) );
  INV_X1 U9553 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7978) );
  OAI21_X1 U9554 ( .B1(n7980), .B2(n7979), .A(n7978), .ZN(n7981) );
  NAND2_X1 U9555 ( .A1(n7981), .A2(n7995), .ZN(n9147) );
  OR2_X1 U9556 ( .A1(n6634), .A2(n9147), .ZN(n7983) );
  INV_X1 U9557 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8759) );
  OR2_X1 U9558 ( .A1(n8121), .A2(n8759), .ZN(n7982) );
  NAND4_X1 U9559 ( .A1(n7985), .A2(n7984), .A3(n7983), .A4(n7982), .ZN(n9168)
         );
  NAND2_X1 U9560 ( .A1(n9168), .A2(n8176), .ZN(n7987) );
  NAND2_X1 U9561 ( .A1(n7986), .A2(n7987), .ZN(n7991) );
  INV_X1 U9562 ( .A(n7986), .ZN(n7989) );
  INV_X1 U9563 ( .A(n7987), .ZN(n7988) );
  NAND2_X1 U9564 ( .A1(n7989), .A2(n7988), .ZN(n7990) );
  NAND2_X1 U9565 ( .A1(n7992), .A2(n8153), .ZN(n7994) );
  OR2_X1 U9566 ( .A1(n8167), .A2(n8364), .ZN(n7993) );
  XNOR2_X1 U9567 ( .A(n9267), .B(n8116), .ZN(n8004) );
  NAND2_X1 U9568 ( .A1(n7995), .A2(n8844), .ZN(n7996) );
  NAND2_X1 U9569 ( .A1(n8009), .A2(n7996), .ZN(n9135) );
  OR2_X1 U9570 ( .A1(n9135), .A2(n6634), .ZN(n8002) );
  INV_X1 U9571 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9136) );
  OR2_X1 U9572 ( .A1(n8083), .A2(n9136), .ZN(n8001) );
  INV_X1 U9573 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n7997) );
  OR2_X1 U9574 ( .A1(n8121), .A2(n7997), .ZN(n8000) );
  INV_X1 U9575 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7998) );
  OR2_X1 U9576 ( .A1(n8162), .A2(n7998), .ZN(n7999) );
  NOR2_X1 U9577 ( .A1(n8790), .A2(n6602), .ZN(n8003) );
  XNOR2_X1 U9578 ( .A(n8004), .B(n8003), .ZN(n8842) );
  NAND2_X1 U9579 ( .A1(n8005), .A2(n8153), .ZN(n8008) );
  OR2_X1 U9580 ( .A1(n8167), .A2(n8006), .ZN(n8007) );
  XNOR2_X1 U9581 ( .A(n9118), .B(n8094), .ZN(n8019) );
  NAND2_X1 U9582 ( .A1(n8009), .A2(n8800), .ZN(n8010) );
  NAND2_X1 U9583 ( .A1(n8025), .A2(n8010), .ZN(n9123) );
  INV_X1 U9584 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8011) );
  OR2_X1 U9585 ( .A1(n8162), .A2(n8011), .ZN(n8013) );
  INV_X1 U9586 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9117) );
  OR2_X1 U9587 ( .A1(n8083), .A2(n9117), .ZN(n8012) );
  AND2_X1 U9588 ( .A1(n8013), .A2(n8012), .ZN(n8016) );
  INV_X1 U9589 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8014) );
  OR2_X1 U9590 ( .A1(n6615), .A2(n8014), .ZN(n8015) );
  OAI211_X1 U9591 ( .C1(n9123), .C2(n6634), .A(n8016), .B(n8015), .ZN(n9131)
         );
  NAND2_X1 U9592 ( .A1(n9131), .A2(n8176), .ZN(n8017) );
  XNOR2_X1 U9593 ( .A(n8019), .B(n8017), .ZN(n8798) );
  INV_X1 U9594 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U9595 ( .A1(n8020), .A2(n8153), .ZN(n8023) );
  OR2_X1 U9596 ( .A1(n8167), .A2(n8021), .ZN(n8022) );
  XNOR2_X1 U9597 ( .A(n9255), .B(n8094), .ZN(n8031) );
  NAND2_X1 U9598 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  AND2_X1 U9599 ( .A1(n8027), .A2(n8026), .ZN(n9099) );
  NAND2_X1 U9600 ( .A1(n9099), .A2(n8099), .ZN(n8030) );
  AOI22_X1 U9601 ( .A1(n8157), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8158), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n8029) );
  INV_X1 U9602 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8579) );
  OR2_X1 U9603 ( .A1(n8162), .A2(n8579), .ZN(n8028) );
  OR2_X1 U9604 ( .A1(n9094), .A2(n6602), .ZN(n8852) );
  INV_X1 U9605 ( .A(n8031), .ZN(n8032) );
  NAND2_X1 U9606 ( .A1(n8035), .A2(n8153), .ZN(n8038) );
  OR2_X1 U9607 ( .A1(n8167), .A2(n8036), .ZN(n8037) );
  XNOR2_X1 U9608 ( .A(n9252), .B(n8094), .ZN(n8055) );
  INV_X1 U9609 ( .A(n8055), .ZN(n8039) );
  NAND2_X1 U9610 ( .A1(n8040), .A2(n8153), .ZN(n8043) );
  OR2_X1 U9611 ( .A1(n8167), .A2(n8041), .ZN(n8042) );
  XNOR2_X1 U9612 ( .A(n9247), .B(n8094), .ZN(n8833) );
  INV_X1 U9613 ( .A(n8833), .ZN(n8057) );
  INV_X1 U9614 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8836) );
  OR2_X2 U9615 ( .A1(n8044), .A2(n8836), .ZN(n8067) );
  NAND2_X1 U9616 ( .A1(n8044), .A2(n8836), .ZN(n8045) );
  AND2_X1 U9617 ( .A1(n8067), .A2(n8045), .ZN(n9072) );
  NAND2_X1 U9618 ( .A1(n9072), .A2(n8099), .ZN(n8052) );
  INV_X1 U9619 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9620 ( .A1(n8046), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8048) );
  INV_X1 U9621 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8705) );
  OR2_X1 U9622 ( .A1(n8121), .A2(n8705), .ZN(n8047) );
  OAI211_X1 U9623 ( .C1(n8083), .C2(n8049), .A(n8048), .B(n8047), .ZN(n8050)
         );
  INV_X1 U9624 ( .A(n8050), .ZN(n8051) );
  NOR2_X1 U9625 ( .A1(n9108), .A2(n6602), .ZN(n8831) );
  NOR2_X1 U9626 ( .A1(n8056), .A2(n8055), .ZN(n8830) );
  NAND2_X1 U9627 ( .A1(n9057), .A2(n8176), .ZN(n8832) );
  NAND2_X1 U9628 ( .A1(n8833), .A2(n8832), .ZN(n8059) );
  INV_X1 U9629 ( .A(n8832), .ZN(n8058) );
  AOI22_X1 U9630 ( .A1(n8830), .A2(n8059), .B1(n8058), .B2(n8057), .ZN(n8060)
         );
  OR2_X1 U9631 ( .A1(n8167), .A2(n8444), .ZN(n8063) );
  XNOR2_X1 U9632 ( .A(n9242), .B(n8116), .ZN(n8808) );
  INV_X1 U9633 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U9634 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9635 ( .A1(n8080), .A2(n8068), .ZN(n9051) );
  OR2_X1 U9636 ( .A1(n9051), .A2(n6634), .ZN(n8073) );
  INV_X1 U9637 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8736) );
  INV_X1 U9638 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8686) );
  OR2_X1 U9639 ( .A1(n8121), .A2(n8686), .ZN(n8070) );
  INV_X1 U9640 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9050) );
  OR2_X1 U9641 ( .A1(n8083), .A2(n9050), .ZN(n8069) );
  OAI211_X1 U9642 ( .C1(n8162), .C2(n8736), .A(n8070), .B(n8069), .ZN(n8071)
         );
  INV_X1 U9643 ( .A(n8071), .ZN(n8072) );
  INV_X1 U9644 ( .A(n9069), .ZN(n8897) );
  NAND2_X1 U9645 ( .A1(n8897), .A2(n8176), .ZN(n8807) );
  INV_X1 U9646 ( .A(n8808), .ZN(n8074) );
  OR2_X1 U9647 ( .A1(n8167), .A2(n8076), .ZN(n8077) );
  XNOR2_X1 U9648 ( .A(n9237), .B(n8094), .ZN(n8088) );
  INV_X1 U9649 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U9650 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  INV_X1 U9651 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U9652 ( .A1(n8158), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8085) );
  INV_X1 U9653 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8082) );
  OR2_X1 U9654 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  OAI211_X1 U9655 ( .C1(n8162), .C2(n8634), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI21_X2 U9656 ( .B1(n9038), .B2(n8099), .A(n8086), .ZN(n9021) );
  OR2_X1 U9657 ( .A1(n9021), .A2(n6602), .ZN(n8087) );
  AOI21_X1 U9658 ( .B1(n8088), .B2(n8087), .A(n8089), .ZN(n8869) );
  INV_X1 U9659 ( .A(n8089), .ZN(n8090) );
  NAND2_X1 U9660 ( .A1(n8091), .A2(n8153), .ZN(n8093) );
  OR2_X1 U9661 ( .A1(n8167), .A2(n8689), .ZN(n8092) );
  XNOR2_X1 U9662 ( .A(n9230), .B(n8094), .ZN(n8101) );
  XNOR2_X1 U9663 ( .A(n8106), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9014) );
  INV_X1 U9664 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U9665 ( .A1(n8157), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9666 ( .A1(n8158), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8095) );
  OAI211_X1 U9667 ( .C1(n8097), .C2(n8162), .A(n8096), .B(n8095), .ZN(n8098)
         );
  OR2_X1 U9668 ( .A1(n9036), .A2(n6602), .ZN(n8100) );
  NOR2_X1 U9669 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  AOI21_X1 U9670 ( .B1(n8101), .B2(n8100), .A(n8102), .ZN(n8419) );
  OR2_X1 U9671 ( .A1(n8167), .A2(n8417), .ZN(n8103) );
  INV_X1 U9672 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8421) );
  INV_X1 U9673 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8105) );
  OAI21_X1 U9674 ( .B1(n8106), .B2(n8421), .A(n8105), .ZN(n8109) );
  INV_X1 U9675 ( .A(n8106), .ZN(n8108) );
  AND2_X1 U9676 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8107) );
  NAND2_X1 U9677 ( .A1(n8108), .A2(n8107), .ZN(n8402) );
  NAND2_X1 U9678 ( .A1(n8109), .A2(n8402), .ZN(n8120) );
  OR2_X1 U9679 ( .A1(n8120), .A2(n6634), .ZN(n8115) );
  INV_X1 U9680 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U9681 ( .A1(n8157), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U9682 ( .A1(n8158), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8110) );
  OAI211_X1 U9683 ( .C1(n8162), .C2(n8112), .A(n8111), .B(n8110), .ZN(n8113)
         );
  INV_X1 U9684 ( .A(n8113), .ZN(n8114) );
  INV_X1 U9685 ( .A(n9022), .ZN(n8896) );
  NAND2_X1 U9686 ( .A1(n8896), .A2(n8176), .ZN(n8117) );
  XNOR2_X1 U9687 ( .A(n8117), .B(n8116), .ZN(n8118) );
  XNOR2_X1 U9688 ( .A(n9226), .B(n8118), .ZN(n8119) );
  INV_X1 U9689 ( .A(n8120), .ZN(n8997) );
  AOI22_X1 U9690 ( .A1(n8997), .A2(n8871), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8128) );
  OR2_X1 U9691 ( .A1(n8402), .A2(n6634), .ZN(n8126) );
  INV_X1 U9692 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U9693 ( .A1(n8157), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8123) );
  INV_X1 U9694 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8718) );
  OR2_X1 U9695 ( .A1(n8121), .A2(n8718), .ZN(n8122) );
  OAI211_X1 U9696 ( .C1(n8162), .C2(n8669), .A(n8123), .B(n8122), .ZN(n8124)
         );
  INV_X1 U9697 ( .A(n8124), .ZN(n8125) );
  NAND2_X1 U9698 ( .A1(n8126), .A2(n8125), .ZN(n9002) );
  NAND2_X1 U9699 ( .A1(n9002), .A2(n8875), .ZN(n8127) );
  OAI211_X1 U9700 ( .C1(n9036), .C2(n8873), .A(n8128), .B(n8127), .ZN(n8129)
         );
  AOI21_X1 U9701 ( .B1(n9226), .B2(n8848), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9702 ( .B1(n8131), .B2(n8866), .A(n8130), .ZN(P2_U3222) );
  NAND2_X1 U9703 ( .A1(n9773), .A2(n9770), .ZN(n8134) );
  NAND2_X1 U9704 ( .A1(n9482), .A2(n8132), .ZN(n9903) );
  NOR2_X1 U9705 ( .A1(n10078), .A2(n9903), .ZN(n9555) );
  AOI21_X1 U9706 ( .B1(n10078), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9555), .ZN(
        n8133) );
  OAI211_X1 U9707 ( .C1(n9775), .C2(n9766), .A(n8134), .B(n8133), .ZN(P1_U3261) );
  INV_X1 U9708 ( .A(n8287), .ZN(n8135) );
  OAI21_X2 U9709 ( .B1(n8136), .B2(n8135), .A(n8286), .ZN(n9194) );
  NAND2_X1 U9710 ( .A1(n9194), .A2(n8290), .ZN(n8137) );
  NAND2_X1 U9711 ( .A1(n9287), .A2(n9181), .ZN(n8289) );
  NAND2_X1 U9712 ( .A1(n8137), .A2(n8289), .ZN(n9178) );
  XNOR2_X1 U9713 ( .A(n9284), .B(n8862), .ZN(n9177) );
  OR2_X1 U9714 ( .A1(n9284), .A2(n8862), .ZN(n8295) );
  INV_X1 U9715 ( .A(n9153), .ZN(n9183) );
  OR2_X1 U9716 ( .A1(n9278), .A2(n9183), .ZN(n8298) );
  NAND2_X1 U9717 ( .A1(n9278), .A2(n9183), .ZN(n8304) );
  INV_X1 U9718 ( .A(n9168), .ZN(n8392) );
  OR2_X1 U9719 ( .A1(n9273), .A2(n8392), .ZN(n8306) );
  NAND2_X1 U9720 ( .A1(n9273), .A2(n8392), .ZN(n9128) );
  NAND2_X1 U9721 ( .A1(n9151), .A2(n9152), .ZN(n9127) );
  NAND2_X1 U9722 ( .A1(n9267), .A2(n8790), .ZN(n8308) );
  NAND2_X1 U9723 ( .A1(n8310), .A2(n8308), .ZN(n9133) );
  INV_X1 U9724 ( .A(n9128), .ZN(n8138) );
  NOR2_X1 U9725 ( .A1(n9133), .A2(n8138), .ZN(n8139) );
  NAND2_X1 U9726 ( .A1(n9127), .A2(n8139), .ZN(n8140) );
  INV_X1 U9727 ( .A(n9131), .ZN(n9107) );
  OR2_X1 U9728 ( .A1(n9260), .A2(n9107), .ZN(n8309) );
  NAND2_X1 U9729 ( .A1(n9260), .A2(n9107), .ZN(n9103) );
  NAND2_X1 U9730 ( .A1(n8309), .A2(n9103), .ZN(n9121) );
  NAND2_X1 U9731 ( .A1(n9255), .A2(n9094), .ZN(n8311) );
  INV_X1 U9732 ( .A(n9103), .ZN(n8143) );
  NOR2_X1 U9733 ( .A1(n9106), .A2(n8143), .ZN(n8144) );
  NAND2_X1 U9734 ( .A1(n9252), .A2(n9108), .ZN(n9065) );
  INV_X1 U9735 ( .A(n9089), .ZN(n8145) );
  NOR2_X1 U9736 ( .A1(n9079), .A2(n8145), .ZN(n8146) );
  NAND2_X1 U9737 ( .A1(n9247), .A2(n9093), .ZN(n8318) );
  INV_X1 U9738 ( .A(n9065), .ZN(n8147) );
  NOR2_X1 U9739 ( .A1(n9066), .A2(n8147), .ZN(n8148) );
  NAND2_X1 U9740 ( .A1(n9064), .A2(n8148), .ZN(n8149) );
  NAND2_X1 U9741 ( .A1(n9242), .A2(n9069), .ZN(n8204) );
  NAND2_X1 U9742 ( .A1(n8206), .A2(n8204), .ZN(n9045) );
  NAND2_X1 U9743 ( .A1(n9230), .A2(n9036), .ZN(n8327) );
  INV_X1 U9744 ( .A(n9019), .ZN(n8151) );
  NOR2_X1 U9745 ( .A1(n9008), .A2(n8151), .ZN(n8152) );
  NAND2_X2 U9746 ( .A1(n9017), .A2(n8152), .ZN(n9024) );
  NAND2_X1 U9747 ( .A1(n9329), .A2(n8153), .ZN(n8155) );
  INV_X1 U9748 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9331) );
  OR2_X1 U9749 ( .A1(n8167), .A2(n9331), .ZN(n8154) );
  INV_X1 U9750 ( .A(n8407), .ZN(n8198) );
  INV_X1 U9751 ( .A(n9002), .ZN(n8332) );
  INV_X1 U9752 ( .A(n8163), .ZN(n8165) );
  INV_X1 U9753 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8381) );
  NOR2_X1 U9754 ( .A1(n8167), .A2(n8381), .ZN(n8156) );
  INV_X1 U9755 ( .A(n8987), .ZN(n9894) );
  INV_X1 U9756 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U9757 ( .A1(n8157), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U9758 ( .A1(n8158), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8159) );
  OAI211_X1 U9759 ( .C1(n8162), .C2(n8161), .A(n8160), .B(n8159), .ZN(n8895)
         );
  AND2_X1 U9760 ( .A1(n8987), .A2(n8895), .ZN(n8199) );
  OAI21_X1 U9761 ( .B1(n8165), .B2(n9894), .A(n8164), .ZN(n8173) );
  NAND2_X1 U9762 ( .A1(n9323), .A2(n8153), .ZN(n8169) );
  OR2_X1 U9763 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  INV_X1 U9764 ( .A(n8982), .ZN(n8172) );
  INV_X1 U9765 ( .A(n8895), .ZN(n8170) );
  NAND2_X1 U9766 ( .A1(n9894), .A2(n8170), .ZN(n8171) );
  INV_X1 U9767 ( .A(n9133), .ZN(n9129) );
  INV_X1 U9768 ( .A(n9166), .ZN(n8193) );
  INV_X1 U9769 ( .A(n9202), .ZN(n8192) );
  NOR4_X1 U9770 ( .A1(n8181), .A2(n8180), .A3(n10204), .A4(n8179), .ZN(n8183)
         );
  NAND4_X1 U9771 ( .A1(n8183), .A2(n8246), .A3(n8259), .A4(n8182), .ZN(n8187)
         );
  INV_X1 U9772 ( .A(n8184), .ZN(n8186) );
  NOR4_X1 U9773 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(n8189)
         );
  NAND4_X1 U9774 ( .A1(n8280), .A2(n8274), .A3(n8190), .A4(n8189), .ZN(n8191)
         );
  NOR4_X1 U9775 ( .A1(n8193), .A2(n8192), .A3(n8281), .A4(n8191), .ZN(n8194)
         );
  INV_X1 U9776 ( .A(n9177), .ZN(n8292) );
  NAND4_X1 U9777 ( .A1(n9129), .A2(n9152), .A3(n8194), .A4(n8292), .ZN(n8195)
         );
  NOR4_X1 U9778 ( .A1(n9079), .A2(n9106), .A3(n9121), .A4(n8195), .ZN(n8196)
         );
  NAND4_X1 U9779 ( .A1(n8150), .A2(n9055), .A3(n8397), .A4(n8196), .ZN(n8197)
         );
  NOR4_X1 U9780 ( .A1(n8198), .A2(n9001), .A3(n9008), .A4(n8197), .ZN(n8201)
         );
  INV_X1 U9781 ( .A(n8199), .ZN(n8340) );
  NAND4_X1 U9782 ( .A1(n8337), .A2(n8201), .A3(n8340), .A4(n8344), .ZN(n8202)
         );
  XNOR2_X1 U9783 ( .A(n8202), .B(n9188), .ZN(n8350) );
  NOR2_X2 U9784 ( .A1(n8203), .A2(n8357), .ZN(n8331) );
  INV_X1 U9785 ( .A(n8331), .ZN(n8343) );
  INV_X1 U9786 ( .A(n8204), .ZN(n8205) );
  OR2_X1 U9787 ( .A1(n9034), .A2(n8205), .ZN(n8208) );
  NAND2_X1 U9788 ( .A1(n8322), .A2(n8206), .ZN(n8207) );
  MUX2_X1 U9789 ( .A(n8208), .B(n8207), .S(n8331), .Z(n8325) );
  AND2_X1 U9790 ( .A1(n8211), .A2(n8262), .ZN(n8209) );
  MUX2_X1 U9791 ( .A(n8250), .B(n8209), .S(n8343), .Z(n8210) );
  AND2_X1 U9792 ( .A1(n8210), .A2(n8254), .ZN(n8252) );
  INV_X1 U9793 ( .A(n8252), .ZN(n8261) );
  OAI211_X1 U9794 ( .C1(n8261), .C2(n8212), .A(n8264), .B(n8211), .ZN(n8257)
         );
  NAND2_X1 U9795 ( .A1(n8240), .A2(n8242), .ZN(n8214) );
  NAND2_X1 U9796 ( .A1(n8216), .A2(n8217), .ZN(n8213) );
  MUX2_X1 U9797 ( .A(n8214), .B(n8213), .S(n8331), .Z(n8244) );
  AND2_X1 U9798 ( .A1(n8216), .A2(n8215), .ZN(n8218) );
  OAI211_X1 U9799 ( .C1(n8244), .C2(n8218), .A(n8217), .B(n8247), .ZN(n8219)
         );
  NAND2_X1 U9800 ( .A1(n8219), .A2(n8343), .ZN(n8228) );
  INV_X1 U9801 ( .A(n8244), .ZN(n8226) );
  AND2_X1 U9802 ( .A1(n8231), .A2(n8220), .ZN(n8221) );
  OAI211_X1 U9803 ( .C1(n8222), .C2(n8221), .A(n8235), .B(n7006), .ZN(n8223)
         );
  NAND3_X1 U9804 ( .A1(n8223), .A2(n8234), .A3(n8343), .ZN(n8224) );
  NAND3_X1 U9805 ( .A1(n8226), .A2(n8225), .A3(n8224), .ZN(n8227) );
  OR2_X1 U9806 ( .A1(n8230), .A2(n8229), .ZN(n8241) );
  NAND2_X1 U9807 ( .A1(n7006), .A2(n8231), .ZN(n8232) );
  NAND3_X1 U9808 ( .A1(n8234), .A2(n8233), .A3(n8232), .ZN(n8236) );
  NAND3_X1 U9809 ( .A1(n8236), .A2(n8331), .A3(n8235), .ZN(n8237) );
  NAND2_X1 U9810 ( .A1(n8910), .A2(n8238), .ZN(n8239) );
  AND2_X1 U9811 ( .A1(n8240), .A2(n8239), .ZN(n8243) );
  OAI211_X1 U9812 ( .C1(n8244), .C2(n8243), .A(n8242), .B(n8241), .ZN(n8245)
         );
  NAND3_X1 U9813 ( .A1(n8260), .A2(n8259), .A3(n8248), .ZN(n8251) );
  NAND3_X1 U9814 ( .A1(n8251), .A2(n8250), .A3(n8249), .ZN(n8253) );
  NAND2_X1 U9815 ( .A1(n8253), .A2(n8252), .ZN(n8255) );
  NAND3_X1 U9816 ( .A1(n8255), .A2(n8265), .A3(n8254), .ZN(n8256) );
  MUX2_X1 U9817 ( .A(n8257), .B(n8256), .S(n8343), .Z(n8271) );
  NAND4_X1 U9818 ( .A1(n8260), .A2(n8259), .A3(n8331), .A4(n8258), .ZN(n8263)
         );
  AOI21_X1 U9819 ( .B1(n8263), .B2(n8262), .A(n8261), .ZN(n8270) );
  NAND2_X1 U9820 ( .A1(n8272), .A2(n8264), .ZN(n8267) );
  NAND2_X1 U9821 ( .A1(n8273), .A2(n8265), .ZN(n8266) );
  MUX2_X1 U9822 ( .A(n8267), .B(n8266), .S(n8331), .Z(n8268) );
  INV_X1 U9823 ( .A(n8268), .ZN(n8269) );
  OAI21_X1 U9824 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8276) );
  MUX2_X1 U9825 ( .A(n8273), .B(n8272), .S(n8331), .Z(n8275) );
  MUX2_X1 U9826 ( .A(n8278), .B(n8277), .S(n8331), .Z(n8279) );
  INV_X1 U9827 ( .A(n8281), .ZN(n8285) );
  MUX2_X1 U9828 ( .A(n8283), .B(n8282), .S(n8331), .Z(n8284) );
  MUX2_X1 U9829 ( .A(n8287), .B(n8286), .S(n8331), .Z(n8288) );
  MUX2_X1 U9830 ( .A(n8290), .B(n8289), .S(n8343), .Z(n8291) );
  NAND2_X1 U9831 ( .A1(n9284), .A2(n8862), .ZN(n8293) );
  AND2_X1 U9832 ( .A1(n8304), .A2(n8293), .ZN(n8294) );
  MUX2_X1 U9833 ( .A(n8295), .B(n8294), .S(n8331), .Z(n8296) );
  NAND3_X1 U9834 ( .A1(n8297), .A2(n8296), .A3(n8298), .ZN(n8305) );
  NAND3_X1 U9835 ( .A1(n8305), .A2(n8298), .A3(n8306), .ZN(n8299) );
  NAND2_X1 U9836 ( .A1(n8299), .A2(n9128), .ZN(n8300) );
  NAND2_X1 U9837 ( .A1(n8300), .A2(n8310), .ZN(n8301) );
  NAND3_X1 U9838 ( .A1(n8301), .A2(n8308), .A3(n9103), .ZN(n8302) );
  NAND3_X1 U9839 ( .A1(n8302), .A2(n8331), .A3(n8309), .ZN(n8303) );
  MUX2_X1 U9840 ( .A(n8331), .B(n8303), .S(n9089), .Z(n8314) );
  NAND2_X1 U9841 ( .A1(n8305), .A2(n8304), .ZN(n8307) );
  MUX2_X1 U9842 ( .A(n8312), .B(n8311), .S(n8331), .Z(n8313) );
  NAND3_X1 U9843 ( .A1(n5027), .A2(n8314), .A3(n8313), .ZN(n8317) );
  MUX2_X1 U9844 ( .A(n9065), .B(n8315), .S(n8331), .Z(n8316) );
  NAND3_X1 U9845 ( .A1(n8397), .A2(n8317), .A3(n8316), .ZN(n8321) );
  MUX2_X1 U9846 ( .A(n8319), .B(n8318), .S(n4630), .Z(n8320) );
  AND3_X1 U9847 ( .A1(n9055), .A2(n8321), .A3(n8320), .ZN(n8324) );
  INV_X1 U9848 ( .A(n9008), .ZN(n9018) );
  MUX2_X1 U9849 ( .A(n9019), .B(n8322), .S(n8343), .Z(n8323) );
  AOI21_X1 U9850 ( .B1(n8329), .B2(n8327), .A(n8331), .ZN(n8328) );
  OAI21_X1 U9851 ( .B1(n8331), .B2(n8330), .A(n8407), .ZN(n8336) );
  NAND2_X1 U9852 ( .A1(n9002), .A2(n8331), .ZN(n8334) );
  NAND2_X1 U9853 ( .A1(n8332), .A2(n8343), .ZN(n8333) );
  MUX2_X1 U9854 ( .A(n8334), .B(n8333), .S(n9220), .Z(n8335) );
  INV_X1 U9855 ( .A(n8337), .ZN(n8338) );
  MUX2_X1 U9856 ( .A(n8339), .B(n8343), .S(n8338), .Z(n8347) );
  NAND2_X1 U9857 ( .A1(n8344), .A2(n8340), .ZN(n8342) );
  NAND3_X1 U9858 ( .A1(n8342), .A2(n8341), .A3(n8343), .ZN(n8346) );
  NOR2_X1 U9859 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  AOI21_X1 U9860 ( .B1(n8351), .B2(n8353), .A(n8352), .ZN(n8348) );
  AOI211_X1 U9861 ( .C1(n8354), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8355)
         );
  NOR4_X1 U9862 ( .A1(n8356), .A2(n10212), .A3(n9182), .A4(n8408), .ZN(n8359)
         );
  OAI21_X1 U9863 ( .B1(n8360), .B2(n8357), .A(P2_B_REG_SCAN_IN), .ZN(n8358) );
  INV_X1 U9864 ( .A(n8361), .ZN(n8416) );
  OAI222_X1 U9865 ( .A1(n9881), .A2(n8416), .B1(n5922), .B2(P1_U3084), .C1(
        n8362), .C2(n8383), .ZN(P1_U3325) );
  OAI222_X1 U9866 ( .A1(n9330), .A2(n8364), .B1(n4490), .B2(n8363), .C1(n6549), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NOR2_X1 U9867 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6557), .ZN(n8369) );
  AOI211_X1 U9868 ( .C1(n8367), .C2(n8366), .A(n8365), .B(n10171), .ZN(n8368)
         );
  AOI211_X1 U9869 ( .C1(n10187), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n8369), .B(
        n8368), .ZN(n8375) );
  AND2_X1 U9870 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8373) );
  MUX2_X1 U9871 ( .A(n8370), .B(P2_REG2_REG_1__SCAN_IN), .S(n8376), .Z(n8372)
         );
  OAI211_X1 U9872 ( .C1(n8373), .C2(n8372), .A(n10185), .B(n8371), .ZN(n8374)
         );
  OAI211_X1 U9873 ( .C1(n10170), .C2(n8376), .A(n8375), .B(n8374), .ZN(
        P2_U3246) );
  OAI222_X1 U9874 ( .A1(n8383), .A2(n8379), .B1(n9881), .B2(n8378), .C1(
        P1_U3084), .C2(n8377), .ZN(P1_U3331) );
  INV_X1 U9875 ( .A(n8380), .ZN(n8386) );
  OAI222_X1 U9876 ( .A1(n8382), .A2(P2_U3152), .B1(n4490), .B2(n8386), .C1(
        n8381), .C2(n9330), .ZN(P2_U3328) );
  INV_X1 U9877 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8384) );
  OAI222_X1 U9878 ( .A1(n9881), .A2(n8386), .B1(n8385), .B2(P1_U3084), .C1(
        n8384), .C2(n8383), .ZN(P1_U3323) );
  INV_X1 U9879 ( .A(n9267), .ZN(n9138) );
  INV_X1 U9880 ( .A(n9273), .ZN(n9150) );
  INV_X1 U9881 ( .A(n9284), .ZN(n8390) );
  INV_X1 U9882 ( .A(n8862), .ZN(n9198) );
  NAND2_X1 U9883 ( .A1(n8390), .A2(n8862), .ZN(n8391) );
  NAND2_X1 U9884 ( .A1(n9174), .A2(n8391), .ZN(n9159) );
  OAI21_X1 U9885 ( .B1(n9138), .B2(n8790), .A(n9265), .ZN(n9114) );
  NAND2_X1 U9886 ( .A1(n9118), .A2(n9107), .ZN(n8393) );
  INV_X1 U9887 ( .A(n9255), .ZN(n9101) );
  INV_X1 U9888 ( .A(n9108), .ZN(n8395) );
  OAI22_X1 U9889 ( .A1(n9063), .A2(n8397), .B1(n9247), .B2(n9057), .ZN(n9046)
         );
  NAND2_X1 U9890 ( .A1(n9046), .A2(n9045), .ZN(n9044) );
  NAND2_X1 U9891 ( .A1(n9044), .A2(n8398), .ZN(n9030) );
  NAND2_X1 U9892 ( .A1(n9030), .A2(n9034), .ZN(n9029) );
  INV_X1 U9893 ( .A(n9021), .ZN(n9058) );
  NAND2_X1 U9894 ( .A1(n8878), .A2(n9021), .ZN(n8399) );
  NAND2_X1 U9895 ( .A1(n9029), .A2(n8399), .ZN(n9009) );
  NAND2_X1 U9896 ( .A1(n9009), .A2(n9008), .ZN(n9007) );
  INV_X1 U9897 ( .A(n9036), .ZN(n9003) );
  NAND2_X1 U9898 ( .A1(n9016), .A2(n9036), .ZN(n8400) );
  NAND2_X1 U9899 ( .A1(n9007), .A2(n8400), .ZN(n8993) );
  NAND2_X1 U9900 ( .A1(n8993), .A2(n9001), .ZN(n8992) );
  OAI21_X1 U9901 ( .B1(n8896), .B2(n9226), .A(n8992), .ZN(n8401) );
  INV_X1 U9902 ( .A(n9287), .ZN(n9207) );
  NAND2_X1 U9903 ( .A1(n9146), .A2(n9138), .ZN(n9140) );
  INV_X1 U9904 ( .A(n9247), .ZN(n9075) );
  INV_X1 U9905 ( .A(n9230), .ZN(n9016) );
  NAND2_X1 U9906 ( .A1(n9037), .A2(n9016), .ZN(n9011) );
  AOI21_X1 U9907 ( .B1(n9220), .B2(n8995), .A(n8986), .ZN(n9221) );
  INV_X1 U9908 ( .A(n9220), .ZN(n8405) );
  INV_X1 U9909 ( .A(n8402), .ZN(n8403) );
  AOI22_X1 U9910 ( .A1(n8403), .A2(n9161), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10210), .ZN(n8404) );
  OAI21_X1 U9911 ( .B1(n8405), .B2(n9164), .A(n8404), .ZN(n8414) );
  XNOR2_X1 U9912 ( .A(n8406), .B(n8407), .ZN(n8412) );
  INV_X1 U9913 ( .A(n8408), .ZN(n8409) );
  AOI21_X1 U9914 ( .B1(n8409), .B2(P2_B_REG_SCAN_IN), .A(n9184), .ZN(n8981) );
  AOI22_X1 U9915 ( .A1(n8896), .A2(n9195), .B1(n8981), .B2(n8895), .ZN(n8410)
         );
  INV_X1 U9916 ( .A(n8410), .ZN(n8411) );
  NOR2_X1 U9917 ( .A1(n9223), .A2(n10210), .ZN(n8413) );
  AOI211_X1 U9918 ( .C1(n9221), .C2(n9211), .A(n8414), .B(n8413), .ZN(n8415)
         );
  OAI21_X1 U9919 ( .B1(n9224), .B2(n9214), .A(n8415), .ZN(P2_U3267) );
  OAI222_X1 U9920 ( .A1(n9330), .A2(n8417), .B1(n4490), .B2(n8416), .C1(n6411), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  OAI211_X1 U9921 ( .C1(n8420), .C2(n8419), .A(n8418), .B(n8882), .ZN(n8425)
         );
  OAI22_X1 U9922 ( .A1(n9021), .A2(n8873), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8421), .ZN(n8423) );
  NOR2_X1 U9923 ( .A1(n9022), .A2(n8887), .ZN(n8422) );
  AOI211_X1 U9924 ( .C1(n8871), .C2(n9014), .A(n8423), .B(n8422), .ZN(n8424)
         );
  OAI211_X1 U9925 ( .C1(n9016), .C2(n8893), .A(n8425), .B(n8424), .ZN(P2_U3216) );
  XNOR2_X1 U9926 ( .A(n8426), .B(n8831), .ZN(n8431) );
  NAND2_X1 U9927 ( .A1(n9057), .A2(n8875), .ZN(n8428) );
  AOI22_X1 U9928 ( .A1(n8394), .A2(n8890), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8427) );
  OAI211_X1 U9929 ( .C1(n8885), .C2(n9085), .A(n8428), .B(n8427), .ZN(n8429)
         );
  AOI21_X1 U9930 ( .B1(n9252), .B2(n8848), .A(n8429), .ZN(n8430) );
  OAI21_X1 U9931 ( .B1(n8431), .B2(n8866), .A(n8430), .ZN(P2_U3218) );
  AOI22_X1 U9932 ( .A1(n6557), .A2(keyinput141), .B1(n8433), .B2(keyinput207), 
        .ZN(n8432) );
  OAI221_X1 U9933 ( .B1(n6557), .B2(keyinput141), .C1(n8433), .C2(keyinput207), 
        .A(n8432), .ZN(n8441) );
  INV_X1 U9934 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U9935 ( .A1(n10217), .A2(keyinput163), .B1(n8705), .B2(keyinput164), 
        .ZN(n8434) );
  OAI221_X1 U9936 ( .B1(n10217), .B2(keyinput163), .C1(n8705), .C2(keyinput164), .A(n8434), .ZN(n8440) );
  AOI22_X1 U9937 ( .A1(n6856), .A2(keyinput159), .B1(n8436), .B2(keyinput152), 
        .ZN(n8435) );
  OAI221_X1 U9938 ( .B1(n6856), .B2(keyinput159), .C1(n8436), .C2(keyinput152), 
        .A(n8435), .ZN(n8439) );
  AOI22_X1 U9939 ( .A1(n6261), .A2(keyinput145), .B1(keyinput169), .B2(n8844), 
        .ZN(n8437) );
  OAI221_X1 U9940 ( .B1(n6261), .B2(keyinput145), .C1(n8844), .C2(keyinput169), 
        .A(n8437), .ZN(n8438) );
  NOR4_X1 U9941 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(n8459)
         );
  AOI22_X1 U9942 ( .A1(n10218), .A2(keyinput184), .B1(n8634), .B2(keyinput234), 
        .ZN(n8442) );
  OAI221_X1 U9943 ( .B1(n10218), .B2(keyinput184), .C1(n8634), .C2(keyinput234), .A(n8442), .ZN(n8448) );
  INV_X1 U9944 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U9945 ( .A1(n10153), .A2(keyinput224), .B1(n8444), .B2(keyinput221), 
        .ZN(n8443) );
  OAI221_X1 U9946 ( .B1(n10153), .B2(keyinput224), .C1(n8444), .C2(keyinput221), .A(n8443), .ZN(n8447) );
  AOI22_X1 U9947 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput188), .B1(
        P1_D_REG_27__SCAN_IN), .B2(keyinput251), .ZN(n8445) );
  OAI221_X1 U9948 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput188), .C1(
        P1_D_REG_27__SCAN_IN), .C2(keyinput251), .A(n8445), .ZN(n8446) );
  NOR3_X1 U9949 ( .A1(n8448), .A2(n8447), .A3(n8446), .ZN(n8458) );
  AOI22_X1 U9950 ( .A1(n10220), .A2(keyinput228), .B1(n8450), .B2(keyinput255), 
        .ZN(n8449) );
  OAI221_X1 U9951 ( .B1(n10220), .B2(keyinput228), .C1(n8450), .C2(keyinput255), .A(n8449), .ZN(n8456) );
  AOI22_X1 U9952 ( .A1(n8662), .A2(keyinput134), .B1(keyinput196), .B2(n8759), 
        .ZN(n8451) );
  OAI221_X1 U9953 ( .B1(n8662), .B2(keyinput134), .C1(n8759), .C2(keyinput196), 
        .A(n8451), .ZN(n8455) );
  AOI22_X1 U9954 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput175), .B1(n8453), 
        .B2(keyinput130), .ZN(n8452) );
  OAI221_X1 U9955 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput175), .C1(n8453), 
        .C2(keyinput130), .A(n8452), .ZN(n8454) );
  NOR3_X1 U9956 ( .A1(n8456), .A2(n8455), .A3(n8454), .ZN(n8457) );
  NAND3_X1 U9957 ( .A1(n8459), .A2(n8458), .A3(n8457), .ZN(n8538) );
  INV_X1 U9958 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10085) );
  INV_X1 U9959 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8648) );
  AOI22_X1 U9960 ( .A1(n10085), .A2(keyinput242), .B1(keyinput227), .B2(n8648), 
        .ZN(n8460) );
  OAI221_X1 U9961 ( .B1(n10085), .B2(keyinput242), .C1(n8648), .C2(keyinput227), .A(n8460), .ZN(n8473) );
  AOI22_X1 U9962 ( .A1(n5274), .A2(keyinput214), .B1(keyinput190), .B2(n8836), 
        .ZN(n8461) );
  OAI221_X1 U9963 ( .B1(n5274), .B2(keyinput214), .C1(n8836), .C2(keyinput190), 
        .A(n8461), .ZN(n8472) );
  XOR2_X1 U9964 ( .A(n5321), .B(keyinput240), .Z(n8465) );
  XNOR2_X1 U9965 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput246), .ZN(n8464) );
  XNOR2_X1 U9966 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput247), .ZN(n8463) );
  NAND3_X1 U9967 ( .A1(n8465), .A2(n8464), .A3(n8463), .ZN(n8471) );
  XNOR2_X1 U9968 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput208), .ZN(n8469) );
  XNOR2_X1 U9969 ( .A(SI_0_), .B(keyinput183), .ZN(n8468) );
  XNOR2_X1 U9970 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput158), .ZN(n8467) );
  XNOR2_X1 U9971 ( .A(SI_3_), .B(keyinput151), .ZN(n8466) );
  NAND4_X1 U9972 ( .A1(n8469), .A2(n8468), .A3(n8467), .A4(n8466), .ZN(n8470)
         );
  NOR4_X1 U9973 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n8489)
         );
  INV_X1 U9974 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10213) );
  XOR2_X1 U9975 ( .A(keyinput155), .B(n10213), .Z(n8488) );
  XOR2_X1 U9976 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput135), .Z(n8479) );
  XNOR2_X1 U9977 ( .A(n8474), .B(keyinput162), .ZN(n8478) );
  XNOR2_X1 U9978 ( .A(n8475), .B(keyinput173), .ZN(n8477) );
  XNOR2_X1 U9979 ( .A(n8670), .B(keyinput167), .ZN(n8476) );
  NOR4_X1 U9980 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n8487)
         );
  XOR2_X1 U9981 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput206), .Z(n8485) );
  XNOR2_X1 U9982 ( .A(n8480), .B(keyinput140), .ZN(n8484) );
  XNOR2_X1 U9983 ( .A(n8481), .B(keyinput132), .ZN(n8483) );
  XNOR2_X1 U9984 ( .A(keyinput187), .B(n7187), .ZN(n8482) );
  NOR4_X1 U9985 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n8486)
         );
  NAND4_X1 U9986 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n8537)
         );
  AOI22_X1 U9987 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput154), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(keyinput209), .ZN(n8490) );
  OAI221_X1 U9988 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput154), .C1(
        P1_DATAO_REG_17__SCAN_IN), .C2(keyinput209), .A(n8490), .ZN(n8497) );
  AOI22_X1 U9989 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput223), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(keyinput198), .ZN(n8491) );
  OAI221_X1 U9990 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput223), .C1(
        P1_REG3_REG_18__SCAN_IN), .C2(keyinput198), .A(n8491), .ZN(n8496) );
  AOI22_X1 U9991 ( .A1(P1_REG2_REG_30__SCAN_IN), .A2(keyinput129), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput171), .ZN(n8492) );
  OAI221_X1 U9992 ( .B1(P1_REG2_REG_30__SCAN_IN), .B2(keyinput129), .C1(
        P1_REG1_REG_24__SCAN_IN), .C2(keyinput171), .A(n8492), .ZN(n8495) );
  AOI22_X1 U9993 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput147), .B1(
        P1_REG1_REG_17__SCAN_IN), .B2(keyinput168), .ZN(n8493) );
  OAI221_X1 U9994 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput147), .C1(
        P1_REG1_REG_17__SCAN_IN), .C2(keyinput168), .A(n8493), .ZN(n8494) );
  NOR4_X1 U9995 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n8525)
         );
  AOI22_X1 U9996 ( .A1(P2_REG0_REG_21__SCAN_IN), .A2(keyinput241), .B1(
        P2_REG1_REG_29__SCAN_IN), .B2(keyinput211), .ZN(n8498) );
  OAI221_X1 U9997 ( .B1(P2_REG0_REG_21__SCAN_IN), .B2(keyinput241), .C1(
        P2_REG1_REG_29__SCAN_IN), .C2(keyinput211), .A(n8498), .ZN(n8505) );
  AOI22_X1 U9998 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput244), .B1(
        P2_REG2_REG_24__SCAN_IN), .B2(keyinput231), .ZN(n8499) );
  OAI221_X1 U9999 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput244), .C1(
        P2_REG2_REG_24__SCAN_IN), .C2(keyinput231), .A(n8499), .ZN(n8504) );
  AOI22_X1 U10000 ( .A1(P2_D_REG_20__SCAN_IN), .A2(keyinput153), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(keyinput215), .ZN(n8500) );
  OAI221_X1 U10001 ( .B1(P2_D_REG_20__SCAN_IN), .B2(keyinput153), .C1(
        P1_DATAO_REG_1__SCAN_IN), .C2(keyinput215), .A(n8500), .ZN(n8503) );
  AOI22_X1 U10002 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput180), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput156), .ZN(n8501) );
  OAI221_X1 U10003 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput180), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput156), .A(n8501), .ZN(n8502) );
  NOR4_X1 U10004 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n8524)
         );
  AOI22_X1 U10005 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput137), .B1(
        P1_REG1_REG_12__SCAN_IN), .B2(keyinput212), .ZN(n8506) );
  OAI221_X1 U10006 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput137), .C1(
        P1_REG1_REG_12__SCAN_IN), .C2(keyinput212), .A(n8506), .ZN(n8513) );
  AOI22_X1 U10007 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput174), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput254), .ZN(n8507) );
  OAI221_X1 U10008 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput174), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput254), .A(n8507), .ZN(n8512) );
  AOI22_X1 U10009 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput136), .B1(
        P2_REG2_REG_26__SCAN_IN), .B2(keyinput191), .ZN(n8508) );
  OAI221_X1 U10010 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput136), .C1(
        P2_REG2_REG_26__SCAN_IN), .C2(keyinput191), .A(n8508), .ZN(n8511) );
  AOI22_X1 U10011 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput197), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput222), .ZN(n8509) );
  OAI221_X1 U10012 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput197), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput222), .A(n8509), .ZN(n8510) );
  NOR4_X1 U10013 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n8523)
         );
  AOI22_X1 U10014 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput230), .B1(
        P1_REG1_REG_21__SCAN_IN), .B2(keyinput203), .ZN(n8514) );
  OAI221_X1 U10015 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput230), .C1(
        P1_REG1_REG_21__SCAN_IN), .C2(keyinput203), .A(n8514), .ZN(n8521) );
  AOI22_X1 U10016 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(keyinput250), .B1(
        P2_ADDR_REG_9__SCAN_IN), .B2(keyinput128), .ZN(n8515) );
  OAI221_X1 U10017 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(keyinput250), .C1(
        P2_ADDR_REG_9__SCAN_IN), .C2(keyinput128), .A(n8515), .ZN(n8520) );
  AOI22_X1 U10018 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(keyinput245), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput172), .ZN(n8516) );
  OAI221_X1 U10019 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(keyinput245), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput172), .A(n8516), .ZN(n8519) );
  AOI22_X1 U10020 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput237), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput200), .ZN(n8517) );
  OAI221_X1 U10021 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput237), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput200), .A(n8517), .ZN(n8518) );
  NOR4_X1 U10022 ( .A1(n8521), .A2(n8520), .A3(n8519), .A4(n8518), .ZN(n8522)
         );
  NAND4_X1 U10023 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n8536)
         );
  INV_X1 U10024 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10083) );
  INV_X1 U10025 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10026 ( .A1(n10083), .A2(keyinput189), .B1(keyinput170), .B2(n9928), .ZN(n8526) );
  OAI221_X1 U10027 ( .B1(n10083), .B2(keyinput189), .C1(n9928), .C2(
        keyinput170), .A(n8526), .ZN(n8534) );
  AOI22_X1 U10028 ( .A1(n8664), .A2(keyinput161), .B1(keyinput192), .B2(n8764), 
        .ZN(n8527) );
  OAI221_X1 U10029 ( .B1(n8664), .B2(keyinput161), .C1(n8764), .C2(keyinput192), .A(n8527), .ZN(n8533) );
  AOI22_X1 U10030 ( .A1(n8529), .A2(keyinput131), .B1(keyinput225), .B2(n7826), 
        .ZN(n8528) );
  OAI221_X1 U10031 ( .B1(n8529), .B2(keyinput131), .C1(n7826), .C2(keyinput225), .A(n8528), .ZN(n8532) );
  AOI22_X1 U10032 ( .A1(n8751), .A2(keyinput226), .B1(keyinput182), .B2(n5296), 
        .ZN(n8530) );
  OAI221_X1 U10033 ( .B1(n8751), .B2(keyinput226), .C1(n5296), .C2(keyinput182), .A(n8530), .ZN(n8531) );
  OR4_X1 U10034 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n8535)
         );
  NOR4_X1 U10035 ( .A1(n8538), .A2(n8537), .A3(n8536), .A4(n8535), .ZN(n8566)
         );
  AOI22_X1 U10036 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(keyinput253), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput219), .ZN(n8539) );
  OAI221_X1 U10037 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(keyinput253), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput219), .A(n8539), .ZN(n8546) );
  AOI22_X1 U10038 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput210), .B1(
        P1_REG2_REG_25__SCAN_IN), .B2(keyinput165), .ZN(n8540) );
  OAI221_X1 U10039 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput210), .C1(
        P1_REG2_REG_25__SCAN_IN), .C2(keyinput165), .A(n8540), .ZN(n8545) );
  AOI22_X1 U10040 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(keyinput233), .B1(
        P2_REG1_REG_12__SCAN_IN), .B2(keyinput243), .ZN(n8541) );
  OAI221_X1 U10041 ( .B1(P2_REG0_REG_4__SCAN_IN), .B2(keyinput233), .C1(
        P2_REG1_REG_12__SCAN_IN), .C2(keyinput243), .A(n8541), .ZN(n8544) );
  AOI22_X1 U10042 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(keyinput235), .B1(
        P1_REG1_REG_4__SCAN_IN), .B2(keyinput229), .ZN(n8542) );
  OAI221_X1 U10043 ( .B1(P2_IR_REG_5__SCAN_IN), .B2(keyinput235), .C1(
        P1_REG1_REG_4__SCAN_IN), .C2(keyinput229), .A(n8542), .ZN(n8543) );
  NOR4_X1 U10044 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(n8565)
         );
  AOI22_X1 U10045 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput252), .B1(
        P2_IR_REG_27__SCAN_IN), .B2(keyinput248), .ZN(n8547) );
  OAI221_X1 U10046 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput252), .C1(
        P2_IR_REG_27__SCAN_IN), .C2(keyinput248), .A(n8547), .ZN(n8554) );
  AOI22_X1 U10047 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(keyinput249), .B1(
        P1_REG3_REG_21__SCAN_IN), .B2(keyinput195), .ZN(n8548) );
  OAI221_X1 U10048 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(keyinput249), .C1(
        P1_REG3_REG_21__SCAN_IN), .C2(keyinput195), .A(n8548), .ZN(n8553) );
  AOI22_X1 U10049 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput178), .B1(
        P1_REG1_REG_23__SCAN_IN), .B2(keyinput181), .ZN(n8549) );
  OAI221_X1 U10050 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput178), .C1(
        P1_REG1_REG_23__SCAN_IN), .C2(keyinput181), .A(n8549), .ZN(n8552) );
  AOI22_X1 U10051 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput216), .B1(
        P1_REG3_REG_10__SCAN_IN), .B2(keyinput139), .ZN(n8550) );
  OAI221_X1 U10052 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput216), .C1(
        P1_REG3_REG_10__SCAN_IN), .C2(keyinput139), .A(n8550), .ZN(n8551) );
  NOR4_X1 U10053 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(n8564)
         );
  AOI22_X1 U10054 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput193), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput238), .ZN(n8555) );
  OAI221_X1 U10055 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput193), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput238), .A(n8555), .ZN(n8562) );
  AOI22_X1 U10056 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput157), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput146), .ZN(n8556) );
  OAI221_X1 U10057 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput157), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput146), .A(n8556), .ZN(n8561) );
  AOI22_X1 U10058 ( .A1(P2_D_REG_27__SCAN_IN), .A2(keyinput213), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput232), .ZN(n8557) );
  OAI221_X1 U10059 ( .B1(P2_D_REG_27__SCAN_IN), .B2(keyinput213), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput232), .A(n8557), .ZN(n8560) );
  AOI22_X1 U10060 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(keyinput144), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput143), .ZN(n8558) );
  OAI221_X1 U10061 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(keyinput144), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput143), .A(n8558), .ZN(n8559) );
  NOR4_X1 U10062 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n8563)
         );
  NAND4_X1 U10063 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n8786)
         );
  INV_X1 U10064 ( .A(SI_18_), .ZN(n8568) );
  AOI22_X1 U10065 ( .A1(n9889), .A2(keyinput177), .B1(n8568), .B2(keyinput138), 
        .ZN(n8567) );
  OAI221_X1 U10066 ( .B1(n9889), .B2(keyinput177), .C1(n8568), .C2(keyinput138), .A(n8567), .ZN(n8576) );
  INV_X1 U10067 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10030) );
  AOI22_X1 U10068 ( .A1(n8712), .A2(keyinput179), .B1(keyinput176), .B2(n10030), .ZN(n8569) );
  OAI221_X1 U10069 ( .B1(n8712), .B2(keyinput179), .C1(n10030), .C2(
        keyinput176), .A(n8569), .ZN(n8575) );
  AOI22_X1 U10070 ( .A1(n5437), .A2(keyinput166), .B1(keyinput194), .B2(n10329), .ZN(n8570) );
  OAI221_X1 U10071 ( .B1(n5437), .B2(keyinput166), .C1(n10329), .C2(
        keyinput194), .A(n8570), .ZN(n8574) );
  AOI22_X1 U10072 ( .A1(n8770), .A2(keyinput205), .B1(keyinput201), .B2(n8572), 
        .ZN(n8571) );
  OAI221_X1 U10073 ( .B1(n8770), .B2(keyinput205), .C1(n8572), .C2(keyinput201), .A(n8571), .ZN(n8573) );
  NOR4_X1 U10074 ( .A1(n8576), .A2(n8575), .A3(n8574), .A4(n8573), .ZN(n8600)
         );
  AOI22_X1 U10075 ( .A1(n8689), .A2(keyinput199), .B1(keyinput185), .B2(n9331), 
        .ZN(n8577) );
  OAI221_X1 U10076 ( .B1(n8689), .B2(keyinput199), .C1(n9331), .C2(keyinput185), .A(n8577), .ZN(n8586) );
  AOI22_X1 U10077 ( .A1(n8579), .A2(keyinput142), .B1(keyinput186), .B2(n6934), 
        .ZN(n8578) );
  OAI221_X1 U10078 ( .B1(n8579), .B2(keyinput142), .C1(n6934), .C2(keyinput186), .A(n8578), .ZN(n8585) );
  INV_X1 U10079 ( .A(SI_6_), .ZN(n8752) );
  AOI22_X1 U10080 ( .A1(n8581), .A2(keyinput204), .B1(n8752), .B2(keyinput133), 
        .ZN(n8580) );
  OAI221_X1 U10081 ( .B1(n8581), .B2(keyinput204), .C1(n8752), .C2(keyinput133), .A(n8580), .ZN(n8584) );
  AOI22_X1 U10082 ( .A1(P1_U3084), .A2(keyinput220), .B1(keyinput202), .B2(
        n8718), .ZN(n8582) );
  OAI221_X1 U10083 ( .B1(P1_U3084), .B2(keyinput220), .C1(n8718), .C2(
        keyinput202), .A(n8582), .ZN(n8583) );
  NOR4_X1 U10084 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n8599)
         );
  AOI22_X1 U10085 ( .A1(n8588), .A2(keyinput160), .B1(keyinput239), .B2(n8636), 
        .ZN(n8587) );
  OAI221_X1 U10086 ( .B1(n8588), .B2(keyinput160), .C1(n8636), .C2(keyinput239), .A(n8587), .ZN(n8597) );
  INV_X1 U10087 ( .A(SI_30_), .ZN(n8590) );
  AOI22_X1 U10088 ( .A1(n5453), .A2(keyinput217), .B1(keyinput148), .B2(n8590), 
        .ZN(n8589) );
  OAI221_X1 U10089 ( .B1(n5453), .B2(keyinput217), .C1(n8590), .C2(keyinput148), .A(n8589), .ZN(n8596) );
  AOI22_X1 U10090 ( .A1(n7265), .A2(keyinput150), .B1(n8592), .B2(keyinput236), 
        .ZN(n8591) );
  OAI221_X1 U10091 ( .B1(n7265), .B2(keyinput150), .C1(n8592), .C2(keyinput236), .A(n8591), .ZN(n8595) );
  AOI22_X1 U10092 ( .A1(n7686), .A2(keyinput218), .B1(n10077), .B2(keyinput149), .ZN(n8593) );
  OAI221_X1 U10093 ( .B1(n7686), .B2(keyinput218), .C1(n10077), .C2(
        keyinput149), .A(n8593), .ZN(n8594) );
  NOR4_X1 U10094 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n8598)
         );
  NAND3_X1 U10095 ( .A1(n8600), .A2(n8599), .A3(n8598), .ZN(n8785) );
  OAI22_X1 U10096 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput46), .B1(
        keyinput0), .B2(P2_ADDR_REG_9__SCAN_IN), .ZN(n8601) );
  AOI221_X1 U10097 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput46), .C1(
        P2_ADDR_REG_9__SCAN_IN), .C2(keyinput0), .A(n8601), .ZN(n8608) );
  OAI22_X1 U10098 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(keyinput45), .B1(
        keyinput94), .B2(P1_REG2_REG_1__SCAN_IN), .ZN(n8602) );
  AOI221_X1 U10099 ( .B1(P1_DATAO_REG_12__SCAN_IN), .B2(keyinput45), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput94), .A(n8602), .ZN(n8607) );
  OAI22_X1 U10100 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(keyinput14), .B1(
        keyinput113), .B2(P2_REG0_REG_21__SCAN_IN), .ZN(n8603) );
  AOI221_X1 U10101 ( .B1(P2_REG1_REG_22__SCAN_IN), .B2(keyinput14), .C1(
        P2_REG0_REG_21__SCAN_IN), .C2(keyinput113), .A(n8603), .ZN(n8606) );
  OAI22_X1 U10102 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(keyinput12), .B1(
        P2_REG1_REG_23__SCAN_IN), .B2(keyinput116), .ZN(n8604) );
  AOI221_X1 U10103 ( .B1(P1_DATAO_REG_0__SCAN_IN), .B2(keyinput12), .C1(
        keyinput116), .C2(P2_REG1_REG_23__SCAN_IN), .A(n8604), .ZN(n8605) );
  NAND4_X1 U10104 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n8660)
         );
  OAI22_X1 U10105 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput112), .B1(
        P2_IR_REG_5__SCAN_IN), .B2(keyinput107), .ZN(n8609) );
  AOI221_X1 U10106 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput112), .C1(
        keyinput107), .C2(P2_IR_REG_5__SCAN_IN), .A(n8609), .ZN(n8616) );
  OAI22_X1 U10107 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput114), .B1(
        keyinput104), .B2(P2_STATE_REG_SCAN_IN), .ZN(n8610) );
  AOI221_X1 U10108 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput114), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput104), .A(n8610), .ZN(n8615) );
  OAI22_X1 U10109 ( .A1(SI_18_), .A2(keyinput10), .B1(P1_DATAO_REG_1__SCAN_IN), 
        .B2(keyinput87), .ZN(n8611) );
  AOI221_X1 U10110 ( .B1(SI_18_), .B2(keyinput10), .C1(keyinput87), .C2(
        P1_DATAO_REG_1__SCAN_IN), .A(n8611), .ZN(n8614) );
  OAI22_X1 U10111 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(keyinput40), .B1(
        keyinput29), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n8612) );
  AOI221_X1 U10112 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(keyinput40), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput29), .A(n8612), .ZN(n8613) );
  NAND4_X1 U10113 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n8659)
         );
  AOI22_X1 U10114 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput17), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput44), .ZN(n8617) );
  OAI221_X1 U10115 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput17), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput44), .A(n8617), .ZN(n8624) );
  AOI22_X1 U10116 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput103), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput91), .ZN(n8618) );
  OAI221_X1 U10117 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput103), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput91), .A(n8618), .ZN(n8623) );
  AOI22_X1 U10118 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput65), .B1(SI_30_), 
        .B2(keyinput20), .ZN(n8619) );
  OAI221_X1 U10119 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput65), .C1(SI_30_), 
        .C2(keyinput20), .A(n8619), .ZN(n8622) );
  AOI22_X1 U10120 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(keyinput79), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(keyinput24), .ZN(n8620) );
  OAI221_X1 U10121 ( .B1(P1_REG0_REG_18__SCAN_IN), .B2(keyinput79), .C1(
        P1_DATAO_REG_14__SCAN_IN), .C2(keyinput24), .A(n8620), .ZN(n8621) );
  NOR4_X1 U10122 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n8657)
         );
  AOI22_X1 U10123 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput9), .B1(
        P1_REG2_REG_16__SCAN_IN), .B2(keyinput38), .ZN(n8625) );
  OAI221_X1 U10124 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput9), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(keyinput38), .A(n8625), .ZN(n8632) );
  AOI22_X1 U10125 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(keyinput122), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput30), .ZN(n8626) );
  OAI221_X1 U10126 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(keyinput122), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput30), .A(n8626), .ZN(n8631) );
  AOI22_X1 U10127 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(keyinput59), .B1(
        P2_REG2_REG_12__SCAN_IN), .B2(keyinput90), .ZN(n8627) );
  OAI221_X1 U10128 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(keyinput59), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput90), .A(n8627), .ZN(n8630) );
  AOI22_X1 U10129 ( .A1(SI_29_), .A2(keyinput86), .B1(P2_IR_REG_14__SCAN_IN), 
        .B2(keyinput108), .ZN(n8628) );
  OAI221_X1 U10130 ( .B1(SI_29_), .B2(keyinput86), .C1(P2_IR_REG_14__SCAN_IN), 
        .C2(keyinput108), .A(n8628), .ZN(n8629) );
  NOR4_X1 U10131 ( .A1(n8632), .A2(n8631), .A3(n8630), .A4(n8629), .ZN(n8656)
         );
  AOI22_X1 U10132 ( .A1(n7756), .A2(keyinput19), .B1(n8634), .B2(keyinput106), 
        .ZN(n8633) );
  OAI221_X1 U10133 ( .B1(n7756), .B2(keyinput19), .C1(n8634), .C2(keyinput106), 
        .A(n8633), .ZN(n8640) );
  AOI22_X1 U10134 ( .A1(n8637), .A2(keyinput70), .B1(keyinput111), .B2(n8636), 
        .ZN(n8635) );
  OAI221_X1 U10135 ( .B1(n8637), .B2(keyinput70), .C1(n8636), .C2(keyinput111), 
        .A(n8635), .ZN(n8639) );
  XOR2_X1 U10136 ( .A(SI_0_), .B(keyinput55), .Z(n8638) );
  OR3_X1 U10137 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8644) );
  AOI22_X1 U10138 ( .A1(n9084), .A2(keyinput8), .B1(keyinput115), .B2(n7476), 
        .ZN(n8641) );
  OAI221_X1 U10139 ( .B1(n9084), .B2(keyinput8), .C1(n7476), .C2(keyinput115), 
        .A(n8641), .ZN(n8643) );
  XNOR2_X1 U10140 ( .A(n10030), .B(keyinput48), .ZN(n8642) );
  NOR3_X1 U10141 ( .A1(n8644), .A2(n8643), .A3(n8642), .ZN(n8655) );
  AOI22_X1 U10142 ( .A1(P1_REG2_REG_30__SCAN_IN), .A2(keyinput1), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput76), .ZN(n8645) );
  OAI221_X1 U10143 ( .B1(P1_REG2_REG_30__SCAN_IN), .B2(keyinput1), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput76), .A(n8645), .ZN(n8653) );
  AOI22_X1 U10144 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput124), .B1(
        P1_REG2_REG_5__SCAN_IN), .B2(keyinput127), .ZN(n8646) );
  OAI221_X1 U10145 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput124), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(keyinput127), .A(n8646), .ZN(n8652) );
  AOI22_X1 U10146 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput109), .B1(n8648), 
        .B2(keyinput99), .ZN(n8647) );
  OAI221_X1 U10147 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput109), .C1(n8648), 
        .C2(keyinput99), .A(n8647), .ZN(n8651) );
  AOI22_X1 U10148 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(keyinput37), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput93), .ZN(n8649) );
  OAI221_X1 U10149 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(keyinput37), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput93), .A(n8649), .ZN(n8650) );
  NOR4_X1 U10150 ( .A1(n8653), .A2(n8652), .A3(n8651), .A4(n8650), .ZN(n8654)
         );
  NAND4_X1 U10151 ( .A1(n8657), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n8658)
         );
  NOR3_X1 U10152 ( .A1(n8660), .A2(n8659), .A3(n8658), .ZN(n8784) );
  AOI22_X1 U10153 ( .A1(n9050), .A2(keyinput95), .B1(n8662), .B2(keyinput6), 
        .ZN(n8661) );
  OAI221_X1 U10154 ( .B1(n9050), .B2(keyinput95), .C1(n8662), .C2(keyinput6), 
        .A(n8661), .ZN(n8674) );
  AOI22_X1 U10155 ( .A1(n8665), .A2(keyinput69), .B1(n8664), .B2(keyinput33), 
        .ZN(n8663) );
  OAI221_X1 U10156 ( .B1(n8665), .B2(keyinput69), .C1(n8664), .C2(keyinput33), 
        .A(n8663), .ZN(n8673) );
  AOI22_X1 U10157 ( .A1(n8667), .A2(keyinput81), .B1(keyinput105), .B2(n6652), 
        .ZN(n8666) );
  OAI221_X1 U10158 ( .B1(n8667), .B2(keyinput81), .C1(n6652), .C2(keyinput105), 
        .A(n8666), .ZN(n8672) );
  AOI22_X1 U10159 ( .A1(n8670), .A2(keyinput39), .B1(keyinput83), .B2(n8669), 
        .ZN(n8668) );
  OAI221_X1 U10160 ( .B1(n8670), .B2(keyinput39), .C1(n8669), .C2(keyinput83), 
        .A(n8668), .ZN(n8671) );
  NOR4_X1 U10161 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n8684)
         );
  AOI22_X1 U10162 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput73), .B1(
        P2_REG2_REG_26__SCAN_IN), .B2(keyinput63), .ZN(n8675) );
  OAI221_X1 U10163 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput73), .C1(
        P2_REG2_REG_26__SCAN_IN), .C2(keyinput63), .A(n8675), .ZN(n8682) );
  AOI22_X1 U10164 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(keyinput49), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(keyinput15), .ZN(n8676) );
  OAI221_X1 U10165 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(keyinput49), .C1(
        P1_REG3_REG_11__SCAN_IN), .C2(keyinput15), .A(n8676), .ZN(n8681) );
  AOI22_X1 U10166 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(keyinput32), .B1(
        P1_D_REG_14__SCAN_IN), .B2(keyinput61), .ZN(n8677) );
  OAI221_X1 U10167 ( .B1(P1_REG3_REG_8__SCAN_IN), .B2(keyinput32), .C1(
        P1_D_REG_14__SCAN_IN), .C2(keyinput61), .A(n8677), .ZN(n8680) );
  AOI22_X1 U10168 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput2), .B1(
        P1_REG1_REG_15__SCAN_IN), .B2(keyinput3), .ZN(n8678) );
  OAI221_X1 U10169 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput2), .C1(
        P1_REG1_REG_15__SCAN_IN), .C2(keyinput3), .A(n8678), .ZN(n8679) );
  NOR4_X1 U10170 ( .A1(n8682), .A2(n8681), .A3(n8680), .A4(n8679), .ZN(n8683)
         );
  AND2_X1 U10171 ( .A1(n8684), .A2(n8683), .ZN(n8782) );
  AOI22_X1 U10172 ( .A1(n10213), .A2(keyinput27), .B1(n8686), .B2(keyinput50), 
        .ZN(n8685) );
  OAI221_X1 U10173 ( .B1(n10213), .B2(keyinput27), .C1(n8686), .C2(keyinput50), 
        .A(n8685), .ZN(n8695) );
  AOI22_X1 U10174 ( .A1(P1_U3084), .A2(keyinput92), .B1(keyinput88), .B2(n6456), .ZN(n8687) );
  OAI221_X1 U10175 ( .B1(P1_U3084), .B2(keyinput92), .C1(n6456), .C2(
        keyinput88), .A(n8687), .ZN(n8694) );
  AOI22_X1 U10176 ( .A1(n8689), .A2(keyinput71), .B1(keyinput60), .B2(n5592), 
        .ZN(n8688) );
  OAI221_X1 U10177 ( .B1(n8689), .B2(keyinput71), .C1(n5592), .C2(keyinput60), 
        .A(n8688), .ZN(n8693) );
  AOI22_X1 U10178 ( .A1(n10217), .A2(keyinput35), .B1(keyinput52), .B2(n8691), 
        .ZN(n8690) );
  OAI221_X1 U10179 ( .B1(n10217), .B2(keyinput35), .C1(n8691), .C2(keyinput52), 
        .A(n8690), .ZN(n8692) );
  NOR4_X1 U10180 ( .A1(n8695), .A2(n8694), .A3(n8693), .A4(n8692), .ZN(n8781)
         );
  AOI22_X1 U10181 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput62), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput18), .ZN(n8696) );
  OAI221_X1 U10182 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput62), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput18), .A(n8696), .ZN(n8703) );
  AOI22_X1 U10183 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput13), .B1(
        P2_REG2_REG_6__SCAN_IN), .B2(keyinput121), .ZN(n8697) );
  OAI221_X1 U10184 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput13), .C1(
        P2_REG2_REG_6__SCAN_IN), .C2(keyinput121), .A(n8697), .ZN(n8702) );
  AOI22_X1 U10185 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput26), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput28), .ZN(n8698) );
  OAI221_X1 U10186 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput26), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput28), .A(n8698), .ZN(n8701) );
  AOI22_X1 U10187 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput78), .B1(
        P1_REG1_REG_2__SCAN_IN), .B2(keyinput96), .ZN(n8699) );
  OAI221_X1 U10188 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput78), .C1(
        P1_REG1_REG_2__SCAN_IN), .C2(keyinput96), .A(n8699), .ZN(n8700) );
  NOR4_X1 U10189 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n8780)
         );
  INV_X1 U10190 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U10191 ( .A1(n8705), .A2(keyinput36), .B1(n10084), .B2(keyinput126), 
        .ZN(n8704) );
  OAI221_X1 U10192 ( .B1(n8705), .B2(keyinput36), .C1(n10084), .C2(keyinput126), .A(n8704), .ZN(n8709) );
  INV_X1 U10193 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8707) );
  AOI22_X1 U10194 ( .A1(n7265), .A2(keyinput22), .B1(n8707), .B2(keyinput53), 
        .ZN(n8706) );
  OAI221_X1 U10195 ( .B1(n7265), .B2(keyinput22), .C1(n8707), .C2(keyinput53), 
        .A(n8706), .ZN(n8708) );
  NOR2_X1 U10196 ( .A1(n8709), .A2(n8708), .ZN(n8716) );
  AOI22_X1 U10197 ( .A1(n10216), .A2(keyinput25), .B1(n9117), .B2(keyinput110), 
        .ZN(n8710) );
  OAI221_X1 U10198 ( .B1(n10216), .B2(keyinput25), .C1(n9117), .C2(keyinput110), .A(n8710), .ZN(n8714) );
  AOI22_X1 U10199 ( .A1(n6856), .A2(keyinput31), .B1(n8712), .B2(keyinput51), 
        .ZN(n8711) );
  OAI221_X1 U10200 ( .B1(n6856), .B2(keyinput31), .C1(n8712), .C2(keyinput51), 
        .A(n8711), .ZN(n8713) );
  NOR2_X1 U10201 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  AND2_X1 U10202 ( .A1(n8716), .A2(n8715), .ZN(n8747) );
  AOI22_X1 U10203 ( .A1(n8718), .A2(keyinput74), .B1(keyinput66), .B2(n10329), 
        .ZN(n8717) );
  OAI221_X1 U10204 ( .B1(n8718), .B2(keyinput74), .C1(n10329), .C2(keyinput66), 
        .A(n8717), .ZN(n8723) );
  INV_X1 U10205 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U10206 ( .A1(n10082), .A2(keyinput123), .B1(keyinput21), .B2(n10077), .ZN(n8719) );
  OAI221_X1 U10207 ( .B1(n10082), .B2(keyinput123), .C1(n10077), .C2(
        keyinput21), .A(n8719), .ZN(n8722) );
  INV_X1 U10208 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U10209 ( .A1(n10081), .A2(keyinput72), .B1(keyinput41), .B2(n8844), 
        .ZN(n8720) );
  OAI221_X1 U10210 ( .B1(n10081), .B2(keyinput72), .C1(n8844), .C2(keyinput41), 
        .A(n8720), .ZN(n8721) );
  NOR3_X1 U10211 ( .A1(n8723), .A2(n8722), .A3(n8721), .ZN(n8746) );
  XNOR2_X1 U10212 ( .A(n9928), .B(keyinput42), .ZN(n8734) );
  XNOR2_X1 U10213 ( .A(SI_3_), .B(keyinput23), .ZN(n8727) );
  XNOR2_X1 U10214 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput120), .ZN(n8726) );
  XNOR2_X1 U10215 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput11), .ZN(n8725) );
  XNOR2_X1 U10216 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput80), .ZN(n8724) );
  NAND4_X1 U10217 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n8733)
         );
  XNOR2_X1 U10218 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput7), .ZN(n8731) );
  XNOR2_X1 U10219 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput100), .ZN(n8730) );
  XNOR2_X1 U10220 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput118), .ZN(n8729) );
  XNOR2_X1 U10221 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput4), .ZN(n8728) );
  NAND4_X1 U10222 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n8732)
         );
  NOR3_X1 U10223 ( .A1(n8734), .A2(n8733), .A3(n8732), .ZN(n8745) );
  AOI22_X1 U10224 ( .A1(n6278), .A2(keyinput84), .B1(keyinput82), .B2(n8736), 
        .ZN(n8735) );
  OAI221_X1 U10225 ( .B1(n6278), .B2(keyinput84), .C1(n8736), .C2(keyinput82), 
        .A(n8735), .ZN(n8743) );
  XNOR2_X1 U10226 ( .A(n10215), .B(keyinput102), .ZN(n8742) );
  XNOR2_X1 U10227 ( .A(P1_REG1_REG_21__SCAN_IN), .B(keyinput75), .ZN(n8740) );
  XNOR2_X1 U10228 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput119), .ZN(n8739) );
  XNOR2_X1 U10229 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput34), .ZN(n8738) );
  XNOR2_X1 U10230 ( .A(keyinput117), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8737)
         );
  NAND4_X1 U10231 ( .A1(n8740), .A2(n8739), .A3(n8738), .A4(n8737), .ZN(n8741)
         );
  NOR3_X1 U10232 ( .A1(n8743), .A2(n8742), .A3(n8741), .ZN(n8744) );
  NAND4_X1 U10233 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n8778)
         );
  INV_X1 U10234 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8749) );
  AOI22_X1 U10235 ( .A1(n8749), .A2(keyinput43), .B1(n5296), .B2(keyinput54), 
        .ZN(n8748) );
  OAI221_X1 U10236 ( .B1(n8749), .B2(keyinput43), .C1(n5296), .C2(keyinput54), 
        .A(n8748), .ZN(n8757) );
  AOI22_X1 U10237 ( .A1(n8752), .A2(keyinput5), .B1(n8751), .B2(keyinput98), 
        .ZN(n8750) );
  OAI221_X1 U10238 ( .B1(n8752), .B2(keyinput5), .C1(n8751), .C2(keyinput98), 
        .A(n8750), .ZN(n8756) );
  XNOR2_X1 U10239 ( .A(keyinput125), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n8754) );
  XNOR2_X1 U10240 ( .A(keyinput16), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U10241 ( .A1(n8754), .A2(n8753), .ZN(n8755) );
  NOR3_X1 U10242 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(n8776) );
  AOI22_X1 U10243 ( .A1(n8759), .A2(keyinput68), .B1(keyinput56), .B2(n10218), 
        .ZN(n8758) );
  OAI221_X1 U10244 ( .B1(n8759), .B2(keyinput68), .C1(n10218), .C2(keyinput56), 
        .A(n8758), .ZN(n8762) );
  AOI22_X1 U10245 ( .A1(n9331), .A2(keyinput57), .B1(keyinput58), .B2(n6934), 
        .ZN(n8760) );
  OAI221_X1 U10246 ( .B1(n9331), .B2(keyinput57), .C1(n6934), .C2(keyinput58), 
        .A(n8760), .ZN(n8761) );
  NOR2_X1 U10247 ( .A1(n8762), .A2(n8761), .ZN(n8775) );
  AOI22_X1 U10248 ( .A1(n8764), .A2(keyinput64), .B1(n5453), .B2(keyinput89), 
        .ZN(n8763) );
  OAI221_X1 U10249 ( .B1(n8764), .B2(keyinput64), .C1(n5453), .C2(keyinput89), 
        .A(n8763), .ZN(n8767) );
  AOI22_X1 U10250 ( .A1(n6806), .A2(keyinput47), .B1(n7826), .B2(keyinput97), 
        .ZN(n8765) );
  OAI221_X1 U10251 ( .B1(n6806), .B2(keyinput47), .C1(n7826), .C2(keyinput97), 
        .A(n8765), .ZN(n8766) );
  NOR2_X1 U10252 ( .A1(n8767), .A2(n8766), .ZN(n8774) );
  AOI22_X1 U10253 ( .A1(n9385), .A2(keyinput67), .B1(keyinput85), .B2(n10214), 
        .ZN(n8768) );
  OAI221_X1 U10254 ( .B1(n9385), .B2(keyinput67), .C1(n10214), .C2(keyinput85), 
        .A(n8768), .ZN(n8772) );
  AOI22_X1 U10255 ( .A1(n8770), .A2(keyinput77), .B1(n10157), .B2(keyinput101), 
        .ZN(n8769) );
  OAI221_X1 U10256 ( .B1(n8770), .B2(keyinput77), .C1(n10157), .C2(keyinput101), .A(n8769), .ZN(n8771) );
  NOR2_X1 U10257 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND4_X1 U10258 ( .A1(n8776), .A2(n8775), .A3(n8774), .A4(n8773), .ZN(n8777)
         );
  NOR2_X1 U10259 ( .A1(n8778), .A2(n8777), .ZN(n8779) );
  AND4_X1 U10260 ( .A1(n8782), .A2(n8781), .A3(n8780), .A4(n8779), .ZN(n8783)
         );
  OAI211_X1 U10261 ( .C1(n8786), .C2(n8785), .A(n8784), .B(n8783), .ZN(n8797)
         );
  OAI21_X1 U10262 ( .B1(n8789), .B2(n8788), .A(n8787), .ZN(n8795) );
  NOR2_X1 U10263 ( .A1(n9150), .A2(n8893), .ZN(n8794) );
  INV_X1 U10264 ( .A(n8790), .ZN(n9154) );
  AOI22_X1 U10265 ( .A1(n9154), .A2(n8875), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8792) );
  NAND2_X1 U10266 ( .A1(n8890), .A2(n9153), .ZN(n8791) );
  OAI211_X1 U10267 ( .C1(n8885), .C2(n9147), .A(n8792), .B(n8791), .ZN(n8793)
         );
  AOI211_X1 U10268 ( .C1(n8795), .C2(n8882), .A(n8794), .B(n8793), .ZN(n8796)
         );
  XOR2_X1 U10269 ( .A(n8797), .B(n8796), .Z(P2_U3221) );
  XNOR2_X1 U10270 ( .A(n8799), .B(n8798), .ZN(n8805) );
  OAI22_X1 U10271 ( .A1(n9094), .A2(n8887), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8800), .ZN(n8801) );
  AOI21_X1 U10272 ( .B1(n8890), .B2(n9154), .A(n8801), .ZN(n8802) );
  OAI21_X1 U10273 ( .B1(n9123), .B2(n8885), .A(n8802), .ZN(n8803) );
  AOI21_X1 U10274 ( .B1(n9260), .B2(n8848), .A(n8803), .ZN(n8804) );
  OAI21_X1 U10275 ( .B1(n8805), .B2(n8866), .A(n8804), .ZN(P2_U3225) );
  XNOR2_X1 U10276 ( .A(n8808), .B(n8807), .ZN(n8809) );
  XNOR2_X1 U10277 ( .A(n8806), .B(n8809), .ZN(n8814) );
  NAND2_X1 U10278 ( .A1(n9058), .A2(n8875), .ZN(n8811) );
  AOI22_X1 U10279 ( .A1(n9057), .A2(n8890), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8810) );
  OAI211_X1 U10280 ( .C1(n8885), .C2(n9051), .A(n8811), .B(n8810), .ZN(n8812)
         );
  AOI21_X1 U10281 ( .B1(n9242), .B2(n8848), .A(n8812), .ZN(n8813) );
  OAI21_X1 U10282 ( .B1(n8814), .B2(n8866), .A(n8813), .ZN(P2_U3227) );
  OAI21_X1 U10283 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8818) );
  NAND2_X1 U10284 ( .A1(n8818), .A2(n8882), .ZN(n8822) );
  NOR2_X1 U10285 ( .A1(n8885), .A2(n9204), .ZN(n8820) );
  NAND2_X1 U10286 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8935) );
  OAI21_X1 U10287 ( .B1(n8887), .B2(n8862), .A(n8935), .ZN(n8819) );
  AOI211_X1 U10288 ( .C1(n8890), .C2(n9196), .A(n8820), .B(n8819), .ZN(n8821)
         );
  OAI211_X1 U10289 ( .C1(n9207), .C2(n8893), .A(n8822), .B(n8821), .ZN(
        P2_U3228) );
  XNOR2_X1 U10290 ( .A(n8823), .B(n8824), .ZN(n8829) );
  OAI22_X1 U10291 ( .A1(n8887), .A2(n9183), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8949), .ZN(n8825) );
  AOI21_X1 U10292 ( .B1(n8890), .B2(n8898), .A(n8825), .ZN(n8826) );
  OAI21_X1 U10293 ( .B1(n9187), .B2(n8885), .A(n8826), .ZN(n8827) );
  AOI21_X1 U10294 ( .B1(n9284), .B2(n8848), .A(n8827), .ZN(n8828) );
  OAI21_X1 U10295 ( .B1(n8829), .B2(n8866), .A(n8828), .ZN(P2_U3230) );
  AOI21_X1 U10296 ( .B1(n8831), .B2(n8426), .A(n8830), .ZN(n8835) );
  XNOR2_X1 U10297 ( .A(n8833), .B(n8832), .ZN(n8834) );
  XNOR2_X1 U10298 ( .A(n8835), .B(n8834), .ZN(n8841) );
  OAI22_X1 U10299 ( .A1(n9108), .A2(n8873), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8836), .ZN(n8837) );
  AOI21_X1 U10300 ( .B1(n9072), .B2(n8871), .A(n8837), .ZN(n8838) );
  OAI21_X1 U10301 ( .B1(n9069), .B2(n8887), .A(n8838), .ZN(n8839) );
  AOI21_X1 U10302 ( .B1(n9247), .B2(n8848), .A(n8839), .ZN(n8840) );
  OAI21_X1 U10303 ( .B1(n8841), .B2(n8866), .A(n8840), .ZN(P2_U3231) );
  XNOR2_X1 U10304 ( .A(n8843), .B(n8842), .ZN(n8850) );
  OAI22_X1 U10305 ( .A1(n8887), .A2(n9107), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8844), .ZN(n8845) );
  AOI21_X1 U10306 ( .B1(n8890), .B2(n9168), .A(n8845), .ZN(n8846) );
  OAI21_X1 U10307 ( .B1(n9135), .B2(n8885), .A(n8846), .ZN(n8847) );
  AOI21_X1 U10308 ( .B1(n9267), .B2(n8848), .A(n8847), .ZN(n8849) );
  OAI21_X1 U10309 ( .B1(n8850), .B2(n8866), .A(n8849), .ZN(P2_U3235) );
  OAI21_X1 U10310 ( .B1(n8853), .B2(n8852), .A(n8851), .ZN(n8854) );
  NAND2_X1 U10311 ( .A1(n8854), .A2(n8882), .ZN(n8858) );
  AOI22_X1 U10312 ( .A1(n8890), .A2(n9131), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8855) );
  OAI21_X1 U10313 ( .B1(n9108), .B2(n8887), .A(n8855), .ZN(n8856) );
  AOI21_X1 U10314 ( .B1(n9099), .B2(n8871), .A(n8856), .ZN(n8857) );
  OAI211_X1 U10315 ( .C1(n9101), .C2(n8893), .A(n8858), .B(n8857), .ZN(
        P2_U3237) );
  XNOR2_X1 U10316 ( .A(n8860), .B(n8859), .ZN(n8867) );
  NAND2_X1 U10317 ( .A1(n8875), .A2(n9168), .ZN(n8861) );
  NAND2_X1 U10318 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n10190)
         );
  OAI211_X1 U10319 ( .C1(n8862), .C2(n8873), .A(n8861), .B(n10190), .ZN(n8864)
         );
  NOR2_X1 U10320 ( .A1(n4739), .A2(n8893), .ZN(n8863) );
  AOI211_X1 U10321 ( .C1(n8871), .C2(n9162), .A(n8864), .B(n8863), .ZN(n8865)
         );
  OAI21_X1 U10322 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(P2_U3240) );
  INV_X1 U10323 ( .A(n9237), .ZN(n8878) );
  OAI211_X1 U10324 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8882), .ZN(n8877)
         );
  AOI22_X1 U10325 ( .A1(n9038), .A2(n8871), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8872) );
  OAI21_X1 U10326 ( .B1(n9069), .B2(n8873), .A(n8872), .ZN(n8874) );
  AOI21_X1 U10327 ( .B1(n9003), .B2(n8875), .A(n8874), .ZN(n8876) );
  OAI211_X1 U10328 ( .C1(n8878), .C2(n8893), .A(n8877), .B(n8876), .ZN(
        P2_U3242) );
  OAI21_X1 U10329 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8883) );
  NAND2_X1 U10330 ( .A1(n8883), .A2(n8882), .ZN(n8892) );
  NOR2_X1 U10331 ( .A1(n8885), .A2(n8884), .ZN(n8889) );
  OAI21_X1 U10332 ( .B1(n8887), .B2(n9181), .A(n8886), .ZN(n8888) );
  AOI211_X1 U10333 ( .C1(n8890), .C2(n8899), .A(n8889), .B(n8888), .ZN(n8891)
         );
  OAI211_X1 U10334 ( .C1(n8894), .C2(n8893), .A(n8892), .B(n8891), .ZN(
        P2_U3243) );
  MUX2_X1 U10335 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8895), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U10336 ( .A(n9002), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8913), .Z(
        P2_U3581) );
  MUX2_X1 U10337 ( .A(n8896), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8913), .Z(
        P2_U3580) );
  MUX2_X1 U10338 ( .A(n9003), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8913), .Z(
        P2_U3579) );
  MUX2_X1 U10339 ( .A(n9058), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8913), .Z(
        P2_U3578) );
  MUX2_X1 U10340 ( .A(n8897), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8913), .Z(
        P2_U3577) );
  MUX2_X1 U10341 ( .A(n9057), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8913), .Z(
        P2_U3576) );
  MUX2_X1 U10342 ( .A(n8394), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8913), .Z(
        P2_U3574) );
  MUX2_X1 U10343 ( .A(n9131), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8913), .Z(
        P2_U3573) );
  MUX2_X1 U10344 ( .A(n9154), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8913), .Z(
        P2_U3572) );
  MUX2_X1 U10345 ( .A(n9168), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8913), .Z(
        P2_U3571) );
  MUX2_X1 U10346 ( .A(n9153), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8913), .Z(
        P2_U3570) );
  MUX2_X1 U10347 ( .A(n9198), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8913), .Z(
        P2_U3569) );
  MUX2_X1 U10348 ( .A(n8898), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8913), .Z(
        P2_U3568) );
  MUX2_X1 U10349 ( .A(n9196), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8913), .Z(
        P2_U3567) );
  MUX2_X1 U10350 ( .A(n8899), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8913), .Z(
        P2_U3566) );
  MUX2_X1 U10351 ( .A(n8900), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8913), .Z(
        P2_U3565) );
  MUX2_X1 U10352 ( .A(n8901), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8913), .Z(
        P2_U3564) );
  MUX2_X1 U10353 ( .A(n8902), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8913), .Z(
        P2_U3563) );
  MUX2_X1 U10354 ( .A(n8903), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8913), .Z(
        P2_U3562) );
  MUX2_X1 U10355 ( .A(n8904), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8913), .Z(
        P2_U3561) );
  MUX2_X1 U10356 ( .A(n8905), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8913), .Z(
        P2_U3560) );
  MUX2_X1 U10357 ( .A(n8906), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8913), .Z(
        P2_U3559) );
  MUX2_X1 U10358 ( .A(n8907), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8913), .Z(
        P2_U3558) );
  MUX2_X1 U10359 ( .A(n8908), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8913), .Z(
        P2_U3557) );
  MUX2_X1 U10360 ( .A(n8909), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8913), .Z(
        P2_U3556) );
  MUX2_X1 U10361 ( .A(n8910), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8913), .Z(
        P2_U3555) );
  MUX2_X1 U10362 ( .A(n8911), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8913), .Z(
        P2_U3554) );
  MUX2_X1 U10363 ( .A(n8912), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8913), .Z(
        P2_U3553) );
  MUX2_X1 U10364 ( .A(n8914), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8913), .Z(
        P2_U3552) );
  AOI211_X1 U10365 ( .C1(n8917), .C2(n8916), .A(n10171), .B(n8915), .ZN(n8918)
         );
  INV_X1 U10366 ( .A(n8918), .ZN(n8928) );
  NOR2_X1 U10367 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8919), .ZN(n8922) );
  NOR2_X1 U10368 ( .A1(n10170), .A2(n8920), .ZN(n8921) );
  AOI211_X1 U10369 ( .C1(n10187), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n8922), .B(
        n8921), .ZN(n8927) );
  OAI211_X1 U10370 ( .C1(n8925), .C2(n8924), .A(n10185), .B(n8923), .ZN(n8926)
         );
  NAND3_X1 U10371 ( .A1(n8928), .A2(n8927), .A3(n8926), .ZN(P2_U3252) );
  NOR2_X1 U10372 ( .A1(n8930), .A2(n8929), .ZN(n8932) );
  NOR2_X1 U10373 ( .A1(n8932), .A2(n8931), .ZN(n8934) );
  MUX2_X1 U10374 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9205), .S(n8955), .Z(n8933) );
  NAND2_X1 U10375 ( .A1(n8933), .A2(n8934), .ZN(n8956) );
  OAI211_X1 U10376 ( .C1(n8934), .C2(n8933), .A(n10185), .B(n8956), .ZN(n8948)
         );
  INV_X1 U10377 ( .A(n8935), .ZN(n8936) );
  AOI21_X1 U10378 ( .B1(n10187), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8936), .ZN(
        n8947) );
  NOR2_X1 U10379 ( .A1(n8938), .A2(n8937), .ZN(n8940) );
  NOR2_X1 U10380 ( .A1(n8940), .A2(n8939), .ZN(n8943) );
  XNOR2_X1 U10381 ( .A(n8955), .B(n8941), .ZN(n8942) );
  NAND2_X1 U10382 ( .A1(n8942), .A2(n8943), .ZN(n8950) );
  OAI21_X1 U10383 ( .B1(n8943), .B2(n8942), .A(n8950), .ZN(n8944) );
  NAND2_X1 U10384 ( .A1(n8944), .A2(n10181), .ZN(n8946) );
  NAND2_X1 U10385 ( .A1(n10183), .A2(n8955), .ZN(n8945) );
  NAND4_X1 U10386 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(
        P2_U3261) );
  NOR2_X1 U10387 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8949), .ZN(n8954) );
  XNOR2_X1 U10388 ( .A(n8971), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8951) );
  AOI211_X1 U10389 ( .C1(n8952), .C2(n8951), .A(n8970), .B(n10171), .ZN(n8953)
         );
  AOI211_X1 U10390 ( .C1(n10187), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8954), .B(
        n8953), .ZN(n8961) );
  XNOR2_X1 U10391 ( .A(n8962), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8959) );
  INV_X1 U10392 ( .A(n8955), .ZN(n8957) );
  OAI21_X1 U10393 ( .B1(n8957), .B2(n9205), .A(n8956), .ZN(n8958) );
  NAND2_X1 U10394 ( .A1(n8959), .A2(n8958), .ZN(n8963) );
  OAI211_X1 U10395 ( .C1(n8959), .C2(n8958), .A(n10185), .B(n8963), .ZN(n8960)
         );
  OAI211_X1 U10396 ( .C1(n10170), .C2(n8962), .A(n8961), .B(n8960), .ZN(
        P2_U3262) );
  NAND2_X1 U10397 ( .A1(n8971), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U10398 ( .A1(n8964), .A2(n8963), .ZN(n8966) );
  XNOR2_X1 U10399 ( .A(n8965), .B(n8966), .ZN(n10186) );
  NAND2_X1 U10400 ( .A1(n10186), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U10401 ( .A1(n8966), .A2(n10182), .ZN(n8967) );
  NAND2_X1 U10402 ( .A1(n10184), .A2(n8967), .ZN(n8968) );
  XOR2_X1 U10403 ( .A(n8968), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8975) );
  XNOR2_X1 U10404 ( .A(n10182), .B(n8969), .ZN(n10179) );
  NOR2_X1 U10405 ( .A1(n10182), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8972) );
  XNOR2_X1 U10406 ( .A(n8973), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8974) );
  AND2_X1 U10407 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8977) );
  AOI21_X1 U10408 ( .B1(n10187), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8977), .ZN(
        n8978) );
  NAND2_X1 U10409 ( .A1(n8979), .A2(n8978), .ZN(P2_U3264) );
  NAND2_X1 U10410 ( .A1(n8987), .A2(n8986), .ZN(n8985) );
  XNOR2_X1 U10411 ( .A(n9217), .B(n8985), .ZN(n9219) );
  NOR2_X1 U10412 ( .A1(n9190), .A2(n8980), .ZN(n8983) );
  NAND2_X1 U10413 ( .A1(n8982), .A2(n8981), .ZN(n9891) );
  NOR2_X1 U10414 ( .A1(n10210), .A2(n9891), .ZN(n8989) );
  AOI211_X1 U10415 ( .C1(n9217), .C2(n10205), .A(n8983), .B(n8989), .ZN(n8984)
         );
  OAI21_X1 U10416 ( .B1(n9219), .B2(n8991), .A(n8984), .ZN(P2_U3265) );
  NOR2_X1 U10417 ( .A1(n8987), .A2(n9164), .ZN(n8988) );
  AOI211_X1 U10418 ( .C1(n10210), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8989), .B(
        n8988), .ZN(n8990) );
  OAI21_X1 U10419 ( .B1(n8991), .B2(n9892), .A(n8990), .ZN(P2_U3266) );
  OAI21_X1 U10420 ( .B1(n8993), .B2(n9001), .A(n8992), .ZN(n8994) );
  INV_X1 U10421 ( .A(n8994), .ZN(n9229) );
  INV_X1 U10422 ( .A(n8995), .ZN(n8996) );
  AOI211_X1 U10423 ( .C1(n9226), .C2(n9011), .A(n10261), .B(n8996), .ZN(n9225)
         );
  INV_X1 U10424 ( .A(n9226), .ZN(n8999) );
  AOI22_X1 U10425 ( .A1(n8997), .A2(n9161), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10210), .ZN(n8998) );
  OAI21_X1 U10426 ( .B1(n8999), .B2(n9164), .A(n8998), .ZN(n9005) );
  XNOR2_X1 U10427 ( .A(n9000), .B(n9001), .ZN(n9004) );
  AOI222_X1 U10428 ( .A1(n10194), .A2(n9004), .B1(n9003), .B2(n9195), .C1(
        n9002), .C2(n9197), .ZN(n9228) );
  OAI21_X1 U10429 ( .B1(n9229), .B2(n9214), .A(n9006), .ZN(P2_U3268) );
  OAI21_X1 U10430 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9010) );
  INV_X1 U10431 ( .A(n9010), .ZN(n9234) );
  INV_X1 U10432 ( .A(n9037), .ZN(n9013) );
  INV_X1 U10433 ( .A(n9011), .ZN(n9012) );
  AOI21_X1 U10434 ( .B1(n9230), .B2(n9013), .A(n9012), .ZN(n9231) );
  AOI22_X1 U10435 ( .A1(n9014), .A2(n9161), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10210), .ZN(n9015) );
  OAI21_X1 U10436 ( .B1(n9016), .B2(n9164), .A(n9015), .ZN(n9027) );
  AOI21_X1 U10437 ( .B1(n9017), .B2(n9019), .A(n9018), .ZN(n9020) );
  NOR2_X1 U10438 ( .A1(n9020), .A2(n9180), .ZN(n9025) );
  OAI22_X1 U10439 ( .A1(n9022), .A2(n9184), .B1(n9021), .B2(n9182), .ZN(n9023)
         );
  AOI21_X1 U10440 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9233) );
  NOR2_X1 U10441 ( .A1(n9233), .A2(n10210), .ZN(n9026) );
  AOI211_X1 U10442 ( .C1(n9231), .C2(n9211), .A(n9027), .B(n9026), .ZN(n9028)
         );
  OAI21_X1 U10443 ( .B1(n9234), .B2(n9214), .A(n9028), .ZN(P2_U3269) );
  OAI21_X1 U10444 ( .B1(n9030), .B2(n9034), .A(n9029), .ZN(n9031) );
  INV_X1 U10445 ( .A(n9031), .ZN(n9239) );
  AOI22_X1 U10446 ( .A1(n9237), .A2(n10205), .B1(n10210), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9043) );
  INV_X1 U10447 ( .A(n9017), .ZN(n9032) );
  OAI222_X1 U10448 ( .A1(n9184), .A2(n9036), .B1(n9182), .B2(n9069), .C1(n9180), .C2(n9035), .ZN(n9235) );
  AOI211_X1 U10449 ( .C1(n9237), .C2(n9048), .A(n10261), .B(n9037), .ZN(n9236)
         );
  INV_X1 U10450 ( .A(n9236), .ZN(n9040) );
  INV_X1 U10451 ( .A(n9038), .ZN(n9039) );
  OAI22_X1 U10452 ( .A1(n9040), .A2(n9188), .B1(n10199), .B2(n9039), .ZN(n9041) );
  OAI21_X1 U10453 ( .B1(n9235), .B2(n9041), .A(n9190), .ZN(n9042) );
  OAI211_X1 U10454 ( .C1(n9239), .C2(n9214), .A(n9043), .B(n9042), .ZN(
        P2_U3270) );
  OAI21_X1 U10455 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9047) );
  INV_X1 U10456 ( .A(n9047), .ZN(n9244) );
  AOI211_X1 U10457 ( .C1(n9242), .C2(n9070), .A(n10261), .B(n4746), .ZN(n9241)
         );
  INV_X1 U10458 ( .A(n9242), .ZN(n9049) );
  NOR2_X1 U10459 ( .A1(n9049), .A2(n9164), .ZN(n9053) );
  OAI22_X1 U10460 ( .A1(n9051), .A2(n10199), .B1(n9050), .B2(n9190), .ZN(n9052) );
  AOI211_X1 U10461 ( .C1(n9241), .C2(n9172), .A(n9053), .B(n9052), .ZN(n9062)
         );
  OAI211_X1 U10462 ( .C1(n9056), .C2(n9055), .A(n9054), .B(n10194), .ZN(n9060)
         );
  AOI22_X1 U10463 ( .A1(n9058), .A2(n9197), .B1(n9195), .B2(n9057), .ZN(n9059)
         );
  NAND2_X1 U10464 ( .A1(n9060), .A2(n9059), .ZN(n9240) );
  NAND2_X1 U10465 ( .A1(n9240), .A2(n9190), .ZN(n9061) );
  OAI211_X1 U10466 ( .C1(n9244), .C2(n9214), .A(n9062), .B(n9061), .ZN(
        P2_U3271) );
  XNOR2_X1 U10467 ( .A(n9063), .B(n9066), .ZN(n9249) );
  NAND2_X1 U10468 ( .A1(n9064), .A2(n9065), .ZN(n9067) );
  XNOR2_X1 U10469 ( .A(n9067), .B(n9066), .ZN(n9068) );
  OAI222_X1 U10470 ( .A1(n9184), .A2(n9069), .B1(n9182), .B2(n9108), .C1(n9068), .C2(n9180), .ZN(n9245) );
  INV_X1 U10471 ( .A(n9081), .ZN(n9071) );
  AOI211_X1 U10472 ( .C1(n9247), .C2(n9071), .A(n10261), .B(n4742), .ZN(n9246)
         );
  NAND2_X1 U10473 ( .A1(n9246), .A2(n9172), .ZN(n9074) );
  AOI22_X1 U10474 ( .A1(n9072), .A2(n9161), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10210), .ZN(n9073) );
  OAI211_X1 U10475 ( .C1(n9075), .C2(n9164), .A(n9074), .B(n9073), .ZN(n9076)
         );
  AOI21_X1 U10476 ( .B1(n9245), .B2(n9190), .A(n9076), .ZN(n9077) );
  OAI21_X1 U10477 ( .B1(n9249), .B2(n9214), .A(n9077), .ZN(P2_U3272) );
  OAI21_X1 U10478 ( .B1(n9080), .B2(n9079), .A(n9078), .ZN(n9254) );
  INV_X1 U10479 ( .A(n9098), .ZN(n9082) );
  AOI211_X1 U10480 ( .C1(n9252), .C2(n9082), .A(n10261), .B(n9081), .ZN(n9251)
         );
  NOR2_X1 U10481 ( .A1(n9083), .A2(n9164), .ZN(n9087) );
  OAI22_X1 U10482 ( .A1(n9085), .A2(n10199), .B1(n9084), .B2(n9190), .ZN(n9086) );
  AOI211_X1 U10483 ( .C1(n9251), .C2(n9172), .A(n9087), .B(n9086), .ZN(n9096)
         );
  INV_X1 U10484 ( .A(n9064), .ZN(n9091) );
  AOI21_X1 U10485 ( .B1(n9088), .B2(n9089), .A(n5027), .ZN(n9090) );
  NOR2_X1 U10486 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  OAI222_X1 U10487 ( .A1(n9182), .A2(n9094), .B1(n9184), .B2(n9093), .C1(n9180), .C2(n9092), .ZN(n9250) );
  NAND2_X1 U10488 ( .A1(n9250), .A2(n9190), .ZN(n9095) );
  OAI211_X1 U10489 ( .C1(n9254), .C2(n9214), .A(n9096), .B(n9095), .ZN(
        P2_U3273) );
  XOR2_X1 U10490 ( .A(n9097), .B(n9106), .Z(n9259) );
  AOI21_X1 U10491 ( .B1(n9255), .B2(n9116), .A(n9098), .ZN(n9256) );
  AOI22_X1 U10492 ( .A1(n10210), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9099), 
        .B2(n9161), .ZN(n9100) );
  OAI21_X1 U10493 ( .B1(n9101), .B2(n9164), .A(n9100), .ZN(n9112) );
  NAND2_X1 U10494 ( .A1(n9102), .A2(n9103), .ZN(n9105) );
  INV_X1 U10495 ( .A(n9088), .ZN(n9104) );
  AOI211_X1 U10496 ( .C1(n9106), .C2(n9105), .A(n9180), .B(n9104), .ZN(n9110)
         );
  OAI22_X1 U10497 ( .A1(n9108), .A2(n9184), .B1(n9107), .B2(n9182), .ZN(n9109)
         );
  NOR2_X1 U10498 ( .A1(n9110), .A2(n9109), .ZN(n9258) );
  NOR2_X1 U10499 ( .A1(n9258), .A2(n10210), .ZN(n9111) );
  AOI211_X1 U10500 ( .C1(n9256), .C2(n9211), .A(n9112), .B(n9111), .ZN(n9113)
         );
  OAI21_X1 U10501 ( .B1(n9259), .B2(n9214), .A(n9113), .ZN(P2_U3274) );
  XNOR2_X1 U10502 ( .A(n9114), .B(n9121), .ZN(n9264) );
  NAND2_X1 U10503 ( .A1(n9140), .A2(n9260), .ZN(n9115) );
  AND2_X1 U10504 ( .A1(n9116), .A2(n9115), .ZN(n9261) );
  OAI22_X1 U10505 ( .A1(n9118), .A2(n9164), .B1(n9190), .B2(n9117), .ZN(n9119)
         );
  AOI21_X1 U10506 ( .B1(n9261), .B2(n9211), .A(n9119), .ZN(n9126) );
  OAI21_X1 U10507 ( .B1(n8142), .B2(n8141), .A(n9102), .ZN(n9122) );
  AOI222_X1 U10508 ( .A1(n10194), .A2(n9122), .B1(n8394), .B2(n9197), .C1(
        n9154), .C2(n9195), .ZN(n9263) );
  OAI21_X1 U10509 ( .B1(n9123), .B2(n10199), .A(n9263), .ZN(n9124) );
  NAND2_X1 U10510 ( .A1(n9124), .A2(n9190), .ZN(n9125) );
  OAI211_X1 U10511 ( .C1(n9264), .C2(n9214), .A(n9126), .B(n9125), .ZN(
        P2_U3275) );
  NAND2_X1 U10512 ( .A1(n9127), .A2(n9128), .ZN(n9130) );
  XNOR2_X1 U10513 ( .A(n9130), .B(n9129), .ZN(n9132) );
  AOI222_X1 U10514 ( .A1(n10194), .A2(n9132), .B1(n9131), .B2(n9197), .C1(
        n9168), .C2(n9195), .ZN(n9270) );
  OR2_X1 U10515 ( .A1(n9134), .A2(n9133), .ZN(n9266) );
  NAND3_X1 U10516 ( .A1(n9266), .A2(n9265), .A3(n10207), .ZN(n9143) );
  OAI22_X1 U10517 ( .A1(n9190), .A2(n9136), .B1(n9135), .B2(n10199), .ZN(n9137) );
  AOI21_X1 U10518 ( .B1(n9267), .B2(n10205), .A(n9137), .ZN(n9142) );
  OR2_X1 U10519 ( .A1(n9146), .A2(n9138), .ZN(n9139) );
  AND2_X1 U10520 ( .A1(n9140), .A2(n9139), .ZN(n9268) );
  NAND2_X1 U10521 ( .A1(n9268), .A2(n9211), .ZN(n9141) );
  AND3_X1 U10522 ( .A1(n9143), .A2(n9142), .A3(n9141), .ZN(n9144) );
  OAI21_X1 U10523 ( .B1(n10210), .B2(n9270), .A(n9144), .ZN(P2_U3276) );
  XOR2_X1 U10524 ( .A(n9145), .B(n9152), .Z(n9276) );
  AOI211_X1 U10525 ( .C1(n9273), .C2(n4741), .A(n10261), .B(n9146), .ZN(n9272)
         );
  INV_X1 U10526 ( .A(n9147), .ZN(n9148) );
  AOI22_X1 U10527 ( .A1(n10210), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9148), 
        .B2(n9161), .ZN(n9149) );
  OAI21_X1 U10528 ( .B1(n9150), .B2(n9164), .A(n9149), .ZN(n9157) );
  OAI21_X1 U10529 ( .B1(n9152), .B2(n9151), .A(n9127), .ZN(n9155) );
  AOI222_X1 U10530 ( .A1(n10194), .A2(n9155), .B1(n9154), .B2(n9197), .C1(
        n9153), .C2(n9195), .ZN(n9275) );
  NOR2_X1 U10531 ( .A1(n9275), .A2(n10210), .ZN(n9156) );
  AOI211_X1 U10532 ( .C1(n9272), .C2(n9172), .A(n9157), .B(n9156), .ZN(n9158)
         );
  OAI21_X1 U10533 ( .B1(n9214), .B2(n9276), .A(n9158), .ZN(P2_U3277) );
  XNOR2_X1 U10534 ( .A(n9159), .B(n9166), .ZN(n9281) );
  AOI211_X1 U10535 ( .C1(n9278), .C2(n9185), .A(n10261), .B(n9160), .ZN(n9277)
         );
  AOI22_X1 U10536 ( .A1(n10210), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9162), 
        .B2(n9161), .ZN(n9163) );
  OAI21_X1 U10537 ( .B1(n4739), .B2(n9164), .A(n9163), .ZN(n9171) );
  OAI21_X1 U10538 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9169) );
  AOI222_X1 U10539 ( .A1(n10194), .A2(n9169), .B1(n9168), .B2(n9197), .C1(
        n9198), .C2(n9195), .ZN(n9280) );
  NOR2_X1 U10540 ( .A1(n9280), .A2(n10210), .ZN(n9170) );
  AOI211_X1 U10541 ( .C1(n9277), .C2(n9172), .A(n9171), .B(n9170), .ZN(n9173)
         );
  OAI21_X1 U10542 ( .B1(n9281), .B2(n9214), .A(n9173), .ZN(P2_U3278) );
  OAI21_X1 U10543 ( .B1(n9175), .B2(n9177), .A(n9174), .ZN(n9176) );
  INV_X1 U10544 ( .A(n9176), .ZN(n9286) );
  AOI22_X1 U10545 ( .A1(n9284), .A2(n10205), .B1(n10210), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n9193) );
  XNOR2_X1 U10546 ( .A(n9178), .B(n9177), .ZN(n9179) );
  OAI222_X1 U10547 ( .A1(n9184), .A2(n9183), .B1(n9182), .B2(n9181), .C1(n9180), .C2(n9179), .ZN(n9282) );
  INV_X1 U10548 ( .A(n9185), .ZN(n9186) );
  AOI211_X1 U10549 ( .C1(n9284), .C2(n9210), .A(n10261), .B(n9186), .ZN(n9283)
         );
  INV_X1 U10550 ( .A(n9283), .ZN(n9189) );
  OAI22_X1 U10551 ( .A1(n9189), .A2(n9188), .B1(n10199), .B2(n9187), .ZN(n9191) );
  OAI21_X1 U10552 ( .B1(n9282), .B2(n9191), .A(n9190), .ZN(n9192) );
  OAI211_X1 U10553 ( .C1(n9286), .C2(n9214), .A(n9193), .B(n9192), .ZN(
        P2_U3279) );
  XNOR2_X1 U10554 ( .A(n9194), .B(n9202), .ZN(n9199) );
  AOI222_X1 U10555 ( .A1(n10194), .A2(n9199), .B1(n9198), .B2(n9197), .C1(
        n9196), .C2(n9195), .ZN(n9290) );
  AOI21_X1 U10556 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(n9203) );
  INV_X1 U10557 ( .A(n9203), .ZN(n9291) );
  OAI22_X1 U10558 ( .A1(n9190), .A2(n9205), .B1(n9204), .B2(n10199), .ZN(n9206) );
  AOI21_X1 U10559 ( .B1(n9287), .B2(n10205), .A(n9206), .ZN(n9213) );
  OR2_X1 U10560 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  AND2_X1 U10561 ( .A1(n9210), .A2(n9209), .ZN(n9288) );
  NAND2_X1 U10562 ( .A1(n9288), .A2(n9211), .ZN(n9212) );
  OAI211_X1 U10563 ( .C1(n9291), .C2(n9214), .A(n9213), .B(n9212), .ZN(n9215)
         );
  INV_X1 U10564 ( .A(n9215), .ZN(n9216) );
  OAI21_X1 U10565 ( .B1(n10210), .B2(n9290), .A(n9216), .ZN(P2_U3280) );
  NAND2_X1 U10566 ( .A1(n9217), .A2(n6570), .ZN(n9218) );
  OAI211_X1 U10567 ( .C1(n9219), .C2(n10261), .A(n9891), .B(n9218), .ZN(n9305)
         );
  MUX2_X1 U10568 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9305), .S(n10295), .Z(
        P2_U3551) );
  AOI22_X1 U10569 ( .A1(n9221), .A2(n10197), .B1(n6570), .B2(n9220), .ZN(n9222) );
  OAI211_X1 U10570 ( .C1(n9224), .C2(n9297), .A(n9223), .B(n9222), .ZN(n9306)
         );
  MUX2_X1 U10571 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9306), .S(n10295), .Z(
        P2_U3549) );
  AOI21_X1 U10572 ( .B1(n6570), .B2(n9226), .A(n9225), .ZN(n9227) );
  OAI211_X1 U10573 ( .C1(n9229), .C2(n9297), .A(n9228), .B(n9227), .ZN(n9307)
         );
  MUX2_X1 U10574 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9307), .S(n10295), .Z(
        P2_U3548) );
  AOI22_X1 U10575 ( .A1(n9231), .A2(n10197), .B1(n6570), .B2(n9230), .ZN(n9232) );
  OAI211_X1 U10576 ( .C1(n9234), .C2(n9297), .A(n9233), .B(n9232), .ZN(n9308)
         );
  MUX2_X1 U10577 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9308), .S(n10295), .Z(
        P2_U3547) );
  AOI211_X1 U10578 ( .C1(n6570), .C2(n9237), .A(n9236), .B(n9235), .ZN(n9238)
         );
  OAI21_X1 U10579 ( .B1(n9239), .B2(n9297), .A(n9238), .ZN(n9309) );
  MUX2_X1 U10580 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9309), .S(n10295), .Z(
        P2_U3546) );
  AOI211_X1 U10581 ( .C1(n6570), .C2(n9242), .A(n9241), .B(n9240), .ZN(n9243)
         );
  OAI21_X1 U10582 ( .B1(n9244), .B2(n9297), .A(n9243), .ZN(n9310) );
  MUX2_X1 U10583 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9310), .S(n10295), .Z(
        P2_U3545) );
  AOI211_X1 U10584 ( .C1(n6570), .C2(n9247), .A(n9246), .B(n9245), .ZN(n9248)
         );
  OAI21_X1 U10585 ( .B1(n9249), .B2(n9297), .A(n9248), .ZN(n9311) );
  MUX2_X1 U10586 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9311), .S(n10295), .Z(
        P2_U3544) );
  AOI211_X1 U10587 ( .C1(n6570), .C2(n9252), .A(n9251), .B(n9250), .ZN(n9253)
         );
  OAI21_X1 U10588 ( .B1(n9254), .B2(n9297), .A(n9253), .ZN(n9312) );
  MUX2_X1 U10589 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9312), .S(n10295), .Z(
        P2_U3543) );
  AOI22_X1 U10590 ( .A1(n9256), .A2(n10197), .B1(n6570), .B2(n9255), .ZN(n9257) );
  OAI211_X1 U10591 ( .C1(n9259), .C2(n9297), .A(n9258), .B(n9257), .ZN(n9313)
         );
  MUX2_X1 U10592 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9313), .S(n10295), .Z(
        P2_U3542) );
  AOI22_X1 U10593 ( .A1(n9261), .A2(n10197), .B1(n6570), .B2(n9260), .ZN(n9262) );
  OAI211_X1 U10594 ( .C1(n9264), .C2(n9297), .A(n9263), .B(n9262), .ZN(n9314)
         );
  MUX2_X1 U10595 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9314), .S(n10295), .Z(
        P2_U3541) );
  NAND3_X1 U10596 ( .A1(n9266), .A2(n9265), .A3(n10279), .ZN(n9271) );
  AOI22_X1 U10597 ( .A1(n9268), .A2(n10197), .B1(n6570), .B2(n9267), .ZN(n9269) );
  NAND3_X1 U10598 ( .A1(n9271), .A2(n9270), .A3(n9269), .ZN(n9315) );
  MUX2_X1 U10599 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9315), .S(n10295), .Z(
        P2_U3540) );
  AOI21_X1 U10600 ( .B1(n6570), .B2(n9273), .A(n9272), .ZN(n9274) );
  OAI211_X1 U10601 ( .C1(n9276), .C2(n9297), .A(n9275), .B(n9274), .ZN(n9316)
         );
  MUX2_X1 U10602 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9316), .S(n10295), .Z(
        P2_U3539) );
  AOI21_X1 U10603 ( .B1(n6570), .B2(n9278), .A(n9277), .ZN(n9279) );
  OAI211_X1 U10604 ( .C1(n9281), .C2(n9297), .A(n9280), .B(n9279), .ZN(n9317)
         );
  MUX2_X1 U10605 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9317), .S(n10295), .Z(
        P2_U3538) );
  AOI211_X1 U10606 ( .C1(n6570), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI21_X1 U10607 ( .B1(n9286), .B2(n9297), .A(n9285), .ZN(n9318) );
  MUX2_X1 U10608 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9318), .S(n10295), .Z(
        P2_U3537) );
  AOI22_X1 U10609 ( .A1(n9288), .A2(n10197), .B1(n6570), .B2(n9287), .ZN(n9289) );
  OAI211_X1 U10610 ( .C1(n9291), .C2(n9297), .A(n9290), .B(n9289), .ZN(n9319)
         );
  MUX2_X1 U10611 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9319), .S(n10295), .Z(
        P2_U3536) );
  INV_X1 U10612 ( .A(n9292), .ZN(n9298) );
  AOI22_X1 U10613 ( .A1(n9294), .A2(n10197), .B1(n6570), .B2(n9293), .ZN(n9295) );
  OAI211_X1 U10614 ( .C1(n9298), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9321)
         );
  MUX2_X1 U10615 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9321), .S(n10295), .Z(
        P2_U3535) );
  NAND2_X1 U10616 ( .A1(n9299), .A2(n6570), .ZN(n9301) );
  OAI211_X1 U10617 ( .C1(n9302), .C2(n10258), .A(n9301), .B(n9300), .ZN(n9303)
         );
  OR2_X1 U10618 ( .A1(n9304), .A2(n9303), .ZN(n9322) );
  MUX2_X1 U10619 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9322), .S(n10295), .Z(
        P2_U3533) );
  MUX2_X1 U10620 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9305), .S(n9320), .Z(
        P2_U3519) );
  MUX2_X1 U10621 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9306), .S(n9320), .Z(
        P2_U3517) );
  MUX2_X1 U10622 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9307), .S(n9320), .Z(
        P2_U3516) );
  MUX2_X1 U10623 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9308), .S(n9320), .Z(
        P2_U3515) );
  MUX2_X1 U10624 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9309), .S(n9320), .Z(
        P2_U3514) );
  MUX2_X1 U10625 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9310), .S(n9320), .Z(
        P2_U3513) );
  MUX2_X1 U10626 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9311), .S(n9320), .Z(
        P2_U3512) );
  MUX2_X1 U10627 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9312), .S(n9320), .Z(
        P2_U3511) );
  MUX2_X1 U10628 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9313), .S(n9320), .Z(
        P2_U3510) );
  MUX2_X1 U10629 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9314), .S(n9320), .Z(
        P2_U3509) );
  MUX2_X1 U10630 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9315), .S(n9320), .Z(
        P2_U3508) );
  MUX2_X1 U10631 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9316), .S(n9320), .Z(
        P2_U3507) );
  MUX2_X1 U10632 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9317), .S(n9320), .Z(
        P2_U3505) );
  MUX2_X1 U10633 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9318), .S(n9320), .Z(
        P2_U3502) );
  MUX2_X1 U10634 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9319), .S(n9320), .Z(
        P2_U3499) );
  MUX2_X1 U10635 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9321), .S(n9320), .Z(
        P2_U3496) );
  MUX2_X1 U10636 ( .A(n9322), .B(P2_REG0_REG_13__SCAN_IN), .S(n10281), .Z(
        P2_U3490) );
  INV_X1 U10637 ( .A(n9323), .ZN(n9877) );
  NOR4_X1 U10638 ( .A1(n9325), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9324), .A4(
        P2_U3152), .ZN(n9326) );
  AOI21_X1 U10639 ( .B1(n9327), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9326), .ZN(
        n9328) );
  OAI21_X1 U10640 ( .B1(n9877), .B2(n4490), .A(n9328), .ZN(P2_U3327) );
  INV_X1 U10641 ( .A(n9329), .ZN(n9880) );
  OAI222_X1 U10642 ( .A1(n9332), .A2(P2_U3152), .B1(n4490), .B2(n9880), .C1(
        n9331), .C2(n9330), .ZN(P2_U3329) );
  MUX2_X1 U10643 ( .A(n9333), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10644 ( .A(n9335), .B(n9334), .ZN(n9336) );
  XNOR2_X1 U10645 ( .A(n9337), .B(n9336), .ZN(n9344) );
  OAI22_X1 U10646 ( .A1(n9464), .A2(n9396), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9338), .ZN(n9342) );
  INV_X1 U10647 ( .A(n9583), .ZN(n9339) );
  OAI22_X1 U10648 ( .A1(n9340), .A2(n9451), .B1(n9453), .B2(n9339), .ZN(n9341)
         );
  AOI211_X1 U10649 ( .C1(n9789), .C2(n9477), .A(n9342), .B(n9341), .ZN(n9343)
         );
  OAI21_X1 U10650 ( .B1(n9344), .B2(n9470), .A(n9343), .ZN(P1_U3212) );
  AOI22_X1 U10651 ( .A1(n9476), .A2(n9736), .B1(n9475), .B2(n9345), .ZN(n9347)
         );
  OAI211_X1 U10652 ( .C1(n9348), .C2(n9464), .A(n9347), .B(n9346), .ZN(n9356)
         );
  INV_X1 U10653 ( .A(n9349), .ZN(n9354) );
  AOI21_X1 U10654 ( .B1(n9353), .B2(n9351), .A(n9350), .ZN(n9352) );
  AOI211_X1 U10655 ( .C1(n9354), .C2(n9353), .A(n9470), .B(n9352), .ZN(n9355)
         );
  AOI211_X1 U10656 ( .C1(n9477), .C2(n9357), .A(n9356), .B(n9355), .ZN(n9358)
         );
  INV_X1 U10657 ( .A(n9358), .ZN(P1_U3213) );
  INV_X1 U10658 ( .A(n9363), .ZN(n9360) );
  NOR2_X1 U10659 ( .A1(n9360), .A2(n9359), .ZN(n9365) );
  AOI21_X1 U10660 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9364) );
  OAI21_X1 U10661 ( .B1(n9365), .B2(n9364), .A(n9428), .ZN(n9371) );
  INV_X1 U10662 ( .A(n9634), .ZN(n9366) );
  OAI22_X1 U10663 ( .A1(n9386), .A2(n9464), .B1(n9453), .B2(n9366), .ZN(n9369)
         );
  OAI22_X1 U10664 ( .A1(n9451), .A2(n9398), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9367), .ZN(n9368) );
  NOR2_X1 U10665 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  OAI211_X1 U10666 ( .C1(n9636), .C2(n9372), .A(n9371), .B(n9370), .ZN(
        P1_U3214) );
  INV_X1 U10667 ( .A(n9373), .ZN(n9374) );
  AOI21_X1 U10668 ( .B1(n9376), .B2(n9375), .A(n9374), .ZN(n9380) );
  NAND2_X1 U10669 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9550) );
  OAI21_X1 U10670 ( .B1(n9451), .B2(n9388), .A(n9550), .ZN(n9378) );
  OAI22_X1 U10671 ( .A1(n9420), .A2(n9464), .B1(n9453), .B2(n9686), .ZN(n9377)
         );
  AOI211_X1 U10672 ( .C1(n9828), .C2(n9477), .A(n9378), .B(n9377), .ZN(n9379)
         );
  OAI21_X1 U10673 ( .B1(n9380), .B2(n9470), .A(n9379), .ZN(P1_U3217) );
  NOR2_X1 U10674 ( .A1(n4759), .A2(n9382), .ZN(n9383) );
  XNOR2_X1 U10675 ( .A(n9384), .B(n9383), .ZN(n9392) );
  OAI22_X1 U10676 ( .A1(n9451), .A2(n9386), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9385), .ZN(n9390) );
  INV_X1 U10677 ( .A(n9660), .ZN(n9387) );
  OAI22_X1 U10678 ( .A1(n9388), .A2(n9464), .B1(n9453), .B2(n9387), .ZN(n9389)
         );
  AOI211_X1 U10679 ( .C1(n9818), .C2(n9477), .A(n9390), .B(n9389), .ZN(n9391)
         );
  OAI21_X1 U10680 ( .B1(n9392), .B2(n9470), .A(n9391), .ZN(P1_U3221) );
  XOR2_X1 U10681 ( .A(n9394), .B(n9393), .Z(n9402) );
  OAI22_X1 U10682 ( .A1(n9451), .A2(n9396), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9395), .ZN(n9400) );
  INV_X1 U10683 ( .A(n9605), .ZN(n9397) );
  OAI22_X1 U10684 ( .A1(n9398), .A2(n9464), .B1(n9453), .B2(n9397), .ZN(n9399)
         );
  AOI211_X1 U10685 ( .C1(n9798), .C2(n9477), .A(n9400), .B(n9399), .ZN(n9401)
         );
  OAI21_X1 U10686 ( .B1(n9402), .B2(n9470), .A(n9401), .ZN(P1_U3223) );
  INV_X1 U10687 ( .A(n9404), .ZN(n9405) );
  AOI21_X1 U10688 ( .B1(n9403), .B2(n9406), .A(n9405), .ZN(n9413) );
  NAND2_X1 U10689 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9509) );
  INV_X1 U10690 ( .A(n9509), .ZN(n9410) );
  INV_X1 U10691 ( .A(n9745), .ZN(n9407) );
  OAI22_X1 U10692 ( .A1(n9408), .A2(n9464), .B1(n9453), .B2(n9407), .ZN(n9409)
         );
  AOI211_X1 U10693 ( .C1(n9476), .C2(n9738), .A(n9410), .B(n9409), .ZN(n9412)
         );
  NAND2_X1 U10694 ( .A1(n9741), .A2(n9477), .ZN(n9411) );
  OAI211_X1 U10695 ( .C1(n9413), .C2(n9470), .A(n9412), .B(n9411), .ZN(
        P1_U3224) );
  INV_X1 U10696 ( .A(n9414), .ZN(n9419) );
  AOI21_X1 U10697 ( .B1(n9416), .B2(n9418), .A(n9415), .ZN(n9417) );
  AOI21_X1 U10698 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9424) );
  NAND2_X1 U10699 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9514) );
  OAI21_X1 U10700 ( .B1(n9464), .B2(n9754), .A(n9514), .ZN(n9422) );
  OAI22_X1 U10701 ( .A1(n9420), .A2(n9451), .B1(n9453), .B2(n9719), .ZN(n9421)
         );
  AOI211_X1 U10702 ( .C1(n9837), .C2(n9477), .A(n9422), .B(n9421), .ZN(n9423)
         );
  OAI21_X1 U10703 ( .B1(n9424), .B2(n9470), .A(n9423), .ZN(P1_U3226) );
  OAI21_X1 U10704 ( .B1(n9427), .B2(n9426), .A(n9425), .ZN(n9429) );
  NAND2_X1 U10705 ( .A1(n9429), .A2(n9428), .ZN(n9433) );
  AOI22_X1 U10706 ( .A1(n9476), .A2(n9627), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9432) );
  AOI22_X1 U10707 ( .A1(n9474), .A2(n9652), .B1(n9475), .B2(n9621), .ZN(n9431)
         );
  NAND2_X1 U10708 ( .A1(n9803), .A2(n9477), .ZN(n9430) );
  NAND4_X1 U10709 ( .A1(n9433), .A2(n9432), .A3(n9431), .A4(n9430), .ZN(
        P1_U3227) );
  XNOR2_X1 U10710 ( .A(n9435), .B(n9434), .ZN(n9436) );
  XNOR2_X1 U10711 ( .A(n9437), .B(n9436), .ZN(n9444) );
  OAI22_X1 U10712 ( .A1(n9451), .A2(n9454), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9438), .ZN(n9442) );
  INV_X1 U10713 ( .A(n9674), .ZN(n9439) );
  OAI22_X1 U10714 ( .A1(n9440), .A2(n9464), .B1(n9453), .B2(n9439), .ZN(n9441)
         );
  AOI211_X1 U10715 ( .C1(n9823), .C2(n9477), .A(n9442), .B(n9441), .ZN(n9443)
         );
  OAI21_X1 U10716 ( .B1(n9444), .B2(n9470), .A(n9443), .ZN(P1_U3231) );
  NAND2_X1 U10717 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  XOR2_X1 U10718 ( .A(n9448), .B(n9447), .Z(n9458) );
  OAI22_X1 U10719 ( .A1(n9451), .A2(n9450), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9449), .ZN(n9456) );
  INV_X1 U10720 ( .A(n9646), .ZN(n9452) );
  OAI22_X1 U10721 ( .A1(n9454), .A2(n9464), .B1(n9453), .B2(n9452), .ZN(n9455)
         );
  AOI211_X1 U10722 ( .C1(n9812), .C2(n9477), .A(n9456), .B(n9455), .ZN(n9457)
         );
  OAI21_X1 U10723 ( .B1(n9458), .B2(n9470), .A(n9457), .ZN(P1_U3233) );
  NAND2_X1 U10724 ( .A1(n9460), .A2(n9459), .ZN(n9461) );
  XOR2_X1 U10725 ( .A(n9462), .B(n9461), .Z(n9468) );
  AOI22_X1 U10726 ( .A1(n9476), .A2(n9710), .B1(n9475), .B2(n9702), .ZN(n9463)
         );
  NAND2_X1 U10727 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10031)
         );
  OAI211_X1 U10728 ( .C1(n9465), .C2(n9464), .A(n9463), .B(n10031), .ZN(n9466)
         );
  AOI21_X1 U10729 ( .B1(n9832), .B2(n9477), .A(n9466), .ZN(n9467) );
  OAI21_X1 U10730 ( .B1(n9468), .B2(n9470), .A(n9467), .ZN(P1_U3236) );
  AOI21_X1 U10731 ( .B1(n9469), .B2(n9471), .A(n9470), .ZN(n9473) );
  NAND2_X1 U10732 ( .A1(n9473), .A2(n9472), .ZN(n9481) );
  AOI22_X1 U10733 ( .A1(n9474), .A2(n9627), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9480) );
  AOI22_X1 U10734 ( .A1(n9476), .A2(n9600), .B1(n9475), .B2(n9591), .ZN(n9479)
         );
  NAND2_X1 U10735 ( .A1(n9792), .A2(n9477), .ZN(n9478) );
  NAND4_X1 U10736 ( .A1(n9481), .A2(n9480), .A3(n9479), .A4(n9478), .ZN(
        P1_U3238) );
  MUX2_X1 U10737 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9482), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10738 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9483), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10739 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9568), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10740 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9576), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10741 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9600), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10742 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9614), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10743 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9627), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10744 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9640), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10745 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9652), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10746 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9665), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10747 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9680), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10748 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9693), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10749 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9710), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10750 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9726), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10751 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9738), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10752 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9727), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10753 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9736), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10754 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9484), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10755 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9485), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10756 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9486), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10757 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9487), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9488), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10759 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9489), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10760 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9490), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10761 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9491), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10762 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9492), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10763 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9493), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10764 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9494), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10765 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9495), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10766 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9496), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10767 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6391), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10768 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n5941), .S(P1_U4006), .Z(
        P1_U3555) );
  NOR2_X1 U10769 ( .A1(n9497), .A2(n9503), .ZN(n9499) );
  NOR2_X1 U10770 ( .A1(n9515), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9500) );
  AOI21_X1 U10771 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9515), .A(n9500), .ZN(
        n9501) );
  AOI211_X1 U10772 ( .C1(n4564), .C2(n9501), .A(n9516), .B(n10032), .ZN(n9513)
         );
  NOR2_X1 U10773 ( .A1(n9503), .A2(n9502), .ZN(n9505) );
  NOR2_X1 U10774 ( .A1(n9505), .A2(n9504), .ZN(n9508) );
  NOR2_X1 U10775 ( .A1(n9515), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9506) );
  AOI21_X1 U10776 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9515), .A(n9506), .ZN(
        n9507) );
  NOR2_X1 U10777 ( .A1(n9508), .A2(n9507), .ZN(n9522) );
  AOI211_X1 U10778 ( .C1(n9508), .C2(n9507), .A(n9522), .B(n9982), .ZN(n9512)
         );
  NAND2_X1 U10779 ( .A1(n9999), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9510) );
  OAI211_X1 U10780 ( .C1(n9515), .C2(n9971), .A(n9510), .B(n9509), .ZN(n9511)
         );
  OR3_X1 U10781 ( .A1(n9513), .A2(n9512), .A3(n9511), .ZN(P1_U3257) );
  INV_X1 U10782 ( .A(n9524), .ZN(n9538) );
  INV_X1 U10783 ( .A(n9514), .ZN(n9521) );
  INV_X1 U10784 ( .A(n9515), .ZN(n9523) );
  AOI21_X1 U10785 ( .B1(n9523), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9516), .ZN(
        n9519) );
  NAND2_X1 U10786 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9538), .ZN(n9517) );
  OAI21_X1 U10787 ( .B1(n9538), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9517), .ZN(
        n9518) );
  NOR2_X1 U10788 ( .A1(n9519), .A2(n9518), .ZN(n9537) );
  AOI211_X1 U10789 ( .C1(n9519), .C2(n9518), .A(n9537), .B(n10032), .ZN(n9520)
         );
  AOI211_X1 U10790 ( .C1(n9538), .C2(n10038), .A(n9521), .B(n9520), .ZN(n9530)
         );
  AOI21_X1 U10791 ( .B1(n9523), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9522), .ZN(
        n9527) );
  MUX2_X1 U10792 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9525), .S(n9524), .Z(n9526) );
  NOR2_X1 U10793 ( .A1(n9527), .A2(n9526), .ZN(n9531) );
  AOI211_X1 U10794 ( .C1(n9527), .C2(n9526), .A(n9531), .B(n9982), .ZN(n9528)
         );
  AOI21_X1 U10795 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n9999), .A(n9528), .ZN(
        n9529) );
  NAND2_X1 U10796 ( .A1(n9530), .A2(n9529), .ZN(P1_U3258) );
  XNOR2_X1 U10797 ( .A(n9539), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10041) );
  AOI21_X1 U10798 ( .B1(n9538), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9531), .ZN(
        n10040) );
  NAND2_X1 U10799 ( .A1(n10041), .A2(n10040), .ZN(n9534) );
  INV_X1 U10800 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U10801 ( .A1(n9539), .A2(n9532), .ZN(n9533) );
  NAND2_X1 U10802 ( .A1(n9534), .A2(n9533), .ZN(n9536) );
  XNOR2_X1 U10803 ( .A(n9536), .B(n9535), .ZN(n9547) );
  INV_X1 U10804 ( .A(n9547), .ZN(n9543) );
  INV_X1 U10805 ( .A(n9539), .ZN(n10039) );
  NAND2_X1 U10806 ( .A1(n10039), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9540) );
  OAI21_X1 U10807 ( .B1(n10039), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9540), .ZN(
        n10034) );
  NOR2_X1 U10808 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U10809 ( .A(n9540), .ZN(n9541) );
  NOR2_X1 U10810 ( .A1(n10033), .A2(n9541), .ZN(n9542) );
  XNOR2_X1 U10811 ( .A(n9542), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9545) );
  INV_X1 U10812 ( .A(n10032), .ZN(n10021) );
  AOI22_X1 U10813 ( .A1(n10043), .A2(n9543), .B1(n9545), .B2(n10021), .ZN(
        n9549) );
  OAI21_X1 U10814 ( .B1(n9545), .B2(n9544), .A(n9971), .ZN(n9546) );
  AOI21_X1 U10815 ( .B1(n10043), .B2(n9547), .A(n9546), .ZN(n9548) );
  MUX2_X1 U10816 ( .A(n9549), .B(n9548), .S(n10054), .Z(n9551) );
  OAI211_X1 U10817 ( .C1(n4877), .C2(n10046), .A(n9551), .B(n9550), .ZN(
        P1_U3260) );
  AOI21_X1 U10818 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9906) );
  NAND2_X1 U10819 ( .A1(n9906), .A2(n9770), .ZN(n9557) );
  AOI21_X1 U10820 ( .B1(n10078), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9555), .ZN(
        n9556) );
  OAI211_X1 U10821 ( .C1(n9904), .C2(n9766), .A(n9557), .B(n9556), .ZN(
        P1_U3262) );
  AOI21_X1 U10822 ( .B1(n9567), .B2(n9559), .A(n9558), .ZN(n9560) );
  INV_X1 U10823 ( .A(n9560), .ZN(n9786) );
  AOI21_X1 U10824 ( .B1(n9782), .B2(n9580), .A(n4789), .ZN(n9783) );
  INV_X1 U10825 ( .A(n9782), .ZN(n9564) );
  AOI22_X1 U10826 ( .A1(n10078), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9562), 
        .B2(n10074), .ZN(n9563) );
  OAI21_X1 U10827 ( .B1(n9564), .B2(n9766), .A(n9563), .ZN(n9571) );
  OAI21_X1 U10828 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9569) );
  AOI222_X1 U10829 ( .A1(n10061), .A2(n9569), .B1(n9568), .B2(n9737), .C1(
        n9600), .C2(n9735), .ZN(n9785) );
  NOR2_X1 U10830 ( .A1(n9785), .A2(n10078), .ZN(n9570) );
  AOI211_X1 U10831 ( .C1(n9783), .C2(n9770), .A(n9571), .B(n9570), .ZN(n9572)
         );
  OAI21_X1 U10832 ( .B1(n9786), .B2(n9750), .A(n9572), .ZN(P1_U3263) );
  XNOR2_X1 U10833 ( .A(n9574), .B(n9573), .ZN(n9791) );
  OAI21_X1 U10834 ( .B1(n4527), .B2(n9575), .A(n10061), .ZN(n9579) );
  AOI22_X1 U10835 ( .A1(n9735), .A2(n9614), .B1(n9576), .B2(n9737), .ZN(n9577)
         );
  OAI21_X1 U10836 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9787) );
  INV_X1 U10837 ( .A(n9590), .ZN(n9582) );
  INV_X1 U10838 ( .A(n9580), .ZN(n9581) );
  AOI211_X1 U10839 ( .C1(n9789), .C2(n9582), .A(n10132), .B(n9581), .ZN(n9788)
         );
  NAND2_X1 U10840 ( .A1(n9788), .A2(n9697), .ZN(n9585) );
  AOI22_X1 U10841 ( .A1(n10078), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9583), 
        .B2(n10074), .ZN(n9584) );
  OAI211_X1 U10842 ( .C1(n9586), .C2(n9766), .A(n9585), .B(n9584), .ZN(n9587)
         );
  AOI21_X1 U10843 ( .B1(n9787), .B2(n10075), .A(n9587), .ZN(n9588) );
  OAI21_X1 U10844 ( .B1(n9791), .B2(n9750), .A(n9588), .ZN(P1_U3264) );
  XOR2_X1 U10845 ( .A(n9598), .B(n9589), .Z(n9796) );
  AOI21_X1 U10846 ( .B1(n9792), .B2(n9604), .A(n9590), .ZN(n9793) );
  AOI22_X1 U10847 ( .A1(n10078), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9591), 
        .B2(n10074), .ZN(n9592) );
  OAI21_X1 U10848 ( .B1(n9593), .B2(n9766), .A(n9592), .ZN(n9602) );
  INV_X1 U10849 ( .A(n9594), .ZN(n9595) );
  NOR2_X1 U10850 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  XOR2_X1 U10851 ( .A(n9598), .B(n9597), .Z(n9599) );
  AOI222_X1 U10852 ( .A1(n9627), .A2(n9735), .B1(n9600), .B2(n9737), .C1(
        n10061), .C2(n9599), .ZN(n9795) );
  NOR2_X1 U10853 ( .A1(n9795), .A2(n10078), .ZN(n9601) );
  AOI211_X1 U10854 ( .C1(n9793), .C2(n9770), .A(n9602), .B(n9601), .ZN(n9603)
         );
  OAI21_X1 U10855 ( .B1(n9750), .B2(n9796), .A(n9603), .ZN(P1_U3265) );
  XOR2_X1 U10856 ( .A(n9612), .B(n4548), .Z(n9801) );
  AOI211_X1 U10857 ( .C1(n9798), .C2(n9619), .A(n10132), .B(n4788), .ZN(n9797)
         );
  INV_X1 U10858 ( .A(n9798), .ZN(n9607) );
  AOI22_X1 U10859 ( .A1(n10078), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9605), 
        .B2(n10074), .ZN(n9606) );
  OAI21_X1 U10860 ( .B1(n9607), .B2(n9766), .A(n9606), .ZN(n9616) );
  INV_X1 U10861 ( .A(n9608), .ZN(n9609) );
  NOR2_X1 U10862 ( .A1(n9610), .A2(n9609), .ZN(n9611) );
  XOR2_X1 U10863 ( .A(n9612), .B(n9611), .Z(n9613) );
  AOI222_X1 U10864 ( .A1(n9640), .A2(n9735), .B1(n9614), .B2(n9737), .C1(
        n10061), .C2(n9613), .ZN(n9800) );
  NOR2_X1 U10865 ( .A1(n9800), .A2(n10078), .ZN(n9615) );
  AOI211_X1 U10866 ( .C1(n9697), .C2(n9797), .A(n9616), .B(n9615), .ZN(n9617)
         );
  OAI21_X1 U10867 ( .B1(n9750), .B2(n9801), .A(n9617), .ZN(P1_U3266) );
  XOR2_X1 U10868 ( .A(n9625), .B(n9618), .Z(n9806) );
  INV_X1 U10869 ( .A(n9632), .ZN(n9620) );
  AOI211_X1 U10870 ( .C1(n9803), .C2(n9620), .A(n10132), .B(n4784), .ZN(n9802)
         );
  AOI22_X1 U10871 ( .A1(n10078), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9621), 
        .B2(n10074), .ZN(n9622) );
  OAI21_X1 U10872 ( .B1(n9623), .B2(n9766), .A(n9622), .ZN(n9629) );
  XOR2_X1 U10873 ( .A(n9625), .B(n9624), .Z(n9626) );
  AOI222_X1 U10874 ( .A1(n9652), .A2(n9735), .B1(n9627), .B2(n9737), .C1(
        n10061), .C2(n9626), .ZN(n9805) );
  NOR2_X1 U10875 ( .A1(n9805), .A2(n10078), .ZN(n9628) );
  AOI211_X1 U10876 ( .C1(n9802), .C2(n9697), .A(n9629), .B(n9628), .ZN(n9630)
         );
  OAI21_X1 U10877 ( .B1(n9750), .B2(n9806), .A(n9630), .ZN(P1_U3267) );
  XNOR2_X1 U10878 ( .A(n9631), .B(n9638), .ZN(n9811) );
  INV_X1 U10879 ( .A(n9645), .ZN(n9633) );
  AOI21_X1 U10880 ( .B1(n9807), .B2(n9633), .A(n9632), .ZN(n9808) );
  AOI22_X1 U10881 ( .A1(n10078), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9634), 
        .B2(n10074), .ZN(n9635) );
  OAI21_X1 U10882 ( .B1(n9636), .B2(n9766), .A(n9635), .ZN(n9642) );
  XOR2_X1 U10883 ( .A(n9638), .B(n9637), .Z(n9639) );
  AOI222_X1 U10884 ( .A1(n9665), .A2(n9735), .B1(n9640), .B2(n9737), .C1(
        n10061), .C2(n9639), .ZN(n9810) );
  NOR2_X1 U10885 ( .A1(n9810), .A2(n10078), .ZN(n9641) );
  AOI211_X1 U10886 ( .C1(n9808), .C2(n9770), .A(n9642), .B(n9641), .ZN(n9643)
         );
  OAI21_X1 U10887 ( .B1(n9750), .B2(n9811), .A(n9643), .ZN(P1_U3268) );
  XNOR2_X1 U10888 ( .A(n9644), .B(n9651), .ZN(n9816) );
  AOI21_X1 U10889 ( .B1(n9812), .B2(n9658), .A(n9645), .ZN(n9813) );
  AOI22_X1 U10890 ( .A1(n10078), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9646), 
        .B2(n10074), .ZN(n9647) );
  OAI21_X1 U10891 ( .B1(n9648), .B2(n9766), .A(n9647), .ZN(n9655) );
  OAI21_X1 U10892 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9653) );
  AOI222_X1 U10893 ( .A1(n10061), .A2(n9653), .B1(n9652), .B2(n9737), .C1(
        n9680), .C2(n9735), .ZN(n9815) );
  NOR2_X1 U10894 ( .A1(n9815), .A2(n10078), .ZN(n9654) );
  AOI211_X1 U10895 ( .C1(n9813), .C2(n9770), .A(n9655), .B(n9654), .ZN(n9656)
         );
  OAI21_X1 U10896 ( .B1(n9750), .B2(n9816), .A(n9656), .ZN(P1_U3269) );
  XNOR2_X1 U10897 ( .A(n9657), .B(n9663), .ZN(n9821) );
  INV_X1 U10898 ( .A(n9658), .ZN(n9659) );
  AOI211_X1 U10899 ( .C1(n9818), .C2(n9671), .A(n10132), .B(n9659), .ZN(n9817)
         );
  INV_X1 U10900 ( .A(n9818), .ZN(n9662) );
  AOI22_X1 U10901 ( .A1(n10078), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9660), 
        .B2(n10074), .ZN(n9661) );
  OAI21_X1 U10902 ( .B1(n9662), .B2(n9766), .A(n9661), .ZN(n9668) );
  XNOR2_X1 U10903 ( .A(n9664), .B(n9663), .ZN(n9666) );
  AOI222_X1 U10904 ( .A1(n10061), .A2(n9666), .B1(n9665), .B2(n9737), .C1(
        n9693), .C2(n9735), .ZN(n9820) );
  NOR2_X1 U10905 ( .A1(n9820), .A2(n10078), .ZN(n9667) );
  AOI211_X1 U10906 ( .C1(n9817), .C2(n9697), .A(n9668), .B(n9667), .ZN(n9669)
         );
  OAI21_X1 U10907 ( .B1(n9750), .B2(n9821), .A(n9669), .ZN(P1_U3270) );
  XOR2_X1 U10908 ( .A(n9670), .B(n9677), .Z(n9826) );
  INV_X1 U10909 ( .A(n9685), .ZN(n9673) );
  INV_X1 U10910 ( .A(n9671), .ZN(n9672) );
  AOI211_X1 U10911 ( .C1(n9823), .C2(n9673), .A(n10132), .B(n9672), .ZN(n9822)
         );
  AOI22_X1 U10912 ( .A1(n10078), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9674), 
        .B2(n10074), .ZN(n9675) );
  OAI21_X1 U10913 ( .B1(n9676), .B2(n9766), .A(n9675), .ZN(n9682) );
  XNOR2_X1 U10914 ( .A(n9678), .B(n9677), .ZN(n9679) );
  AOI222_X1 U10915 ( .A1(n9710), .A2(n9735), .B1(n9680), .B2(n9737), .C1(
        n10061), .C2(n9679), .ZN(n9825) );
  NOR2_X1 U10916 ( .A1(n9825), .A2(n10078), .ZN(n9681) );
  AOI211_X1 U10917 ( .C1(n9822), .C2(n9697), .A(n9682), .B(n9681), .ZN(n9683)
         );
  OAI21_X1 U10918 ( .B1(n9750), .B2(n9826), .A(n9683), .ZN(P1_U3271) );
  XNOR2_X1 U10919 ( .A(n9684), .B(n9692), .ZN(n9831) );
  AOI211_X1 U10920 ( .C1(n9828), .C2(n9700), .A(n10132), .B(n9685), .ZN(n9827)
         );
  INV_X1 U10921 ( .A(n9686), .ZN(n9687) );
  AOI22_X1 U10922 ( .A1(n10078), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9687), 
        .B2(n10074), .ZN(n9688) );
  OAI21_X1 U10923 ( .B1(n9689), .B2(n9766), .A(n9688), .ZN(n9696) );
  OAI21_X1 U10924 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9694) );
  AOI222_X1 U10925 ( .A1(n10061), .A2(n9694), .B1(n9693), .B2(n9737), .C1(
        n9726), .C2(n9735), .ZN(n9830) );
  NOR2_X1 U10926 ( .A1(n9830), .A2(n10078), .ZN(n9695) );
  AOI211_X1 U10927 ( .C1(n9827), .C2(n9697), .A(n9696), .B(n9695), .ZN(n9698)
         );
  OAI21_X1 U10928 ( .B1(n9750), .B2(n9831), .A(n9698), .ZN(P1_U3272) );
  XNOR2_X1 U10929 ( .A(n9699), .B(n9709), .ZN(n9836) );
  INV_X1 U10930 ( .A(n9700), .ZN(n9701) );
  AOI21_X1 U10931 ( .B1(n9832), .B2(n9717), .A(n9701), .ZN(n9833) );
  INV_X1 U10932 ( .A(n9832), .ZN(n9704) );
  AOI22_X1 U10933 ( .A1(n10078), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9702), 
        .B2(n10074), .ZN(n9703) );
  OAI21_X1 U10934 ( .B1(n9704), .B2(n9766), .A(n9703), .ZN(n9713) );
  INV_X1 U10935 ( .A(n9705), .ZN(n9706) );
  NOR2_X1 U10936 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  XOR2_X1 U10937 ( .A(n9709), .B(n9708), .Z(n9711) );
  AOI222_X1 U10938 ( .A1(n10061), .A2(n9711), .B1(n9710), .B2(n9737), .C1(
        n9738), .C2(n9735), .ZN(n9835) );
  NOR2_X1 U10939 ( .A1(n9835), .A2(n10078), .ZN(n9712) );
  AOI211_X1 U10940 ( .C1(n9833), .C2(n9770), .A(n9713), .B(n9712), .ZN(n9714)
         );
  OAI21_X1 U10941 ( .B1(n9750), .B2(n9836), .A(n9714), .ZN(P1_U3273) );
  XNOR2_X1 U10942 ( .A(n9715), .B(n9723), .ZN(n9841) );
  INV_X1 U10943 ( .A(n9716), .ZN(n9742) );
  INV_X1 U10944 ( .A(n9717), .ZN(n9718) );
  AOI21_X1 U10945 ( .B1(n9837), .B2(n9742), .A(n9718), .ZN(n9838) );
  INV_X1 U10946 ( .A(n9719), .ZN(n9720) );
  AOI22_X1 U10947 ( .A1(n10078), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10074), 
        .B2(n9720), .ZN(n9721) );
  OAI21_X1 U10948 ( .B1(n9722), .B2(n9766), .A(n9721), .ZN(n9729) );
  XNOR2_X1 U10949 ( .A(n9724), .B(n9723), .ZN(n9725) );
  AOI222_X1 U10950 ( .A1(n9727), .A2(n9735), .B1(n9726), .B2(n9737), .C1(
        n10061), .C2(n9725), .ZN(n9840) );
  NOR2_X1 U10951 ( .A1(n9840), .A2(n10078), .ZN(n9728) );
  AOI211_X1 U10952 ( .C1(n9838), .C2(n9770), .A(n9729), .B(n9728), .ZN(n9730)
         );
  OAI21_X1 U10953 ( .B1(n9750), .B2(n9841), .A(n9730), .ZN(P1_U3274) );
  XNOR2_X1 U10954 ( .A(n9731), .B(n4926), .ZN(n9912) );
  INV_X1 U10955 ( .A(n9912), .ZN(n9751) );
  OAI21_X1 U10956 ( .B1(n4926), .B2(n9733), .A(n9732), .ZN(n9734) );
  NAND2_X1 U10957 ( .A1(n9734), .A2(n10061), .ZN(n9740) );
  AOI22_X1 U10958 ( .A1(n9738), .A2(n9737), .B1(n9736), .B2(n9735), .ZN(n9739)
         );
  NAND2_X1 U10959 ( .A1(n9740), .A2(n9739), .ZN(n9911) );
  INV_X1 U10960 ( .A(n9741), .ZN(n9909) );
  INV_X1 U10961 ( .A(n9763), .ZN(n9743) );
  OAI211_X1 U10962 ( .C1(n9909), .C2(n9743), .A(n9742), .B(n10140), .ZN(n9908)
         );
  NOR2_X1 U10963 ( .A1(n9908), .A2(n9744), .ZN(n9748) );
  AOI22_X1 U10964 ( .A1(n10078), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9745), 
        .B2(n10074), .ZN(n9746) );
  OAI21_X1 U10965 ( .B1(n9909), .B2(n9766), .A(n9746), .ZN(n9747) );
  AOI211_X1 U10966 ( .C1(n9911), .C2(n10075), .A(n9748), .B(n9747), .ZN(n9749)
         );
  OAI21_X1 U10967 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(P1_U3275) );
  XNOR2_X1 U10968 ( .A(n9752), .B(n9755), .ZN(n9759) );
  OAI22_X1 U10969 ( .A1(n9754), .A2(n10058), .B1(n9753), .B2(n10056), .ZN(
        n9758) );
  XNOR2_X1 U10970 ( .A(n9756), .B(n9755), .ZN(n9847) );
  NOR2_X1 U10971 ( .A1(n9847), .A2(n10064), .ZN(n9757) );
  AOI211_X1 U10972 ( .C1(n9759), .C2(n10061), .A(n9758), .B(n9757), .ZN(n9846)
         );
  NAND2_X1 U10973 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  NAND2_X1 U10974 ( .A1(n9763), .A2(n9762), .ZN(n9843) );
  INV_X1 U10975 ( .A(n9843), .ZN(n9771) );
  AOI22_X1 U10976 ( .A1(n10078), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9764), 
        .B2(n10074), .ZN(n9765) );
  OAI21_X1 U10977 ( .B1(n9842), .B2(n9766), .A(n9765), .ZN(n9769) );
  NOR2_X1 U10978 ( .A1(n9847), .A2(n9767), .ZN(n9768) );
  AOI211_X1 U10979 ( .C1(n9771), .C2(n9770), .A(n9769), .B(n9768), .ZN(n9772)
         );
  OAI21_X1 U10980 ( .B1(n9846), .B2(n10078), .A(n9772), .ZN(P1_U3276) );
  NAND2_X1 U10981 ( .A1(n9773), .A2(n10140), .ZN(n9774) );
  OAI211_X1 U10982 ( .C1(n10130), .C2(n9775), .A(n9774), .B(n9903), .ZN(n9855)
         );
  AND2_X2 U10983 ( .A1(n9776), .A2(n9871), .ZN(n10169) );
  MUX2_X1 U10984 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9855), .S(n10169), .Z(
        P1_U3554) );
  AOI22_X1 U10985 ( .A1(n9778), .A2(n10140), .B1(n10139), .B2(n9777), .ZN(
        n9779) );
  MUX2_X1 U10986 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9856), .S(n10169), .Z(
        P1_U3552) );
  AOI22_X1 U10987 ( .A1(n9783), .A2(n10140), .B1(n10139), .B2(n9782), .ZN(
        n9784) );
  OAI211_X1 U10988 ( .C1(n9786), .C2(n9883), .A(n9785), .B(n9784), .ZN(n9857)
         );
  MUX2_X1 U10989 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9857), .S(n10169), .Z(
        P1_U3551) );
  AOI211_X1 U10990 ( .C1(n10139), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9790)
         );
  OAI21_X1 U10991 ( .B1(n9791), .B2(n9883), .A(n9790), .ZN(n9858) );
  MUX2_X1 U10992 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9858), .S(n10169), .Z(
        P1_U3550) );
  AOI22_X1 U10993 ( .A1(n9793), .A2(n10140), .B1(n10139), .B2(n9792), .ZN(
        n9794) );
  OAI211_X1 U10994 ( .C1(n9796), .C2(n9883), .A(n9795), .B(n9794), .ZN(n9859)
         );
  MUX2_X1 U10995 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9859), .S(n10169), .Z(
        P1_U3549) );
  AOI21_X1 U10996 ( .B1(n10139), .B2(n9798), .A(n9797), .ZN(n9799) );
  OAI211_X1 U10997 ( .C1(n9801), .C2(n9883), .A(n9800), .B(n9799), .ZN(n9860)
         );
  MUX2_X1 U10998 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9860), .S(n10169), .Z(
        P1_U3548) );
  AOI21_X1 U10999 ( .B1(n10139), .B2(n9803), .A(n9802), .ZN(n9804) );
  OAI211_X1 U11000 ( .C1(n9806), .C2(n9883), .A(n9805), .B(n9804), .ZN(n9861)
         );
  MUX2_X1 U11001 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9861), .S(n10169), .Z(
        P1_U3547) );
  AOI22_X1 U11002 ( .A1(n9808), .A2(n10140), .B1(n10139), .B2(n9807), .ZN(
        n9809) );
  OAI211_X1 U11003 ( .C1(n9811), .C2(n9883), .A(n9810), .B(n9809), .ZN(n9862)
         );
  MUX2_X1 U11004 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9862), .S(n10169), .Z(
        P1_U3546) );
  AOI22_X1 U11005 ( .A1(n9813), .A2(n10140), .B1(n10139), .B2(n9812), .ZN(
        n9814) );
  OAI211_X1 U11006 ( .C1(n9816), .C2(n9883), .A(n9815), .B(n9814), .ZN(n9863)
         );
  MUX2_X1 U11007 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9863), .S(n10169), .Z(
        P1_U3545) );
  AOI21_X1 U11008 ( .B1(n10139), .B2(n9818), .A(n9817), .ZN(n9819) );
  OAI211_X1 U11009 ( .C1(n9821), .C2(n9883), .A(n9820), .B(n9819), .ZN(n9864)
         );
  MUX2_X1 U11010 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9864), .S(n10169), .Z(
        P1_U3544) );
  AOI21_X1 U11011 ( .B1(n10139), .B2(n9823), .A(n9822), .ZN(n9824) );
  OAI211_X1 U11012 ( .C1(n9826), .C2(n9883), .A(n9825), .B(n9824), .ZN(n9865)
         );
  MUX2_X1 U11013 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9865), .S(n10169), .Z(
        P1_U3543) );
  AOI21_X1 U11014 ( .B1(n10139), .B2(n9828), .A(n9827), .ZN(n9829) );
  OAI211_X1 U11015 ( .C1(n9831), .C2(n9883), .A(n9830), .B(n9829), .ZN(n9866)
         );
  MUX2_X1 U11016 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9866), .S(n10169), .Z(
        P1_U3542) );
  AOI22_X1 U11017 ( .A1(n9833), .A2(n10140), .B1(n10139), .B2(n9832), .ZN(
        n9834) );
  OAI211_X1 U11018 ( .C1(n9836), .C2(n9883), .A(n9835), .B(n9834), .ZN(n9867)
         );
  MUX2_X1 U11019 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9867), .S(n10169), .Z(
        P1_U3541) );
  AOI22_X1 U11020 ( .A1(n9838), .A2(n10140), .B1(n10139), .B2(n9837), .ZN(
        n9839) );
  OAI211_X1 U11021 ( .C1(n9841), .C2(n9883), .A(n9840), .B(n9839), .ZN(n9868)
         );
  MUX2_X1 U11022 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9868), .S(n10169), .Z(
        P1_U3540) );
  OAI22_X1 U11023 ( .A1(n9843), .A2(n10132), .B1(n9842), .B2(n10130), .ZN(
        n9844) );
  INV_X1 U11024 ( .A(n9844), .ZN(n9845) );
  OAI211_X1 U11025 ( .C1(n10145), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9869)
         );
  MUX2_X1 U11026 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9869), .S(n10169), .Z(
        P1_U3538) );
  AOI22_X1 U11027 ( .A1(n9849), .A2(n10140), .B1(n10139), .B2(n9848), .ZN(
        n9850) );
  OAI211_X1 U11028 ( .C1(n10145), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9870)
         );
  MUX2_X1 U11029 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9870), .S(n10169), .Z(
        P1_U3536) );
  MUX2_X1 U11030 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9853), .S(n10169), .Z(
        P1_U3534) );
  MUX2_X1 U11031 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9854), .S(n10169), .Z(
        P1_U3523) );
  MUX2_X1 U11032 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9855), .S(n10150), .Z(
        P1_U3522) );
  MUX2_X1 U11033 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9856), .S(n10150), .Z(
        P1_U3520) );
  MUX2_X1 U11034 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9857), .S(n10150), .Z(
        P1_U3519) );
  MUX2_X1 U11035 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9858), .S(n10150), .Z(
        P1_U3518) );
  MUX2_X1 U11036 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9859), .S(n10150), .Z(
        P1_U3517) );
  MUX2_X1 U11037 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9860), .S(n10150), .Z(
        P1_U3516) );
  MUX2_X1 U11038 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9861), .S(n10150), .Z(
        P1_U3515) );
  MUX2_X1 U11039 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9862), .S(n10150), .Z(
        P1_U3514) );
  MUX2_X1 U11040 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9863), .S(n10150), .Z(
        P1_U3513) );
  MUX2_X1 U11041 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9864), .S(n10150), .Z(
        P1_U3512) );
  MUX2_X1 U11042 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9865), .S(n10150), .Z(
        P1_U3511) );
  MUX2_X1 U11043 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9866), .S(n10150), .Z(
        P1_U3510) );
  MUX2_X1 U11044 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9867), .S(n10150), .Z(
        P1_U3508) );
  MUX2_X1 U11045 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9868), .S(n10150), .Z(
        P1_U3505) );
  MUX2_X1 U11046 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9869), .S(n10150), .Z(
        P1_U3499) );
  MUX2_X1 U11047 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9870), .S(n10150), .Z(
        P1_U3493) );
  MUX2_X1 U11048 ( .A(n9871), .B(P1_D_REG_0__SCAN_IN), .S(n10090), .Z(P1_U3440) );
  NOR4_X1 U11049 ( .A1(n9873), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9872), .ZN(n9874) );
  AOI21_X1 U11050 ( .B1(n9875), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9874), .ZN(
        n9876) );
  OAI21_X1 U11051 ( .B1(n9877), .B2(n9881), .A(n9876), .ZN(P1_U3322) );
  INV_X1 U11052 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9878) );
  OAI222_X1 U11053 ( .A1(n9881), .A2(n9880), .B1(n9879), .B2(P1_U3084), .C1(
        n9878), .C2(n8383), .ZN(P1_U3324) );
  MUX2_X1 U11054 ( .A(n9882), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11055 ( .A(n9883), .ZN(n10136) );
  NAND3_X1 U11056 ( .A1(n9886), .A2(n9885), .A3(n9884), .ZN(n9887) );
  AOI21_X1 U11057 ( .B1(n10136), .B2(n9888), .A(n9887), .ZN(n9890) );
  AOI22_X1 U11058 ( .A1(n10150), .A2(n9890), .B1(n5576), .B2(n10149), .ZN(
        P1_U3484) );
  AOI22_X1 U11059 ( .A1(n10169), .A2(n9890), .B1(n9889), .B2(n10166), .ZN(
        P1_U3533) );
  INV_X1 U11060 ( .A(n9891), .ZN(n9893) );
  AOI22_X1 U11061 ( .A1(n10295), .A2(n9900), .B1(n8161), .B2(n10293), .ZN(
        P2_U3550) );
  OAI22_X1 U11062 ( .A1(n9896), .A2(n10261), .B1(n9895), .B2(n10275), .ZN(
        n9898) );
  AOI211_X1 U11063 ( .C1(n9899), .C2(n10279), .A(n9898), .B(n9897), .ZN(n9902)
         );
  AOI22_X1 U11064 ( .A1(n10295), .A2(n9902), .B1(n7625), .B2(n10293), .ZN(
        P2_U3534) );
  INV_X1 U11065 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U11066 ( .A1(n9320), .A2(n9902), .B1(n9901), .B2(n10281), .ZN(
        P2_U3493) );
  OAI21_X1 U11067 ( .B1(n9904), .B2(n10130), .A(n9903), .ZN(n9905) );
  AOI21_X1 U11068 ( .B1(n9906), .B2(n10140), .A(n9905), .ZN(n9924) );
  INV_X1 U11069 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9907) );
  AOI22_X1 U11070 ( .A1(n10169), .A2(n9924), .B1(n9907), .B2(n10166), .ZN(
        P1_U3553) );
  OAI21_X1 U11071 ( .B1(n9909), .B2(n10130), .A(n9908), .ZN(n9910) );
  AOI211_X1 U11072 ( .C1(n9912), .C2(n10136), .A(n9911), .B(n9910), .ZN(n9925)
         );
  INV_X1 U11073 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U11074 ( .A1(n10169), .A2(n9925), .B1(n9913), .B2(n10166), .ZN(
        P1_U3539) );
  OAI21_X1 U11075 ( .B1(n9915), .B2(n10130), .A(n9914), .ZN(n9916) );
  AOI211_X1 U11076 ( .C1(n9918), .C2(n10136), .A(n9917), .B(n9916), .ZN(n9926)
         );
  AOI22_X1 U11077 ( .A1(n10169), .A2(n9926), .B1(n6276), .B2(n10166), .ZN(
        P1_U3537) );
  OAI21_X1 U11078 ( .B1(n9920), .B2(n10130), .A(n9919), .ZN(n9921) );
  AOI211_X1 U11079 ( .C1(n9923), .C2(n10136), .A(n9922), .B(n9921), .ZN(n9927)
         );
  AOI22_X1 U11080 ( .A1(n10169), .A2(n9927), .B1(n6278), .B2(n10166), .ZN(
        P1_U3535) );
  AOI22_X1 U11081 ( .A1(n10150), .A2(n9924), .B1(n5269), .B2(n10149), .ZN(
        P1_U3521) );
  AOI22_X1 U11082 ( .A1(n10150), .A2(n9925), .B1(n5436), .B2(n10149), .ZN(
        P1_U3502) );
  AOI22_X1 U11083 ( .A1(n10150), .A2(n9926), .B1(n5452), .B2(n10149), .ZN(
        P1_U3496) );
  AOI22_X1 U11084 ( .A1(n10150), .A2(n9927), .B1(n5483), .B2(n10149), .ZN(
        P1_U3490) );
  XOR2_X1 U11085 ( .A(n9928), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11086 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11087 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10301) );
  OAI21_X1 U11088 ( .B1(n5925), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9929), .ZN(
        n9958) );
  AOI21_X1 U11089 ( .B1(n5925), .B2(n9930), .A(n9958), .ZN(n9931) );
  XNOR2_X1 U11090 ( .A(n9931), .B(n9957), .ZN(n9933) );
  AND2_X1 U11091 ( .A1(n9933), .A2(n9932), .ZN(n9934) );
  AOI21_X1 U11092 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .A(n9934), 
        .ZN(n9935) );
  OAI21_X1 U11093 ( .B1(n10301), .B2(n10046), .A(n9935), .ZN(P1_U3241) );
  AOI22_X1 U11094 ( .A1(n10038), .A2(n9936), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        P1_U3084), .ZN(n9945) );
  NAND2_X1 U11095 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9939) );
  AOI211_X1 U11096 ( .C1(n9939), .C2(n9938), .A(n9937), .B(n9982), .ZN(n9943)
         );
  AOI211_X1 U11097 ( .C1(n9956), .C2(n9941), .A(n9940), .B(n10032), .ZN(n9942)
         );
  AOI211_X1 U11098 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9999), .A(n9943), .B(
        n9942), .ZN(n9944) );
  NAND2_X1 U11099 ( .A1(n9945), .A2(n9944), .ZN(P1_U3242) );
  AOI22_X1 U11100 ( .A1(n10038), .A2(n9946), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n9962) );
  AOI211_X1 U11101 ( .C1(n9949), .C2(n9948), .A(n9947), .B(n9982), .ZN(n9954)
         );
  AOI211_X1 U11102 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n10032), .ZN(n9953)
         );
  AOI211_X1 U11103 ( .C1(P1_ADDR_REG_2__SCAN_IN), .C2(n9999), .A(n9954), .B(
        n9953), .ZN(n9961) );
  MUX2_X1 U11104 ( .A(n9956), .B(n9955), .S(n5925), .Z(n9960) );
  NAND2_X1 U11105 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  OAI211_X1 U11106 ( .C1(n9960), .C2(n5922), .A(P1_U4006), .B(n9959), .ZN(
        n9975) );
  NAND3_X1 U11107 ( .A1(n9962), .A2(n9961), .A3(n9975), .ZN(P1_U3243) );
  OAI21_X1 U11108 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9966) );
  AOI22_X1 U11109 ( .A1(n9999), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(n10021), .B2(
        n9966), .ZN(n9977) );
  OAI21_X1 U11110 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9974) );
  NOR2_X1 U11111 ( .A1(n9971), .A2(n9970), .ZN(n9972) );
  AOI211_X1 U11112 ( .C1(n10043), .C2(n9974), .A(n9973), .B(n9972), .ZN(n9976)
         );
  NAND3_X1 U11113 ( .A1(n9977), .A2(n9976), .A3(n9975), .ZN(P1_U3245) );
  AOI22_X1 U11114 ( .A1(n9999), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9978), .B2(
        n10038), .ZN(n9990) );
  OAI21_X1 U11115 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9988) );
  AOI211_X1 U11116 ( .C1(n9985), .C2(n9984), .A(n9983), .B(n9982), .ZN(n9986)
         );
  AOI211_X1 U11117 ( .C1(n10021), .C2(n9988), .A(n9987), .B(n9986), .ZN(n9989)
         );
  NAND2_X1 U11118 ( .A1(n9990), .A2(n9989), .ZN(P1_U3246) );
  AOI211_X1 U11119 ( .C1(n9993), .C2(n9992), .A(n10032), .B(n9991), .ZN(n9994)
         );
  AOI211_X1 U11120 ( .C1(n10038), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10002) );
  XNOR2_X1 U11121 ( .A(n9998), .B(n9997), .ZN(n10000) );
  AOI22_X1 U11122 ( .A1(n10043), .A2(n10000), .B1(n9999), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U11123 ( .A1(n10002), .A2(n10001), .ZN(P1_U3247) );
  AOI21_X1 U11124 ( .B1(n10038), .B2(n10004), .A(n10003), .ZN(n10014) );
  OAI21_X1 U11125 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(n10012) );
  OAI21_X1 U11126 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n10011) );
  AOI22_X1 U11127 ( .A1(n10012), .A2(n10021), .B1(n10043), .B2(n10011), .ZN(
        n10013) );
  OAI211_X1 U11128 ( .C1(n10046), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        P1_U3248) );
  OAI21_X1 U11129 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(n10022) );
  INV_X1 U11130 ( .A(n10019), .ZN(n10020) );
  AOI21_X1 U11131 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10029) );
  OAI21_X1 U11132 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10027) );
  AOI22_X1 U11133 ( .A1(n10027), .A2(n10043), .B1(n10026), .B2(n10038), .ZN(
        n10028) );
  OAI211_X1 U11134 ( .C1(n10030), .C2(n10046), .A(n10029), .B(n10028), .ZN(
        P1_U3252) );
  INV_X1 U11135 ( .A(n10031), .ZN(n10037) );
  AOI211_X1 U11136 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10036) );
  AOI211_X1 U11137 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10045) );
  XNOR2_X1 U11138 ( .A(n10041), .B(n10040), .ZN(n10042) );
  NAND2_X1 U11139 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  OAI211_X1 U11140 ( .C1(n10046), .C2(n10336), .A(n10045), .B(n10044), .ZN(
        P1_U3259) );
  XOR2_X1 U11141 ( .A(n6816), .B(n10047), .Z(n10065) );
  INV_X1 U11142 ( .A(n10065), .ZN(n10095) );
  INV_X1 U11143 ( .A(n10048), .ZN(n10049) );
  OAI211_X1 U11144 ( .C1(n10092), .C2(n10050), .A(n10049), .B(n10140), .ZN(
        n10091) );
  AOI22_X1 U11145 ( .A1(n10074), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n10052), 
        .B2(n10051), .ZN(n10053) );
  OAI21_X1 U11146 ( .B1(n10091), .B2(n10054), .A(n10053), .ZN(n10066) );
  XNOR2_X1 U11147 ( .A(n6816), .B(n10055), .ZN(n10062) );
  OAI22_X1 U11148 ( .A1(n10059), .A2(n10058), .B1(n10057), .B2(n10056), .ZN(
        n10060) );
  AOI21_X1 U11149 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10063) );
  OAI21_X1 U11150 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(n10093) );
  AOI211_X1 U11151 ( .C1(n10067), .C2(n10095), .A(n10066), .B(n10093), .ZN(
        n10068) );
  AOI22_X1 U11152 ( .A1(n10078), .A2(n5500), .B1(n10068), .B2(n10075), .ZN(
        P1_U3290) );
  NOR2_X1 U11153 ( .A1(n10070), .A2(n10069), .ZN(n10073) );
  INV_X1 U11154 ( .A(n10071), .ZN(n10072) );
  AOI211_X1 U11155 ( .C1(n10074), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10073), .B(
        n10072), .ZN(n10076) );
  AOI22_X1 U11156 ( .A1(n10078), .A2(n10077), .B1(n10076), .B2(n10075), .ZN(
        P1_U3291) );
  AND2_X1 U11157 ( .A1(n10080), .A2(n10079), .ZN(n10086) );
  INV_X1 U11158 ( .A(n10086), .ZN(n10087) );
  AND2_X1 U11159 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10087), .ZN(P1_U3292) );
  AND2_X1 U11160 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10087), .ZN(P1_U3293) );
  NOR2_X1 U11161 ( .A1(n10086), .A2(n10081), .ZN(P1_U3294) );
  AND2_X1 U11162 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10087), .ZN(P1_U3295) );
  NOR2_X1 U11163 ( .A1(n10086), .A2(n10082), .ZN(P1_U3296) );
  AND2_X1 U11164 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10087), .ZN(P1_U3297) );
  AND2_X1 U11165 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10087), .ZN(P1_U3298) );
  AND2_X1 U11166 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10087), .ZN(P1_U3299) );
  AND2_X1 U11167 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10087), .ZN(P1_U3300) );
  AND2_X1 U11168 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10087), .ZN(P1_U3301) );
  AND2_X1 U11169 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10087), .ZN(P1_U3302) );
  AND2_X1 U11170 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10087), .ZN(P1_U3303) );
  AND2_X1 U11171 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10087), .ZN(P1_U3304) );
  AND2_X1 U11172 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10087), .ZN(P1_U3305) );
  AND2_X1 U11173 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10087), .ZN(P1_U3306) );
  AND2_X1 U11174 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10087), .ZN(P1_U3307) );
  AND2_X1 U11175 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10087), .ZN(P1_U3308) );
  NOR2_X1 U11176 ( .A1(n10086), .A2(n10083), .ZN(P1_U3309) );
  AND2_X1 U11177 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10087), .ZN(P1_U3310) );
  NOR2_X1 U11178 ( .A1(n10086), .A2(n10084), .ZN(P1_U3311) );
  AND2_X1 U11179 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10087), .ZN(P1_U3312) );
  AND2_X1 U11180 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10087), .ZN(P1_U3313) );
  AND2_X1 U11181 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10087), .ZN(P1_U3314) );
  NOR2_X1 U11182 ( .A1(n10086), .A2(n10085), .ZN(P1_U3315) );
  AND2_X1 U11183 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10087), .ZN(P1_U3316) );
  AND2_X1 U11184 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10087), .ZN(P1_U3317) );
  AND2_X1 U11185 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10087), .ZN(P1_U3318) );
  AND2_X1 U11186 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10087), .ZN(P1_U3319) );
  AND2_X1 U11187 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10087), .ZN(P1_U3320) );
  AND2_X1 U11188 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10087), .ZN(P1_U3321) );
  INV_X1 U11189 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10089) );
  AOI21_X1 U11190 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(P1_U3441) );
  INV_X1 U11191 ( .A(n10145), .ZN(n10101) );
  OAI21_X1 U11192 ( .B1(n10092), .B2(n10130), .A(n10091), .ZN(n10094) );
  AOI211_X1 U11193 ( .C1(n10101), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10152) );
  AOI22_X1 U11194 ( .A1(n10150), .A2(n10152), .B1(n5499), .B2(n10149), .ZN(
        P1_U3457) );
  OAI22_X1 U11195 ( .A1(n10097), .A2(n10132), .B1(n10096), .B2(n10130), .ZN(
        n10099) );
  AOI211_X1 U11196 ( .C1(n10101), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10154) );
  AOI22_X1 U11197 ( .A1(n10150), .A2(n10154), .B1(n5508), .B2(n10149), .ZN(
        P1_U3460) );
  INV_X1 U11198 ( .A(n10102), .ZN(n10108) );
  NOR2_X1 U11199 ( .A1(n10102), .A2(n10145), .ZN(n10107) );
  OAI211_X1 U11200 ( .C1(n10132), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10106) );
  AOI211_X1 U11201 ( .C1(n10108), .C2(n10148), .A(n10107), .B(n10106), .ZN(
        n10156) );
  AOI22_X1 U11202 ( .A1(n10150), .A2(n10156), .B1(n5555), .B2(n10149), .ZN(
        P1_U3463) );
  OAI211_X1 U11203 ( .C1(n10132), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10112) );
  AOI21_X1 U11204 ( .B1(n10136), .B2(n10113), .A(n10112), .ZN(n10158) );
  AOI22_X1 U11205 ( .A1(n10150), .A2(n10158), .B1(n5489), .B2(n10149), .ZN(
        P1_U3466) );
  NAND3_X1 U11206 ( .A1(n10115), .A2(n10114), .A3(n10136), .ZN(n10116) );
  AND4_X1 U11207 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10160) );
  AOI22_X1 U11208 ( .A1(n10150), .A2(n10160), .B1(n5523), .B2(n10149), .ZN(
        P1_U3469) );
  OAI22_X1 U11209 ( .A1(n10120), .A2(n10132), .B1(n4781), .B2(n10130), .ZN(
        n10122) );
  AOI211_X1 U11210 ( .C1(n10123), .C2(n10136), .A(n10122), .B(n10121), .ZN(
        n10162) );
  AOI22_X1 U11211 ( .A1(n10150), .A2(n10162), .B1(n5539), .B2(n10149), .ZN(
        P1_U3472) );
  OAI21_X1 U11212 ( .B1(n10125), .B2(n10130), .A(n10124), .ZN(n10127) );
  AOI211_X1 U11213 ( .C1(n10136), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10164) );
  INV_X1 U11214 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U11215 ( .A1(n10150), .A2(n10164), .B1(n10129), .B2(n10149), .ZN(
        P1_U3475) );
  OAI22_X1 U11216 ( .A1(n10133), .A2(n10132), .B1(n10131), .B2(n10130), .ZN(
        n10135) );
  AOI211_X1 U11217 ( .C1(n10137), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10165) );
  AOI22_X1 U11218 ( .A1(n10150), .A2(n10165), .B1(n5615), .B2(n10149), .ZN(
        P1_U3478) );
  INV_X1 U11219 ( .A(n10144), .ZN(n10147) );
  AOI22_X1 U11220 ( .A1(n10141), .A2(n10140), .B1(n10139), .B2(n10138), .ZN(
        n10142) );
  OAI211_X1 U11221 ( .C1(n10145), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10146) );
  AOI21_X1 U11222 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(n10168) );
  AOI22_X1 U11223 ( .A1(n10150), .A2(n10168), .B1(n5592), .B2(n10149), .ZN(
        P1_U3481) );
  INV_X1 U11224 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U11225 ( .A1(n10169), .A2(n10152), .B1(n10151), .B2(n10166), .ZN(
        P1_U3524) );
  AOI22_X1 U11226 ( .A1(n10169), .A2(n10154), .B1(n10153), .B2(n10166), .ZN(
        P1_U3525) );
  INV_X1 U11227 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11228 ( .A1(n10169), .A2(n10156), .B1(n10155), .B2(n10166), .ZN(
        P1_U3526) );
  AOI22_X1 U11229 ( .A1(n10169), .A2(n10158), .B1(n10157), .B2(n10166), .ZN(
        P1_U3527) );
  INV_X1 U11230 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U11231 ( .A1(n10169), .A2(n10160), .B1(n10159), .B2(n10166), .ZN(
        P1_U3528) );
  INV_X1 U11232 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U11233 ( .A1(n10169), .A2(n10162), .B1(n10161), .B2(n10166), .ZN(
        P1_U3529) );
  INV_X1 U11234 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11235 ( .A1(n10169), .A2(n10164), .B1(n10163), .B2(n10166), .ZN(
        P1_U3530) );
  AOI22_X1 U11236 ( .A1(n10169), .A2(n10165), .B1(n6286), .B2(n10166), .ZN(
        P1_U3531) );
  AOI22_X1 U11237 ( .A1(n10169), .A2(n10168), .B1(n10167), .B2(n10166), .ZN(
        P1_U3532) );
  AOI22_X1 U11238 ( .A1(n10185), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10181), .ZN(n10177) );
  AOI22_X1 U11239 ( .A1(n10187), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10176) );
  OAI21_X1 U11240 ( .B1(n10171), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10170), .ZN(
        n10174) );
  NOR2_X1 U11241 ( .A1(n10172), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10173) );
  OAI21_X1 U11242 ( .B1(n10174), .B2(n10173), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10175) );
  OAI211_X1 U11243 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10177), .A(n10176), .B(
        n10175), .ZN(P2_U3245) );
  XNOR2_X1 U11244 ( .A(n10179), .B(n10178), .ZN(n10180) );
  AOI22_X1 U11245 ( .A1(n10183), .A2(n10182), .B1(n10181), .B2(n10180), .ZN(
        n10191) );
  OAI211_X1 U11246 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n10186), .A(n10185), 
        .B(n10184), .ZN(n10189) );
  NAND2_X1 U11247 ( .A1(n10187), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n10188) );
  NAND4_X1 U11248 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        P2_U3263) );
  XOR2_X1 U11249 ( .A(n10192), .B(n10204), .Z(n10195) );
  AOI21_X1 U11250 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10248) );
  OAI211_X1 U11251 ( .C1(n10198), .C2(n10249), .A(n10197), .B(n10196), .ZN(
        n10247) );
  OAI22_X1 U11252 ( .A1(n10247), .A2(n10201), .B1(n10200), .B2(n10199), .ZN(
        n10202) );
  INV_X1 U11253 ( .A(n10202), .ZN(n10209) );
  XNOR2_X1 U11254 ( .A(n10203), .B(n10204), .ZN(n10251) );
  AOI222_X1 U11255 ( .A1(n10251), .A2(n10207), .B1(P2_REG2_REG_4__SCAN_IN), 
        .B2(n10210), .C1(n10206), .C2(n10205), .ZN(n10208) );
  OAI211_X1 U11256 ( .C1(n10210), .C2(n10248), .A(n10209), .B(n10208), .ZN(
        P2_U3292) );
  NOR2_X1 U11257 ( .A1(n10212), .A2(n10211), .ZN(n10219) );
  INV_X1 U11258 ( .A(n10219), .ZN(n10223) );
  AND2_X1 U11259 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10223), .ZN(P2_U3297) );
  AND2_X1 U11260 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10223), .ZN(P2_U3298) );
  AND2_X1 U11261 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10223), .ZN(P2_U3299) );
  NOR2_X1 U11262 ( .A1(n10219), .A2(n10213), .ZN(P2_U3300) );
  NOR2_X1 U11263 ( .A1(n10219), .A2(n10214), .ZN(P2_U3301) );
  AND2_X1 U11264 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10223), .ZN(P2_U3302) );
  AND2_X1 U11265 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10223), .ZN(P2_U3303) );
  AND2_X1 U11266 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10223), .ZN(P2_U3304) );
  NOR2_X1 U11267 ( .A1(n10219), .A2(n10215), .ZN(P2_U3305) );
  AND2_X1 U11268 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10223), .ZN(P2_U3306) );
  AND2_X1 U11269 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10223), .ZN(P2_U3307) );
  NOR2_X1 U11270 ( .A1(n10219), .A2(n10216), .ZN(P2_U3308) );
  AND2_X1 U11271 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10223), .ZN(P2_U3309) );
  AND2_X1 U11272 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10223), .ZN(P2_U3310) );
  AND2_X1 U11273 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10223), .ZN(P2_U3311) );
  NOR2_X1 U11274 ( .A1(n10219), .A2(n10217), .ZN(P2_U3312) );
  AND2_X1 U11275 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10223), .ZN(P2_U3313) );
  AND2_X1 U11276 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10223), .ZN(P2_U3314) );
  AND2_X1 U11277 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10223), .ZN(P2_U3315) );
  AND2_X1 U11278 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10223), .ZN(P2_U3316) );
  AND2_X1 U11279 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10223), .ZN(P2_U3317) );
  AND2_X1 U11280 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10223), .ZN(P2_U3318) );
  AND2_X1 U11281 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10223), .ZN(P2_U3319) );
  AND2_X1 U11282 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10223), .ZN(P2_U3320) );
  AND2_X1 U11283 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10223), .ZN(P2_U3321) );
  NOR2_X1 U11284 ( .A1(n10219), .A2(n10218), .ZN(P2_U3322) );
  AND2_X1 U11285 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10223), .ZN(P2_U3323) );
  AND2_X1 U11286 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10223), .ZN(P2_U3324) );
  AND2_X1 U11287 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10223), .ZN(P2_U3325) );
  AND2_X1 U11288 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10223), .ZN(P2_U3326) );
  AOI22_X1 U11289 ( .A1(n10225), .A2(n10221), .B1(n10220), .B2(n10223), .ZN(
        P2_U3437) );
  INV_X1 U11290 ( .A(n10222), .ZN(n10224) );
  AOI22_X1 U11291 ( .A1(n10225), .A2(n10224), .B1(n6532), .B2(n10223), .ZN(
        P2_U3438) );
  INV_X1 U11292 ( .A(n10226), .ZN(n10227) );
  OAI21_X1 U11293 ( .B1(n10228), .B2(n10275), .A(n10227), .ZN(n10231) );
  INV_X1 U11294 ( .A(n10229), .ZN(n10230) );
  AOI211_X1 U11295 ( .C1(n10279), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        n10283) );
  AOI22_X1 U11296 ( .A1(n9320), .A2(n10283), .B1(n6558), .B2(n10281), .ZN(
        P2_U3454) );
  INV_X1 U11297 ( .A(n10233), .ZN(n10237) );
  OAI211_X1 U11298 ( .C1(n4489), .C2(n10275), .A(n10235), .B(n10234), .ZN(
        n10236) );
  AOI21_X1 U11299 ( .B1(n10279), .B2(n10237), .A(n10236), .ZN(n10285) );
  INV_X1 U11300 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U11301 ( .A1(n9320), .A2(n10285), .B1(n10238), .B2(n10281), .ZN(
        P2_U3457) );
  INV_X1 U11302 ( .A(n10243), .ZN(n10245) );
  AOI211_X1 U11303 ( .C1(n6570), .C2(n10241), .A(n10240), .B(n10239), .ZN(
        n10242) );
  OAI21_X1 U11304 ( .B1(n10258), .B2(n10243), .A(n10242), .ZN(n10244) );
  AOI21_X1 U11305 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(n10286) );
  AOI22_X1 U11306 ( .A1(n9320), .A2(n10286), .B1(n6614), .B2(n10281), .ZN(
        P2_U3460) );
  OAI211_X1 U11307 ( .C1(n10249), .C2(n10275), .A(n10248), .B(n10247), .ZN(
        n10250) );
  AOI21_X1 U11308 ( .B1(n10279), .B2(n10251), .A(n10250), .ZN(n10288) );
  AOI22_X1 U11309 ( .A1(n9320), .A2(n10288), .B1(n6652), .B2(n10281), .ZN(
        P2_U3463) );
  AND2_X1 U11310 ( .A1(n10252), .A2(n10279), .ZN(n10256) );
  OAI22_X1 U11311 ( .A1(n10254), .A2(n10261), .B1(n10253), .B2(n10275), .ZN(
        n10255) );
  NOR3_X1 U11312 ( .A1(n10257), .A2(n10256), .A3(n10255), .ZN(n10290) );
  AOI22_X1 U11313 ( .A1(n9320), .A2(n10290), .B1(n6856), .B2(n10281), .ZN(
        P2_U3469) );
  INV_X1 U11314 ( .A(n10258), .ZN(n10272) );
  INV_X1 U11315 ( .A(n10259), .ZN(n10265) );
  OAI22_X1 U11316 ( .A1(n10262), .A2(n10261), .B1(n10260), .B2(n10275), .ZN(
        n10264) );
  AOI211_X1 U11317 ( .C1(n10272), .C2(n10265), .A(n10264), .B(n10263), .ZN(
        n10291) );
  AOI22_X1 U11318 ( .A1(n9320), .A2(n10291), .B1(n6964), .B2(n10281), .ZN(
        P2_U3475) );
  INV_X1 U11319 ( .A(n10266), .ZN(n10271) );
  OAI21_X1 U11320 ( .B1(n10268), .B2(n10275), .A(n10267), .ZN(n10270) );
  AOI211_X1 U11321 ( .C1(n10272), .C2(n10271), .A(n10270), .B(n10269), .ZN(
        n10292) );
  INV_X1 U11322 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U11323 ( .A1(n9320), .A2(n10292), .B1(n10273), .B2(n10281), .ZN(
        P2_U3481) );
  OAI21_X1 U11324 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(n10278) );
  AOI211_X1 U11325 ( .C1(n10280), .C2(n10279), .A(n10278), .B(n10277), .ZN(
        n10294) );
  INV_X1 U11326 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U11327 ( .A1(n9320), .A2(n10294), .B1(n10282), .B2(n10281), .ZN(
        P2_U3487) );
  AOI22_X1 U11328 ( .A1(n10295), .A2(n10283), .B1(n4688), .B2(n10293), .ZN(
        P2_U3521) );
  INV_X1 U11329 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U11330 ( .A1(n10295), .A2(n10285), .B1(n10284), .B2(n10293), .ZN(
        P2_U3522) );
  AOI22_X1 U11331 ( .A1(n10295), .A2(n10286), .B1(n6414), .B2(n10293), .ZN(
        P2_U3523) );
  INV_X1 U11332 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11333 ( .A1(n10295), .A2(n10288), .B1(n10287), .B2(n10293), .ZN(
        P2_U3524) );
  INV_X1 U11334 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U11335 ( .A1(n10295), .A2(n10290), .B1(n10289), .B2(n10293), .ZN(
        P2_U3526) );
  AOI22_X1 U11336 ( .A1(n10295), .A2(n10291), .B1(n6667), .B2(n10293), .ZN(
        P2_U3528) );
  AOI22_X1 U11337 ( .A1(n10295), .A2(n10292), .B1(n7228), .B2(n10293), .ZN(
        P2_U3530) );
  AOI22_X1 U11338 ( .A1(n10295), .A2(n10294), .B1(n7476), .B2(n10293), .ZN(
        P2_U3532) );
  INV_X1 U11339 ( .A(n10296), .ZN(n10297) );
  NAND2_X1 U11340 ( .A1(n10298), .A2(n10297), .ZN(n10299) );
  XOR2_X1 U11341 ( .A(n10300), .B(n10299), .Z(ADD_1071_U5) );
  INV_X1 U11342 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U11343 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10302), .B2(n10301), .ZN(ADD_1071_U46) );
  OAI21_X1 U11344 ( .B1(n10305), .B2(n10304), .A(n10303), .ZN(ADD_1071_U56) );
  OAI21_X1 U11345 ( .B1(n10308), .B2(n10307), .A(n10306), .ZN(ADD_1071_U57) );
  OAI21_X1 U11346 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(ADD_1071_U58) );
  OAI21_X1 U11347 ( .B1(n10314), .B2(n10313), .A(n10312), .ZN(ADD_1071_U59) );
  OAI21_X1 U11348 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(ADD_1071_U60) );
  OAI21_X1 U11349 ( .B1(n10320), .B2(n10319), .A(n10318), .ZN(ADD_1071_U61) );
  AOI21_X1 U11350 ( .B1(n10323), .B2(n10322), .A(n10321), .ZN(ADD_1071_U62) );
  AOI21_X1 U11351 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(ADD_1071_U63) );
  AOI21_X1 U11352 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(ADD_1071_U48) );
  XOR2_X1 U11353 ( .A(n10330), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11354 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  XOR2_X1 U11355 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10333), .Z(ADD_1071_U51) );
  OAI21_X1 U11356 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(n10337) );
  XNOR2_X1 U11357 ( .A(n10337), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11358 ( .B1(n10340), .B2(n10339), .A(n10338), .ZN(ADD_1071_U47) );
  XOR2_X1 U11359 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10341), .Z(ADD_1071_U49) );
  XOR2_X1 U11360 ( .A(n10343), .B(n10342), .Z(ADD_1071_U54) );
  XOR2_X1 U11361 ( .A(n10345), .B(n10344), .Z(ADD_1071_U53) );
  XNOR2_X1 U11362 ( .A(n10347), .B(n10346), .ZN(ADD_1071_U52) );
  NOR2_X1 U4994 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5243) );
  CLKBUF_X1 U5003 ( .A(n5992), .Z(n6165) );
  CLKBUF_X1 U5015 ( .A(n5563), .Z(n5684) );
  NAND2_X2 U5034 ( .A1(n6549), .A2(n8976), .ZN(n8356) );
  CLKBUF_X1 U5204 ( .A(n6615), .Z(n8121) );
  CLKBUF_X1 U5836 ( .A(n5409), .Z(n5546) );
  OR3_X1 U6031 ( .A1(n7781), .A2(n7508), .A3(n7727), .ZN(n5930) );
endmodule

