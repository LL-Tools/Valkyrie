

module b15_C_SARLock_k_64_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703;

  AOI21_X1 U3409 ( .B1(n5221), .B2(n5202), .A(n5226), .ZN(n4131) );
  INV_X1 U3410 ( .A(n4080), .ZN(n4120) );
  CLKBUF_X2 U3411 ( .A(n4471), .Z(n2979) );
  AND2_X1 U3412 ( .A1(n4399), .A2(n3954), .ZN(n3973) );
  CLKBUF_X2 U3413 ( .A(n3782), .Z(n3663) );
  CLKBUF_X2 U3414 ( .A(n3195), .Z(n2973) );
  CLKBUF_X2 U3415 ( .A(n3207), .Z(n3906) );
  INV_X1 U3416 ( .A(n4278), .ZN(n3946) );
  AND4_X1 U3417 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3125)
         );
  AND2_X1 U3418 ( .A1(n4436), .A2(n4797), .ZN(n3207) );
  AND2_X1 U3419 ( .A1(n3119), .A2(n3118), .ZN(n3184) );
  AND2_X1 U3420 ( .A1(n4436), .A2(n3118), .ZN(n3186) );
  CLKBUF_X2 U3421 ( .A(n3904), .Z(n2977) );
  CLKBUF_X1 U3422 ( .A(n3187), .Z(n2965) );
  BUF_X1 U3423 ( .A(n3224), .Z(n3257) );
  AOI22_X1 U3425 ( .A1(n6631), .A2(keyinput44), .B1(keyinput18), .B2(n6630), 
        .ZN(n6629) );
  AND2_X1 U3426 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4797) );
  OAI221_X1 U3427 ( .B1(n6631), .B2(keyinput44), .C1(n6630), .C2(keyinput18), 
        .A(n6629), .ZN(n6644) );
  INV_X1 U3428 ( .A(n5912), .ZN(n5883) );
  AND2_X2 U3429 ( .A1(n4443), .A2(n4799), .ZN(n3904) );
  OR4_X1 U3431 ( .A1(n3067), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4347), .ZN(n2960) );
  AOI21_X2 U3432 ( .B1(n4532), .B2(n4533), .A(n4155), .ZN(n6083) );
  NAND2_X2 U3433 ( .A1(n5015), .A2(n4215), .ZN(n5055) );
  NAND2_X2 U3434 ( .A1(n3219), .A2(n3218), .ZN(n3255) );
  NAND2_X2 U3435 ( .A1(n3006), .A2(n2994), .ZN(n6414) );
  AND2_X4 U3436 ( .A1(n3112), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5145)
         );
  OAI21_X1 U3437 ( .B1(n3079), .B2(n3001), .A(n4219), .ZN(n3029) );
  INV_X4 U3438 ( .A(n4219), .ZN(n2967) );
  AND2_X1 U3439 ( .A1(n5382), .A2(n3045), .ZN(n5575) );
  XNOR2_X1 U3440 ( .A(n3294), .B(n3293), .ZN(n3435) );
  OR2_X1 U3441 ( .A1(n5283), .A2(n5282), .ZN(n5285) );
  CLKBUF_X2 U3442 ( .A(n4469), .Z(n2978) );
  NAND3_X1 U3443 ( .A1(n4401), .A2(n4256), .A3(n3222), .ZN(n4275) );
  CLKBUF_X2 U3444 ( .A(n4018), .Z(n4119) );
  NOR2_X2 U34450 ( .A1(n4278), .A2(n3253), .ZN(n4256) );
  NAND2_X1 U34460 ( .A1(n3220), .A2(n3256), .ZN(n4142) );
  CLKBUF_X2 U34470 ( .A(n3335), .Z(n3907) );
  BUF_X2 U34480 ( .A(n3184), .Z(n3905) );
  BUF_X2 U3449 ( .A(n3185), .Z(n3624) );
  CLKBUF_X2 U3450 ( .A(n3284), .Z(n3897) );
  INV_X2 U34510 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3110) );
  OR2_X1 U34520 ( .A1(n5518), .A2(n6065), .ZN(n4349) );
  NOR2_X1 U34530 ( .A1(n5420), .A2(n5519), .ZN(n4351) );
  AND2_X1 U3454 ( .A1(n3067), .A2(n2989), .ZN(n5409) );
  INV_X1 U34550 ( .A(n5427), .ZN(n5670) );
  INV_X1 U34560 ( .A(n5673), .ZN(n5435) );
  NAND2_X1 U3457 ( .A1(n5237), .A2(n3099), .ZN(n5423) );
  INV_X1 U3458 ( .A(n5447), .ZN(n5404) );
  NOR2_X1 U34590 ( .A1(n4355), .A2(n4354), .ZN(n3930) );
  AND2_X1 U34600 ( .A1(n5334), .A2(n5342), .ZN(n5673) );
  OR2_X1 U34610 ( .A1(n5336), .A2(n5250), .ZN(n5427) );
  OR2_X1 U34620 ( .A1(n5238), .A2(n4344), .ZN(n4345) );
  NAND2_X1 U34630 ( .A1(n3101), .A2(n3100), .ZN(n3099) );
  NAND2_X1 U34640 ( .A1(n4343), .A2(n4344), .ZN(n4355) );
  CLKBUF_X1 U34650 ( .A(n4343), .Z(n5238) );
  NOR2_X1 U3466 ( .A1(n3063), .A2(n3023), .ZN(n3022) );
  INV_X1 U3467 ( .A(n3080), .ZN(n3079) );
  NOR2_X1 U34680 ( .A1(n4221), .A2(n4220), .ZN(n4222) );
  NOR2_X1 U34690 ( .A1(n4230), .A2(n3083), .ZN(n3082) );
  INV_X1 U34700 ( .A(n5093), .ZN(n3064) );
  AND2_X2 U34710 ( .A1(n4206), .A2(n4209), .ZN(n4219) );
  NAND2_X1 U34720 ( .A1(n3392), .A2(n3425), .ZN(n3479) );
  AND2_X1 U34730 ( .A1(n3470), .A2(n3471), .ZN(n4512) );
  NAND2_X1 U34740 ( .A1(n3058), .A2(n3057), .ZN(n3056) );
  AND2_X1 U3475 ( .A1(n4393), .A2(n4394), .ZN(n3465) );
  AND2_X1 U3476 ( .A1(n3378), .A2(n3377), .ZN(n4539) );
  NAND2_X1 U3477 ( .A1(n3455), .A2(n3454), .ZN(n4824) );
  NAND2_X1 U3478 ( .A1(n3450), .A2(n3353), .ZN(n3439) );
  AND2_X1 U3479 ( .A1(n6414), .A2(n6429), .ZN(n4657) );
  NAND2_X1 U3480 ( .A1(n3364), .A2(n3363), .ZN(n4513) );
  CLKBUF_X1 U3481 ( .A(n3266), .Z(n3360) );
  AOI21_X1 U3482 ( .B1(n3250), .B2(n3249), .A(n3248), .ZN(n4272) );
  AND3_X1 U3483 ( .A1(n3261), .A2(n3260), .A3(n3259), .ZN(n3262) );
  NOR2_X1 U3484 ( .A1(n3350), .A2(n6419), .ZN(n3451) );
  INV_X2 U3485 ( .A(n4020), .ZN(n4406) );
  NAND2_X1 U3486 ( .A1(n2981), .A2(n5211), .ZN(n3232) );
  OR2_X1 U3487 ( .A1(n3366), .A2(n3318), .ZN(n3306) );
  NAND2_X4 U3488 ( .A1(n3215), .A2(n3420), .ZN(n3217) );
  OR2_X1 U3489 ( .A1(n3341), .A2(n3340), .ZN(n4148) );
  NAND2_X1 U3490 ( .A1(n3221), .A2(n3237), .ZN(n4398) );
  OR2_X1 U3491 ( .A1(n3317), .A2(n3316), .ZN(n4211) );
  CLKBUF_X1 U3492 ( .A(n3221), .Z(n3222) );
  INV_X1 U3493 ( .A(n3247), .ZN(n4399) );
  INV_X1 U3494 ( .A(n3220), .ZN(n4265) );
  NAND2_X2 U3495 ( .A1(n3135), .A2(n3134), .ZN(n3237) );
  OR2_X1 U3496 ( .A1(n3176), .A2(n3175), .ZN(n3256) );
  NOR2_X1 U3497 ( .A1(n3003), .A2(n2986), .ZN(n3002) );
  OR2_X2 U3498 ( .A1(n3155), .A2(n3154), .ZN(n5211) );
  OR2_X2 U3499 ( .A1(n3193), .A2(n3192), .ZN(n4278) );
  AND3_X2 U3500 ( .A1(n3165), .A2(n3107), .A3(n3106), .ZN(n3247) );
  AND4_X1 U3501 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3108)
         );
  AND4_X1 U3502 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3145)
         );
  AND4_X1 U3503 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3124)
         );
  AND4_X1 U3504 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3134)
         );
  AND4_X1 U3505 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3213)
         );
  AND4_X1 U3506 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3212)
         );
  AND4_X1 U3507 ( .A1(n3208), .A2(n3209), .A3(n3211), .A4(n3005), .ZN(n3004)
         );
  BUF_X2 U3508 ( .A(n2966), .Z(n3898) );
  AND2_X1 U3509 ( .A1(n3210), .A2(n3202), .ZN(n3005) );
  BUF_X2 U3510 ( .A(n3329), .Z(n3903) );
  INV_X2 U3511 ( .A(n6063), .ZN(n6075) );
  BUF_X2 U3512 ( .A(n3328), .Z(n3307) );
  BUF_X2 U3513 ( .A(n3904), .Z(n2976) );
  BUF_X2 U3514 ( .A(n3904), .Z(n2974) );
  BUF_X2 U3515 ( .A(n3186), .Z(n3753) );
  AND2_X1 U3516 ( .A1(n3031), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3119)
         );
  NOR2_X1 U3517 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3118) );
  NOR2_X1 U3518 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3111) );
  AND2_X2 U3519 ( .A1(n2961), .A2(n3541), .ZN(n5051) );
  NOR2_X1 U3520 ( .A1(n5052), .A2(n5034), .ZN(n2961) );
  CLKBUF_X1 U3521 ( .A(n6396), .Z(n2962) );
  AND2_X2 U3522 ( .A1(n3420), .A2(n5211), .ZN(n3456) );
  INV_X1 U3523 ( .A(n2963), .ZN(n4318) );
  INV_X2 U3524 ( .A(n3140), .ZN(n3161) );
  AND2_X2 U3525 ( .A1(n3253), .A2(n3946), .ZN(n4136) );
  NAND3_X4 U3526 ( .A1(n3002), .A2(n3213), .A3(n2982), .ZN(n3253) );
  AND2_X2 U3527 ( .A1(n4319), .A2(n4320), .ZN(n2963) );
  AND2_X1 U3528 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4442) );
  AND2_X2 U3529 ( .A1(n3178), .A2(n3177), .ZN(n3986) );
  AND2_X1 U3530 ( .A1(n3216), .A2(n4438), .ZN(n3261) );
  AND2_X2 U3531 ( .A1(n4398), .A2(n3247), .ZN(n2981) );
  AND2_X2 U3532 ( .A1(n3212), .A2(n3004), .ZN(n2982) );
  NAND2_X1 U3533 ( .A1(n3265), .A2(n3245), .ZN(n3295) );
  NAND2_X1 U3534 ( .A1(n4568), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3365) );
  INV_X2 U3535 ( .A(n3237), .ZN(n3420) );
  AND2_X1 U3536 ( .A1(n3119), .A2(n4797), .ZN(n2964) );
  BUF_X4 U3537 ( .A(n3187), .Z(n2966) );
  AND2_X2 U3538 ( .A1(n3019), .A2(n3017), .ZN(n2983) );
  NAND2_X1 U3539 ( .A1(n3014), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3241) );
  NOR2_X4 U3540 ( .A1(n5377), .A2(n3677), .ZN(n5365) );
  INV_X2 U3541 ( .A(n3221), .ZN(n3215) );
  XNOR2_X1 U3542 ( .A(n4355), .B(n4354), .ZN(n5217) );
  NAND2_X2 U3543 ( .A1(n3435), .A2(n3436), .ZN(n3469) );
  NAND3_X2 U3544 ( .A1(n3027), .A2(n2987), .A3(n3026), .ZN(n5472) );
  NOR2_X2 U3545 ( .A1(n5359), .A2(n3094), .ZN(n4319) );
  NAND2_X2 U3546 ( .A1(n5365), .A2(n5366), .ZN(n5359) );
  NOR2_X1 U3547 ( .A1(n3110), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3117)
         );
  AND2_X2 U3548 ( .A1(n3110), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4443)
         );
  OR2_X2 U3549 ( .A1(n5122), .A2(n3091), .ZN(n5377) );
  NAND2_X1 U3550 ( .A1(n3541), .A2(n3540), .ZN(n5035) );
  AND2_X1 U3551 ( .A1(n5145), .A2(n4797), .ZN(n3334) );
  AND2_X2 U3552 ( .A1(n5145), .A2(n4797), .ZN(n2971) );
  AOI211_X2 U3553 ( .C1(n6059), .C2(n5621), .A(n5437), .B(n5436), .ZN(n5438)
         );
  NOR2_X2 U3554 ( .A1(n4422), .A2(n4429), .ZN(n4428) );
  NAND2_X2 U3555 ( .A1(n3279), .A2(n4800), .ZN(n4470) );
  NAND2_X2 U3556 ( .A1(n3056), .A2(n3469), .ZN(n4468) );
  AND2_X1 U3557 ( .A1(n3117), .A2(n5145), .ZN(n2968) );
  INV_X1 U3558 ( .A(n3140), .ZN(n2969) );
  INV_X2 U3559 ( .A(n3140), .ZN(n3896) );
  AND2_X1 U3560 ( .A1(n5145), .A2(n4797), .ZN(n2970) );
  AND2_X4 U3562 ( .A1(n4797), .A2(n4799), .ZN(n3879) );
  NOR2_X4 U3563 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4799) );
  AND2_X1 U3564 ( .A1(n3119), .A2(n4797), .ZN(n3195) );
  XNOR2_X1 U3565 ( .A(n3441), .B(n3440), .ZN(n4469) );
  AND2_X4 U3566 ( .A1(n4442), .A2(n3111), .ZN(n3862) );
  AND2_X1 U3567 ( .A1(n3253), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3954) );
  AOI21_X1 U3568 ( .B1(n3940), .B2(n4187), .A(n3939), .ZN(n3975) );
  AOI22_X1 U3569 ( .A1(n3983), .A2(n3973), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6419), .ZN(n3974) );
  NOR2_X1 U3570 ( .A1(n5335), .A2(n5341), .ZN(n3104) );
  INV_X1 U3571 ( .A(n3890), .ZN(n3922) );
  NOR2_X1 U3572 ( .A1(n5139), .A2(n6419), .ZN(n3890) );
  NOR2_X1 U3573 ( .A1(n3077), .A2(n3072), .ZN(n3071) );
  INV_X1 U3574 ( .A(n4224), .ZN(n3072) );
  NAND2_X1 U3575 ( .A1(n3079), .A2(n3078), .ZN(n3077) );
  AOI21_X1 U3576 ( .B1(n3079), .B2(n3076), .A(n3075), .ZN(n3074) );
  INV_X1 U3577 ( .A(n5481), .ZN(n3075) );
  NOR2_X1 U3578 ( .A1(n3082), .A2(n4231), .ZN(n3076) );
  INV_X1 U3579 ( .A(n3029), .ZN(n3028) );
  INV_X1 U3580 ( .A(n3065), .ZN(n3062) );
  INV_X1 U3581 ( .A(n4217), .ZN(n3023) );
  NAND2_X1 U3582 ( .A1(n4222), .A2(n3064), .ZN(n3063) );
  NOR2_X1 U3583 ( .A1(n3043), .A2(n5062), .ZN(n3042) );
  INV_X1 U3584 ( .A(n4066), .ZN(n3043) );
  NAND2_X1 U3585 ( .A1(n5055), .A2(n4216), .ZN(n3024) );
  AND2_X1 U3586 ( .A1(n6525), .A2(n3991), .ZN(n5888) );
  NOR2_X1 U3587 ( .A1(n5888), .A2(n6279), .ZN(n5028) );
  NAND2_X1 U3588 ( .A1(n3093), .A2(n5273), .ZN(n3091) );
  NAND2_X1 U3589 ( .A1(n4657), .A2(n4417), .ZN(n6004) );
  INV_X1 U3590 ( .A(n3792), .ZN(n3927) );
  INV_X1 U3591 ( .A(n3087), .ZN(n3086) );
  OAI21_X1 U3592 ( .B1(n3088), .B2(n5061), .A(n5084), .ZN(n3087) );
  INV_X1 U3593 ( .A(n4903), .ZN(n3524) );
  NOR2_X1 U3594 ( .A1(n5432), .A2(n3069), .ZN(n3068) );
  INV_X1 U3595 ( .A(n4235), .ZN(n3069) );
  NOR2_X1 U3596 ( .A1(n4094), .A2(n3048), .ZN(n3047) );
  NAND2_X1 U3597 ( .A1(n4254), .A2(n4253), .ZN(n4291) );
  AND2_X1 U3598 ( .A1(n6418), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3979) );
  OR2_X1 U3599 ( .A1(n5331), .A2(n5874), .ZN(n3032) );
  NAND2_X1 U3600 ( .A1(n3934), .A2(n3933), .ZN(n3942) );
  INV_X1 U3601 ( .A(n4227), .ZN(n3083) );
  NAND2_X1 U3602 ( .A1(n3417), .A2(n3416), .ZN(n3487) );
  AND2_X1 U3603 ( .A1(n3231), .A2(n3230), .ZN(n3242) );
  NOR2_X1 U3604 ( .A1(n3938), .A2(n6182), .ZN(n3983) );
  NAND2_X1 U3605 ( .A1(n5252), .A2(n3050), .ZN(n3049) );
  INV_X1 U3606 ( .A(n3051), .ZN(n3050) );
  AOI22_X1 U3607 ( .A1(n3335), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U3608 ( .A1(n3782), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U3609 ( .A1(n3334), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3132) );
  INV_X1 U3610 ( .A(n5239), .ZN(n3103) );
  INV_X1 U3611 ( .A(n5359), .ZN(n3096) );
  AND2_X1 U3612 ( .A1(n4240), .A2(n4241), .ZN(n4257) );
  NOR2_X1 U3613 ( .A1(n5466), .A2(n3018), .ZN(n3017) );
  OAI21_X1 U3614 ( .B1(n4230), .B2(n3081), .A(n4229), .ZN(n3080) );
  NAND2_X1 U3615 ( .A1(n4228), .A2(n4227), .ZN(n3081) );
  NAND2_X1 U3616 ( .A1(n5496), .A2(n3082), .ZN(n3073) );
  AND2_X1 U3617 ( .A1(n4257), .A2(n4256), .ZN(n4409) );
  NAND2_X1 U3618 ( .A1(n3016), .A2(n3236), .ZN(n3015) );
  CLKBUF_X1 U3619 ( .A(n4248), .Z(n4451) );
  INV_X1 U3620 ( .A(n4539), .ZN(n3379) );
  AOI22_X1 U3621 ( .A1(n3328), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3120) );
  AOI21_X1 U3622 ( .B1(n6434), .B2(n4822), .A(n5186), .ZN(n4480) );
  AND2_X1 U3623 ( .A1(n3986), .A2(n3988), .ZN(n6397) );
  INV_X1 U3624 ( .A(n5888), .ZN(n5064) );
  AND2_X1 U3625 ( .A1(n3676), .A2(n3675), .ZN(n5379) );
  OAI21_X1 U3626 ( .B1(n4386), .B2(n3919), .A(n3457), .ZN(n4394) );
  NAND2_X1 U3627 ( .A1(n3838), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3857)
         );
  NAND2_X1 U3628 ( .A1(n3095), .A2(n5351), .ZN(n3094) );
  NOR2_X1 U3629 ( .A1(n6631), .A2(n3641), .ZN(n3674) );
  INV_X1 U3630 ( .A(n3640), .ZN(n3641) );
  NAND2_X1 U3631 ( .A1(n3622), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3623)
         );
  NOR2_X1 U3632 ( .A1(n6637), .A2(n3623), .ZN(n3640) );
  AND3_X1 U3633 ( .A1(n3621), .A2(n3620), .A3(n3619), .ZN(n5128) );
  NOR2_X1 U3634 ( .A1(n3579), .A2(n3090), .ZN(n3089) );
  INV_X1 U3635 ( .A(n5061), .ZN(n3090) );
  NAND2_X1 U3636 ( .A1(n3085), .A2(n3579), .ZN(n3084) );
  NAND2_X1 U3637 ( .A1(n5051), .A2(n5061), .ZN(n3085) );
  NOR2_X1 U3638 ( .A1(n3558), .A2(n5840), .ZN(n3574) );
  INV_X1 U3639 ( .A(n4503), .ZN(n3485) );
  INV_X1 U3640 ( .A(n5453), .ZN(n5440) );
  NOR2_X1 U3641 ( .A1(n3046), .A2(n5572), .ZN(n3045) );
  INV_X1 U3642 ( .A(n3047), .ZN(n3046) );
  NAND2_X1 U3643 ( .A1(n3021), .A2(n3020), .ZN(n3019) );
  INV_X1 U3644 ( .A(n5686), .ZN(n3020) );
  INV_X1 U3645 ( .A(n5688), .ZN(n3021) );
  AND2_X1 U3646 ( .A1(n3061), .A2(n5091), .ZN(n3060) );
  NAND2_X1 U3647 ( .A1(n3024), .A2(n3022), .ZN(n3025) );
  AND2_X1 U3648 ( .A1(n4071), .A2(n4070), .ZN(n5062) );
  INV_X1 U3649 ( .A(n5586), .ZN(n6106) );
  OR3_X1 U3650 ( .A1(n4441), .A2(n4786), .A3(n4276), .ZN(n4277) );
  NAND2_X1 U3651 ( .A1(n4291), .A2(n6399), .ZN(n5585) );
  NAND2_X1 U3652 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  NAND2_X1 U3653 ( .A1(n3351), .A2(n3347), .ZN(n3348) );
  NAND2_X1 U3654 ( .A1(n3346), .A2(n4148), .ZN(n3349) );
  NOR2_X1 U3655 ( .A1(n4512), .A2(n4597), .ZN(n4603) );
  NAND2_X1 U3656 ( .A1(n3010), .A2(n3007), .ZN(n3006) );
  INV_X1 U3657 ( .A(n3008), .ZN(n3007) );
  INV_X1 U3658 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U3659 ( .A1(n2984), .A2(n3035), .ZN(n3034) );
  NAND2_X1 U3660 ( .A1(n4138), .A2(n4137), .ZN(n3035) );
  INV_X1 U3661 ( .A(n5633), .ZN(n5622) );
  OR2_X1 U3662 ( .A1(n5826), .A2(n4002), .ZN(n5296) );
  XNOR2_X1 U3663 ( .A(n4131), .B(n3033), .ZN(n5331) );
  INV_X1 U3664 ( .A(n4132), .ZN(n3033) );
  INV_X1 U3665 ( .A(n5251), .ZN(n3100) );
  INV_X1 U3666 ( .A(n5250), .ZN(n3101) );
  NOR2_X2 U3667 ( .A1(n5944), .A2(n5210), .ZN(n5941) );
  OAI21_X1 U3668 ( .B1(n4456), .B2(n4416), .A(n6429), .ZN(n4418) );
  XNOR2_X1 U3669 ( .A(n3995), .B(n3994), .ZN(n4339) );
  INV_X1 U3670 ( .A(n5423), .ZN(n3098) );
  INV_X1 U3671 ( .A(n6090), .ZN(n6059) );
  INV_X1 U3672 ( .A(n5483), .ZN(n6080) );
  NAND2_X2 U3673 ( .A1(n4657), .A2(n4331), .ZN(n6065) );
  XNOR2_X1 U3674 ( .A(n3055), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4341)
         );
  NAND2_X1 U3675 ( .A1(n4239), .A2(n2960), .ZN(n3055) );
  AND2_X1 U3676 ( .A1(n5717), .A2(n4303), .ZN(n5532) );
  AND2_X1 U3677 ( .A1(n5560), .A2(n4299), .ZN(n5710) );
  INV_X1 U3678 ( .A(n4733), .ZN(n4689) );
  AOI21_X1 U3679 ( .B1(n6390), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3936), 
        .ZN(n3937) );
  INV_X1 U3680 ( .A(n3942), .ZN(n3935) );
  INV_X1 U3681 ( .A(n4231), .ZN(n3078) );
  OR2_X1 U3682 ( .A1(n3402), .A2(n3401), .ZN(n4188) );
  OR2_X1 U3683 ( .A1(n3415), .A2(n3414), .ZN(n4199) );
  OR2_X1 U3684 ( .A1(n3305), .A2(n3304), .ZN(n4141) );
  OR2_X1 U3685 ( .A1(n3290), .A2(n3289), .ZN(n3291) );
  OR2_X1 U3686 ( .A1(n3376), .A2(n3375), .ZN(n4171) );
  AOI22_X1 U3687 ( .A1(n2969), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3688 ( .A1(n3366), .A2(n3365), .ZN(n3976) );
  NAND2_X1 U3689 ( .A1(n3201), .A2(n3200), .ZN(n3003) );
  NOR2_X1 U3690 ( .A1(n3748), .A2(n5360), .ZN(n3095) );
  OR2_X1 U3691 ( .A1(n5467), .A2(n5262), .ZN(n3748) );
  OR2_X1 U3692 ( .A1(n5343), .A2(n3054), .ZN(n3051) );
  INV_X1 U3693 ( .A(n5337), .ZN(n3054) );
  NOR2_X1 U3694 ( .A1(n3066), .A2(n4223), .ZN(n3065) );
  INV_X1 U3695 ( .A(n5075), .ZN(n3066) );
  INV_X1 U3696 ( .A(n4035), .ZN(n3039) );
  NOR2_X1 U3697 ( .A1(n4266), .A2(n4020), .ZN(n4126) );
  INV_X1 U3698 ( .A(n3291), .ZN(n4164) );
  NAND2_X1 U3699 ( .A1(n4211), .A2(n3247), .ZN(n3351) );
  INV_X1 U3700 ( .A(n4141), .ZN(n3318) );
  NAND2_X1 U3701 ( .A1(n3247), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U3702 ( .A1(n3220), .A2(n3252), .ZN(n4273) );
  AND2_X1 U3703 ( .A1(n3228), .A2(n3268), .ZN(n4947) );
  INV_X1 U3704 ( .A(n2978), .ZN(n4699) );
  AOI22_X1 U3705 ( .A1(n3195), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3706 ( .A1(n3973), .A2(n4187), .ZN(n3978) );
  OAI21_X1 U3707 ( .B1(n3974), .B2(n3975), .A(n3009), .ZN(n3008) );
  NAND2_X1 U3708 ( .A1(n3976), .A2(n3977), .ZN(n3009) );
  OR2_X1 U3709 ( .A1(n3973), .A2(n3980), .ZN(n3012) );
  NAND2_X1 U3710 ( .A1(n3974), .A2(n3975), .ZN(n3011) );
  INV_X1 U3711 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6665) );
  INV_X1 U3712 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6631) );
  INV_X1 U3713 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5812) );
  INV_X1 U3714 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U3715 ( .A1(n4407), .A2(n4406), .ZN(n4405) );
  NOR3_X1 U3716 ( .A1(n5242), .A2(n4130), .A3(n4129), .ZN(n5224) );
  NAND2_X1 U3717 ( .A1(n3053), .A2(n3052), .ZN(n5242) );
  INV_X1 U3718 ( .A(n5240), .ZN(n3052) );
  INV_X1 U3719 ( .A(n3053), .ZN(n5254) );
  OR2_X1 U3720 ( .A1(n3840), .A2(n3839), .ZN(n5335) );
  INV_X1 U3721 ( .A(n4273), .ZN(n4401) );
  AOI22_X1 U3722 ( .A1(n3334), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U3723 ( .A1(n3856), .A2(n3855), .B1(n3893), .B2(n5425), .ZN(n5251)
         );
  NAND2_X1 U3724 ( .A1(n4413), .A2(n4412), .ZN(n4456) );
  OR2_X1 U3725 ( .A1(n5770), .A2(n4411), .ZN(n4412) );
  AOI22_X1 U3726 ( .A1(n3328), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3131) );
  AND2_X1 U3727 ( .A1(n4660), .A2(n4659), .ZN(n5948) );
  NAND2_X1 U3728 ( .A1(n6052), .A2(n4658), .ZN(n4660) );
  OR2_X1 U3729 ( .A1(n3924), .A2(n5205), .ZN(n3992) );
  AOI22_X1 U3730 ( .A1(n3895), .A2(n3894), .B1(n3893), .B2(n5203), .ZN(n4344)
         );
  NAND2_X1 U3731 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3924)
         );
  AND2_X1 U3732 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n3837), .ZN(n3838)
         );
  NOR2_X1 U3733 ( .A1(n3791), .A2(n5638), .ZN(n3813) );
  AND2_X1 U3734 ( .A1(n5628), .A2(n3990), .ZN(n3773) );
  AND2_X1 U3735 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3744), .ZN(n3745)
         );
  NAND2_X1 U3736 ( .A1(n3745), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3791)
         );
  NOR2_X1 U3737 ( .A1(n3694), .A2(n5653), .ZN(n3695) );
  AND2_X1 U3738 ( .A1(n3693), .A2(n3692), .ZN(n5366) );
  INV_X1 U3739 ( .A(n5379), .ZN(n3677) );
  NAND2_X1 U3740 ( .A1(n3674), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3694)
         );
  AND2_X1 U3741 ( .A1(n3639), .A2(n3638), .ZN(n5281) );
  NOR2_X1 U3742 ( .A1(n3618), .A2(n5812), .ZN(n3622) );
  AND2_X1 U3743 ( .A1(n3574), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3575)
         );
  NAND2_X1 U3744 ( .A1(n3575), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3618)
         );
  NAND2_X1 U3745 ( .A1(n3573), .A2(n3572), .ZN(n5061) );
  NAND2_X1 U3746 ( .A1(n3542), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3558)
         );
  NAND2_X1 U3747 ( .A1(n3508), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3525)
         );
  AND2_X1 U3748 ( .A1(n3503), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3508)
         );
  NOR2_X1 U3749 ( .A1(n3481), .A2(n4910), .ZN(n3489) );
  AOI21_X1 U3750 ( .B1(n4178), .B2(n3615), .A(n3484), .ZN(n4503) );
  NOR2_X1 U3751 ( .A1(n6591), .A2(n3473), .ZN(n3472) );
  NAND2_X1 U3752 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3473) );
  INV_X1 U3753 ( .A(n3465), .ZN(n4425) );
  AND2_X1 U3754 ( .A1(n4257), .A2(n4255), .ZN(n4331) );
  NOR2_X1 U3755 ( .A1(n5344), .A2(n3051), .ZN(n5339) );
  NOR2_X1 U3756 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  OR2_X1 U3757 ( .A1(n5356), .A2(n4322), .ZN(n5344) );
  OR2_X1 U3758 ( .A1(n5097), .A2(n5100), .ZN(n4301) );
  NAND2_X1 U3759 ( .A1(n5354), .A2(n5353), .ZN(n5356) );
  NAND2_X1 U3760 ( .A1(n3019), .A2(n2993), .ZN(n5453) );
  AOI21_X1 U3761 ( .B1(n2967), .B2(n6670), .A(n2983), .ZN(n5460) );
  AND2_X1 U3762 ( .A1(n5575), .A2(n5268), .ZN(n5354) );
  NAND2_X1 U3763 ( .A1(n5382), .A2(n5371), .ZN(n5370) );
  NAND2_X1 U3764 ( .A1(n3028), .A2(n3001), .ZN(n3026) );
  NAND2_X1 U3765 ( .A1(n3073), .A2(n3028), .ZN(n3027) );
  OR2_X1 U3766 ( .A1(n4290), .A2(n6137), .ZN(n5584) );
  OR2_X1 U3767 ( .A1(n2967), .A2(n5693), .ZN(n5481) );
  OR2_X1 U3768 ( .A1(n2967), .A2(n4226), .ZN(n4227) );
  OR2_X1 U3769 ( .A1(n5131), .A2(n5130), .ZN(n5283) );
  NOR2_X1 U3770 ( .A1(n5861), .A2(n3041), .ZN(n5763) );
  NAND2_X1 U3771 ( .A1(n3042), .A2(n5761), .ZN(n3041) );
  NAND2_X1 U3772 ( .A1(n5763), .A2(n5125), .ZN(n5131) );
  INV_X1 U3773 ( .A(n3042), .ZN(n3040) );
  NOR2_X1 U3774 ( .A1(n2967), .A2(n6685), .ZN(n4220) );
  INV_X1 U3775 ( .A(n6054), .ZN(n4221) );
  NAND2_X1 U3776 ( .A1(n5074), .A2(n3065), .ZN(n3059) );
  NAND2_X1 U3777 ( .A1(n5859), .A2(n5858), .ZN(n5861) );
  NAND2_X1 U3778 ( .A1(n3044), .A2(n4066), .ZN(n5833) );
  INV_X1 U3779 ( .A(n5861), .ZN(n3044) );
  AND2_X1 U3780 ( .A1(n4056), .A2(n4055), .ZN(n4364) );
  NOR2_X1 U3781 ( .A1(n4746), .A2(n4364), .ZN(n5859) );
  NAND2_X1 U3782 ( .A1(n3038), .A2(n3036), .ZN(n4748) );
  INV_X1 U3783 ( .A(n4043), .ZN(n3038) );
  NOR2_X1 U3784 ( .A1(n4432), .A2(n3037), .ZN(n3036) );
  NAND2_X1 U3785 ( .A1(n3039), .A2(n4499), .ZN(n3037) );
  NAND2_X1 U3786 ( .A1(n4052), .A2(n4051), .ZN(n4746) );
  INV_X1 U3787 ( .A(n4749), .ZN(n4051) );
  INV_X1 U3788 ( .A(n4748), .ZN(n4052) );
  OR2_X1 U3789 ( .A1(n4432), .A2(n4035), .ZN(n5885) );
  OR2_X1 U3790 ( .A1(n4451), .A2(n4020), .ZN(n4454) );
  AND2_X1 U3791 ( .A1(n4080), .A2(n4119), .ZN(n4379) );
  NAND2_X1 U3792 ( .A1(n3244), .A2(n2995), .ZN(n3245) );
  INV_X1 U3793 ( .A(n3241), .ZN(n3244) );
  NAND2_X1 U3794 ( .A1(n3263), .A2(n3321), .ZN(n3326) );
  AND2_X1 U3795 ( .A1(n3454), .A2(n4208), .ZN(n3353) );
  INV_X1 U3796 ( .A(n3436), .ZN(n3057) );
  INV_X1 U3797 ( .A(n3435), .ZN(n3058) );
  INV_X1 U3798 ( .A(n3469), .ZN(n3030) );
  INV_X1 U3799 ( .A(n6270), .ZN(n6274) );
  OR2_X1 U3800 ( .A1(n3251), .A2(n3222), .ZN(n5139) );
  NAND2_X1 U3801 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6414), .ZN(n5190) );
  INV_X1 U3802 ( .A(n4256), .ZN(n3948) );
  NOR2_X1 U3803 ( .A1(n6274), .A2(n2978), .ZN(n4592) );
  AND2_X1 U3804 ( .A1(n2978), .A2(n4824), .ZN(n6183) );
  AND2_X1 U3805 ( .A1(n4512), .A2(n4468), .ZN(n6270) );
  AND2_X1 U3806 ( .A1(n2978), .A2(n4700), .ZN(n6269) );
  OR2_X1 U3807 ( .A1(n6512), .A2(n4480), .ZN(n4580) );
  OR2_X1 U3808 ( .A1(n6398), .A2(n3989), .ZN(n4370) );
  NAND2_X1 U3809 ( .A1(n4657), .A2(n3016), .ZN(n5969) );
  AND2_X1 U3810 ( .A1(n5969), .A2(n4370), .ZN(n6525) );
  AND2_X1 U3811 ( .A1(n5640), .A2(n4007), .ZN(n5633) );
  INV_X1 U3812 ( .A(n5301), .ZN(n5892) );
  NAND2_X1 U3813 ( .A1(n5028), .A2(n3999), .ZN(n5826) );
  INV_X1 U3814 ( .A(n5903), .ZN(n5864) );
  INV_X1 U3815 ( .A(n5874), .ZN(n5906) );
  NAND2_X1 U3816 ( .A1(n5826), .A2(n5064), .ZN(n5886) );
  AND2_X1 U3817 ( .A1(n5384), .A2(n5383), .ZN(n5806) );
  INV_X1 U3818 ( .A(n5925), .ZN(n5930) );
  NAND2_X1 U3819 ( .A1(n4404), .A2(n5934), .ZN(n5925) );
  AND2_X1 U3820 ( .A1(n5392), .A2(n5212), .ZN(n5945) );
  AND2_X1 U3821 ( .A1(n5392), .A2(n4420), .ZN(n5134) );
  INV_X1 U3822 ( .A(n5134), .ZN(n5083) );
  INV_X1 U3823 ( .A(n6527), .ZN(n5966) );
  INV_X1 U3824 ( .A(n6412), .ZN(n4656) );
  CLKBUF_X1 U3825 ( .A(n6043), .Z(n6050) );
  AND2_X1 U3826 ( .A1(n3643), .A2(n3642), .ZN(n5703) );
  AND2_X1 U3827 ( .A1(n5127), .A2(n5129), .ZN(n5493) );
  CLKBUF_X1 U3828 ( .A(n5120), .Z(n5121) );
  AND2_X1 U3829 ( .A1(n5087), .A2(n5086), .ZN(n5919) );
  NAND2_X1 U3830 ( .A1(n5074), .A2(n5075), .ZN(n6055) );
  CLKBUF_X1 U3831 ( .A(n4901), .Z(n4902) );
  INV_X1 U3832 ( .A(n6065), .ZN(n6085) );
  NAND2_X1 U3833 ( .A1(n5382), .A2(n3047), .ZN(n5573) );
  NAND2_X1 U3834 ( .A1(n3019), .A2(n5685), .ZN(n5465) );
  AND2_X1 U3835 ( .A1(n4295), .A2(n4294), .ZN(n5735) );
  NAND2_X1 U3836 ( .A1(n5584), .A2(n4282), .ZN(n5739) );
  OR2_X1 U3837 ( .A1(n5585), .A2(n4289), .ZN(n4282) );
  INV_X1 U3838 ( .A(n5585), .ZN(n6172) );
  INV_X1 U3839 ( .A(n5100), .ZN(n5594) );
  INV_X1 U3840 ( .A(n6094), .ZN(n6169) );
  INV_X1 U3841 ( .A(n6318), .ZN(n6272) );
  AND2_X1 U3842 ( .A1(n2978), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6271) );
  INV_X1 U3843 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6390) );
  INV_X1 U3844 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U3845 ( .A1(n4805), .A2(n4804), .ZN(n6181) );
  INV_X1 U3846 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4461) );
  NOR2_X1 U3847 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5194) );
  INV_X1 U3848 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5774) );
  NOR2_X1 U3849 ( .A1(n4602), .A2(n4700), .ZN(n4733) );
  NAND2_X1 U3850 ( .A1(n4544), .A2(n6269), .ZN(n4760) );
  AND2_X1 U3851 ( .A1(n6184), .A2(n6269), .ZN(n6262) );
  INV_X1 U3852 ( .A(n4837), .ZN(n4861) );
  INV_X1 U3853 ( .A(n5009), .ZN(n4727) );
  NAND2_X1 U3854 ( .A1(n4592), .A2(n4700), .ZN(n5009) );
  OAI211_X1 U3855 ( .C1(n6368), .C2(n6514), .A(n6327), .B(n6326), .ZN(n6374)
         );
  INV_X1 U3856 ( .A(n5153), .ZN(n5180) );
  INV_X1 U3857 ( .A(n4643), .ZN(n4931) );
  INV_X1 U3858 ( .A(n5152), .ZN(n5179) );
  AND2_X1 U3859 ( .A1(n3979), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6429) );
  AND2_X1 U3860 ( .A1(n6448), .A2(STATE_REG_1__SCAN_IN), .ZN(n6537) );
  AOI21_X1 U3861 ( .B1(n5232), .B2(REIP_REG_31__SCAN_IN), .A(n3013), .ZN(n4139) );
  NAND2_X1 U3862 ( .A1(n3034), .A2(n3032), .ZN(n3013) );
  NOR2_X1 U3863 ( .A1(n5944), .A2(n5211), .ZN(n5393) );
  OAI21_X1 U3864 ( .B1(n4341), .B2(n6065), .A(n4342), .ZN(U2955) );
  OAI211_X1 U3865 ( .C1(n5538), .C2(n6065), .A(n3102), .B(n3097), .ZN(U2959)
         );
  AOI21_X1 U3866 ( .B1(n6059), .B2(n5425), .A(n5424), .ZN(n3102) );
  NAND2_X1 U3867 ( .A1(n3098), .A2(n6075), .ZN(n3097) );
  NOR3_X1 U3868 ( .A1(n4308), .A2(n4307), .A3(n4306), .ZN(n4309) );
  AND2_X1 U3869 ( .A1(n4305), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4306)
         );
  INV_X1 U3870 ( .A(n4080), .ZN(n4121) );
  AND2_X2 U3871 ( .A1(n4436), .A2(n4443), .ZN(n3328) );
  INV_X1 U3872 ( .A(n4080), .ZN(n4266) );
  NAND2_X1 U3873 ( .A1(n3096), .A2(n3712), .ZN(n5261) );
  NOR2_X1 U3874 ( .A1(n5122), .A2(n3092), .ZN(n2980) );
  NOR2_X1 U3875 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3893) );
  INV_X1 U3876 ( .A(n3893), .ZN(n3919) );
  AND2_X1 U3877 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4436) );
  AND2_X1 U3878 ( .A1(n4278), .A2(n3256), .ZN(n4015) );
  INV_X1 U3879 ( .A(n4015), .ZN(n4080) );
  NAND2_X1 U3880 ( .A1(n4436), .A2(n3117), .ZN(n3140) );
  OR2_X1 U3881 ( .A1(n5122), .A2(n5128), .ZN(n5127) );
  NAND2_X1 U3882 ( .A1(n4345), .A2(n4355), .ZN(n5199) );
  AND2_X1 U3883 ( .A1(n4799), .A2(n3118), .ZN(n3284) );
  AND2_X1 U3884 ( .A1(n3145), .A2(n3108), .ZN(n3220) );
  NOR3_X1 U3885 ( .A1(n5219), .A2(REIP_REG_31__SCAN_IN), .A3(n4012), .ZN(n2984) );
  INV_X1 U3886 ( .A(n3256), .ZN(n3252) );
  NAND2_X1 U3887 ( .A1(n4236), .A2(n3068), .ZN(n3067) );
  OR2_X1 U3888 ( .A1(n5199), .A2(n6063), .ZN(n2985) );
  AND2_X1 U3889 ( .A1(n3185), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n2986) );
  AND2_X1 U3890 ( .A1(n3070), .A2(n3074), .ZN(n2987) );
  NAND2_X1 U3891 ( .A1(n3073), .A2(n3079), .ZN(n5449) );
  AND2_X1 U3892 ( .A1(n3096), .A2(n3095), .ZN(n2988) );
  OAI21_X1 U3893 ( .B1(n5496), .B2(n4228), .A(n4227), .ZN(n5488) );
  NAND2_X1 U3894 ( .A1(n3030), .A2(n3379), .ZN(n3470) );
  INV_X1 U3895 ( .A(n3833), .ZN(n3928) );
  INV_X1 U3897 ( .A(n6396), .ZN(n3016) );
  NAND2_X1 U3898 ( .A1(n3024), .A2(n4217), .ZN(n5074) );
  INV_X1 U3899 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U3900 ( .A1(n3025), .A2(n3060), .ZN(n5706) );
  NAND2_X1 U3901 ( .A1(n3059), .A2(n4222), .ZN(n5090) );
  NAND2_X1 U3902 ( .A1(n2967), .A2(n5716), .ZN(n2989) );
  AND2_X1 U3903 ( .A1(n5251), .A2(n3104), .ZN(n2990) );
  NOR2_X1 U3904 ( .A1(n3255), .A2(n4142), .ZN(n4240) );
  NAND2_X1 U3905 ( .A1(n5051), .A2(n3089), .ZN(n3591) );
  INV_X1 U3906 ( .A(n5685), .ZN(n3018) );
  NAND2_X1 U3907 ( .A1(n3591), .A2(n3084), .ZN(n2991) );
  INV_X1 U3908 ( .A(n5360), .ZN(n3712) );
  AND2_X1 U3909 ( .A1(n4743), .A2(n4744), .ZN(n2992) );
  AND2_X1 U3910 ( .A1(n3017), .A2(n5458), .ZN(n2993) );
  INV_X1 U3911 ( .A(n4187), .ZN(n4207) );
  AND2_X1 U3912 ( .A1(n4278), .A2(n3215), .ZN(n4187) );
  OR2_X1 U3913 ( .A1(n3985), .A2(n3978), .ZN(n2994) );
  OR2_X1 U3914 ( .A1(n3243), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2995)
         );
  AND2_X1 U3915 ( .A1(n4074), .A2(n4073), .ZN(n5761) );
  INV_X1 U3916 ( .A(n5341), .ZN(n3816) );
  INV_X1 U3917 ( .A(n3093), .ZN(n3092) );
  NOR2_X1 U3918 ( .A1(n5281), .A2(n5128), .ZN(n3093) );
  AND2_X1 U3919 ( .A1(n3524), .A2(n4362), .ZN(n2996) );
  AND2_X1 U3920 ( .A1(n2990), .A2(n3103), .ZN(n2997) );
  AND2_X1 U3921 ( .A1(n2989), .A2(n3109), .ZN(n2998) );
  NOR2_X1 U3922 ( .A1(n5861), .A2(n3040), .ZN(n2999) );
  NAND2_X1 U3923 ( .A1(n3420), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3606) );
  INV_X1 U3924 ( .A(n3606), .ZN(n3615) );
  NOR2_X1 U3925 ( .A1(n4043), .A2(n5885), .ZN(n3000) );
  INV_X1 U3926 ( .A(n3579), .ZN(n3088) );
  INV_X1 U3927 ( .A(n5371), .ZN(n3048) );
  OR2_X1 U3928 ( .A1(n6435), .A2(n6318), .ZN(n6063) );
  OR2_X1 U3929 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3001) );
  INV_X1 U3930 ( .A(n5211), .ZN(n4404) );
  NAND3_X1 U3931 ( .A1(n3972), .A2(n3012), .A3(n3011), .ZN(n3010) );
  NAND3_X1 U3932 ( .A1(n4258), .A2(n5770), .A3(n3015), .ZN(n3014) );
  NAND2_X1 U3933 ( .A1(n3239), .A2(n3986), .ZN(n5770) );
  NAND2_X1 U3934 ( .A1(n3238), .A2(n3429), .ZN(n4258) );
  NAND2_X1 U3935 ( .A1(n5706), .A2(n5707), .ZN(n4225) );
  NAND3_X1 U3936 ( .A1(n3470), .A2(n3471), .A3(n4187), .ZN(n4168) );
  INV_X2 U3937 ( .A(n3253), .ZN(n4568) );
  INV_X1 U3938 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3031) );
  NOR2_X2 U3939 ( .A1(n5344), .A2(n3049), .ZN(n3053) );
  OAI21_X2 U3940 ( .B1(n4468), .B2(n4207), .A(n4159), .ZN(n6082) );
  NAND3_X1 U3941 ( .A1(n3062), .A2(n4222), .A3(n3064), .ZN(n3061) );
  NAND2_X1 U3942 ( .A1(n3067), .A2(n2998), .ZN(n5420) );
  NAND2_X1 U3943 ( .A1(n4236), .A2(n4235), .ZN(n5410) );
  INV_X1 U3944 ( .A(n3067), .ZN(n5431) );
  NAND2_X1 U3945 ( .A1(n4225), .A2(n4224), .ZN(n5496) );
  NAND2_X1 U3946 ( .A1(n4225), .A2(n3071), .ZN(n3070) );
  OAI211_X1 U3947 ( .C1(n5051), .C2(n3088), .A(n3591), .B(n3086), .ZN(n5086)
         );
  NAND3_X1 U3948 ( .A1(n4744), .A2(n4743), .A3(n4362), .ZN(n4361) );
  NAND3_X1 U3949 ( .A1(n4744), .A2(n4743), .A3(n2996), .ZN(n4901) );
  NAND2_X1 U3950 ( .A1(n2963), .A2(n2990), .ZN(n5237) );
  AND2_X1 U3951 ( .A1(n2963), .A2(n3104), .ZN(n5250) );
  NAND2_X1 U3952 ( .A1(n2963), .A2(n3816), .ZN(n5334) );
  AND2_X2 U3953 ( .A1(n2963), .A2(n2997), .ZN(n4343) );
  OR2_X1 U3954 ( .A1(n5217), .A2(n6063), .ZN(n3105) );
  NAND2_X1 U3955 ( .A1(n5394), .A2(n5393), .ZN(n5396) );
  XNOR2_X1 U3956 ( .A(n3930), .B(n3929), .ZN(n5394) );
  NOR2_X1 U3957 ( .A1(n4468), .A2(n3379), .ZN(n6184) );
  AND2_X1 U3958 ( .A1(n4240), .A2(n3223), .ZN(n3226) );
  AND3_X1 U3959 ( .A1(n3164), .A2(n3163), .A3(n3162), .ZN(n3106) );
  AND4_X1 U3960 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3107)
         );
  AND2_X1 U3961 ( .A1(n2967), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3109)
         );
  INV_X1 U3962 ( .A(n3429), .ZN(n5210) );
  AND2_X1 U3963 ( .A1(n5211), .A2(n3237), .ZN(n3429) );
  INV_X1 U3964 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6637) );
  AND2_X1 U3965 ( .A1(n5934), .A2(n5211), .ZN(n5931) );
  AND2_X1 U3966 ( .A1(n3976), .A2(n3982), .ZN(n3965) );
  AND2_X1 U3967 ( .A1(n3948), .A2(n3947), .ZN(n3970) );
  INV_X1 U3968 ( .A(n4148), .ZN(n3347) );
  OR2_X1 U3969 ( .A1(n3389), .A2(n3388), .ZN(n4189) );
  NOR2_X1 U3970 ( .A1(n3935), .A2(n3941), .ZN(n3936) );
  AOI22_X1 U3971 ( .A1(n3328), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3171) );
  XNOR2_X1 U3972 ( .A(n4461), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3941)
         );
  AND2_X1 U3973 ( .A1(n6188), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3951)
         );
  NOR2_X1 U3974 ( .A1(n5211), .A2(n6279), .ZN(n3480) );
  INV_X1 U3975 ( .A(n3743), .ZN(n3744) );
  INV_X1 U3976 ( .A(n3480), .ZN(n3833) );
  INV_X1 U3977 ( .A(n5034), .ZN(n3540) );
  NAND2_X1 U3978 ( .A1(n4437), .A2(n6419), .ZN(n3378) );
  NOR2_X1 U3979 ( .A1(n4004), .A2(n5296), .ZN(n5656) );
  NOR2_X1 U3980 ( .A1(n3857), .A2(n5422), .ZN(n3858) );
  NOR2_X1 U3981 ( .A1(n3525), .A2(n5863), .ZN(n3542) );
  OR2_X1 U3982 ( .A1(n4166), .A2(n6531), .ZN(n4167) );
  OR3_X1 U3983 ( .A1(n2967), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5520), 
        .ZN(n4347) );
  NOR2_X1 U3984 ( .A1(n5831), .A2(n5832), .ZN(n4066) );
  NAND2_X1 U3985 ( .A1(n4034), .A2(n4033), .ZN(n4035) );
  INV_X1 U3986 ( .A(n4876), .ZN(n4870) );
  INV_X1 U3987 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5653) );
  INV_X1 U3988 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5840) );
  INV_X1 U3989 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4910) );
  AND3_X1 U3990 ( .A1(n6092), .A2(n6423), .A3(n6430), .ZN(n3991) );
  AND2_X1 U3991 ( .A1(n4406), .A2(n5216), .ZN(n4129) );
  AOI21_X1 U3992 ( .B1(n4186), .B2(n3615), .A(n3492), .ZN(n4497) );
  OR2_X1 U3993 ( .A1(n4451), .A2(n6531), .ZN(n6412) );
  INV_X1 U3994 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6591) );
  INV_X1 U3995 ( .A(n4301), .ZN(n6137) );
  NAND2_X1 U3996 ( .A1(n4291), .A2(n4262), .ZN(n6094) );
  INV_X1 U3997 ( .A(n4512), .ZN(n4806) );
  NAND2_X1 U3998 ( .A1(n4544), .A2(n6183), .ZN(n4971) );
  INV_X1 U3999 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4595) );
  INV_X1 U4000 ( .A(n6262), .ZN(n4860) );
  INV_X1 U4001 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4986) );
  INV_X1 U4002 ( .A(n4824), .ZN(n4700) );
  INV_X1 U4003 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6279) );
  INV_X1 U4004 ( .A(n4136), .ZN(n6531) );
  AND2_X1 U4005 ( .A1(n4310), .A2(n4001), .ZN(n5259) );
  NAND2_X1 U4006 ( .A1(n5028), .A2(n4135), .ZN(n5874) );
  INV_X1 U4007 ( .A(n5659), .ZN(n5879) );
  NOR2_X2 U4008 ( .A1(n5888), .A2(n4316), .ZN(n5912) );
  AND2_X1 U4009 ( .A1(n4065), .A2(n4064), .ZN(n5832) );
  INV_X1 U4010 ( .A(n5934), .ZN(n5386) );
  INV_X1 U4011 ( .A(n5669), .ZN(n5942) );
  INV_X2 U4012 ( .A(n5392), .ZN(n5944) );
  OAI21_X1 U4013 ( .B1(n4136), .B2(n4249), .A(n5970), .ZN(n6043) );
  NAND2_X1 U4014 ( .A1(n3695), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3743)
         );
  INV_X1 U4015 ( .A(n5696), .ZN(n5935) );
  AND2_X1 U4016 ( .A1(n3489), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3503)
         );
  NAND2_X1 U4017 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3472), .ZN(n3481)
         );
  NAND2_X1 U4018 ( .A1(n6065), .A2(n4333), .ZN(n5483) );
  AND2_X1 U4019 ( .A1(n5373), .A2(n5372), .ZN(n5657) );
  AND2_X1 U4020 ( .A1(n4291), .A2(n5141), .ZN(n5100) );
  OR2_X1 U4021 ( .A1(n5103), .A2(n6172), .ZN(n5586) );
  INV_X1 U4022 ( .A(n6095), .ZN(n6175) );
  AND2_X1 U4023 ( .A1(n6397), .A2(n4278), .ZN(n5141) );
  INV_X1 U4024 ( .A(n5190), .ZN(n5186) );
  OAI21_X1 U4025 ( .B1(n4642), .B2(n4641), .A(n4640), .ZN(n4688) );
  INV_X1 U4026 ( .A(n4972), .ZN(n4942) );
  OAI221_X1 U4027 ( .B1(n4974), .B2(n6514), .C1(n4974), .C2(n4948), .A(n4985), 
        .ZN(n4970) );
  OAI21_X1 U4028 ( .B1(n4519), .B2(n4518), .A(n4517), .ZN(n4627) );
  INV_X1 U4029 ( .A(n6190), .ZN(n6217) );
  INV_X1 U4030 ( .A(n6187), .ZN(n6216) );
  INV_X1 U4031 ( .A(n6221), .ZN(n6259) );
  OAI21_X1 U4032 ( .B1(n4836), .B2(n4835), .A(n4834), .ZN(n4859) );
  AND2_X1 U4033 ( .A1(n4592), .A2(n4824), .ZN(n4837) );
  OAI211_X1 U4034 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4986), .A(n4985), .B(n4984), .ZN(n5008) );
  INV_X1 U4035 ( .A(n6377), .ZN(n6319) );
  NOR2_X2 U4036 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4480), .ZN(n4946) );
  INV_X1 U4037 ( .A(n3919), .ZN(n3990) );
  INV_X1 U4038 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6418) );
  INV_X1 U4039 ( .A(n5905), .ZN(n5889) );
  NAND2_X1 U4040 ( .A1(n5064), .A2(n3996), .ZN(n5659) );
  AND2_X1 U4041 ( .A1(n4906), .A2(n5659), .ZN(n5910) );
  AND2_X2 U4042 ( .A1(n4403), .A2(n6429), .ZN(n5934) );
  INV_X1 U4043 ( .A(n5493), .ZN(n5300) );
  INV_X1 U4044 ( .A(n4899), .ZN(n5311) );
  NAND2_X1 U4045 ( .A1(n5392), .A2(n4419), .ZN(n5669) );
  NAND2_X1 U4046 ( .A1(n4418), .A2(n6004), .ZN(n5392) );
  INV_X1 U4047 ( .A(n5948), .ZN(n5968) );
  NAND2_X2 U4048 ( .A1(n4657), .A2(n4656), .ZN(n6052) );
  NAND2_X1 U4049 ( .A1(n5483), .A2(n4336), .ZN(n6090) );
  AND2_X1 U4050 ( .A1(n5571), .A2(n4302), .ZN(n5717) );
  AND2_X1 U4051 ( .A1(n5564), .A2(n5578), .ZN(n5571) );
  OR2_X1 U4052 ( .A1(n6526), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U4053 ( .A1(n4291), .A2(n4261), .ZN(n6095) );
  INV_X1 U4054 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U4055 ( .A1(n6184), .A2(n6183), .ZN(n6221) );
  NAND2_X1 U4056 ( .A1(n6270), .A2(n6183), .ZN(n6307) );
  NAND2_X1 U4057 ( .A1(n6270), .A2(n6269), .ZN(n6377) );
  INV_X1 U4058 ( .A(n4698), .ZN(n4783) );
  INV_X1 U4059 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6514) );
  INV_X1 U4060 ( .A(n6701), .ZN(n6438) );
  INV_X1 U4061 ( .A(n6501), .ZN(n6508) );
  AND2_X2 U4062 ( .A1(n3117), .A2(n4799), .ZN(n3335) );
  AOI22_X1 U4063 ( .A1(n3335), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4064 ( .A1(n2977), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4065 ( .A1(n3329), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3114) );
  AND2_X4 U4066 ( .A1(n4443), .A2(n5145), .ZN(n3782) );
  AOI22_X1 U4067 ( .A1(n3782), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3123) );
  AND2_X2 U4068 ( .A1(n4443), .A2(n3119), .ZN(n3187) );
  AOI22_X1 U4069 ( .A1(n2965), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3122) );
  AND2_X2 U4070 ( .A1(n3117), .A2(n5145), .ZN(n3185) );
  AOI22_X1 U4071 ( .A1(n2968), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3121) );
  AND2_X2 U4072 ( .A1(n3125), .A2(n3124), .ZN(n3221) );
  AOI22_X1 U4073 ( .A1(n2976), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4074 ( .A1(n2964), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3126) );
  AND4_X2 U4075 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n3135)
         );
  AOI22_X1 U4076 ( .A1(n3161), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4077 ( .A1(n3185), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4078 ( .A1(n3185), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4079 ( .A1(n3335), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4080 ( .A1(n3328), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4081 ( .A1(n3782), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4082 ( .A1(n2969), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4083 ( .A1(n3184), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4084 ( .A1(n2974), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4085 ( .A1(n4398), .A2(n3220), .ZN(n3156) );
  AOI22_X1 U4086 ( .A1(n2968), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4087 ( .A1(n3335), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4088 ( .A1(n3328), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4089 ( .A1(n3184), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3146) );
  NAND4_X1 U4090 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3155)
         );
  AOI22_X1 U4091 ( .A1(n3161), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4092 ( .A1(n3782), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4093 ( .A1(n2964), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3150) );
  NAND4_X1 U4094 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3154)
         );
  NAND2_X1 U4095 ( .A1(n3156), .A2(n5211), .ZN(n3166) );
  AOI22_X1 U4096 ( .A1(n3329), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4097 ( .A1(n2966), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4098 ( .A1(n3782), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4099 ( .A1(n2968), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4100 ( .A1(n3328), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4101 ( .A1(n2975), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4102 ( .A1(n3335), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4103 ( .A1(n2969), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U4104 ( .A1(n3456), .A2(n4399), .ZN(n3251) );
  NAND2_X1 U4105 ( .A1(n3166), .A2(n3251), .ZN(n3178) );
  AOI22_X1 U4106 ( .A1(n3329), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4107 ( .A1(n3161), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4108 ( .A1(n3335), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4109 ( .A1(n2976), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U4110 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3176)
         );
  AOI22_X1 U4111 ( .A1(n3185), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4112 ( .A1(n3782), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4113 ( .A1(n2966), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3172) );
  NAND4_X1 U4114 ( .A1(n3174), .A2(n3173), .A3(n3172), .A4(n3171), .ZN(n3175)
         );
  NAND2_X1 U4115 ( .A1(n3217), .A2(n3256), .ZN(n3177) );
  INV_X1 U4116 ( .A(n3456), .ZN(n3179) );
  NAND2_X1 U4117 ( .A1(n2981), .A2(n3179), .ZN(n3987) );
  AOI22_X1 U4118 ( .A1(n2969), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4119 ( .A1(n3329), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4120 ( .A1(n3335), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4121 ( .A1(n3904), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3180) );
  NAND4_X1 U4122 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3193)
         );
  AOI22_X1 U4123 ( .A1(n3185), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4124 ( .A1(n3782), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3284), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4125 ( .A1(n2966), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3186), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4126 ( .A1(n3328), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3188) );
  NAND4_X1 U4127 ( .A1(n3191), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3192)
         );
  AOI21_X1 U4128 ( .B1(n3987), .B2(n4265), .A(n4278), .ZN(n3194) );
  NAND2_X1 U4129 ( .A1(n3986), .A2(n3194), .ZN(n3214) );
  NAND2_X1 U4130 ( .A1(n3161), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4131 ( .A1(n3329), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3198) );
  NAND2_X1 U4132 ( .A1(n2964), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4133 ( .A1(n3862), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4134 ( .A1(n3782), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4135 ( .A1(n2966), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3201)
         );
  NAND2_X1 U4136 ( .A1(n3284), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4137 ( .A1(n3334), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3206)
         );
  NAND2_X1 U4138 ( .A1(n2977), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4139 ( .A1(n3184), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4140 ( .A1(n3879), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3203)
         );
  NAND2_X1 U4141 ( .A1(n3335), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4142 ( .A1(n3328), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3210)
         );
  NAND2_X1 U4143 ( .A1(n3207), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3209)
         );
  NAND2_X1 U4144 ( .A1(n3186), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4145 ( .A1(n3214), .A2(n4568), .ZN(n3246) );
  NAND2_X1 U4146 ( .A1(n3232), .A2(n4136), .ZN(n3216) );
  AND2_X1 U4147 ( .A1(n3247), .A2(n3215), .ZN(n4255) );
  NAND2_X1 U4148 ( .A1(n4255), .A2(n4015), .ZN(n4438) );
  INV_X1 U4149 ( .A(n3217), .ZN(n3224) );
  NAND2_X1 U4150 ( .A1(n3224), .A2(n3247), .ZN(n3219) );
  AND2_X1 U4151 ( .A1(n4398), .A2(n5211), .ZN(n3218) );
  NAND2_X1 U4152 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6440) );
  OAI21_X1 U4153 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6440), .ZN(n3997) );
  NAND2_X1 U4154 ( .A1(n3946), .A2(n3997), .ZN(n3236) );
  NAND2_X1 U4155 ( .A1(n3236), .A2(n3222), .ZN(n3223) );
  NOR2_X1 U4156 ( .A1(n3257), .A2(n4568), .ZN(n3225) );
  NAND2_X1 U4157 ( .A1(n3232), .A2(n3225), .ZN(n4269) );
  NAND4_X1 U4158 ( .A1(n3246), .A2(n3261), .A3(n3226), .A4(n4269), .ZN(n3227)
         );
  AND2_X2 U4159 ( .A1(n3227), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3266) );
  INV_X1 U4160 ( .A(n3266), .ZN(n3240) );
  NAND2_X1 U4161 ( .A1(n5194), .A2(n6419), .ZN(n6526) );
  INV_X1 U4162 ( .A(n6526), .ZN(n3270) );
  NAND2_X1 U4163 ( .A1(n6188), .A2(n4595), .ZN(n3228) );
  NAND2_X1 U4164 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4165 ( .A1(n3270), .A2(n4947), .ZN(n3231) );
  INV_X1 U4166 ( .A(n3979), .ZN(n3229) );
  NAND2_X1 U4167 ( .A1(n3229), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3230) );
  INV_X1 U4168 ( .A(n3232), .ZN(n3234) );
  NOR2_X1 U4169 ( .A1(n4142), .A2(n3215), .ZN(n3233) );
  NAND2_X1 U4170 ( .A1(n3234), .A2(n3233), .ZN(n4248) );
  INV_X1 U4171 ( .A(n4248), .ZN(n3235) );
  NAND2_X1 U4172 ( .A1(n3235), .A2(n3253), .ZN(n6396) );
  INV_X1 U4173 ( .A(n4275), .ZN(n3238) );
  NOR2_X1 U4174 ( .A1(n3987), .A2(n3948), .ZN(n3239) );
  OAI211_X2 U4175 ( .C1(n3240), .C2(n3112), .A(n3242), .B(n3241), .ZN(n3265)
         );
  INV_X1 U4176 ( .A(n3242), .ZN(n3243) );
  INV_X1 U4177 ( .A(n3295), .ZN(n3264) );
  NAND2_X1 U4178 ( .A1(n3266), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3324) );
  MUX2_X1 U4179 ( .A(n3979), .B(n6526), .S(n6188), .Z(n3323) );
  NAND2_X1 U4180 ( .A1(n3324), .A2(n3323), .ZN(n3263) );
  INV_X1 U4181 ( .A(n3246), .ZN(n3250) );
  NAND2_X1 U4182 ( .A1(n4187), .A2(n3247), .ZN(n3249) );
  NAND2_X1 U4183 ( .A1(n3257), .A2(n4136), .ZN(n4242) );
  OAI21_X1 U4184 ( .B1(n4568), .B2(n3220), .A(n4242), .ZN(n3248) );
  NAND2_X1 U4185 ( .A1(n5194), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5780) );
  INV_X1 U4186 ( .A(n5780), .ZN(n6428) );
  NAND2_X1 U4187 ( .A1(n3252), .A2(n3253), .ZN(n4018) );
  OAI211_X1 U4188 ( .C1(n3251), .C2(n4273), .A(n6428), .B(n4018), .ZN(n3254)
         );
  INV_X1 U4189 ( .A(n3254), .ZN(n3260) );
  OAI21_X1 U4190 ( .B1(n3257), .B2(n3247), .A(n3256), .ZN(n3258) );
  OAI21_X1 U4191 ( .B1(n3255), .B2(n3258), .A(n4278), .ZN(n3259) );
  NAND2_X1 U4192 ( .A1(n4272), .A2(n3262), .ZN(n3321) );
  NAND2_X1 U4193 ( .A1(n3264), .A2(n3326), .ZN(n3278) );
  BUF_X1 U4194 ( .A(n3265), .Z(n3275) );
  NAND2_X1 U4195 ( .A1(n3278), .A2(n3275), .ZN(n3273) );
  INV_X1 U4196 ( .A(n3268), .ZN(n3267) );
  NAND2_X1 U4197 ( .A1(n3267), .A2(n6665), .ZN(n6268) );
  NAND2_X1 U4198 ( .A1(n3268), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4199 ( .A1(n6268), .A2(n3269), .ZN(n4515) );
  NAND2_X1 U4200 ( .A1(n3270), .A2(n4515), .ZN(n3271) );
  OAI21_X1 U4201 ( .B1(n3979), .B2(n6665), .A(n3271), .ZN(n3272) );
  AOI21_X2 U4202 ( .B1(n3360), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3272), 
        .ZN(n3274) );
  NAND2_X1 U4203 ( .A1(n3273), .A2(n3274), .ZN(n3279) );
  INV_X1 U4204 ( .A(n3274), .ZN(n3276) );
  AND2_X2 U4205 ( .A1(n3276), .A2(n3275), .ZN(n3277) );
  NAND2_X2 U4206 ( .A1(n3278), .A2(n3277), .ZN(n4800) );
  AOI22_X1 U4207 ( .A1(n3896), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3283) );
  INV_X1 U4208 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6639) );
  AOI22_X1 U4209 ( .A1(n3903), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4210 ( .A1(n3907), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4211 ( .A1(n2977), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3280) );
  NAND4_X1 U4212 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3290)
         );
  AOI22_X1 U4213 ( .A1(n3185), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4214 ( .A1(n3663), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4215 ( .A1(n3898), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4216 ( .A1(n3307), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4217 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  OAI22_X2 U4218 ( .A1(n4470), .A2(STATE2_REG_0__SCAN_IN), .B1(n4164), .B2(
        n3366), .ZN(n3294) );
  INV_X1 U4219 ( .A(n3365), .ZN(n3292) );
  AOI22_X1 U4220 ( .A1(n3973), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3292), 
        .B2(n3291), .ZN(n3293) );
  XNOR2_X1 U4221 ( .A(n3295), .B(n3326), .ZN(n4471) );
  AOI22_X1 U4222 ( .A1(n3663), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4223 ( .A1(n3329), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4224 ( .A1(n2973), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4225 ( .A1(n3879), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3296) );
  NAND4_X1 U4226 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3305)
         );
  AOI22_X1 U4227 ( .A1(n3185), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4228 ( .A1(n3896), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4229 ( .A1(n3907), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4230 ( .A1(n3905), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4231 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  OAI21_X2 U4232 ( .B1(n2979), .B2(STATE2_REG_0__SCAN_IN), .A(n3306), .ZN(
        n3440) );
  AOI22_X1 U4233 ( .A1(n2968), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4234 ( .A1(n2974), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4235 ( .A1(n3334), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4236 ( .A1(n3905), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3308) );
  NAND4_X1 U4237 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3317)
         );
  AOI22_X1 U4238 ( .A1(n3896), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3329), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4239 ( .A1(n3335), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4240 ( .A1(n3663), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4241 ( .A1(n2973), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3312) );
  NAND4_X1 U4242 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3316)
         );
  NAND2_X1 U4243 ( .A1(n3973), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3320) );
  OR2_X1 U4244 ( .A1(n3365), .A2(n3318), .ZN(n3319) );
  OAI211_X1 U4245 ( .C1(n3366), .C2(n4211), .A(n3320), .B(n3319), .ZN(n3438)
         );
  NAND2_X1 U4246 ( .A1(n3440), .A2(n3438), .ZN(n3355) );
  INV_X1 U4247 ( .A(n3321), .ZN(n3322) );
  AND2_X1 U4248 ( .A1(n3323), .A2(n3322), .ZN(n3325) );
  NAND2_X1 U4249 ( .A1(n3325), .A2(n3324), .ZN(n3327) );
  AND2_X2 U4250 ( .A1(n3327), .A2(n3326), .ZN(n3446) );
  NAND2_X1 U4251 ( .A1(n3446), .A2(n6419), .ZN(n3450) );
  NAND2_X1 U4252 ( .A1(n3973), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4253 ( .A1(n2975), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4254 ( .A1(n3185), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4255 ( .A1(n3307), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4256 ( .A1(n3329), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3330) );
  NAND4_X1 U4257 ( .A1(n3333), .A2(n3332), .A3(n3331), .A4(n3330), .ZN(n3341)
         );
  AOI22_X1 U4258 ( .A1(n3896), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4259 ( .A1(n2971), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4260 ( .A1(n3898), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4261 ( .A1(n3907), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3336) );
  NAND4_X1 U4262 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3340)
         );
  AOI21_X1 U4263 ( .B1(n4568), .B2(n4148), .A(n6419), .ZN(n3342) );
  AND2_X1 U4264 ( .A1(n3342), .A2(n3351), .ZN(n3343) );
  NAND2_X1 U4265 ( .A1(n3344), .A2(n3343), .ZN(n3449) );
  INV_X1 U4266 ( .A(n4211), .ZN(n3345) );
  NAND2_X1 U4267 ( .A1(n3345), .A2(n3247), .ZN(n3346) );
  NAND2_X1 U4268 ( .A1(n3449), .A2(n3451), .ZN(n3454) );
  INV_X1 U4269 ( .A(n3351), .ZN(n3352) );
  NAND2_X1 U4270 ( .A1(n3352), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4208) );
  INV_X1 U4271 ( .A(n3439), .ZN(n3354) );
  NAND2_X1 U4272 ( .A1(n3355), .A2(n3354), .ZN(n3359) );
  INV_X1 U4273 ( .A(n3440), .ZN(n3357) );
  INV_X1 U4274 ( .A(n3438), .ZN(n3356) );
  NAND2_X1 U4275 ( .A1(n3357), .A2(n3356), .ZN(n3358) );
  AND2_X2 U4276 ( .A1(n3359), .A2(n3358), .ZN(n3436) );
  NAND2_X1 U4277 ( .A1(n3360), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3364) );
  NOR3_X1 U4278 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6665), .A3(n4595), 
        .ZN(n6233) );
  NAND2_X1 U4279 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6233), .ZN(n6224) );
  NAND2_X1 U4280 ( .A1(n6390), .A2(n6224), .ZN(n3361) );
  NAND3_X1 U4281 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5150) );
  INV_X1 U4282 ( .A(n5150), .ZN(n4874) );
  NAND2_X1 U4283 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4874), .ZN(n4932) );
  NAND2_X1 U4284 ( .A1(n3361), .A2(n4932), .ZN(n4830) );
  OAI22_X1 U4285 ( .A1(n6526), .A2(n4830), .B1(n3979), .B2(n6390), .ZN(n3362)
         );
  INV_X1 U4286 ( .A(n3362), .ZN(n3363) );
  XNOR2_X2 U4287 ( .A(n4800), .B(n4513), .ZN(n4437) );
  AOI22_X1 U4288 ( .A1(n3896), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4289 ( .A1(n3898), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4290 ( .A1(n3903), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4291 ( .A1(n3907), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4292 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3376)
         );
  AOI22_X1 U4293 ( .A1(n3624), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4294 ( .A1(n2974), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4295 ( .A1(n3897), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4296 ( .A1(n2971), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4297 ( .A1(n3374), .A2(n3373), .A3(n3372), .A4(n3371), .ZN(n3375)
         );
  AOI22_X1 U4298 ( .A1(n3976), .A2(n4171), .B1(n3973), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3377) );
  INV_X1 U4299 ( .A(n3470), .ZN(n3392) );
  AOI22_X1 U4300 ( .A1(n3896), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4301 ( .A1(n3903), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4302 ( .A1(n3907), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4303 ( .A1(n2975), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3380) );
  NAND4_X1 U4304 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3389)
         );
  AOI22_X1 U4305 ( .A1(n3624), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4306 ( .A1(n3663), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4307 ( .A1(n3898), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4308 ( .A1(n3307), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3384) );
  NAND4_X1 U4309 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3388)
         );
  NAND2_X1 U4310 ( .A1(n3976), .A2(n4189), .ZN(n3391) );
  NAND2_X1 U4311 ( .A1(n3973), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4312 ( .A1(n3391), .A2(n3390), .ZN(n3425) );
  INV_X1 U4313 ( .A(n3479), .ZN(n3405) );
  AOI22_X1 U4314 ( .A1(n3663), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4315 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3307), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4316 ( .A1(n3907), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4317 ( .A1(n3903), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4318 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3402)
         );
  AOI22_X1 U4319 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n3624), .B1(n2971), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4320 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n3898), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4321 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n3896), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4322 ( .A1(n2974), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4323 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  NAND2_X1 U4324 ( .A1(n3976), .A2(n4188), .ZN(n3404) );
  NAND2_X1 U4325 ( .A1(n3973), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4326 ( .A1(n3404), .A2(n3403), .ZN(n3478) );
  NAND2_X1 U4327 ( .A1(n3405), .A2(n3478), .ZN(n3488) );
  INV_X1 U4328 ( .A(n3488), .ZN(n3418) );
  AOI22_X1 U4329 ( .A1(n3896), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4330 ( .A1(n3903), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4331 ( .A1(n3907), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4332 ( .A1(n2975), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3406) );
  NAND4_X1 U4333 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n3415)
         );
  AOI22_X1 U4334 ( .A1(n3624), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4335 ( .A1(n3663), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4336 ( .A1(n3898), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3411) );
  INV_X1 U4337 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U4338 ( .A1(n3307), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3410) );
  NAND4_X1 U4339 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n3414)
         );
  NAND2_X1 U4340 ( .A1(n3976), .A2(n4199), .ZN(n3417) );
  NAND2_X1 U4341 ( .A1(n3973), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3416) );
  NAND2_X1 U4342 ( .A1(n3418), .A2(n3487), .ZN(n4206) );
  AOI22_X1 U4343 ( .A1(n3976), .A2(n4211), .B1(n3973), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3419) );
  XNOR2_X1 U4344 ( .A(n4206), .B(n3419), .ZN(n4197) );
  INV_X1 U4345 ( .A(n4197), .ZN(n3421) );
  NAND2_X1 U4346 ( .A1(n3421), .A2(n3615), .ZN(n3424) );
  INV_X1 U4347 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4897) );
  XNOR2_X1 U4348 ( .A(n3503), .B(n4897), .ZN(n5303) );
  NAND2_X1 U4349 ( .A1(n4986), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3792) );
  OAI22_X1 U4350 ( .A1(n5303), .A2(n3919), .B1(n3792), .B2(n4897), .ZN(n3422)
         );
  AOI21_X1 U4351 ( .B1(n3928), .B2(EAX_REG_7__SCAN_IN), .A(n3422), .ZN(n3423)
         );
  NAND2_X1 U4352 ( .A1(n3424), .A2(n3423), .ZN(n4743) );
  INV_X1 U4353 ( .A(n3425), .ZN(n3426) );
  NAND2_X1 U4354 ( .A1(n3470), .A2(n3426), .ZN(n3427) );
  NAND2_X1 U4355 ( .A1(n3427), .A2(n3479), .ZN(n4175) );
  INV_X1 U4356 ( .A(n4175), .ZN(n3428) );
  NAND2_X1 U4357 ( .A1(n3428), .A2(n3615), .ZN(n3434) );
  OAI21_X1 U4358 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3472), .A(n3481), 
        .ZN(n6079) );
  AND2_X1 U4359 ( .A1(n3429), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3458) );
  INV_X1 U4360 ( .A(n3458), .ZN(n3476) );
  INV_X1 U4361 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5890) );
  AOI21_X1 U4362 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5890), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3430) );
  AOI21_X1 U4363 ( .B1(n3928), .B2(EAX_REG_4__SCAN_IN), .A(n3430), .ZN(n3431)
         );
  OAI21_X1 U4364 ( .B1(n5774), .B2(n3476), .A(n3431), .ZN(n3432) );
  OAI21_X1 U4365 ( .B1(n3919), .B2(n6079), .A(n3432), .ZN(n3433) );
  NAND2_X1 U4366 ( .A1(n3434), .A2(n3433), .ZN(n4494) );
  NOR2_X1 U4367 ( .A1(n4468), .A2(n3606), .ZN(n3437) );
  NOR2_X1 U4368 ( .A1(n3437), .A2(n3927), .ZN(n4423) );
  XNOR2_X1 U4369 ( .A(n3439), .B(n3438), .ZN(n3441) );
  NAND2_X1 U4370 ( .A1(n4469), .A2(n3615), .ZN(n3445) );
  AOI22_X1 U4371 ( .A1(n3928), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6279), .ZN(n3443) );
  NAND2_X1 U4372 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3442) );
  AND2_X1 U4373 ( .A1(n3443), .A2(n3442), .ZN(n3444) );
  NAND2_X1 U4374 ( .A1(n3445), .A2(n3444), .ZN(n4393) );
  INV_X1 U4375 ( .A(n3446), .ZN(n5322) );
  AOI22_X1 U4376 ( .A1(n3928), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6279), .ZN(n3448) );
  NAND2_X1 U4377 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3447) );
  OAI211_X1 U4378 ( .C1(n5322), .C2(n3606), .A(n3448), .B(n3447), .ZN(n4386)
         );
  NAND2_X1 U4379 ( .A1(n3450), .A2(n3449), .ZN(n3453) );
  INV_X1 U4380 ( .A(n3451), .ZN(n3452) );
  NAND2_X1 U4381 ( .A1(n3453), .A2(n3452), .ZN(n3455) );
  AOI21_X1 U4382 ( .B1(n4824), .B2(n3456), .A(n6279), .ZN(n4387) );
  NAND2_X1 U4383 ( .A1(n4387), .A2(n4386), .ZN(n3457) );
  NAND2_X1 U4384 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3463) );
  INV_X1 U4385 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3460) );
  OAI21_X1 U4386 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3473), .ZN(n6089) );
  NAND2_X1 U4387 ( .A1(n3893), .A2(n6089), .ZN(n3459) );
  OAI21_X1 U4388 ( .B1(n3792), .B2(n3460), .A(n3459), .ZN(n3461) );
  AOI21_X1 U4389 ( .B1(n3928), .B2(EAX_REG_2__SCAN_IN), .A(n3461), .ZN(n3462)
         );
  NAND2_X1 U4390 ( .A1(n3463), .A2(n3462), .ZN(n3466) );
  NAND2_X1 U4391 ( .A1(n3465), .A2(n3466), .ZN(n3464) );
  NAND2_X1 U4392 ( .A1(n4423), .A2(n3464), .ZN(n3468) );
  INV_X1 U4393 ( .A(n3466), .ZN(n4424) );
  NAND2_X1 U4394 ( .A1(n4425), .A2(n4424), .ZN(n3467) );
  NAND2_X1 U4395 ( .A1(n3468), .A2(n3467), .ZN(n4422) );
  NAND2_X1 U4396 ( .A1(n3469), .A2(n4539), .ZN(n3471) );
  AOI21_X1 U4397 ( .B1(n6591), .B2(n3473), .A(n3472), .ZN(n5913) );
  OAI22_X1 U4398 ( .A1(n5913), .A2(n3919), .B1(n3792), .B2(n6591), .ZN(n3474)
         );
  AOI21_X1 U4399 ( .B1(n3928), .B2(EAX_REG_3__SCAN_IN), .A(n3474), .ZN(n3475)
         );
  OAI21_X1 U4400 ( .B1(n4461), .B2(n3476), .A(n3475), .ZN(n3477) );
  AOI21_X1 U4401 ( .B1(n4512), .B2(n3615), .A(n3477), .ZN(n4429) );
  NAND2_X1 U4402 ( .A1(n4494), .A2(n4428), .ZN(n4502) );
  INV_X1 U4403 ( .A(n4502), .ZN(n3486) );
  XNOR2_X1 U4404 ( .A(n3479), .B(n3478), .ZN(n4178) );
  INV_X1 U4405 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3483) );
  XNOR2_X1 U4406 ( .A(n3481), .B(n4910), .ZN(n4907) );
  AOI22_X1 U4407 ( .A1(n4907), .A2(n3990), .B1(n3927), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3482) );
  OAI21_X1 U4408 ( .B1(n3833), .B2(n3483), .A(n3482), .ZN(n3484) );
  NAND2_X1 U4409 ( .A1(n3486), .A2(n3485), .ZN(n4498) );
  XNOR2_X1 U4410 ( .A(n3488), .B(n3487), .ZN(n4186) );
  INV_X1 U4411 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4828) );
  NOR2_X1 U4412 ( .A1(n3489), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3490)
         );
  OR2_X1 U4413 ( .A1(n3503), .A2(n3490), .ZN(n6070) );
  AOI22_X1 U4414 ( .A1(n6070), .A2(n3990), .B1(n3927), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3491) );
  OAI21_X1 U4415 ( .B1(n3833), .B2(n4828), .A(n3491), .ZN(n3492) );
  NOR2_X2 U4416 ( .A1(n4498), .A2(n4497), .ZN(n4744) );
  AOI22_X1 U4417 ( .A1(n3896), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4418 ( .A1(n3663), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4419 ( .A1(n3307), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4420 ( .A1(n2977), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4421 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3502)
         );
  AOI22_X1 U4422 ( .A1(n3903), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4423 ( .A1(n3905), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4424 ( .A1(n3624), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4425 ( .A1(n3907), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4426 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  OAI21_X1 U4427 ( .B1(n3502), .B2(n3501), .A(n3615), .ZN(n3507) );
  NAND2_X1 U4428 ( .A1(n3928), .A2(EAX_REG_8__SCAN_IN), .ZN(n3506) );
  XNOR2_X1 U4429 ( .A(n3508), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U4430 ( .A1(n5020), .A2(n3990), .ZN(n3505) );
  NAND2_X1 U4431 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3504)
         );
  NAND4_X1 U4432 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n4362)
         );
  XNOR2_X1 U4433 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3525), .ZN(n5867) );
  INV_X1 U4434 ( .A(n5867), .ZN(n3523) );
  AOI22_X1 U4435 ( .A1(n3896), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4436 ( .A1(n3905), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4437 ( .A1(n3907), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4438 ( .A1(n3903), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4439 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3518)
         );
  AOI22_X1 U4440 ( .A1(n3663), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4441 ( .A1(n3624), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4442 ( .A1(n2976), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4443 ( .A1(n3307), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4444 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3517)
         );
  OAI21_X1 U4445 ( .B1(n3518), .B2(n3517), .A(n3615), .ZN(n3521) );
  NAND2_X1 U4446 ( .A1(n3928), .A2(EAX_REG_9__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4447 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3519)
         );
  NAND3_X1 U4448 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3522) );
  AOI21_X1 U4449 ( .B1(n3523), .B2(n3990), .A(n3522), .ZN(n4903) );
  INV_X1 U4450 ( .A(n4901), .ZN(n3541) );
  XNOR2_X1 U4451 ( .A(n3542), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5850)
         );
  AOI22_X1 U4452 ( .A1(n3307), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4453 ( .A1(n2973), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4454 ( .A1(n2971), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4455 ( .A1(n3898), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4456 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3535)
         );
  AOI22_X1 U4457 ( .A1(n3624), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2974), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4458 ( .A1(n3896), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4459 ( .A1(n3907), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4460 ( .A1(n3663), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4461 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3534)
         );
  OAI21_X1 U4462 ( .B1(n3535), .B2(n3534), .A(n3615), .ZN(n3538) );
  NAND2_X1 U4463 ( .A1(n3928), .A2(EAX_REG_10__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4464 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3536)
         );
  NAND3_X1 U4465 ( .A1(n3538), .A2(n3537), .A3(n3536), .ZN(n3539) );
  AOI21_X1 U4466 ( .B1(n5850), .B2(n3990), .A(n3539), .ZN(n5034) );
  XNOR2_X1 U4467 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3558), .ZN(n6058)
         );
  INV_X1 U4468 ( .A(n6058), .ZN(n3557) );
  AOI22_X1 U4469 ( .A1(n3898), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4470 ( .A1(n2971), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4471 ( .A1(n3907), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4472 ( .A1(n3663), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4473 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3552)
         );
  AOI22_X1 U4474 ( .A1(n3896), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2975), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4475 ( .A1(n3903), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4476 ( .A1(n3307), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4477 ( .A1(n3624), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4478 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3551)
         );
  OAI21_X1 U4479 ( .B1(n3552), .B2(n3551), .A(n3615), .ZN(n3555) );
  NAND2_X1 U4480 ( .A1(n3928), .A2(EAX_REG_11__SCAN_IN), .ZN(n3554) );
  NAND2_X1 U4481 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3553)
         );
  NAND3_X1 U4482 ( .A1(n3555), .A2(n3554), .A3(n3553), .ZN(n3556) );
  AOI21_X1 U4483 ( .B1(n3557), .B2(n3990), .A(n3556), .ZN(n5052) );
  XNOR2_X1 U4484 ( .A(n3574), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5115)
         );
  NAND2_X1 U4485 ( .A1(n5115), .A2(n3990), .ZN(n3573) );
  INV_X1 U4486 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5081) );
  INV_X1 U4487 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3559) );
  OAI22_X1 U4488 ( .A1(n3833), .A2(n5081), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3559), .ZN(n3571) );
  AOI22_X1 U4489 ( .A1(n3896), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4490 ( .A1(n3307), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4491 ( .A1(n3663), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4492 ( .A1(n2974), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4493 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3569)
         );
  AOI22_X1 U4494 ( .A1(n2971), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4495 ( .A1(n3624), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4496 ( .A1(n3903), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4497 ( .A1(n3898), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3564) );
  NAND4_X1 U4498 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3568)
         );
  OR2_X1 U4499 ( .A1(n3569), .A2(n3568), .ZN(n3570) );
  AOI22_X1 U4500 ( .A1(n3571), .A2(n3919), .B1(n3615), .B2(n3570), .ZN(n3572)
         );
  INV_X1 U4501 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3577) );
  OAI21_X1 U4502 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3575), .A(n3618), 
        .ZN(n5830) );
  NAND2_X1 U4503 ( .A1(n5830), .A2(n3990), .ZN(n3576) );
  OAI21_X1 U4504 ( .B1(n3577), .B2(n3792), .A(n3576), .ZN(n3578) );
  AOI21_X1 U4505 ( .B1(n3928), .B2(EAX_REG_13__SCAN_IN), .A(n3578), .ZN(n3579)
         );
  AOI22_X1 U4506 ( .A1(n3896), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4507 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n3624), .B1(n3307), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4508 ( .A1(n3903), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4509 ( .A1(n3907), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        INSTQUEUE_REG_8__5__SCAN_IN), .B2(n3862), .ZN(n3580) );
  NAND4_X1 U4510 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3589)
         );
  AOI22_X1 U4511 ( .A1(n2973), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4512 ( .A1(n2975), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4513 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3898), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4514 ( .A1(n2971), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3584) );
  NAND4_X1 U4515 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3588)
         );
  OR2_X1 U4516 ( .A1(n3589), .A2(n3588), .ZN(n3590) );
  AND2_X1 U4517 ( .A1(n3615), .A2(n3590), .ZN(n5084) );
  NAND2_X1 U4518 ( .A1(n5086), .A2(n3591), .ZN(n5120) );
  AOI22_X1 U4519 ( .A1(n3624), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4520 ( .A1(n3307), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4521 ( .A1(n3898), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4522 ( .A1(n3907), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4523 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  AOI22_X1 U4524 ( .A1(n3896), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4525 ( .A1(n2975), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4526 ( .A1(n3905), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4527 ( .A1(n2971), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4528 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  NOR2_X1 U4529 ( .A1(n3601), .A2(n3600), .ZN(n3605) );
  XNOR2_X1 U4530 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3618), .ZN(n5815)
         );
  INV_X1 U4531 ( .A(n5815), .ZN(n3602) );
  AOI22_X1 U4532 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3990), 
        .B2(n3602), .ZN(n3604) );
  NAND2_X1 U4533 ( .A1(n3928), .A2(EAX_REG_14__SCAN_IN), .ZN(n3603) );
  OAI211_X1 U4534 ( .C1(n3606), .C2(n3605), .A(n3604), .B(n3603), .ZN(n5123)
         );
  NAND2_X1 U4535 ( .A1(n5120), .A2(n5123), .ZN(n5122) );
  AOI22_X1 U4536 ( .A1(n3903), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4537 ( .A1(n3896), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4538 ( .A1(n2974), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4539 ( .A1(n3898), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4540 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3617)
         );
  AOI22_X1 U4541 ( .A1(n3624), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4542 ( .A1(n3907), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4543 ( .A1(n3663), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4544 ( .A1(n3879), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4545 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3616)
         );
  OAI21_X1 U4546 ( .B1(n3617), .B2(n3616), .A(n3615), .ZN(n3621) );
  XNOR2_X1 U4547 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3622), .ZN(n5491)
         );
  AOI22_X1 U4548 ( .A1(n3990), .A2(n5491), .B1(n3927), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4549 ( .A1(n3928), .A2(EAX_REG_15__SCAN_IN), .ZN(n3619) );
  AOI21_X1 U4550 ( .B1(n6637), .B2(n3623), .A(n3640), .ZN(n5485) );
  OR2_X1 U4551 ( .A1(n5485), .A2(n3919), .ZN(n3639) );
  AOI22_X1 U4552 ( .A1(n3624), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4553 ( .A1(n3663), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4554 ( .A1(n3307), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4555 ( .A1(n3905), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4556 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3634)
         );
  AOI22_X1 U4557 ( .A1(n3896), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4558 ( .A1(n2971), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4559 ( .A1(n3903), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4560 ( .A1(n2977), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4561 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  OR2_X1 U4562 ( .A1(n3634), .A2(n3633), .ZN(n3637) );
  INV_X1 U4563 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3635) );
  OAI22_X1 U4564 ( .A1(n3833), .A2(n3635), .B1(n3792), .B2(n6637), .ZN(n3636)
         );
  AOI21_X1 U4565 ( .B1(n3890), .B2(n3637), .A(n3636), .ZN(n3638) );
  OR2_X1 U4566 ( .A1(n3640), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3643)
         );
  INV_X1 U4567 ( .A(n3674), .ZN(n3642) );
  AOI22_X1 U4568 ( .A1(n3896), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4569 ( .A1(n3903), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4570 ( .A1(n3907), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4571 ( .A1(n2974), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4572 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3653)
         );
  AOI22_X1 U4573 ( .A1(n3624), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4574 ( .A1(n3782), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4575 ( .A1(n3898), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4576 ( .A1(n3307), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4577 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3652)
         );
  OR2_X1 U4578 ( .A1(n3653), .A2(n3652), .ZN(n3657) );
  INV_X1 U4579 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3655) );
  INV_X1 U4580 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5784) );
  OAI21_X1 U4581 ( .B1(n5784), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6279), 
        .ZN(n3654) );
  OAI21_X1 U4582 ( .B1(n3833), .B2(n3655), .A(n3654), .ZN(n3656) );
  AOI21_X1 U4583 ( .B1(n3890), .B2(n3657), .A(n3656), .ZN(n3658) );
  AOI21_X1 U4584 ( .B1(n5703), .B2(n3990), .A(n3658), .ZN(n5273) );
  AOI22_X1 U4585 ( .A1(n2975), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4586 ( .A1(n2971), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4587 ( .A1(n2973), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4588 ( .A1(n3624), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4589 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3669)
         );
  AOI22_X1 U4590 ( .A1(n3663), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4591 ( .A1(n3896), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4592 ( .A1(n3907), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4593 ( .A1(n3898), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4594 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3668)
         );
  NOR2_X1 U4595 ( .A1(n3669), .A2(n3668), .ZN(n3673) );
  NAND2_X1 U4596 ( .A1(n6279), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3670)
         );
  NAND2_X1 U4597 ( .A1(n3919), .A2(n3670), .ZN(n3671) );
  AOI21_X1 U4598 ( .B1(n3480), .B2(EAX_REG_18__SCAN_IN), .A(n3671), .ZN(n3672)
         );
  OAI21_X1 U4599 ( .B1(n3922), .B2(n3673), .A(n3672), .ZN(n3676) );
  OAI21_X1 U4600 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3674), .A(n3694), 
        .ZN(n5809) );
  OR2_X1 U4601 ( .A1(n3919), .A2(n5809), .ZN(n3675) );
  AOI22_X1 U4602 ( .A1(n3907), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2975), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4603 ( .A1(n2971), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4604 ( .A1(n2973), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4605 ( .A1(n3879), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4606 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3687)
         );
  AOI22_X1 U4607 ( .A1(n3624), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4608 ( .A1(n3663), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4609 ( .A1(n3903), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4610 ( .A1(n3896), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4611 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  NOR2_X1 U4612 ( .A1(n3687), .A2(n3686), .ZN(n3691) );
  NAND2_X1 U4613 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3688)
         );
  NAND2_X1 U4614 ( .A1(n3919), .A2(n3688), .ZN(n3689) );
  AOI21_X1 U4615 ( .B1(n3480), .B2(EAX_REG_19__SCAN_IN), .A(n3689), .ZN(n3690)
         );
  OAI21_X1 U4616 ( .B1(n3922), .B2(n3691), .A(n3690), .ZN(n3693) );
  XNOR2_X1 U4617 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3694), .ZN(n5663)
         );
  NAND2_X1 U4618 ( .A1(n5663), .A2(n3990), .ZN(n3692) );
  OR2_X1 U4619 ( .A1(n3695), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3696)
         );
  NAND2_X1 U4620 ( .A1(n3696), .A2(n3743), .ZN(n5692) );
  AOI22_X1 U4621 ( .A1(n3663), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4622 ( .A1(n3896), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4623 ( .A1(n2977), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4624 ( .A1(n2973), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4625 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3706)
         );
  AOI22_X1 U4626 ( .A1(n3624), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4627 ( .A1(n3907), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4628 ( .A1(n3905), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4629 ( .A1(n3307), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4630 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3705)
         );
  NOR2_X1 U4631 ( .A1(n3706), .A2(n3705), .ZN(n3707) );
  NOR2_X1 U4632 ( .A1(n3922), .A2(n3707), .ZN(n3711) );
  INV_X1 U4633 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4634 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3708)
         );
  OAI211_X1 U4635 ( .C1(n3833), .C2(n3709), .A(n3919), .B(n3708), .ZN(n3710)
         );
  OAI22_X1 U4636 ( .A1(n5692), .A2(n3919), .B1(n3711), .B2(n3710), .ZN(n5360)
         );
  AOI22_X1 U4637 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n3907), .B1(n2974), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4638 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n3663), .B1(n3903), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4639 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n3307), .B1(n3879), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4640 ( .A1(n3898), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4641 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3722)
         );
  AOI22_X1 U4642 ( .A1(n2971), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4643 ( .A1(n3896), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4644 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n3624), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4645 ( .A1(n2973), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3717) );
  NAND4_X1 U4646 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3721)
         );
  NOR2_X1 U4647 ( .A1(n3722), .A2(n3721), .ZN(n3726) );
  NAND2_X1 U4648 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3723)
         );
  NAND2_X1 U4649 ( .A1(n3919), .A2(n3723), .ZN(n3724) );
  AOI21_X1 U4650 ( .B1(n3480), .B2(EAX_REG_21__SCAN_IN), .A(n3724), .ZN(n3725)
         );
  OAI21_X1 U4651 ( .B1(n3922), .B2(n3726), .A(n3725), .ZN(n3728) );
  XNOR2_X1 U4652 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3743), .ZN(n5639)
         );
  NAND2_X1 U4653 ( .A1(n5639), .A2(n3990), .ZN(n3727) );
  NAND2_X1 U4654 ( .A1(n3728), .A2(n3727), .ZN(n5467) );
  AOI22_X1 U4655 ( .A1(n3907), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4656 ( .A1(n3903), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4657 ( .A1(n3896), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4658 ( .A1(n3753), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4659 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3738)
         );
  AOI22_X1 U4660 ( .A1(n3624), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3898), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4661 ( .A1(n2974), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4662 ( .A1(n3905), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4663 ( .A1(n3663), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4664 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3737)
         );
  NOR2_X1 U4665 ( .A1(n3738), .A2(n3737), .ZN(n3742) );
  NAND2_X1 U4666 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3739)
         );
  NAND2_X1 U4667 ( .A1(n3919), .A2(n3739), .ZN(n3740) );
  AOI21_X1 U4668 ( .B1(n3480), .B2(EAX_REG_22__SCAN_IN), .A(n3740), .ZN(n3741)
         );
  OAI21_X1 U4669 ( .B1(n3922), .B2(n3742), .A(n3741), .ZN(n3747) );
  OAI21_X1 U4670 ( .B1(n3745), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3791), 
        .ZN(n5461) );
  OR2_X1 U4671 ( .A1(n5461), .A2(n3919), .ZN(n3746) );
  NAND2_X1 U4672 ( .A1(n3747), .A2(n3746), .ZN(n5262) );
  AOI22_X1 U4673 ( .A1(n3896), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2975), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4674 ( .A1(n3907), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4675 ( .A1(n2971), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4676 ( .A1(n3663), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4677 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3759)
         );
  AOI22_X1 U4678 ( .A1(n3624), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4679 ( .A1(n3898), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4680 ( .A1(n3897), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4681 ( .A1(n3307), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4682 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4683 ( .A1(n3759), .A2(n3758), .ZN(n3777) );
  AOI22_X1 U4684 ( .A1(n3624), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4685 ( .A1(n3905), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4686 ( .A1(n3663), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4687 ( .A1(n2971), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4688 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4689 ( .A1(n3896), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4690 ( .A1(n3903), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4691 ( .A1(n3907), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4692 ( .A1(n3897), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4693 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  NOR2_X1 U4694 ( .A1(n3769), .A2(n3768), .ZN(n3776) );
  XOR2_X1 U4695 ( .A(n3777), .B(n3776), .Z(n3770) );
  NAND2_X1 U4696 ( .A1(n3890), .A2(n3770), .ZN(n3775) );
  NAND2_X1 U4697 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3771)
         );
  NAND2_X1 U4698 ( .A1(n3919), .A2(n3771), .ZN(n3772) );
  AOI21_X1 U4699 ( .B1(n3480), .B2(EAX_REG_23__SCAN_IN), .A(n3772), .ZN(n3774)
         );
  XNOR2_X1 U4700 ( .A(n3791), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5628)
         );
  AOI21_X1 U4701 ( .B1(n3775), .B2(n3774), .A(n3773), .ZN(n5351) );
  NOR2_X1 U4702 ( .A1(n3777), .A2(n3776), .ZN(n3808) );
  AOI22_X1 U4703 ( .A1(n3896), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4704 ( .A1(n3903), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4705 ( .A1(n3907), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4706 ( .A1(n2976), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4707 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3788)
         );
  AOI22_X1 U4708 ( .A1(n3624), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4709 ( .A1(n3782), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4710 ( .A1(n2966), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4711 ( .A1(n3307), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3783) );
  NAND4_X1 U4712 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3787)
         );
  OR2_X1 U4713 ( .A1(n3788), .A2(n3787), .ZN(n3807) );
  INV_X1 U4714 ( .A(n3807), .ZN(n3789) );
  XNOR2_X1 U4715 ( .A(n3808), .B(n3789), .ZN(n3790) );
  NAND2_X1 U4716 ( .A1(n3790), .A2(n3890), .ZN(n3796) );
  INV_X1 U4717 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5638) );
  XNOR2_X1 U4718 ( .A(n3813), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5445)
         );
  AND2_X1 U4719 ( .A1(n5445), .A2(n3893), .ZN(n3794) );
  INV_X1 U4720 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4314) );
  NOR2_X1 U4721 ( .A1(n3792), .A2(n4314), .ZN(n3793) );
  AOI211_X1 U4722 ( .C1(n3480), .C2(EAX_REG_24__SCAN_IN), .A(n3794), .B(n3793), 
        .ZN(n3795) );
  NAND2_X1 U4723 ( .A1(n3796), .A2(n3795), .ZN(n4320) );
  AOI22_X1 U4724 ( .A1(n3896), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4725 ( .A1(n2971), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4726 ( .A1(n2966), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4727 ( .A1(n2973), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4728 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3806)
         );
  AOI22_X1 U4729 ( .A1(n3907), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2977), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4730 ( .A1(n3903), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4731 ( .A1(n3905), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4732 ( .A1(n3624), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4733 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  NOR2_X1 U4734 ( .A1(n3806), .A2(n3805), .ZN(n3818) );
  NAND2_X1 U4735 ( .A1(n3808), .A2(n3807), .ZN(n3817) );
  XOR2_X1 U4736 ( .A(n3818), .B(n3817), .Z(n3809) );
  NAND2_X1 U4737 ( .A1(n3809), .A2(n3890), .ZN(n3812) );
  INV_X1 U4738 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5434) );
  AOI21_X1 U4739 ( .B1(n5434), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3810) );
  AOI21_X1 U4740 ( .B1(n3480), .B2(EAX_REG_25__SCAN_IN), .A(n3810), .ZN(n3811)
         );
  NAND2_X1 U4741 ( .A1(n3812), .A2(n3811), .ZN(n3815) );
  NAND2_X1 U4742 ( .A1(n3813), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3836)
         );
  XNOR2_X1 U4743 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n3836), .ZN(n5621)
         );
  NAND2_X1 U4744 ( .A1(n5621), .A2(n3990), .ZN(n3814) );
  NAND2_X1 U4745 ( .A1(n3815), .A2(n3814), .ZN(n5341) );
  NOR2_X1 U4746 ( .A1(n3818), .A2(n3817), .ZN(n3842) );
  AOI22_X1 U4747 ( .A1(n3896), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4748 ( .A1(n3903), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4749 ( .A1(n3907), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3819), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4750 ( .A1(n2975), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4751 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4752 ( .A1(n3624), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4753 ( .A1(n3663), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4754 ( .A1(n2966), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4755 ( .A1(n3307), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4756 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  OR2_X1 U4757 ( .A1(n3829), .A2(n3828), .ZN(n3841) );
  INV_X1 U4758 ( .A(n3841), .ZN(n3830) );
  XNOR2_X1 U4759 ( .A(n3842), .B(n3830), .ZN(n3835) );
  INV_X1 U4760 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4761 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3831)
         );
  OAI211_X1 U4762 ( .C1(n3833), .C2(n3832), .A(n3919), .B(n3831), .ZN(n3834)
         );
  AOI21_X1 U4763 ( .B1(n3835), .B2(n3890), .A(n3834), .ZN(n3840) );
  INV_X1 U4764 ( .A(n3836), .ZN(n3837) );
  OAI21_X1 U4765 ( .B1(n3838), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n3857), 
        .ZN(n5619) );
  NOR2_X1 U4766 ( .A1(n5619), .A2(n3919), .ZN(n3839) );
  NAND2_X1 U4767 ( .A1(n3842), .A2(n3841), .ZN(n3860) );
  AOI22_X1 U4768 ( .A1(n3907), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4769 ( .A1(n2966), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4770 ( .A1(n3307), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4771 ( .A1(n3897), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4772 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3852)
         );
  AOI22_X1 U4773 ( .A1(n3896), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4774 ( .A1(n3663), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4775 ( .A1(n2973), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4776 ( .A1(n3624), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4777 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  NOR2_X1 U4778 ( .A1(n3852), .A2(n3851), .ZN(n3861) );
  XOR2_X1 U4779 ( .A(n3860), .B(n3861), .Z(n3853) );
  NAND2_X1 U4780 ( .A1(n3853), .A2(n3890), .ZN(n3856) );
  INV_X1 U4781 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5422) );
  AOI21_X1 U4782 ( .B1(n5422), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3854) );
  AOI21_X1 U4783 ( .B1(n3480), .B2(EAX_REG_27__SCAN_IN), .A(n3854), .ZN(n3855)
         );
  XNOR2_X1 U4784 ( .A(n3857), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5425)
         );
  OR2_X1 U4785 ( .A1(n3858), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U4786 ( .A1(n3924), .A2(n3859), .ZN(n5415) );
  NOR2_X1 U4787 ( .A1(n3861), .A2(n3860), .ZN(n3878) );
  AOI22_X1 U4788 ( .A1(n3896), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4789 ( .A1(n3903), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4790 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n3907), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4791 ( .A1(n2974), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4792 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3872)
         );
  AOI22_X1 U4793 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n3624), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4794 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n3663), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4795 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n3898), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4796 ( .A1(n3307), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4797 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  OR2_X1 U4798 ( .A1(n3872), .A2(n3871), .ZN(n3877) );
  XNOR2_X1 U4799 ( .A(n3878), .B(n3877), .ZN(n3875) );
  AOI21_X1 U4800 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6279), .A(n3893), 
        .ZN(n3874) );
  NAND2_X1 U4801 ( .A1(n3928), .A2(EAX_REG_28__SCAN_IN), .ZN(n3873) );
  OAI211_X1 U4802 ( .C1(n3875), .C2(n3922), .A(n3874), .B(n3873), .ZN(n3876)
         );
  OAI21_X1 U4803 ( .B1(n3919), .B2(n5415), .A(n3876), .ZN(n5239) );
  NAND2_X1 U4804 ( .A1(n3878), .A2(n3877), .ZN(n3914) );
  AOI22_X1 U4805 ( .A1(n3907), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4806 ( .A1(n3663), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4807 ( .A1(n3905), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4808 ( .A1(n2966), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4809 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  AOI22_X1 U4810 ( .A1(n3161), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4811 ( .A1(n3624), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4812 ( .A1(n2974), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4813 ( .A1(n2973), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4814 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  NOR2_X1 U4815 ( .A1(n3889), .A2(n3888), .ZN(n3915) );
  XOR2_X1 U4816 ( .A(n3914), .B(n3915), .Z(n3891) );
  NAND2_X1 U4817 ( .A1(n3891), .A2(n3890), .ZN(n3895) );
  INV_X1 U4818 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5205) );
  NOR2_X1 U4819 ( .A1(n5205), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3892) );
  AOI211_X1 U4820 ( .C1(n3480), .C2(EAX_REG_29__SCAN_IN), .A(n3893), .B(n3892), 
        .ZN(n3894) );
  XNOR2_X1 U4821 ( .A(n3924), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5203)
         );
  AOI22_X1 U4822 ( .A1(n3161), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4823 ( .A1(n3663), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4824 ( .A1(n3307), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4825 ( .A1(n3898), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3753), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4826 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3913)
         );
  AOI22_X1 U4827 ( .A1(n2975), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4828 ( .A1(n3624), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4829 ( .A1(n2973), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3862), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4830 ( .A1(n3907), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3906), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4831 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3912)
         );
  NOR2_X1 U4832 ( .A1(n3913), .A2(n3912), .ZN(n3917) );
  NOR2_X1 U4833 ( .A1(n3915), .A2(n3914), .ZN(n3916) );
  XOR2_X1 U4834 ( .A(n3917), .B(n3916), .Z(n3923) );
  NAND2_X1 U4835 ( .A1(n4986), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3918)
         );
  NAND2_X1 U4836 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  AOI21_X1 U4837 ( .B1(n3928), .B2(EAX_REG_30__SCAN_IN), .A(n3920), .ZN(n3921)
         );
  OAI21_X1 U4838 ( .B1(n3923), .B2(n3922), .A(n3921), .ZN(n3926) );
  XNOR2_X1 U4839 ( .A(n3992), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5227)
         );
  NAND2_X1 U4840 ( .A1(n5227), .A2(n3990), .ZN(n3925) );
  NAND2_X1 U4841 ( .A1(n3926), .A2(n3925), .ZN(n4354) );
  AOI22_X1 U4842 ( .A1(n3928), .A2(EAX_REG_31__SCAN_IN), .B1(n3927), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3929) );
  XNOR2_X1 U4843 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3949) );
  NAND2_X1 U4844 ( .A1(n3951), .A2(n3949), .ZN(n3932) );
  NAND2_X1 U4845 ( .A1(n4595), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4846 ( .A1(n3932), .A2(n3931), .ZN(n3945) );
  XNOR2_X1 U4847 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3943) );
  NAND2_X1 U4848 ( .A1(n3945), .A2(n3943), .ZN(n3934) );
  NAND2_X1 U4849 ( .A1(n6665), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3933) );
  OAI222_X1 U4850 ( .A1(n5774), .A2(n3937), .B1(n5774), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3937), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3977) );
  INV_X1 U4851 ( .A(n3976), .ZN(n3940) );
  NAND2_X1 U4852 ( .A1(n3937), .A2(n5774), .ZN(n3938) );
  INV_X1 U4853 ( .A(n3983), .ZN(n3939) );
  XNOR2_X1 U4854 ( .A(n3942), .B(n3941), .ZN(n3980) );
  INV_X1 U4855 ( .A(n3943), .ZN(n3944) );
  XNOR2_X1 U4856 ( .A(n3945), .B(n3944), .ZN(n3982) );
  INV_X1 U4857 ( .A(n3965), .ZN(n3971) );
  NAND2_X1 U4858 ( .A1(n3946), .A2(n3215), .ZN(n3947) );
  AOI21_X1 U4859 ( .B1(n3976), .B2(n4278), .A(n3222), .ZN(n3962) );
  INV_X1 U4860 ( .A(n3949), .ZN(n3950) );
  XNOR2_X1 U4861 ( .A(n3950), .B(n3951), .ZN(n3981) );
  NAND2_X1 U4862 ( .A1(n3981), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3961) );
  INV_X1 U4863 ( .A(n3951), .ZN(n3953) );
  NAND2_X1 U4864 ( .A1(n3031), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3952) );
  NAND2_X1 U4865 ( .A1(n3953), .A2(n3952), .ZN(n3957) );
  OAI21_X1 U4866 ( .B1(n4255), .B2(n3957), .A(n3954), .ZN(n3955) );
  AOI22_X1 U4867 ( .A1(n3962), .A2(n3961), .B1(n3970), .B2(n3955), .ZN(n3959)
         );
  INV_X1 U4868 ( .A(n3959), .ZN(n3956) );
  AOI21_X1 U4869 ( .B1(n3956), .B2(n3981), .A(n3978), .ZN(n3964) );
  INV_X1 U4870 ( .A(n3957), .ZN(n3958) );
  NAND3_X1 U4871 ( .A1(n3959), .A2(n3958), .A3(n3976), .ZN(n3960) );
  OAI21_X1 U4872 ( .B1(n3962), .B2(n3961), .A(n3960), .ZN(n3963) );
  NOR2_X1 U4873 ( .A1(n3964), .A2(n3963), .ZN(n3969) );
  INV_X1 U4874 ( .A(n3982), .ZN(n3967) );
  INV_X1 U4875 ( .A(n3970), .ZN(n3966) );
  AOI211_X1 U4876 ( .C1(n3973), .C2(n3967), .A(n3966), .B(n3965), .ZN(n3968)
         );
  OAI222_X1 U4877 ( .A1(n3971), .A2(n3970), .B1(n4207), .B2(n3980), .C1(n3969), 
        .C2(n3968), .ZN(n3972) );
  INV_X1 U4878 ( .A(n3977), .ZN(n3985) );
  NAND3_X1 U4879 ( .A1(n3982), .A2(n3981), .A3(n3980), .ZN(n3984) );
  AOI21_X1 U4880 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n6398) );
  NOR2_X1 U4881 ( .A1(n3987), .A2(n3253), .ZN(n3988) );
  NAND2_X1 U4882 ( .A1(n6397), .A2(n6429), .ZN(n3989) );
  NOR2_X1 U4883 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6532) );
  NAND3_X1 U4884 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6532), .ZN(n6423) );
  AND2_X1 U4885 ( .A1(n6419), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U4886 ( .A1(n4330), .A2(n3990), .ZN(n6430) );
  INV_X1 U4887 ( .A(n3992), .ZN(n3993) );
  NAND2_X1 U4888 ( .A1(n3993), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3995)
         );
  INV_X1 U4889 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3994) );
  NOR2_X1 U4890 ( .A1(n4339), .A2(n6418), .ZN(n3996) );
  NAND2_X1 U4891 ( .A1(n5394), .A2(n5879), .ZN(n4140) );
  AND2_X1 U4892 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4011) );
  NAND3_X1 U4893 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4006) );
  INV_X1 U4894 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6487) );
  NAND3_X1 U4895 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4004) );
  OR2_X1 U4896 ( .A1(n3997), .A2(STATE_REG_0__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U4897 ( .A1(n3946), .A2(n6445), .ZN(n4250) );
  INV_X1 U4898 ( .A(READY_N), .ZN(n4249) );
  NAND2_X1 U4899 ( .A1(n4249), .A2(n5784), .ZN(n4133) );
  INV_X1 U4900 ( .A(n4133), .ZN(n3998) );
  AND3_X1 U4901 ( .A1(n4250), .A2(n3253), .A3(n3998), .ZN(n3999) );
  INV_X1 U4902 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6475) );
  INV_X1 U4903 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6471) );
  INV_X1 U4904 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6465) );
  INV_X1 U4905 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6584) );
  INV_X1 U4906 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6461) );
  INV_X1 U4907 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6459) );
  NOR3_X1 U4908 ( .A1(n6584), .A2(n6461), .A3(n6459), .ZN(n5896) );
  NAND2_X1 U4909 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5896), .ZN(n4913) );
  NOR2_X1 U4910 ( .A1(n6465), .A2(n4913), .ZN(n4914) );
  NAND3_X1 U4911 ( .A1(n4914), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n4363) );
  NOR2_X1 U4912 ( .A1(n6471), .A2(n4363), .ZN(n5847) );
  NAND3_X1 U4913 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n5847), .ZN(n5835) );
  NOR2_X1 U4914 ( .A1(n6475), .A2(n5835), .ZN(n5836) );
  NAND2_X1 U4915 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5836), .ZN(n5810) );
  INV_X1 U4916 ( .A(n5810), .ZN(n4000) );
  NAND3_X1 U4917 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n4000), .ZN(n4002) );
  NAND2_X1 U4918 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5656), .ZN(n5654) );
  NOR2_X1 U4919 ( .A1(n6487), .A2(n5654), .ZN(n5649) );
  NAND2_X1 U4920 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5649), .ZN(n5641) );
  NOR2_X1 U4921 ( .A1(n4006), .A2(n5641), .ZN(n4310) );
  AND3_X1 U4922 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4001) );
  AND2_X1 U4923 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4009) );
  NAND2_X1 U4924 ( .A1(n5259), .A2(n4009), .ZN(n5219) );
  NAND3_X1 U4925 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4008) );
  NAND3_X1 U4926 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4005) );
  OAI21_X1 U4927 ( .B1(n5888), .B2(n4002), .A(n5886), .ZN(n5819) );
  INV_X1 U4928 ( .A(n5819), .ZN(n4003) );
  AOI21_X1 U4929 ( .B1(n5886), .B2(n4004), .A(n4003), .ZN(n5804) );
  INV_X1 U4930 ( .A(n5804), .ZN(n5277) );
  AOI21_X1 U4931 ( .B1(n5886), .B2(n4005), .A(n5277), .ZN(n5640) );
  NAND2_X1 U4932 ( .A1(n5886), .A2(n4006), .ZN(n4007) );
  AOI21_X1 U4933 ( .B1(n4008), .B2(n5886), .A(n5622), .ZN(n5615) );
  OAI21_X1 U4934 ( .B1(n4009), .B2(n5826), .A(n5615), .ZN(n5248) );
  INV_X1 U4935 ( .A(n5248), .ZN(n4010) );
  OAI21_X1 U4936 ( .B1(n4011), .B2(n5219), .A(n4010), .ZN(n5232) );
  INV_X1 U4937 ( .A(n4011), .ZN(n4012) );
  INV_X1 U4938 ( .A(n4379), .ZN(n4124) );
  NAND2_X1 U4939 ( .A1(n4278), .A2(n3253), .ZN(n4020) );
  OAI22_X1 U4940 ( .A1(n4124), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4020), .ZN(n4132) );
  AND2_X1 U4941 ( .A1(n4020), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4013)
         );
  AOI21_X1 U4942 ( .B1(n4124), .B2(EBX_REG_30__SCAN_IN), .A(n4013), .ZN(n5221)
         );
  INV_X1 U4943 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U4944 ( .A1(n4119), .A2(n5137), .ZN(n4014) );
  OAI211_X1 U4945 ( .C1(EBX_REG_1__SCAN_IN), .C2(n4020), .A(n4014), .B(n4080), 
        .ZN(n4017) );
  INV_X1 U4946 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U4947 ( .A1(n4266), .A2(n4408), .ZN(n4016) );
  NAND2_X1 U4948 ( .A1(n4017), .A2(n4016), .ZN(n4021) );
  NAND2_X1 U4949 ( .A1(n4119), .A2(EBX_REG_0__SCAN_IN), .ZN(n4019) );
  OAI21_X1 U4950 ( .B1(n4120), .B2(EBX_REG_0__SCAN_IN), .A(n4019), .ZN(n4380)
         );
  XNOR2_X1 U4951 ( .A(n4021), .B(n4380), .ZN(n4407) );
  INV_X1 U4952 ( .A(n4021), .ZN(n4022) );
  NAND2_X1 U4953 ( .A1(n4022), .A2(n4380), .ZN(n4023) );
  NAND2_X1 U4954 ( .A1(n4405), .A2(n4023), .ZN(n4432) );
  INV_X1 U4955 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U4956 ( .B1(n4120), .B2(n6179), .A(n4119), .ZN(n4025) );
  INV_X1 U4957 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4026) );
  NAND2_X1 U4958 ( .A1(n4406), .A2(n4026), .ZN(n4024) );
  NAND2_X1 U4959 ( .A1(n4025), .A2(n4024), .ZN(n4028) );
  NAND2_X1 U4960 ( .A1(n4121), .A2(n4026), .ZN(n4027) );
  AND2_X1 U4961 ( .A1(n4028), .A2(n4027), .ZN(n4431) );
  INV_X1 U4962 ( .A(n4431), .ZN(n4034) );
  INV_X1 U4963 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U4964 ( .A1(n4126), .A2(n4029), .ZN(n4032) );
  INV_X1 U4965 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U4966 ( .A1(n4406), .A2(n4029), .ZN(n4030) );
  OAI211_X1 U4967 ( .C1(n4121), .C2(n6164), .A(n4030), .B(n4119), .ZN(n4031)
         );
  NAND2_X1 U4968 ( .A1(n4032), .A2(n4031), .ZN(n4430) );
  INV_X1 U4969 ( .A(n4430), .ZN(n4033) );
  INV_X1 U4970 ( .A(n4126), .ZN(n4116) );
  MUX2_X1 U4971 ( .A(n4116), .B(n4080), .S(EBX_REG_5__SCAN_IN), .Z(n4037) );
  INV_X1 U4972 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U4973 ( .A1(n4379), .A2(n6136), .ZN(n4036) );
  NAND2_X1 U4974 ( .A1(n4037), .A2(n4036), .ZN(n4504) );
  INV_X1 U4975 ( .A(n4504), .ZN(n4042) );
  INV_X1 U4976 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U4977 ( .A1(n4119), .A2(n6155), .ZN(n4039) );
  INV_X1 U4978 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U4979 ( .A1(n4406), .A2(n5933), .ZN(n4038) );
  NAND3_X1 U4980 ( .A1(n4039), .A2(n4080), .A3(n4038), .ZN(n4041) );
  NAND2_X1 U4981 ( .A1(n4121), .A2(n5933), .ZN(n4040) );
  NAND2_X1 U4982 ( .A1(n4041), .A2(n4040), .ZN(n5884) );
  NAND2_X1 U4983 ( .A1(n4042), .A2(n5884), .ZN(n4043) );
  INV_X1 U4984 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U4985 ( .A1(n4119), .A2(n6650), .ZN(n4045) );
  INV_X1 U4986 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U4987 ( .A1(n4406), .A2(n4046), .ZN(n4044) );
  NAND3_X1 U4988 ( .A1(n4045), .A2(n4080), .A3(n4044), .ZN(n4048) );
  NAND2_X1 U4989 ( .A1(n4121), .A2(n4046), .ZN(n4047) );
  NAND2_X1 U4990 ( .A1(n4048), .A2(n4047), .ZN(n4499) );
  MUX2_X1 U4991 ( .A(n4116), .B(n4080), .S(EBX_REG_7__SCAN_IN), .Z(n4050) );
  INV_X1 U4992 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U4993 ( .A1(n4379), .A2(n6134), .ZN(n4049) );
  NAND2_X1 U4994 ( .A1(n4050), .A2(n4049), .ZN(n4749) );
  INV_X1 U4995 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U4996 ( .A1(n4119), .A2(n6125), .ZN(n4054) );
  INV_X1 U4997 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U4998 ( .A1(n4406), .A2(n4360), .ZN(n4053) );
  NAND3_X1 U4999 ( .A1(n4054), .A2(n4080), .A3(n4053), .ZN(n4056) );
  NAND2_X1 U5000 ( .A1(n4121), .A2(n4360), .ZN(n4055) );
  INV_X1 U5001 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U5002 ( .A1(n4126), .A2(n5929), .ZN(n4059) );
  INV_X1 U5003 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5004 ( .A1(n4406), .A2(n5929), .ZN(n4057) );
  OAI211_X1 U5005 ( .C1(n4120), .C2(n6103), .A(n4057), .B(n4119), .ZN(n4058)
         );
  AND2_X1 U5006 ( .A1(n4059), .A2(n4058), .ZN(n5858) );
  INV_X1 U5007 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U5008 ( .A1(n4126), .A2(n6662), .ZN(n4062) );
  INV_X1 U5009 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U5010 ( .A1(n4406), .A2(n6662), .ZN(n4060) );
  OAI211_X1 U5011 ( .C1(n4120), .C2(n6685), .A(n4060), .B(n4119), .ZN(n4061)
         );
  NAND2_X1 U5012 ( .A1(n4062), .A2(n4061), .ZN(n5831) );
  INV_X1 U5013 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U5014 ( .A1(n4119), .A2(n4218), .ZN(n4063) );
  OAI211_X1 U5015 ( .C1(EBX_REG_10__SCAN_IN), .C2(n4020), .A(n4063), .B(n4080), 
        .ZN(n4065) );
  INV_X1 U5016 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U5017 ( .A1(n4121), .A2(n5037), .ZN(n4064) );
  INV_X1 U5018 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U5019 ( .A1(n4119), .A2(n5108), .ZN(n4068) );
  INV_X1 U5020 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4069) );
  NAND2_X1 U5021 ( .A1(n4406), .A2(n4069), .ZN(n4067) );
  NAND3_X1 U5022 ( .A1(n4068), .A2(n4080), .A3(n4067), .ZN(n4071) );
  NAND2_X1 U5023 ( .A1(n4121), .A2(n4069), .ZN(n4070) );
  INV_X1 U5024 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5025 ( .A1(n4126), .A2(n5921), .ZN(n4074) );
  INV_X1 U5026 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U5027 ( .A1(n4406), .A2(n5921), .ZN(n4072) );
  OAI211_X1 U5028 ( .C1(n4120), .C2(n6618), .A(n4072), .B(n4119), .ZN(n4073)
         );
  INV_X1 U5029 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4226) );
  OAI21_X1 U5030 ( .B1(n4120), .B2(n4226), .A(n4119), .ZN(n4076) );
  INV_X1 U5031 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5032 ( .A1(n4406), .A2(n4077), .ZN(n4075) );
  NAND2_X1 U5033 ( .A1(n4076), .A2(n4075), .ZN(n4079) );
  NAND2_X1 U5034 ( .A1(n4121), .A2(n4077), .ZN(n4078) );
  NAND2_X1 U5035 ( .A1(n4079), .A2(n4078), .ZN(n5125) );
  MUX2_X1 U5036 ( .A(n4116), .B(n4080), .S(EBX_REG_15__SCAN_IN), .Z(n4082) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5038 ( .A1(n4379), .A2(n5756), .ZN(n4081) );
  NAND2_X1 U5039 ( .A1(n4082), .A2(n4081), .ZN(n5130) );
  INV_X1 U5040 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U5041 ( .B1(n4120), .B2(n5693), .A(n4119), .ZN(n4084) );
  INV_X1 U5042 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U5043 ( .A1(n4406), .A2(n5389), .ZN(n4083) );
  AOI22_X1 U5044 ( .A1(n4084), .A2(n4083), .B1(n4121), .B2(n5389), .ZN(n5282)
         );
  INV_X1 U5045 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U5046 ( .A1(n4126), .A2(n5274), .ZN(n4087) );
  INV_X1 U5047 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5738) );
  NAND2_X1 U5048 ( .A1(n4406), .A2(n5274), .ZN(n4085) );
  OAI211_X1 U5049 ( .C1(n4120), .C2(n5738), .A(n4085), .B(n4119), .ZN(n4086)
         );
  NAND2_X1 U5050 ( .A1(n4087), .A2(n4086), .ZN(n5278) );
  NOR2_X4 U5051 ( .A1(n5285), .A2(n5278), .ZN(n5382) );
  INV_X1 U5052 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U5053 ( .A1(n4119), .A2(n5474), .ZN(n4089) );
  INV_X1 U5054 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U5055 ( .A1(n4406), .A2(n5374), .ZN(n4088) );
  NAND3_X1 U5056 ( .A1(n4089), .A2(n4080), .A3(n4088), .ZN(n4091) );
  NAND2_X1 U5057 ( .A1(n4266), .A2(n5374), .ZN(n4090) );
  NAND2_X1 U5058 ( .A1(n4091), .A2(n4090), .ZN(n5371) );
  INV_X1 U5059 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5730) );
  NOR2_X1 U5060 ( .A1(n4020), .A2(EBX_REG_18__SCAN_IN), .ZN(n5368) );
  AOI21_X1 U5061 ( .B1(n4379), .B2(n5730), .A(n5368), .ZN(n5367) );
  OAI22_X1 U5062 ( .A1(n4124), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4020), .ZN(n5362) );
  NAND2_X1 U5063 ( .A1(n5367), .A2(n5362), .ZN(n4093) );
  NAND2_X1 U5064 ( .A1(n4266), .A2(EBX_REG_20__SCAN_IN), .ZN(n4092) );
  OAI211_X1 U5065 ( .C1(n5367), .C2(n4266), .A(n4093), .B(n4092), .ZN(n4094)
         );
  INV_X1 U5066 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U5067 ( .A1(n4126), .A2(n5668), .ZN(n4097) );
  INV_X1 U5068 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U5069 ( .A1(n4406), .A2(n5668), .ZN(n4095) );
  OAI211_X1 U5070 ( .C1(n4121), .C2(n6670), .A(n4095), .B(n4119), .ZN(n4096)
         );
  NAND2_X1 U5071 ( .A1(n4097), .A2(n4096), .ZN(n5572) );
  INV_X1 U5072 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5073 ( .A1(n4119), .A2(n5570), .ZN(n4099) );
  INV_X1 U5074 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U5075 ( .A1(n4406), .A2(n4100), .ZN(n4098) );
  NAND3_X1 U5076 ( .A1(n4099), .A2(n4080), .A3(n4098), .ZN(n4102) );
  NAND2_X1 U5077 ( .A1(n4266), .A2(n4100), .ZN(n4101) );
  NAND2_X1 U5078 ( .A1(n4102), .A2(n4101), .ZN(n5268) );
  MUX2_X1 U5079 ( .A(n4116), .B(n4080), .S(EBX_REG_23__SCAN_IN), .Z(n4104) );
  INV_X1 U5080 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U5081 ( .A1(n4379), .A2(n5559), .ZN(n4103) );
  AND2_X1 U5082 ( .A1(n4104), .A2(n4103), .ZN(n5353) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U5084 ( .A1(n4119), .A2(n5550), .ZN(n4106) );
  INV_X1 U5085 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U5086 ( .A1(n4406), .A2(n6647), .ZN(n4105) );
  NAND3_X1 U5087 ( .A1(n4106), .A2(n4080), .A3(n4105), .ZN(n4108) );
  NAND2_X1 U5088 ( .A1(n4121), .A2(n6647), .ZN(n4107) );
  AND2_X1 U5089 ( .A1(n4108), .A2(n4107), .ZN(n4322) );
  INV_X1 U5090 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U5091 ( .A1(n4126), .A2(n5348), .ZN(n4111) );
  INV_X1 U5092 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5093 ( .A1(n4406), .A2(n5348), .ZN(n4109) );
  OAI211_X1 U5094 ( .C1(n4121), .C2(n5716), .A(n4109), .B(n4119), .ZN(n4110)
         );
  NAND2_X1 U5095 ( .A1(n4111), .A2(n4110), .ZN(n5343) );
  INV_X1 U5096 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U5097 ( .B1(n4120), .B2(n6613), .A(n4119), .ZN(n4113) );
  INV_X1 U5098 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U5099 ( .A1(n4406), .A2(n5340), .ZN(n4112) );
  NAND2_X1 U5100 ( .A1(n4113), .A2(n4112), .ZN(n4115) );
  NAND2_X1 U5101 ( .A1(n4266), .A2(n5340), .ZN(n4114) );
  NAND2_X1 U5102 ( .A1(n4115), .A2(n4114), .ZN(n5337) );
  MUX2_X1 U5103 ( .A(n4116), .B(n4080), .S(EBX_REG_27__SCAN_IN), .Z(n4118) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U5105 ( .A1(n4379), .A2(n5535), .ZN(n4117) );
  AND2_X1 U5106 ( .A1(n4118), .A2(n4117), .ZN(n5252) );
  INV_X1 U5107 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4238) );
  OAI21_X1 U5108 ( .B1(n4120), .B2(n4238), .A(n4119), .ZN(n4123) );
  INV_X1 U5109 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U5110 ( .A1(n4406), .A2(n5332), .ZN(n4122) );
  AOI22_X1 U5111 ( .A1(n4123), .A2(n4122), .B1(n4121), .B2(n5332), .ZN(n5240)
         );
  NOR2_X1 U5112 ( .A1(n4124), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4130)
         );
  INV_X1 U5113 ( .A(n4130), .ZN(n4125) );
  INV_X1 U5114 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5216) );
  MUX2_X1 U5115 ( .A(n4125), .B(n5216), .S(n4121), .Z(n4128) );
  NAND2_X1 U5116 ( .A1(n4126), .A2(n5216), .ZN(n4127) );
  NAND2_X1 U5117 ( .A1(n4128), .A2(n4127), .ZN(n5200) );
  NOR2_X1 U5118 ( .A1(n5242), .A2(n5200), .ZN(n5202) );
  NOR2_X1 U5119 ( .A1(n5224), .A2(n4266), .ZN(n5226) );
  NAND2_X1 U5120 ( .A1(n3253), .A2(n4133), .ZN(n4312) );
  NAND2_X1 U5121 ( .A1(n4278), .A2(EBX_REG_31__SCAN_IN), .ZN(n4134) );
  NOR2_X1 U5122 ( .A1(n4312), .A2(n4134), .ZN(n4135) );
  NOR2_X2 U5123 ( .A1(n5888), .A2(n6514), .ZN(n5905) );
  NAND2_X1 U5124 ( .A1(n5905), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4138)
         );
  INV_X1 U5125 ( .A(n6445), .ZN(n4659) );
  NAND3_X1 U5126 ( .A1(n4659), .A2(n4249), .A3(n5784), .ZN(n6411) );
  NAND4_X1 U5127 ( .A1(n5028), .A2(n4136), .A3(EBX_REG_31__SCAN_IN), .A4(n6411), .ZN(n4137) );
  NAND2_X1 U5128 ( .A1(n4140), .A2(n4139), .ZN(U2796) );
  NAND2_X1 U5129 ( .A1(n2978), .A2(n4187), .ZN(n4147) );
  NAND2_X1 U5130 ( .A1(n4141), .A2(n4148), .ZN(n4165) );
  OAI21_X1 U5131 ( .B1(n4148), .B2(n4141), .A(n4165), .ZN(n4144) );
  INV_X1 U5132 ( .A(n4142), .ZN(n4143) );
  OAI211_X1 U5133 ( .C1(n4144), .C2(n6531), .A(n4143), .B(n3215), .ZN(n4145)
         );
  INV_X1 U5134 ( .A(n4145), .ZN(n4146) );
  NAND2_X1 U5135 ( .A1(n4147), .A2(n4146), .ZN(n4532) );
  NAND2_X1 U5136 ( .A1(n4568), .A2(n3256), .ZN(n4156) );
  OAI21_X1 U5137 ( .B1(n6531), .B2(n4148), .A(n4156), .ZN(n4149) );
  INV_X1 U5138 ( .A(n4149), .ZN(n4150) );
  OAI21_X1 U5139 ( .B1(n4824), .B2(n4207), .A(n4150), .ZN(n4376) );
  NAND2_X1 U5140 ( .A1(n4376), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4151)
         );
  NAND2_X1 U5141 ( .A1(n4151), .A2(n5137), .ZN(n4153) );
  AND2_X1 U5142 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4152) );
  NAND2_X1 U5143 ( .A1(n4376), .A2(n4152), .ZN(n4154) );
  AND2_X1 U5144 ( .A1(n4153), .A2(n4154), .ZN(n4533) );
  INV_X1 U5145 ( .A(n4154), .ZN(n4155) );
  XNOR2_X1 U5146 ( .A(n4165), .B(n4164), .ZN(n4158) );
  INV_X1 U5147 ( .A(n4156), .ZN(n4157) );
  AOI21_X1 U5148 ( .B1(n4158), .B2(n4136), .A(n4157), .ZN(n4159) );
  NAND2_X1 U5149 ( .A1(n6082), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4160)
         );
  NAND2_X1 U5150 ( .A1(n6083), .A2(n4160), .ZN(n4163) );
  INV_X1 U5151 ( .A(n6082), .ZN(n4161) );
  NAND2_X1 U5152 ( .A1(n4161), .A2(n6179), .ZN(n4162) );
  AND2_X2 U5153 ( .A1(n4163), .A2(n4162), .ZN(n4665) );
  NAND2_X1 U5154 ( .A1(n4165), .A2(n4164), .ZN(n4172) );
  XNOR2_X1 U5155 ( .A(n4172), .B(n4171), .ZN(n4166) );
  NAND2_X1 U5156 ( .A1(n4168), .A2(n4167), .ZN(n4169) );
  XNOR2_X1 U5157 ( .A(n4169), .B(n6164), .ZN(n4666) );
  NAND2_X1 U5158 ( .A1(n4665), .A2(n4666), .ZN(n4664) );
  NAND2_X1 U5159 ( .A1(n4169), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4170)
         );
  NAND2_X1 U5160 ( .A1(n4664), .A2(n4170), .ZN(n6071) );
  NAND2_X1 U5161 ( .A1(n4172), .A2(n4171), .ZN(n4191) );
  XNOR2_X1 U5162 ( .A(n4191), .B(n4189), .ZN(n4173) );
  NAND2_X1 U5163 ( .A1(n4173), .A2(n4136), .ZN(n4174) );
  OAI21_X2 U5164 ( .B1(n4175), .B2(n4207), .A(n4174), .ZN(n4176) );
  XNOR2_X1 U5165 ( .A(n4176), .B(n6155), .ZN(n6072) );
  NAND2_X1 U5166 ( .A1(n6071), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U5167 ( .A1(n4176), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4177)
         );
  NAND2_X1 U5168 ( .A1(n6074), .A2(n4177), .ZN(n4562) );
  NAND2_X1 U5169 ( .A1(n4178), .A2(n4187), .ZN(n4183) );
  INV_X1 U5170 ( .A(n4191), .ZN(n4179) );
  NAND2_X1 U5171 ( .A1(n4179), .A2(n4189), .ZN(n4180) );
  XNOR2_X1 U5172 ( .A(n4180), .B(n4188), .ZN(n4181) );
  NAND2_X1 U5173 ( .A1(n4181), .A2(n4136), .ZN(n4182) );
  NAND2_X1 U5174 ( .A1(n4183), .A2(n4182), .ZN(n4184) );
  XNOR2_X1 U5175 ( .A(n4184), .B(n6136), .ZN(n4561) );
  NAND2_X1 U5176 ( .A1(n4562), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U5177 ( .A1(n4184), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4185)
         );
  NAND2_X1 U5178 ( .A1(n4560), .A2(n4185), .ZN(n4811) );
  NAND2_X1 U5179 ( .A1(n4186), .A2(n4187), .ZN(n4194) );
  NAND2_X1 U5180 ( .A1(n4189), .A2(n4188), .ZN(n4190) );
  OR2_X1 U5181 ( .A1(n4191), .A2(n4190), .ZN(n4198) );
  XNOR2_X1 U5182 ( .A(n4198), .B(n4199), .ZN(n4192) );
  NAND2_X1 U5183 ( .A1(n4192), .A2(n4136), .ZN(n4193) );
  NAND2_X1 U5184 ( .A1(n4194), .A2(n4193), .ZN(n4195) );
  XNOR2_X1 U5185 ( .A(n4195), .B(n6650), .ZN(n4810) );
  NAND2_X1 U5186 ( .A1(n4811), .A2(n4810), .ZN(n4813) );
  NAND2_X1 U5187 ( .A1(n4195), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4196)
         );
  NAND2_X1 U5188 ( .A1(n4813), .A2(n4196), .ZN(n4895) );
  OR2_X1 U5189 ( .A1(n4197), .A2(n4207), .ZN(n4203) );
  INV_X1 U5190 ( .A(n4198), .ZN(n4200) );
  NAND2_X1 U5191 ( .A1(n4200), .A2(n4199), .ZN(n4210) );
  XNOR2_X1 U5192 ( .A(n4210), .B(n4211), .ZN(n4201) );
  NAND2_X1 U5193 ( .A1(n4201), .A2(n4136), .ZN(n4202) );
  NAND2_X1 U5194 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  XNOR2_X1 U5195 ( .A(n4204), .B(n6134), .ZN(n4894) );
  NAND2_X1 U5196 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  NAND2_X1 U5197 ( .A1(n4204), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4205)
         );
  NAND2_X1 U5198 ( .A1(n4893), .A2(n4205), .ZN(n5017) );
  NOR2_X1 U5199 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  INV_X1 U5200 ( .A(n4210), .ZN(n4212) );
  NAND3_X1 U5201 ( .A1(n4212), .A2(n4136), .A3(n4211), .ZN(n4213) );
  NAND2_X1 U5202 ( .A1(n2967), .A2(n4213), .ZN(n4214) );
  XNOR2_X1 U5203 ( .A(n4214), .B(n6125), .ZN(n5016) );
  NAND2_X1 U5204 ( .A1(n5017), .A2(n5016), .ZN(n5015) );
  NAND2_X1 U5205 ( .A1(n4214), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4215)
         );
  NAND2_X1 U5206 ( .A1(n2967), .A2(n6103), .ZN(n4216) );
  OR2_X1 U5207 ( .A1(n2967), .A2(n6103), .ZN(n4217) );
  NAND2_X1 U5208 ( .A1(n2967), .A2(n4218), .ZN(n5075) );
  AND2_X1 U5209 ( .A1(n2967), .A2(n6685), .ZN(n4223) );
  OR2_X1 U5210 ( .A1(n2967), .A2(n4218), .ZN(n6054) );
  NOR2_X1 U5211 ( .A1(n2967), .A2(n5108), .ZN(n5093) );
  NAND2_X1 U5212 ( .A1(n2967), .A2(n5108), .ZN(n5091) );
  XNOR2_X1 U5213 ( .A(n2967), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5707)
         );
  NAND2_X1 U5214 ( .A1(n2967), .A2(n6618), .ZN(n4224) );
  AND2_X1 U5215 ( .A1(n2967), .A2(n4226), .ZN(n4228) );
  NOR2_X1 U5216 ( .A1(n2967), .A2(n5756), .ZN(n4230) );
  NAND2_X1 U5217 ( .A1(n2967), .A2(n5756), .ZN(n4229) );
  AND2_X1 U5218 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U5219 ( .A1(n5583), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4231) );
  AND2_X1 U5220 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5451) );
  AND2_X1 U5221 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4299) );
  AND2_X1 U5222 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5450) );
  NAND3_X1 U5223 ( .A1(n5451), .A2(n4299), .A3(n5450), .ZN(n4232) );
  NAND2_X1 U5224 ( .A1(n2967), .A2(n4232), .ZN(n4233) );
  NAND2_X1 U5225 ( .A1(n5472), .A2(n4233), .ZN(n4236) );
  NOR2_X1 U5226 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U5227 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5548) );
  NAND4_X1 U5228 ( .A1(n5719), .A2(n5548), .A3(n6670), .A4(n5570), .ZN(n4234)
         );
  NAND2_X1 U5229 ( .A1(n4219), .A2(n4234), .ZN(n4235) );
  XOR2_X1 U5230 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n2967), .Z(n5432) );
  NAND2_X1 U5231 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5519) );
  INV_X1 U5232 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5511) );
  INV_X1 U5233 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4285) );
  NOR2_X1 U5234 ( .A1(n5511), .A2(n4285), .ZN(n4237) );
  NAND2_X1 U5235 ( .A1(n4351), .A2(n4237), .ZN(n4239) );
  NAND2_X1 U5236 ( .A1(n5535), .A2(n4238), .ZN(n5520) );
  INV_X1 U5237 ( .A(n5139), .ZN(n4464) );
  NAND2_X1 U5238 ( .A1(n4464), .A2(n4278), .ZN(n4244) );
  NAND2_X1 U5239 ( .A1(n5139), .A2(n4568), .ZN(n4241) );
  NAND3_X1 U5240 ( .A1(n4257), .A2(n4269), .A3(n4242), .ZN(n4243) );
  INV_X1 U5241 ( .A(n6397), .ZN(n5777) );
  NAND2_X1 U5242 ( .A1(n4243), .A2(n5777), .ZN(n4280) );
  OAI21_X1 U5243 ( .B1(n6414), .B2(n4244), .A(n4280), .ZN(n4457) );
  NAND2_X1 U5244 ( .A1(n4278), .A2(n6445), .ZN(n4245) );
  NOR2_X1 U5245 ( .A1(n6398), .A2(READY_N), .ZN(n4410) );
  AND3_X1 U5246 ( .A1(n4245), .A2(n4410), .A3(n4265), .ZN(n4246) );
  OR2_X1 U5247 ( .A1(n4457), .A2(n4246), .ZN(n4247) );
  NAND2_X1 U5248 ( .A1(n4247), .A2(n6429), .ZN(n4254) );
  NAND2_X1 U5249 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  OAI211_X1 U5250 ( .C1(n4451), .C2(n4251), .A(n3253), .B(n5210), .ZN(n4252)
         );
  NAND3_X1 U5251 ( .A1(n4657), .A2(n3220), .A3(n4252), .ZN(n4253) );
  INV_X1 U5252 ( .A(n4331), .ZN(n6406) );
  INV_X1 U5253 ( .A(n4409), .ZN(n6395) );
  OAI211_X1 U5254 ( .C1(n3247), .C2(n4258), .A(n4454), .B(n5770), .ZN(n4259)
         );
  INV_X1 U5255 ( .A(n4259), .ZN(n4260) );
  NAND3_X1 U5256 ( .A1(n6406), .A2(n6395), .A3(n4260), .ZN(n4261) );
  OAI21_X1 U5257 ( .B1(n4258), .B2(n4399), .A(n6412), .ZN(n4262) );
  INV_X1 U5258 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6509) );
  OR2_X1 U5259 ( .A1(n6092), .A2(n6509), .ZN(n4338) );
  OAI21_X1 U5260 ( .B1(n5331), .B2(n6094), .A(n4338), .ZN(n4308) );
  NAND4_X1 U5261 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U5262 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4263) );
  OR2_X1 U5263 ( .A1(n6138), .A2(n4263), .ZN(n5102) );
  NOR2_X1 U5264 ( .A1(n6134), .A2(n6125), .ZN(n6121) );
  NAND3_X1 U5265 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6121), .ZN(n5107) );
  NOR2_X1 U5266 ( .A1(n5102), .A2(n5107), .ZN(n5099) );
  NAND2_X1 U5267 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U5268 ( .A1(n6618), .A2(n5592), .ZN(n5599) );
  NAND2_X1 U5269 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5599), .ZN(n5747) );
  NAND2_X1 U5270 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5748) );
  NOR2_X1 U5271 ( .A1(n5747), .A2(n5748), .ZN(n4281) );
  NAND2_X1 U5272 ( .A1(n5099), .A2(n4281), .ZN(n4290) );
  NAND2_X1 U5273 ( .A1(n4568), .A2(n4278), .ZN(n5029) );
  OR2_X1 U5274 ( .A1(n5029), .A2(n4265), .ZN(n4455) );
  NAND2_X1 U5275 ( .A1(n4379), .A2(n4455), .ZN(n4264) );
  NAND2_X1 U5276 ( .A1(n4264), .A2(n4142), .ZN(n4270) );
  NAND2_X1 U5277 ( .A1(n5210), .A2(n4265), .ZN(n4268) );
  NAND2_X1 U5278 ( .A1(n3255), .A2(n4266), .ZN(n4267) );
  AND4_X1 U5279 ( .A1(n4270), .A2(n4269), .A3(n4268), .A4(n4267), .ZN(n4271)
         );
  NAND2_X1 U5280 ( .A1(n4272), .A2(n4271), .ZN(n4441) );
  OR2_X1 U5281 ( .A1(n4273), .A2(n3253), .ZN(n4274) );
  NOR2_X1 U5282 ( .A1(n5139), .A2(n4274), .ZN(n4786) );
  OAI22_X1 U5283 ( .A1(n4275), .A2(n3179), .B1(n4438), .B2(n3253), .ZN(n4276)
         );
  NAND2_X1 U5284 ( .A1(n4291), .A2(n4277), .ZN(n4377) );
  INV_X1 U5285 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5189) );
  NOR2_X1 U5286 ( .A1(n4377), .A2(n5189), .ZN(n5097) );
  NOR2_X1 U5287 ( .A1(n5139), .A2(n4568), .ZN(n4279) );
  NAND2_X1 U5288 ( .A1(n4280), .A2(n4279), .ZN(n4435) );
  INV_X1 U5289 ( .A(n4435), .ZN(n6399) );
  AOI21_X1 U5290 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6166) );
  NAND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6151) );
  NOR2_X1 U5292 ( .A1(n6166), .A2(n6151), .ZN(n6140) );
  NAND3_X1 U5293 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6140), .ZN(n6102) );
  NOR2_X1 U5294 ( .A1(n5107), .A2(n6102), .ZN(n5096) );
  NAND2_X1 U5295 ( .A1(n4281), .A2(n5096), .ZN(n4289) );
  NAND2_X1 U5296 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5720) );
  INV_X1 U5297 ( .A(n5720), .ZN(n4283) );
  AND2_X1 U5298 ( .A1(n5583), .A2(n4283), .ZN(n4296) );
  NAND2_X1 U5299 ( .A1(n5739), .A2(n4296), .ZN(n4287) );
  INV_X1 U5300 ( .A(n5451), .ZN(n4288) );
  NOR2_X1 U5301 ( .A1(n4287), .A2(n4288), .ZN(n5560) );
  NAND2_X1 U5302 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5540) );
  INV_X1 U5303 ( .A(n5540), .ZN(n4284) );
  NAND2_X1 U5304 ( .A1(n5710), .A2(n4284), .ZN(n5529) );
  NOR3_X1 U5305 ( .A1(n5519), .A2(n5511), .A3(n4285), .ZN(n4304) );
  INV_X1 U5306 ( .A(n4304), .ZN(n4286) );
  NOR3_X1 U5307 ( .A1(n5529), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4286), 
        .ZN(n4307) );
  NAND2_X1 U5308 ( .A1(n5594), .A2(n4377), .ZN(n5103) );
  INV_X1 U5309 ( .A(n4287), .ZN(n5580) );
  NAND2_X1 U5310 ( .A1(n5580), .A2(n4288), .ZN(n5564) );
  AOI22_X1 U5311 ( .A1(n5103), .A2(n4290), .B1(n4289), .B2(n6172), .ZN(n4295)
         );
  OR2_X1 U5312 ( .A1(n4377), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4293)
         );
  INV_X1 U5313 ( .A(n4291), .ZN(n4292) );
  NAND2_X1 U5314 ( .A1(n4292), .A2(n6092), .ZN(n4671) );
  NAND2_X1 U5315 ( .A1(n4293), .A2(n4671), .ZN(n5101) );
  INV_X1 U5316 ( .A(n5101), .ZN(n4294) );
  INV_X1 U5317 ( .A(n4296), .ZN(n4297) );
  NAND2_X1 U5318 ( .A1(n5586), .A2(n4297), .ZN(n4298) );
  AND2_X1 U5319 ( .A1(n5735), .A2(n4298), .ZN(n5578) );
  INV_X1 U5320 ( .A(n4299), .ZN(n4300) );
  OAI21_X1 U5321 ( .B1(n4301), .B2(n6172), .A(n4300), .ZN(n4302) );
  NAND2_X1 U5322 ( .A1(n5586), .A2(n5540), .ZN(n4303) );
  OAI21_X1 U5323 ( .B1(n6106), .B2(n4304), .A(n5532), .ZN(n4305) );
  OAI21_X1 U5324 ( .B1(n4341), .B2(n6095), .A(n4309), .ZN(U2987) );
  INV_X1 U5325 ( .A(n4310), .ZN(n5612) );
  NOR2_X1 U5326 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5612), .ZN(n5623) );
  INV_X1 U5327 ( .A(n5623), .ZN(n4329) );
  NAND2_X1 U5328 ( .A1(n4136), .A2(n6411), .ZN(n4311) );
  OAI21_X1 U5329 ( .B1(EBX_REG_31__SCAN_IN), .B2(n4312), .A(n4311), .ZN(n4313)
         );
  AND2_X2 U5330 ( .A1(n5028), .A2(n4313), .ZN(n5903) );
  OAI22_X1 U5331 ( .A1(n6647), .A2(n5864), .B1(n4314), .B2(n5889), .ZN(n4315)
         );
  INV_X1 U5332 ( .A(n4315), .ZN(n4328) );
  INV_X1 U5333 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U5334 ( .A1(n4339), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4316) );
  OAI22_X1 U5335 ( .A1(n5633), .A2(n6494), .B1(n5445), .B2(n5883), .ZN(n4317)
         );
  INV_X1 U5336 ( .A(n4317), .ZN(n4327) );
  OR2_X1 U5337 ( .A1(n4319), .A2(n4320), .ZN(n4321) );
  AND2_X1 U5338 ( .A1(n4318), .A2(n4321), .ZN(n5447) );
  NAND2_X1 U5339 ( .A1(n5356), .A2(n4322), .ZN(n4323) );
  AND2_X1 U5340 ( .A1(n5344), .A2(n4323), .ZN(n5553) );
  INV_X1 U5341 ( .A(n5553), .ZN(n4324) );
  OAI22_X1 U5342 ( .A1(n5404), .A2(n5659), .B1(n4324), .B2(n5874), .ZN(n4325)
         );
  INV_X1 U5343 ( .A(n4325), .ZN(n4326) );
  NAND4_X1 U5344 ( .A1(n4329), .A2(n4328), .A3(n4327), .A4(n4326), .ZN(U2803)
         );
  NAND2_X1 U5345 ( .A1(n4330), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6435) );
  NAND2_X2 U5346 ( .A1(n4986), .A2(n6514), .ZN(n6318) );
  NAND2_X1 U5347 ( .A1(n6526), .A2(n6318), .ZN(n4332) );
  NAND2_X1 U5348 ( .A1(n4332), .A2(n6419), .ZN(n4333) );
  NAND2_X1 U5349 ( .A1(n6419), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4335) );
  NAND2_X1 U5350 ( .A1(n5784), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4334) );
  AND2_X1 U5351 ( .A1(n4335), .A2(n4334), .ZN(n4385) );
  INV_X1 U5352 ( .A(n4385), .ZN(n4336) );
  NAND2_X1 U5353 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4337)
         );
  OAI211_X1 U5354 ( .C1(n6090), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4340)
         );
  AOI21_X1 U5355 ( .B1(n5394), .B2(n6075), .A(n4340), .ZN(n4342) );
  INV_X2 U5356 ( .A(n6092), .ZN(n6171) );
  NAND2_X1 U5357 ( .A1(n6171), .A2(REIP_REG_29__SCAN_IN), .ZN(n5512) );
  OAI21_X1 U5358 ( .B1(n5483), .B2(n5205), .A(n5512), .ZN(n4346) );
  AOI21_X1 U5359 ( .B1(n6059), .B2(n5203), .A(n4346), .ZN(n4350) );
  NOR2_X1 U5360 ( .A1(n5409), .A2(n4347), .ZN(n4352) );
  NOR2_X1 U5361 ( .A1(n4351), .A2(n4352), .ZN(n4348) );
  XNOR2_X1 U5362 ( .A(n4348), .B(n5511), .ZN(n5518) );
  NAND3_X1 U5363 ( .A1(n2985), .A2(n4350), .A3(n4349), .ZN(U2957) );
  MUX2_X1 U5364 ( .A(n4352), .B(n4351), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n4353) );
  XNOR2_X1 U5365 ( .A(n4353), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5510)
         );
  INV_X1 U5366 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U5367 ( .A1(n6171), .A2(REIP_REG_30__SCAN_IN), .ZN(n5503) );
  OAI21_X1 U5368 ( .B1(n5483), .B2(n4356), .A(n5503), .ZN(n4357) );
  AOI21_X1 U5369 ( .B1(n6059), .B2(n5227), .A(n4357), .ZN(n4358) );
  OAI211_X1 U5370 ( .C1(n5510), .C2(n6065), .A(n3105), .B(n4358), .ZN(U2956)
         );
  OAI21_X1 U5371 ( .B1(n5826), .B2(n5847), .A(n5064), .ZN(n5866) );
  AOI22_X1 U5372 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5905), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5866), .ZN(n4359) );
  NOR2_X1 U5373 ( .A1(n6318), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U5374 ( .A1(n5064), .A2(n4374), .ZN(n5301) );
  OAI211_X1 U5375 ( .C1(n5864), .C2(n4360), .A(n4359), .B(n5301), .ZN(n4369)
         );
  OAI21_X1 U5376 ( .B1(n2992), .B2(n4362), .A(n4361), .ZN(n5018) );
  NOR2_X1 U5377 ( .A1(n5018), .A2(n5659), .ZN(n4368) );
  NOR3_X1 U5378 ( .A1(n5826), .A2(n5847), .A3(n4363), .ZN(n4367) );
  AOI21_X1 U5379 ( .B1(n4364), .B2(n4746), .A(n5859), .ZN(n6120) );
  INV_X1 U5380 ( .A(n6120), .ZN(n4365) );
  OAI22_X1 U5381 ( .A1(n5020), .A2(n5883), .B1(n5874), .B2(n4365), .ZN(n4366)
         );
  OR4_X1 U5382 ( .A1(n4369), .A2(n4368), .A3(n4367), .A4(n4366), .ZN(U2819) );
  INV_X1 U5383 ( .A(n4370), .ZN(n4373) );
  INV_X1 U5384 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4372) );
  INV_X1 U5385 ( .A(n4374), .ZN(n4371) );
  OAI211_X1 U5386 ( .C1(n4373), .C2(n4372), .A(n5969), .B(n4371), .ZN(U2788)
         );
  NAND2_X1 U5387 ( .A1(n6531), .A2(n5029), .ZN(n5785) );
  OAI21_X1 U5388 ( .B1(n4374), .B2(READREQUEST_REG_SCAN_IN), .A(n6525), .ZN(
        n4375) );
  OAI21_X1 U5389 ( .B1(n6525), .B2(n5785), .A(n4375), .ZN(U3474) );
  XNOR2_X1 U5390 ( .A(n4376), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4392)
         );
  NAND2_X1 U5391 ( .A1(n5585), .A2(n4377), .ZN(n5591) );
  AOI21_X1 U5392 ( .B1(n5594), .B2(n4671), .A(n5189), .ZN(n4378) );
  AOI21_X1 U5393 ( .B1(n5189), .B2(n5591), .A(n4378), .ZN(n4384) );
  NAND2_X1 U5394 ( .A1(n4379), .A2(n5189), .ZN(n4381) );
  AND2_X1 U5395 ( .A1(n4381), .A2(n4380), .ZN(n5325) );
  INV_X1 U5396 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4382) );
  NOR2_X1 U5397 ( .A1(n6092), .A2(n4382), .ZN(n4389) );
  AOI21_X1 U5398 ( .B1(n6169), .B2(n5325), .A(n4389), .ZN(n4383) );
  OAI211_X1 U5399 ( .C1(n4392), .C2(n6095), .A(n4384), .B(n4383), .ZN(U3018)
         );
  NAND2_X1 U5400 ( .A1(n4385), .A2(n5483), .ZN(n4390) );
  XNOR2_X1 U5401 ( .A(n4387), .B(n4386), .ZN(n5329) );
  NOR2_X1 U5402 ( .A1(n5329), .A2(n6063), .ZN(n4388) );
  AOI211_X1 U5403 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4390), .A(n4389), 
        .B(n4388), .ZN(n4391) );
  OAI21_X1 U5404 ( .B1(n4392), .B2(n6065), .A(n4391), .ZN(U2986) );
  INV_X1 U5405 ( .A(n4393), .ZN(n4396) );
  INV_X1 U5406 ( .A(n4394), .ZN(n4395) );
  NAND2_X1 U5407 ( .A1(n4396), .A2(n4395), .ZN(n4397) );
  NAND2_X1 U5408 ( .A1(n4425), .A2(n4397), .ZN(n5320) );
  INV_X1 U5409 ( .A(n4398), .ZN(n4400) );
  NOR2_X1 U5410 ( .A1(n5211), .A2(n4399), .ZN(n4414) );
  NAND4_X1 U5411 ( .A1(n4401), .A2(n4400), .A3(n4406), .A4(n4414), .ZN(n4402)
         );
  OAI21_X1 U5412 ( .B1(n6414), .B2(n4435), .A(n4402), .ZN(n4403) );
  INV_X2 U5413 ( .A(n5931), .ZN(n5390) );
  OAI21_X1 U5414 ( .B1(n4407), .B2(n4406), .A(n4405), .ZN(n5317) );
  INV_X1 U5415 ( .A(n5317), .ZN(n4673) );
  OAI222_X1 U5416 ( .A1(n5320), .A2(n5390), .B1(n4408), .B2(n5934), .C1(n5925), 
        .C2(n4673), .ZN(U2858) );
  NAND2_X1 U5417 ( .A1(n6414), .A2(n4409), .ZN(n4413) );
  INV_X1 U5418 ( .A(n4410), .ZN(n4411) );
  NAND2_X1 U5419 ( .A1(n4414), .A2(n3237), .ZN(n4415) );
  NOR2_X1 U5420 ( .A1(n4275), .A2(n4415), .ZN(n4416) );
  NOR2_X1 U5421 ( .A1(n4454), .A2(READY_N), .ZN(n4417) );
  NAND2_X1 U5422 ( .A1(n3217), .A2(n5211), .ZN(n4419) );
  INV_X1 U5423 ( .A(n4419), .ZN(n4420) );
  AOI22_X1 U5424 ( .A1(n5134), .A2(DATAI_1_), .B1(n5944), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4421) );
  OAI21_X1 U5425 ( .B1(n5669), .B2(n5320), .A(n4421), .ZN(U2890) );
  NAND3_X1 U5426 ( .A1(n4425), .A2(n4424), .A3(n4423), .ZN(n4426) );
  NAND2_X1 U5427 ( .A1(n4422), .A2(n4426), .ZN(n6081) );
  XOR2_X1 U5428 ( .A(n4431), .B(n4432), .Z(n6170) );
  AOI22_X1 U5429 ( .A1(n5930), .A2(n6170), .B1(EBX_REG_2__SCAN_IN), .B2(n5386), 
        .ZN(n4427) );
  OAI21_X1 U5430 ( .B1(n5390), .B2(n6081), .A(n4427), .ZN(U2857) );
  AOI21_X1 U5431 ( .B1(n4429), .B2(n4422), .A(n4428), .ZN(n4668) );
  INV_X1 U5432 ( .A(n4668), .ZN(n5909) );
  OAI21_X1 U5433 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(n4433) );
  AND2_X1 U5434 ( .A1(n4433), .A2(n5885), .ZN(n6157) );
  AOI22_X1 U5435 ( .A1(n5930), .A2(n6157), .B1(EBX_REG_3__SCAN_IN), .B2(n5386), 
        .ZN(n4434) );
  OAI21_X1 U5436 ( .B1(n5909), .B2(n5390), .A(n4434), .ZN(U2856) );
  NAND2_X1 U5437 ( .A1(n4435), .A2(n6395), .ZN(n4794) );
  INV_X1 U5438 ( .A(n4794), .ZN(n4449) );
  INV_X1 U5439 ( .A(n4436), .ZN(n5191) );
  NAND2_X1 U5440 ( .A1(n5191), .A2(n3110), .ZN(n4785) );
  XNOR2_X1 U5441 ( .A(n4785), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4448)
         );
  INV_X1 U5442 ( .A(n5770), .ZN(n4440) );
  NAND3_X1 U5443 ( .A1(n4451), .A2(n4275), .A3(n4438), .ZN(n4439) );
  OR3_X1 U5444 ( .A1(n4441), .A2(n4440), .A3(n4439), .ZN(n4790) );
  NAND2_X1 U5445 ( .A1(n4437), .A2(n4790), .ZN(n4447) );
  XNOR2_X1 U5446 ( .A(n4442), .B(n4461), .ZN(n4445) );
  AOI21_X1 U5447 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n5191), .A(n4443), 
        .ZN(n4444) );
  NAND2_X1 U5448 ( .A1(n3140), .A2(n4444), .ZN(n4450) );
  AOI22_X1 U5449 ( .A1(n5141), .A2(n4445), .B1(n4786), .B2(n4450), .ZN(n4446)
         );
  OAI211_X1 U5450 ( .C1(n4449), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4796)
         );
  AOI22_X1 U5451 ( .A1(n4796), .A2(n5194), .B1(n4450), .B2(n5186), .ZN(n4460)
         );
  OAI21_X1 U5452 ( .B1(n5141), .B2(n3235), .A(n4659), .ZN(n4453) );
  INV_X1 U5453 ( .A(n6414), .ZN(n4452) );
  AOI211_X1 U5454 ( .C1(n4454), .C2(n4453), .A(READY_N), .B(n4452), .ZN(n4459)
         );
  INV_X1 U5455 ( .A(n4455), .ZN(n4458) );
  NOR4_X1 U5456 ( .A1(n4459), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(n4795)
         );
  INV_X1 U5457 ( .A(n4795), .ZN(n6382) );
  NAND2_X1 U5458 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4822) );
  NOR2_X1 U5459 ( .A1(n6419), .A2(n4822), .ZN(n6433) );
  AOI22_X1 U5460 ( .A1(n6382), .A2(n6429), .B1(FLUSH_REG_SCAN_IN), .B2(n6433), 
        .ZN(n5772) );
  NAND2_X1 U5461 ( .A1(n6419), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U5462 ( .A1(n5772), .A2(n6512), .ZN(n5775) );
  MUX2_X1 U5463 ( .A(n4461), .B(n4460), .S(n5775), .Z(n4462) );
  INV_X1 U5464 ( .A(n4462), .ZN(U3456) );
  INV_X1 U5465 ( .A(n5325), .ZN(n4463) );
  INV_X1 U5466 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5321) );
  OAI222_X1 U5467 ( .A1(n4463), .A2(n5925), .B1(n5321), .B2(n5934), .C1(n5390), 
        .C2(n5329), .ZN(U2859) );
  NAND2_X1 U5468 ( .A1(n5141), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6379) );
  INV_X1 U5469 ( .A(n5194), .ZN(n5771) );
  OAI21_X1 U5470 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5190), .A(n5775), 
        .ZN(n5136) );
  AOI22_X1 U5471 ( .A1(n3446), .A2(n4790), .B1(n4464), .B2(n3031), .ZN(n6380)
         );
  OAI22_X1 U5472 ( .A1(n6380), .A2(n5771), .B1(n6418), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4465) );
  OAI22_X1 U5473 ( .A1(n5136), .A2(n4465), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5775), .ZN(n4466) );
  OAI21_X1 U5474 ( .B1(n6379), .B2(n5771), .A(n4466), .ZN(U3461) );
  INV_X1 U5475 ( .A(DATAI_2_), .ZN(n6570) );
  INV_X1 U5476 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6014) );
  OAI222_X1 U5477 ( .A1(n6081), .A2(n5669), .B1(n5083), .B2(n6570), .C1(n5392), 
        .C2(n6014), .ZN(U2889) );
  INV_X1 U5478 ( .A(DATAI_3_), .ZN(n4467) );
  INV_X1 U5479 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6017) );
  OAI222_X1 U5480 ( .A1(n5909), .A2(n5669), .B1(n5083), .B2(n4467), .C1(n5392), 
        .C2(n6017), .ZN(U2888) );
  INV_X1 U5481 ( .A(n6532), .ZN(n6434) );
  NAND2_X1 U5482 ( .A1(DATAI_3_), .A2(n4946), .ZN(n6248) );
  NAND2_X1 U5483 ( .A1(n6184), .A2(n4699), .ZN(n4478) );
  OAI21_X1 U5484 ( .B1(n4478), .B2(n5784), .A(n6272), .ZN(n4519) );
  INV_X1 U5485 ( .A(n4519), .ZN(n4474) );
  INV_X1 U5486 ( .A(n2979), .ZN(n5316) );
  OR2_X1 U5487 ( .A1(n4470), .A2(n5316), .ZN(n6320) );
  INV_X1 U5488 ( .A(n4513), .ZN(n6321) );
  NAND2_X1 U5489 ( .A1(n3446), .A2(n6321), .ZN(n6223) );
  NAND2_X1 U5490 ( .A1(n4595), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4696) );
  OR2_X1 U5491 ( .A1(n4696), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4514)
         );
  NOR2_X1 U5492 ( .A1(n6188), .A2(n4514), .ZN(n4581) );
  INV_X1 U5493 ( .A(n4581), .ZN(n4472) );
  OAI21_X1 U5494 ( .B1(n6320), .B2(n6223), .A(n4472), .ZN(n4476) );
  INV_X1 U5495 ( .A(n4514), .ZN(n4473) );
  AOI22_X1 U5496 ( .A1(n4474), .A2(n4476), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4473), .ZN(n4584) );
  OAI21_X1 U5497 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6514), .A(n4946), 
        .ZN(n6276) );
  AOI21_X1 U5498 ( .B1(n6318), .B2(n4514), .A(n6276), .ZN(n4475) );
  OAI21_X1 U5499 ( .B1(n4519), .B2(n4476), .A(n4475), .ZN(n4579) );
  NAND2_X1 U5500 ( .A1(n6075), .A2(DATAI_27_), .ZN(n6349) );
  INV_X1 U5501 ( .A(n4478), .ZN(n4477) );
  NAND2_X1 U5502 ( .A1(n4477), .A2(n4824), .ZN(n4628) );
  OR2_X1 U5503 ( .A1(n4478), .A2(n4824), .ZN(n6190) );
  NAND2_X1 U5504 ( .A1(n6075), .A2(DATAI_19_), .ZN(n6207) );
  OAI22_X1 U5505 ( .A1(n6349), .A2(n4628), .B1(n6190), .B2(n6207), .ZN(n4479)
         );
  AOI21_X1 U5506 ( .B1(n4579), .B2(INSTQUEUE_REG_5__3__SCAN_IN), .A(n4479), 
        .ZN(n4482) );
  NOR2_X2 U5507 ( .A1(n4580), .A2(n3252), .ZN(n6344) );
  NAND2_X1 U5508 ( .A1(n6344), .A2(n4581), .ZN(n4481) );
  OAI211_X1 U5509 ( .C1(n6248), .C2(n4584), .A(n4482), .B(n4481), .ZN(U3063)
         );
  NAND2_X1 U5510 ( .A1(DATAI_2_), .A2(n4946), .ZN(n6244) );
  INV_X1 U5511 ( .A(DATAI_26_), .ZN(n4483) );
  NOR2_X1 U5512 ( .A1(n6063), .A2(n4483), .ZN(n6241) );
  INV_X1 U5513 ( .A(n6241), .ZN(n6343) );
  NAND2_X1 U5514 ( .A1(n6075), .A2(DATAI_18_), .ZN(n6204) );
  OAI22_X1 U5515 ( .A1(n6343), .A2(n4628), .B1(n6190), .B2(n6204), .ZN(n4484)
         );
  AOI21_X1 U5516 ( .B1(n4579), .B2(INSTQUEUE_REG_5__2__SCAN_IN), .A(n4484), 
        .ZN(n4486) );
  NOR2_X2 U5517 ( .A1(n4580), .A2(n3220), .ZN(n6338) );
  NAND2_X1 U5518 ( .A1(n6338), .A2(n4581), .ZN(n4485) );
  OAI211_X1 U5519 ( .C1(n6244), .C2(n4584), .A(n4486), .B(n4485), .ZN(U3062)
         );
  NAND2_X1 U5520 ( .A1(DATAI_7_), .A2(n4946), .ZN(n6266) );
  NAND2_X1 U5521 ( .A1(n6075), .A2(DATAI_31_), .ZN(n6378) );
  NAND2_X1 U5522 ( .A1(n6075), .A2(DATAI_23_), .ZN(n6222) );
  OAI22_X1 U5523 ( .A1(n6378), .A2(n4628), .B1(n6190), .B2(n6222), .ZN(n4487)
         );
  AOI21_X1 U5524 ( .B1(n4579), .B2(INSTQUEUE_REG_5__7__SCAN_IN), .A(n4487), 
        .ZN(n4489) );
  NOR2_X2 U5525 ( .A1(n4580), .A2(n4404), .ZN(n6369) );
  NAND2_X1 U5526 ( .A1(n6369), .A2(n4581), .ZN(n4488) );
  OAI211_X1 U5527 ( .C1(n6266), .C2(n4584), .A(n4489), .B(n4488), .ZN(U3067)
         );
  NAND2_X1 U5528 ( .A1(DATAI_6_), .A2(n4946), .ZN(n6258) );
  INV_X1 U5529 ( .A(DATAI_30_), .ZN(n4490) );
  NOR2_X1 U5530 ( .A1(n6063), .A2(n4490), .ZN(n6297) );
  INV_X1 U5531 ( .A(n6297), .ZN(n6367) );
  NAND2_X1 U5532 ( .A1(n6075), .A2(DATAI_22_), .ZN(n6301) );
  OAI22_X1 U5533 ( .A1(n6367), .A2(n4628), .B1(n6190), .B2(n6301), .ZN(n4491)
         );
  AOI21_X1 U5534 ( .B1(n4579), .B2(INSTQUEUE_REG_5__6__SCAN_IN), .A(n4491), 
        .ZN(n4493) );
  NOR2_X2 U5535 ( .A1(n4580), .A2(n3420), .ZN(n6362) );
  NAND2_X1 U5536 ( .A1(n6362), .A2(n4581), .ZN(n4492) );
  OAI211_X1 U5537 ( .C1(n6258), .C2(n4584), .A(n4493), .B(n4492), .ZN(U3066)
         );
  XOR2_X1 U5538 ( .A(n4494), .B(n4428), .Z(n6076) );
  INV_X1 U5539 ( .A(n6076), .ZN(n4496) );
  INV_X1 U5540 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6020) );
  INV_X1 U5541 ( .A(DATAI_4_), .ZN(n4495) );
  OAI222_X1 U5542 ( .A1(n5669), .A2(n4496), .B1(n5392), .B2(n6020), .C1(n5083), 
        .C2(n4495), .ZN(U2887) );
  XNOR2_X1 U5543 ( .A(n4497), .B(n4498), .ZN(n6064) );
  OAI21_X1 U5544 ( .B1(n3000), .B2(n4499), .A(n4748), .ZN(n5875) );
  INV_X1 U5545 ( .A(n5875), .ZN(n4819) );
  AOI22_X1 U5546 ( .A1(n5930), .A2(n4819), .B1(EBX_REG_6__SCAN_IN), .B2(n5386), 
        .ZN(n4500) );
  OAI21_X1 U5547 ( .B1(n6064), .B2(n5390), .A(n4500), .ZN(U2853) );
  INV_X1 U5548 ( .A(n4498), .ZN(n4501) );
  AOI21_X1 U5549 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4565) );
  INV_X1 U5550 ( .A(n4565), .ZN(n4918) );
  INV_X1 U5551 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4508) );
  INV_X1 U5552 ( .A(n5884), .ZN(n4505) );
  OAI21_X1 U5553 ( .B1(n5885), .B2(n4505), .A(n4504), .ZN(n4506) );
  INV_X1 U5554 ( .A(n4506), .ZN(n4507) );
  OR2_X1 U5555 ( .A1(n4507), .A2(n3000), .ZN(n4908) );
  OAI222_X1 U5556 ( .A1(n4918), .A2(n5390), .B1(n4508), .B2(n5934), .C1(n4908), 
        .C2(n5925), .ZN(U2854) );
  INV_X1 U5557 ( .A(DATAI_5_), .ZN(n4509) );
  OAI222_X1 U5558 ( .A1(n4918), .A2(n5669), .B1(n5083), .B2(n4509), .C1(n5392), 
        .C2(n3483), .ZN(U2886) );
  NOR2_X1 U5559 ( .A1(n6320), .A2(n6318), .ZN(n6308) );
  INV_X1 U5560 ( .A(n4437), .ZN(n6313) );
  INV_X1 U5561 ( .A(n4830), .ZN(n4510) );
  NOR2_X1 U5562 ( .A1(n4510), .A2(n4947), .ZN(n4634) );
  INV_X1 U5563 ( .A(n4515), .ZN(n4511) );
  NOR2_X1 U5564 ( .A1(n4511), .A2(n6279), .ZN(n6309) );
  AOI22_X1 U5565 ( .A1(n6308), .A2(n6313), .B1(n4634), .B2(n6309), .ZN(n4633)
         );
  INV_X1 U5566 ( .A(n4468), .ZN(n5608) );
  NOR2_X1 U5567 ( .A1(n4512), .A2(n5608), .ZN(n4544) );
  NAND2_X1 U5568 ( .A1(n6272), .A2(n5784), .ZN(n4940) );
  INV_X1 U5569 ( .A(n4940), .ZN(n6322) );
  OAI22_X1 U5570 ( .A1(n4760), .A2(n6322), .B1(n4513), .B2(n6320), .ZN(n4518)
         );
  NOR2_X1 U5571 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4514), .ZN(n4630)
         );
  INV_X1 U5572 ( .A(n4630), .ZN(n4516) );
  NOR2_X1 U5573 ( .A1(n4515), .A2(n6279), .ZN(n6325) );
  OAI21_X1 U5574 ( .B1(n4634), .B2(n4986), .A(n4946), .ZN(n4638) );
  AOI211_X1 U5575 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4516), .A(n6325), .B(
        n4638), .ZN(n4517) );
  NAND2_X1 U5576 ( .A1(n4627), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4522) );
  OAI22_X1 U5577 ( .A1(n6349), .A2(n4760), .B1(n4628), .B2(n6207), .ZN(n4520)
         );
  AOI21_X1 U5578 ( .B1(n6344), .B2(n4630), .A(n4520), .ZN(n4521) );
  OAI211_X1 U5579 ( .C1(n4633), .C2(n6248), .A(n4522), .B(n4521), .ZN(U3055)
         );
  NAND2_X1 U5580 ( .A1(n4627), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4525) );
  OAI22_X1 U5581 ( .A1(n6343), .A2(n4760), .B1(n4628), .B2(n6204), .ZN(n4523)
         );
  AOI21_X1 U5582 ( .B1(n6338), .B2(n4630), .A(n4523), .ZN(n4524) );
  OAI211_X1 U5583 ( .C1(n4633), .C2(n6244), .A(n4525), .B(n4524), .ZN(U3054)
         );
  NAND2_X1 U5584 ( .A1(n4627), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4528) );
  OAI22_X1 U5585 ( .A1(n6378), .A2(n4760), .B1(n4628), .B2(n6222), .ZN(n4526)
         );
  AOI21_X1 U5586 ( .B1(n6369), .B2(n4630), .A(n4526), .ZN(n4527) );
  OAI211_X1 U5587 ( .C1(n4633), .C2(n6266), .A(n4528), .B(n4527), .ZN(U3059)
         );
  NAND2_X1 U5588 ( .A1(n4627), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4531) );
  OAI22_X1 U5589 ( .A1(n6367), .A2(n4760), .B1(n4628), .B2(n6301), .ZN(n4529)
         );
  AOI21_X1 U5590 ( .B1(n6362), .B2(n4630), .A(n4529), .ZN(n4530) );
  OAI211_X1 U5591 ( .C1(n4633), .C2(n6258), .A(n4531), .B(n4530), .ZN(U3058)
         );
  XOR2_X1 U5592 ( .A(n4533), .B(n4532), .Z(n4676) );
  INV_X1 U5593 ( .A(n4676), .ZN(n4537) );
  OAI22_X1 U5594 ( .A1(n5320), .A2(n6063), .B1(n6092), .B2(n6584), .ZN(n4534)
         );
  AOI21_X1 U5595 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6080), .A(n4534), 
        .ZN(n4536) );
  INV_X1 U5596 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U5597 ( .A1(n6059), .A2(n5312), .ZN(n4535) );
  OAI211_X1 U5598 ( .C1(n4537), .C2(n6065), .A(n4536), .B(n4535), .ZN(U2985)
         );
  INV_X1 U5599 ( .A(n6268), .ZN(n4538) );
  NAND2_X1 U5600 ( .A1(n4538), .A2(n6390), .ZN(n4766) );
  INV_X1 U5601 ( .A(n6369), .ZN(n4877) );
  NAND2_X1 U5602 ( .A1(n6184), .A2(n6271), .ZN(n6230) );
  OR2_X1 U5603 ( .A1(n4468), .A2(n4539), .ZN(n4876) );
  NOR2_X1 U5604 ( .A1(n2978), .A2(n5784), .ZN(n4585) );
  NAND2_X1 U5605 ( .A1(n4870), .A2(n4585), .ZN(n4702) );
  NAND3_X1 U5606 ( .A1(n6274), .A2(n6230), .A3(n4702), .ZN(n4540) );
  AND2_X1 U5607 ( .A1(n4540), .A2(n6272), .ZN(n4808) );
  AOI21_X1 U5608 ( .B1(n4468), .B2(n6271), .A(n6318), .ZN(n4541) );
  NOR2_X1 U5609 ( .A1(n4808), .A2(n4541), .ZN(n4548) );
  AND2_X1 U5610 ( .A1(n4470), .A2(n5316), .ZN(n4979) );
  AND2_X1 U5611 ( .A1(n6313), .A2(n4979), .ZN(n4943) );
  NAND2_X1 U5612 ( .A1(n4943), .A2(n3446), .ZN(n4542) );
  NAND2_X1 U5613 ( .A1(n4542), .A2(n4766), .ZN(n4546) );
  NAND3_X1 U5614 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6390), .A3(n6665), .ZN(n4939) );
  AOI21_X1 U5615 ( .B1(n6318), .B2(n4939), .A(n6276), .ZN(n4543) );
  OAI21_X1 U5616 ( .B1(n4548), .B2(n4546), .A(n4543), .ZN(n4762) );
  OAI22_X1 U5617 ( .A1(n6378), .A2(n4971), .B1(n4760), .B2(n6222), .ZN(n4545)
         );
  AOI21_X1 U5618 ( .B1(n4762), .B2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4545), 
        .ZN(n4550) );
  INV_X1 U5619 ( .A(n4546), .ZN(n4547) );
  OAI22_X1 U5620 ( .A1(n4548), .A2(n4547), .B1(n4939), .B2(n6279), .ZN(n4763)
         );
  INV_X1 U5621 ( .A(n6266), .ZN(n6371) );
  NAND2_X1 U5622 ( .A1(n4763), .A2(n6371), .ZN(n4549) );
  OAI211_X1 U5623 ( .C1(n4766), .C2(n4877), .A(n4550), .B(n4549), .ZN(U3051)
         );
  INV_X1 U5624 ( .A(n6362), .ZN(n4889) );
  OAI22_X1 U5625 ( .A1(n6367), .A2(n4971), .B1(n4760), .B2(n6301), .ZN(n4551)
         );
  AOI21_X1 U5626 ( .B1(n4762), .B2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n4551), 
        .ZN(n4553) );
  INV_X1 U5627 ( .A(n6258), .ZN(n6363) );
  NAND2_X1 U5628 ( .A1(n4763), .A2(n6363), .ZN(n4552) );
  OAI211_X1 U5629 ( .C1(n4766), .C2(n4889), .A(n4553), .B(n4552), .ZN(U3050)
         );
  INV_X1 U5630 ( .A(n6338), .ZN(n4885) );
  OAI22_X1 U5631 ( .A1(n6343), .A2(n4971), .B1(n4760), .B2(n6204), .ZN(n4554)
         );
  AOI21_X1 U5632 ( .B1(n4762), .B2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4554), 
        .ZN(n4556) );
  INV_X1 U5633 ( .A(n6244), .ZN(n6339) );
  NAND2_X1 U5634 ( .A1(n4763), .A2(n6339), .ZN(n4555) );
  OAI211_X1 U5635 ( .C1(n4766), .C2(n4885), .A(n4556), .B(n4555), .ZN(U3046)
         );
  INV_X1 U5636 ( .A(n6344), .ZN(n4881) );
  OAI22_X1 U5637 ( .A1(n6349), .A2(n4971), .B1(n4760), .B2(n6207), .ZN(n4557)
         );
  AOI21_X1 U5638 ( .B1(n4762), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4557), 
        .ZN(n4559) );
  INV_X1 U5639 ( .A(n6248), .ZN(n6345) );
  NAND2_X1 U5640 ( .A1(n4763), .A2(n6345), .ZN(n4558) );
  OAI211_X1 U5641 ( .C1(n4766), .C2(n4881), .A(n4559), .B(n4558), .ZN(U3047)
         );
  OAI21_X1 U5642 ( .B1(n4562), .B2(n4561), .A(n4560), .ZN(n6141) );
  AOI22_X1 U5643 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6171), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4563) );
  OAI21_X1 U5644 ( .B1(n4907), .B2(n6090), .A(n4563), .ZN(n4564) );
  AOI21_X1 U5645 ( .B1(n4565), .B2(n6075), .A(n4564), .ZN(n4566) );
  OAI21_X1 U5646 ( .B1(n6065), .B2(n6141), .A(n4566), .ZN(U2981) );
  NAND2_X1 U5647 ( .A1(DATAI_0_), .A2(n4946), .ZN(n6236) );
  NAND2_X1 U5648 ( .A1(n6075), .A2(DATAI_24_), .ZN(n6331) );
  NAND2_X1 U5649 ( .A1(n6075), .A2(DATAI_16_), .ZN(n6198) );
  OAI22_X1 U5650 ( .A1(n6331), .A2(n4628), .B1(n6190), .B2(n6198), .ZN(n4567)
         );
  AOI21_X1 U5651 ( .B1(n4579), .B2(INSTQUEUE_REG_5__0__SCAN_IN), .A(n4567), 
        .ZN(n4570) );
  NOR2_X2 U5652 ( .A1(n4580), .A2(n4568), .ZN(n6316) );
  NAND2_X1 U5653 ( .A1(n6316), .A2(n4581), .ZN(n4569) );
  OAI211_X1 U5654 ( .C1(n6236), .C2(n4584), .A(n4570), .B(n4569), .ZN(U3060)
         );
  NAND2_X1 U5655 ( .A1(DATAI_4_), .A2(n4946), .ZN(n6251) );
  INV_X1 U5656 ( .A(DATAI_28_), .ZN(n4571) );
  NOR2_X1 U5657 ( .A1(n6063), .A2(n4571), .ZN(n6291) );
  INV_X1 U5658 ( .A(n6291), .ZN(n6355) );
  NAND2_X1 U5659 ( .A1(n6075), .A2(DATAI_20_), .ZN(n6294) );
  OAI22_X1 U5660 ( .A1(n6355), .A2(n4628), .B1(n6190), .B2(n6294), .ZN(n4572)
         );
  AOI21_X1 U5661 ( .B1(n4579), .B2(INSTQUEUE_REG_5__4__SCAN_IN), .A(n4572), 
        .ZN(n4574) );
  NOR2_X2 U5662 ( .A1(n4580), .A2(n3247), .ZN(n6350) );
  NAND2_X1 U5663 ( .A1(n6350), .A2(n4581), .ZN(n4573) );
  OAI211_X1 U5664 ( .C1(n6251), .C2(n4584), .A(n4574), .B(n4573), .ZN(U3064)
         );
  NAND2_X1 U5665 ( .A1(DATAI_1_), .A2(n4946), .ZN(n6240) );
  NAND2_X1 U5666 ( .A1(n6075), .A2(DATAI_25_), .ZN(n6337) );
  NAND2_X1 U5667 ( .A1(n6075), .A2(DATAI_17_), .ZN(n6201) );
  OAI22_X1 U5668 ( .A1(n6337), .A2(n4628), .B1(n6190), .B2(n6201), .ZN(n4575)
         );
  AOI21_X1 U5669 ( .B1(n4579), .B2(INSTQUEUE_REG_5__1__SCAN_IN), .A(n4575), 
        .ZN(n4577) );
  NOR2_X2 U5670 ( .A1(n4580), .A2(n3946), .ZN(n6332) );
  NAND2_X1 U5671 ( .A1(n6332), .A2(n4581), .ZN(n4576) );
  OAI211_X1 U5672 ( .C1(n6240), .C2(n4584), .A(n4577), .B(n4576), .ZN(U3061)
         );
  NAND2_X1 U5673 ( .A1(DATAI_5_), .A2(n4946), .ZN(n6255) );
  NAND2_X1 U5674 ( .A1(n6075), .A2(DATAI_29_), .ZN(n6361) );
  NAND2_X1 U5675 ( .A1(n6075), .A2(DATAI_21_), .ZN(n6212) );
  OAI22_X1 U5676 ( .A1(n6361), .A2(n4628), .B1(n6190), .B2(n6212), .ZN(n4578)
         );
  AOI21_X1 U5677 ( .B1(n4579), .B2(INSTQUEUE_REG_5__5__SCAN_IN), .A(n4578), 
        .ZN(n4583) );
  NOR2_X2 U5678 ( .A1(n4580), .A2(n3222), .ZN(n6356) );
  NAND2_X1 U5679 ( .A1(n6356), .A2(n4581), .ZN(n4582) );
  OAI211_X1 U5680 ( .C1(n6255), .C2(n4584), .A(n4583), .B(n4582), .ZN(U3065)
         );
  NAND3_X1 U5681 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6665), .A3(n4595), .ZN(n4832) );
  NOR2_X1 U5682 ( .A1(n6188), .A2(n4832), .ZN(n4586) );
  INV_X1 U5683 ( .A(n4586), .ZN(n4730) );
  INV_X1 U5684 ( .A(n6276), .ZN(n6231) );
  AOI21_X1 U5685 ( .B1(n6270), .B2(n4585), .A(n6318), .ZN(n4589) );
  AND2_X1 U5686 ( .A1(n4437), .A2(n3446), .ZN(n4868) );
  NAND2_X1 U5687 ( .A1(n4470), .A2(n2979), .ZN(n4829) );
  INV_X1 U5688 ( .A(n4829), .ZN(n4587) );
  AOI21_X1 U5689 ( .B1(n4868), .B2(n4587), .A(n4586), .ZN(n4591) );
  AOI22_X1 U5690 ( .A1(n4589), .A2(n4591), .B1(n6318), .B2(n4832), .ZN(n4588)
         );
  NAND2_X1 U5691 ( .A1(n6231), .A2(n4588), .ZN(n4726) );
  INV_X1 U5692 ( .A(n4589), .ZN(n4590) );
  OAI22_X1 U5693 ( .A1(n4591), .A2(n4590), .B1(n4986), .B2(n4832), .ZN(n4725)
         );
  AOI22_X1 U5694 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4726), .B1(n6363), 
        .B2(n4725), .ZN(n4594) );
  INV_X1 U5695 ( .A(n6301), .ZN(n6364) );
  AOI22_X1 U5696 ( .A1(n4727), .A2(n6364), .B1(n4837), .B2(n6297), .ZN(n4593)
         );
  OAI211_X1 U5697 ( .C1(n4889), .C2(n4730), .A(n4594), .B(n4593), .ZN(U3098)
         );
  NAND3_X1 U5698 ( .A1(n6390), .A2(n6665), .A3(n4595), .ZN(n4637) );
  NOR2_X1 U5699 ( .A1(n6188), .A2(n4637), .ZN(n4596) );
  INV_X1 U5700 ( .A(n4596), .ZN(n4736) );
  NOR2_X1 U5701 ( .A1(n4437), .A2(n4829), .ZN(n4642) );
  AOI21_X1 U5702 ( .B1(n4642), .B2(n3446), .A(n4596), .ZN(n4600) );
  NAND2_X1 U5703 ( .A1(n4468), .A2(n4699), .ZN(n4597) );
  AOI21_X1 U5704 ( .B1(n4603), .B2(STATEBS16_REG_SCAN_IN), .A(n6318), .ZN(
        n4599) );
  AOI22_X1 U5705 ( .A1(n4600), .A2(n4599), .B1(n6318), .B2(n4637), .ZN(n4598)
         );
  NAND2_X1 U5706 ( .A1(n6231), .A2(n4598), .ZN(n4732) );
  INV_X1 U5707 ( .A(n4599), .ZN(n4601) );
  OAI22_X1 U5708 ( .A1(n4601), .A2(n4600), .B1(n4986), .B2(n4637), .ZN(n4731)
         );
  AOI22_X1 U5709 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4732), .B1(n6363), 
        .B2(n4731), .ZN(n4605) );
  INV_X1 U5710 ( .A(n4603), .ZN(n4602) );
  NAND2_X1 U5711 ( .A1(n4603), .A2(n4700), .ZN(n4972) );
  AOI22_X1 U5712 ( .A1(n4733), .A2(n6297), .B1(n6364), .B2(n4942), .ZN(n4604)
         );
  OAI211_X1 U5713 ( .C1(n4889), .C2(n4736), .A(n4605), .B(n4604), .ZN(U3034)
         );
  AOI22_X1 U5714 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4732), .B1(n6339), 
        .B2(n4731), .ZN(n4607) );
  INV_X1 U5715 ( .A(n6204), .ZN(n6340) );
  AOI22_X1 U5716 ( .A1(n4733), .A2(n6241), .B1(n6340), .B2(n4942), .ZN(n4606)
         );
  OAI211_X1 U5717 ( .C1(n4885), .C2(n4736), .A(n4607), .B(n4606), .ZN(U3030)
         );
  AOI22_X1 U5718 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4726), .B1(n6371), 
        .B2(n4725), .ZN(n4609) );
  INV_X1 U5719 ( .A(n6222), .ZN(n6373) );
  INV_X1 U5720 ( .A(n6378), .ZN(n6260) );
  AOI22_X1 U5721 ( .A1(n4727), .A2(n6373), .B1(n4837), .B2(n6260), .ZN(n4608)
         );
  OAI211_X1 U5722 ( .C1(n4877), .C2(n4730), .A(n4609), .B(n4608), .ZN(U3099)
         );
  AOI22_X1 U5723 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4726), .B1(n6345), 
        .B2(n4725), .ZN(n4611) );
  INV_X1 U5724 ( .A(n6207), .ZN(n6346) );
  INV_X1 U5725 ( .A(n6349), .ZN(n6245) );
  AOI22_X1 U5726 ( .A1(n4727), .A2(n6346), .B1(n4837), .B2(n6245), .ZN(n4610)
         );
  OAI211_X1 U5727 ( .C1(n4881), .C2(n4730), .A(n4611), .B(n4610), .ZN(U3095)
         );
  AOI22_X1 U5728 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4732), .B1(n6371), 
        .B2(n4731), .ZN(n4613) );
  AOI22_X1 U5729 ( .A1(n4733), .A2(n6260), .B1(n6373), .B2(n4942), .ZN(n4612)
         );
  OAI211_X1 U5730 ( .C1(n4877), .C2(n4736), .A(n4613), .B(n4612), .ZN(U3035)
         );
  AOI22_X1 U5731 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4726), .B1(n6339), 
        .B2(n4725), .ZN(n4615) );
  AOI22_X1 U5732 ( .A1(n4727), .A2(n6340), .B1(n4837), .B2(n6241), .ZN(n4614)
         );
  OAI211_X1 U5733 ( .C1(n4885), .C2(n4730), .A(n4615), .B(n4614), .ZN(U3094)
         );
  AOI22_X1 U5734 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4732), .B1(n6345), 
        .B2(n4731), .ZN(n4617) );
  AOI22_X1 U5735 ( .A1(n4733), .A2(n6245), .B1(n6346), .B2(n4942), .ZN(n4616)
         );
  OAI211_X1 U5736 ( .C1(n4881), .C2(n4736), .A(n4617), .B(n4616), .ZN(U3031)
         );
  NAND2_X1 U5737 ( .A1(n4627), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4620) );
  OAI22_X1 U5738 ( .A1(n6337), .A2(n4760), .B1(n4628), .B2(n6201), .ZN(n4618)
         );
  AOI21_X1 U5739 ( .B1(n6332), .B2(n4630), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5740 ( .C1(n4633), .C2(n6240), .A(n4620), .B(n4619), .ZN(U3053)
         );
  NAND2_X1 U5741 ( .A1(n4627), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4623) );
  OAI22_X1 U5742 ( .A1(n6361), .A2(n4760), .B1(n4628), .B2(n6212), .ZN(n4621)
         );
  AOI21_X1 U5743 ( .B1(n6356), .B2(n4630), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5744 ( .C1(n4633), .C2(n6255), .A(n4623), .B(n4622), .ZN(U3057)
         );
  NAND2_X1 U5745 ( .A1(n4627), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5746 ( .A1(n6355), .A2(n4760), .B1(n4628), .B2(n6294), .ZN(n4624)
         );
  AOI21_X1 U5747 ( .B1(n6350), .B2(n4630), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5748 ( .C1(n4633), .C2(n6251), .A(n4626), .B(n4625), .ZN(U3056)
         );
  NAND2_X1 U5749 ( .A1(n4627), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5750 ( .A1(n6331), .A2(n4760), .B1(n4628), .B2(n6198), .ZN(n4629)
         );
  AOI21_X1 U5751 ( .B1(n6316), .B2(n4630), .A(n4629), .ZN(n4631) );
  OAI211_X1 U5752 ( .C1(n4633), .C2(n6236), .A(n4632), .B(n4631), .ZN(U3052)
         );
  AOI22_X1 U5753 ( .A1(n4642), .A2(n6272), .B1(n6325), .B2(n4634), .ZN(n4694)
         );
  INV_X1 U5754 ( .A(n6269), .ZN(n4635) );
  NOR2_X1 U5755 ( .A1(n4876), .A2(n4635), .ZN(n4643) );
  NOR3_X1 U5756 ( .A1(n4733), .A2(n4643), .A3(n6318), .ZN(n4636) );
  NOR2_X1 U5757 ( .A1(n4636), .A2(n6322), .ZN(n4641) );
  NOR2_X1 U5758 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4637), .ZN(n4691)
         );
  INV_X1 U5759 ( .A(n4691), .ZN(n4639) );
  AOI211_X1 U5760 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4639), .A(n6309), .B(
        n4638), .ZN(n4640) );
  NAND2_X1 U5761 ( .A1(n4688), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4646) );
  OAI22_X1 U5762 ( .A1(n4689), .A2(n6204), .B1(n6343), .B2(n4931), .ZN(n4644)
         );
  AOI21_X1 U5763 ( .B1(n6338), .B2(n4691), .A(n4644), .ZN(n4645) );
  OAI211_X1 U5764 ( .C1(n4694), .C2(n6244), .A(n4646), .B(n4645), .ZN(U3022)
         );
  NAND2_X1 U5765 ( .A1(n4688), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4649) );
  OAI22_X1 U5766 ( .A1(n4689), .A2(n6222), .B1(n6378), .B2(n4931), .ZN(n4647)
         );
  AOI21_X1 U5767 ( .B1(n6369), .B2(n4691), .A(n4647), .ZN(n4648) );
  OAI211_X1 U5768 ( .C1(n4694), .C2(n6266), .A(n4649), .B(n4648), .ZN(U3027)
         );
  NAND2_X1 U5769 ( .A1(n4688), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4652) );
  OAI22_X1 U5770 ( .A1(n4689), .A2(n6301), .B1(n6367), .B2(n4931), .ZN(n4650)
         );
  AOI21_X1 U5771 ( .B1(n6362), .B2(n4691), .A(n4650), .ZN(n4651) );
  OAI211_X1 U5772 ( .C1(n4694), .C2(n6258), .A(n4652), .B(n4651), .ZN(U3026)
         );
  NAND2_X1 U5773 ( .A1(n4688), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4655) );
  OAI22_X1 U5774 ( .A1(n4689), .A2(n6207), .B1(n6349), .B2(n4931), .ZN(n4653)
         );
  AOI21_X1 U5775 ( .B1(n6344), .B2(n4691), .A(n4653), .ZN(n4654) );
  OAI211_X1 U5776 ( .C1(n4694), .C2(n6248), .A(n4655), .B(n4654), .ZN(U3023)
         );
  INV_X1 U5777 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U5778 ( .A1(n4657), .A2(n5141), .ZN(n4658) );
  NAND2_X1 U5779 ( .A1(n5948), .A2(n3253), .ZN(n5050) );
  NOR2_X1 U5780 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4822), .ZN(n5956) );
  INV_X1 U5781 ( .A(n5956), .ZN(n6527) );
  NOR2_X4 U5782 ( .A1(n5948), .A2(n5966), .ZN(n5960) );
  AOI22_X1 U5783 ( .A1(n5966), .A2(UWORD_REG_9__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4661) );
  OAI21_X1 U5784 ( .B1(n5992), .B2(n5050), .A(n4661), .ZN(U2898) );
  INV_X1 U5785 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5997) );
  AOI22_X1 U5786 ( .A1(n5966), .A2(UWORD_REG_11__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5787 ( .B1(n5997), .B2(n5050), .A(n4662), .ZN(U2896) );
  INV_X1 U5788 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6002) );
  AOI22_X1 U5789 ( .A1(n5966), .A2(UWORD_REG_13__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4663) );
  OAI21_X1 U5790 ( .B1(n6002), .B2(n5050), .A(n4663), .ZN(U2894) );
  OAI21_X1 U5791 ( .B1(n4666), .B2(n4665), .A(n4664), .ZN(n6159) );
  NOR2_X1 U5792 ( .A1(n6092), .A2(n6461), .ZN(n6156) );
  NOR2_X1 U5793 ( .A1(n5483), .A2(n6591), .ZN(n4667) );
  AOI211_X1 U5794 ( .C1(n6059), .C2(n5913), .A(n6156), .B(n4667), .ZN(n4670)
         );
  NAND2_X1 U5795 ( .A1(n4668), .A2(n6075), .ZN(n4669) );
  OAI211_X1 U5796 ( .C1(n6159), .C2(n6065), .A(n4670), .B(n4669), .ZN(U2983)
         );
  INV_X1 U5797 ( .A(n4671), .ZN(n4672) );
  AOI21_X1 U5798 ( .B1(n5189), .B2(n5591), .A(n4672), .ZN(n4678) );
  OAI22_X1 U5799 ( .A1(n6094), .A2(n4673), .B1(n6584), .B2(n6092), .ZN(n4675)
         );
  AOI211_X1 U5800 ( .C1(n5189), .C2(n5594), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n6106), .ZN(n4674) );
  AOI211_X1 U5801 ( .C1(n6175), .C2(n4676), .A(n4675), .B(n4674), .ZN(n4677)
         );
  OAI21_X1 U5802 ( .B1(n4678), .B2(n5137), .A(n4677), .ZN(U3017) );
  NAND2_X1 U5803 ( .A1(n4688), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4681) );
  OAI22_X1 U5804 ( .A1(n4689), .A2(n6294), .B1(n6355), .B2(n4931), .ZN(n4679)
         );
  AOI21_X1 U5805 ( .B1(n6350), .B2(n4691), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5806 ( .C1(n4694), .C2(n6251), .A(n4681), .B(n4680), .ZN(U3024)
         );
  NAND2_X1 U5807 ( .A1(n4688), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4684) );
  OAI22_X1 U5808 ( .A1(n4689), .A2(n6201), .B1(n6337), .B2(n4931), .ZN(n4682)
         );
  AOI21_X1 U5809 ( .B1(n6332), .B2(n4691), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5810 ( .C1(n4694), .C2(n6240), .A(n4684), .B(n4683), .ZN(U3021)
         );
  NAND2_X1 U5811 ( .A1(n4688), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4687) );
  OAI22_X1 U5812 ( .A1(n4689), .A2(n6212), .B1(n6361), .B2(n4931), .ZN(n4685)
         );
  AOI21_X1 U5813 ( .B1(n6356), .B2(n4691), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5814 ( .C1(n4694), .C2(n6255), .A(n4687), .B(n4686), .ZN(U3025)
         );
  NAND2_X1 U5815 ( .A1(n4688), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4693) );
  OAI22_X1 U5816 ( .A1(n4689), .A2(n6198), .B1(n6331), .B2(n4931), .ZN(n4690)
         );
  AOI21_X1 U5817 ( .B1(n6316), .B2(n4691), .A(n4690), .ZN(n4692) );
  OAI211_X1 U5818 ( .C1(n4694), .C2(n6236), .A(n4693), .B(n4692), .ZN(U3020)
         );
  INV_X1 U5819 ( .A(n6320), .ZN(n4695) );
  NOR2_X1 U5820 ( .A1(n6390), .A2(n4696), .ZN(n4704) );
  INV_X1 U5821 ( .A(n4704), .ZN(n6315) );
  NOR2_X1 U5822 ( .A1(n6188), .A2(n6315), .ZN(n4781) );
  AOI21_X1 U5823 ( .B1(n4868), .B2(n4695), .A(n4781), .ZN(n4703) );
  NAND2_X1 U5824 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4697) );
  OAI22_X1 U5825 ( .A1(n4703), .A2(n6318), .B1(n4697), .B2(n4696), .ZN(n4698)
         );
  NAND2_X1 U5826 ( .A1(n4870), .A2(n4699), .ZN(n4701) );
  NOR2_X1 U5827 ( .A1(n4701), .A2(n4824), .ZN(n5153) );
  NOR2_X2 U5828 ( .A1(n4701), .A2(n4700), .ZN(n6372) );
  NAND2_X1 U5829 ( .A1(n4703), .A2(n4702), .ZN(n4706) );
  OR2_X1 U5830 ( .A1(n6272), .A2(n4704), .ZN(n4705) );
  OAI211_X1 U5831 ( .C1(n4706), .C2(n6318), .A(n4705), .B(n6231), .ZN(n4778)
         );
  AOI22_X1 U5832 ( .A1(n6372), .A2(n6245), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4778), .ZN(n4707) );
  OAI21_X1 U5833 ( .B1(n5180), .B2(n6207), .A(n4707), .ZN(n4708) );
  AOI21_X1 U5834 ( .B1(n6344), .B2(n4781), .A(n4708), .ZN(n4709) );
  OAI21_X1 U5835 ( .B1(n6248), .B2(n4783), .A(n4709), .ZN(U3127) );
  AOI22_X1 U5836 ( .A1(n6372), .A2(n6241), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4778), .ZN(n4710) );
  OAI21_X1 U5837 ( .B1(n5180), .B2(n6204), .A(n4710), .ZN(n4711) );
  AOI21_X1 U5838 ( .B1(n6338), .B2(n4781), .A(n4711), .ZN(n4712) );
  OAI21_X1 U5839 ( .B1(n6244), .B2(n4783), .A(n4712), .ZN(U3126) );
  INV_X1 U5840 ( .A(n6316), .ZN(n4927) );
  INV_X1 U5841 ( .A(n6236), .ZN(n6317) );
  AOI22_X1 U5842 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4726), .B1(n6317), 
        .B2(n4725), .ZN(n4714) );
  INV_X1 U5843 ( .A(n6198), .ZN(n6328) );
  INV_X1 U5844 ( .A(n6331), .ZN(n6228) );
  AOI22_X1 U5845 ( .A1(n4727), .A2(n6328), .B1(n4837), .B2(n6228), .ZN(n4713)
         );
  OAI211_X1 U5846 ( .C1(n4927), .C2(n4730), .A(n4714), .B(n4713), .ZN(U3092)
         );
  INV_X1 U5847 ( .A(n6350), .ZN(n4933) );
  INV_X1 U5848 ( .A(n6251), .ZN(n6351) );
  AOI22_X1 U5849 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4732), .B1(n6351), 
        .B2(n4731), .ZN(n4716) );
  INV_X1 U5850 ( .A(n6294), .ZN(n6352) );
  AOI22_X1 U5851 ( .A1(n4733), .A2(n6291), .B1(n6352), .B2(n4942), .ZN(n4715)
         );
  OAI211_X1 U5852 ( .C1(n4933), .C2(n4736), .A(n4716), .B(n4715), .ZN(U3032)
         );
  INV_X1 U5853 ( .A(n6356), .ZN(n4919) );
  INV_X1 U5854 ( .A(n6255), .ZN(n6357) );
  AOI22_X1 U5855 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4732), .B1(n6357), 
        .B2(n4731), .ZN(n4718) );
  INV_X1 U5856 ( .A(n6361), .ZN(n6252) );
  INV_X1 U5857 ( .A(n6212), .ZN(n6358) );
  AOI22_X1 U5858 ( .A1(n4733), .A2(n6252), .B1(n6358), .B2(n4942), .ZN(n4717)
         );
  OAI211_X1 U5859 ( .C1(n4919), .C2(n4736), .A(n4718), .B(n4717), .ZN(U3033)
         );
  INV_X1 U5860 ( .A(n6332), .ZN(n4923) );
  INV_X1 U5861 ( .A(n6240), .ZN(n6333) );
  AOI22_X1 U5862 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4726), .B1(n6333), 
        .B2(n4725), .ZN(n4720) );
  INV_X1 U5863 ( .A(n6201), .ZN(n6334) );
  INV_X1 U5864 ( .A(n6337), .ZN(n6237) );
  AOI22_X1 U5865 ( .A1(n4727), .A2(n6334), .B1(n4837), .B2(n6237), .ZN(n4719)
         );
  OAI211_X1 U5866 ( .C1(n4923), .C2(n4730), .A(n4720), .B(n4719), .ZN(U3093)
         );
  AOI22_X1 U5867 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4726), .B1(n6351), 
        .B2(n4725), .ZN(n4722) );
  AOI22_X1 U5868 ( .A1(n4727), .A2(n6352), .B1(n4837), .B2(n6291), .ZN(n4721)
         );
  OAI211_X1 U5869 ( .C1(n4933), .C2(n4730), .A(n4722), .B(n4721), .ZN(U3096)
         );
  AOI22_X1 U5870 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4732), .B1(n6317), 
        .B2(n4731), .ZN(n4724) );
  AOI22_X1 U5871 ( .A1(n4733), .A2(n6228), .B1(n6328), .B2(n4942), .ZN(n4723)
         );
  OAI211_X1 U5872 ( .C1(n4927), .C2(n4736), .A(n4724), .B(n4723), .ZN(U3028)
         );
  AOI22_X1 U5873 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4726), .B1(n6357), 
        .B2(n4725), .ZN(n4729) );
  AOI22_X1 U5874 ( .A1(n4727), .A2(n6358), .B1(n4837), .B2(n6252), .ZN(n4728)
         );
  OAI211_X1 U5875 ( .C1(n4919), .C2(n4730), .A(n4729), .B(n4728), .ZN(U3097)
         );
  AOI22_X1 U5876 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4732), .B1(n6333), 
        .B2(n4731), .ZN(n4735) );
  AOI22_X1 U5877 ( .A1(n4733), .A2(n6237), .B1(n6334), .B2(n4942), .ZN(n4734)
         );
  OAI211_X1 U5878 ( .C1(n4923), .C2(n4736), .A(n4735), .B(n4734), .ZN(U3029)
         );
  AOI22_X1 U5879 ( .A1(n6372), .A2(n6260), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4778), .ZN(n4737) );
  OAI21_X1 U5880 ( .B1(n5180), .B2(n6222), .A(n4737), .ZN(n4738) );
  AOI21_X1 U5881 ( .B1(n6369), .B2(n4781), .A(n4738), .ZN(n4739) );
  OAI21_X1 U5882 ( .B1(n6266), .B2(n4783), .A(n4739), .ZN(U3131) );
  AOI22_X1 U5883 ( .A1(n6372), .A2(n6297), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4778), .ZN(n4740) );
  OAI21_X1 U5884 ( .B1(n5180), .B2(n6301), .A(n4740), .ZN(n4741) );
  AOI21_X1 U5885 ( .B1(n6362), .B2(n4781), .A(n4741), .ZN(n4742) );
  OAI21_X1 U5886 ( .B1(n6258), .B2(n4783), .A(n4742), .ZN(U3130) );
  XOR2_X1 U5887 ( .A(n4743), .B(n4744), .Z(n4899) );
  AOI22_X1 U5888 ( .A1(n5134), .A2(DATAI_7_), .B1(n5944), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4745) );
  OAI21_X1 U5889 ( .B1(n5311), .B2(n5669), .A(n4745), .ZN(U2884) );
  INV_X1 U5890 ( .A(n4746), .ZN(n4747) );
  AOI21_X1 U5891 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n6128) );
  AOI22_X1 U5892 ( .A1(n5930), .A2(n6128), .B1(EBX_REG_7__SCAN_IN), .B2(n5386), 
        .ZN(n4750) );
  OAI21_X1 U5893 ( .B1(n5311), .B2(n5390), .A(n4750), .ZN(U2852) );
  OAI22_X1 U5894 ( .A1(n6355), .A2(n4971), .B1(n4760), .B2(n6294), .ZN(n4751)
         );
  AOI21_X1 U5895 ( .B1(n4762), .B2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n4751), 
        .ZN(n4753) );
  NAND2_X1 U5896 ( .A1(n4763), .A2(n6351), .ZN(n4752) );
  OAI211_X1 U5897 ( .C1(n4766), .C2(n4933), .A(n4753), .B(n4752), .ZN(U3048)
         );
  OAI22_X1 U5898 ( .A1(n6331), .A2(n4971), .B1(n4760), .B2(n6198), .ZN(n4754)
         );
  AOI21_X1 U5899 ( .B1(n4762), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4754), 
        .ZN(n4756) );
  NAND2_X1 U5900 ( .A1(n4763), .A2(n6317), .ZN(n4755) );
  OAI211_X1 U5901 ( .C1(n4766), .C2(n4927), .A(n4756), .B(n4755), .ZN(U3044)
         );
  OAI22_X1 U5902 ( .A1(n6361), .A2(n4971), .B1(n4760), .B2(n6212), .ZN(n4757)
         );
  AOI21_X1 U5903 ( .B1(n4762), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4757), 
        .ZN(n4759) );
  NAND2_X1 U5904 ( .A1(n4763), .A2(n6357), .ZN(n4758) );
  OAI211_X1 U5905 ( .C1(n4766), .C2(n4919), .A(n4759), .B(n4758), .ZN(U3049)
         );
  OAI22_X1 U5906 ( .A1(n6337), .A2(n4971), .B1(n4760), .B2(n6201), .ZN(n4761)
         );
  AOI21_X1 U5907 ( .B1(n4762), .B2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4761), 
        .ZN(n4765) );
  NAND2_X1 U5908 ( .A1(n4763), .A2(n6333), .ZN(n4764) );
  OAI211_X1 U5909 ( .C1(n4766), .C2(n4923), .A(n4765), .B(n4764), .ZN(U3045)
         );
  AOI22_X1 U5910 ( .A1(n5930), .A2(n6120), .B1(EBX_REG_8__SCAN_IN), .B2(n5386), 
        .ZN(n4767) );
  OAI21_X1 U5911 ( .B1(n5018), .B2(n5390), .A(n4767), .ZN(U2851) );
  AOI22_X1 U5912 ( .A1(n5134), .A2(DATAI_8_), .B1(n5944), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4768) );
  OAI21_X1 U5913 ( .B1(n5018), .B2(n5669), .A(n4768), .ZN(U2883) );
  AOI22_X1 U5914 ( .A1(n6372), .A2(n6228), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4778), .ZN(n4769) );
  OAI21_X1 U5915 ( .B1(n5180), .B2(n6198), .A(n4769), .ZN(n4770) );
  AOI21_X1 U5916 ( .B1(n6316), .B2(n4781), .A(n4770), .ZN(n4771) );
  OAI21_X1 U5917 ( .B1(n6236), .B2(n4783), .A(n4771), .ZN(U3124) );
  AOI22_X1 U5918 ( .A1(n6372), .A2(n6237), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4778), .ZN(n4772) );
  OAI21_X1 U5919 ( .B1(n5180), .B2(n6201), .A(n4772), .ZN(n4773) );
  AOI21_X1 U5920 ( .B1(n6332), .B2(n4781), .A(n4773), .ZN(n4774) );
  OAI21_X1 U5921 ( .B1(n6240), .B2(n4783), .A(n4774), .ZN(U3125) );
  AOI22_X1 U5922 ( .A1(n6372), .A2(n6291), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4778), .ZN(n4775) );
  OAI21_X1 U5923 ( .B1(n5180), .B2(n6294), .A(n4775), .ZN(n4776) );
  AOI21_X1 U5924 ( .B1(n6350), .B2(n4781), .A(n4776), .ZN(n4777) );
  OAI21_X1 U5925 ( .B1(n6251), .B2(n4783), .A(n4777), .ZN(U3128) );
  AOI22_X1 U5926 ( .A1(n6372), .A2(n6252), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4778), .ZN(n4779) );
  OAI21_X1 U5927 ( .B1(n5180), .B2(n6212), .A(n4779), .ZN(n4780) );
  AOI21_X1 U5928 ( .B1(n6356), .B2(n4781), .A(n4780), .ZN(n4782) );
  OAI21_X1 U5929 ( .B1(n6255), .B2(n4783), .A(n4782), .ZN(U3129) );
  NAND2_X1 U5930 ( .A1(n4436), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5931 ( .A1(n4785), .A2(n4784), .ZN(n4793) );
  INV_X1 U5932 ( .A(n5141), .ZN(n4789) );
  XNOR2_X1 U5933 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4788) );
  INV_X1 U5934 ( .A(n4786), .ZN(n4787) );
  OAI22_X1 U5935 ( .A1(n4789), .A2(n4788), .B1(n4787), .B2(n4793), .ZN(n4792)
         );
  INV_X1 U5936 ( .A(n4790), .ZN(n5143) );
  NOR2_X1 U5937 ( .A1(n4470), .A2(n5143), .ZN(n4791) );
  AOI211_X1 U5938 ( .C1(n4794), .C2(n4793), .A(n4792), .B(n4791), .ZN(n5187)
         );
  MUX2_X1 U5939 ( .A(n5187), .B(n3110), .S(n4795), .Z(n6388) );
  NOR2_X1 U5940 ( .A1(n6388), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4798) );
  MUX2_X1 U5941 ( .A(n4796), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4795), 
        .Z(n6391) );
  INV_X1 U5942 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6572) );
  AND2_X1 U5943 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6572), .ZN(n4802) );
  AOI22_X1 U5944 ( .A1(n4798), .A2(n6391), .B1(n4797), .B2(n4802), .ZN(n6394)
         );
  OR2_X1 U5945 ( .A1(n4800), .A2(n6321), .ZN(n4801) );
  XNOR2_X1 U5946 ( .A(n4801), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5893)
         );
  INV_X1 U5947 ( .A(n5893), .ZN(n5769) );
  OAI22_X1 U5948 ( .A1(n6382), .A2(n5774), .B1(n5770), .B2(n5769), .ZN(n4803)
         );
  AOI22_X1 U5949 ( .A1(n4803), .A2(n6418), .B1(n4802), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U5950 ( .B1(n6394), .B2(n4799), .A(n6407), .ZN(n4823) );
  OAI21_X1 U5951 ( .B1(n4823), .B2(FLUSH_REG_SCAN_IN), .A(n6433), .ZN(n4805)
         );
  INV_X1 U5952 ( .A(n4946), .ZN(n4804) );
  AND2_X1 U5953 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6514), .ZN(n5609) );
  OAI22_X1 U5954 ( .A1(n4806), .A2(n4940), .B1(n6313), .B2(n5609), .ZN(n4807)
         );
  OAI21_X1 U5955 ( .B1(n4808), .B2(n4807), .A(n6181), .ZN(n4809) );
  OAI21_X1 U5956 ( .B1(n6181), .B2(n6390), .A(n4809), .ZN(U3462) );
  OR2_X1 U5957 ( .A1(n4811), .A2(n4810), .ZN(n4812) );
  NAND2_X1 U5958 ( .A1(n4813), .A2(n4812), .ZN(n6066) );
  NOR2_X1 U5959 ( .A1(n6137), .A2(n5137), .ZN(n6176) );
  AOI21_X1 U5960 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6176), .A(n6172), 
        .ZN(n6158) );
  NAND2_X1 U5961 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6140), .ZN(n4815)
         );
  NOR2_X1 U5962 ( .A1(n6158), .A2(n4815), .ZN(n4817) );
  NAND2_X1 U5963 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4814) );
  AOI21_X1 U5964 ( .B1(n5103), .B2(n4814), .A(n5101), .ZN(n6180) );
  INV_X1 U5965 ( .A(n6180), .ZN(n6148) );
  AOI21_X1 U5966 ( .B1(n5586), .B2(n4815), .A(n6148), .ZN(n6147) );
  INV_X1 U5967 ( .A(n6147), .ZN(n4816) );
  MUX2_X1 U5968 ( .A(n4817), .B(n4816), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4818) );
  INV_X1 U5969 ( .A(n4818), .ZN(n4821) );
  AOI22_X1 U5970 ( .A1(n6169), .A2(n4819), .B1(n6171), .B2(REIP_REG_6__SCAN_IN), .ZN(n4820) );
  OAI211_X1 U5971 ( .C1(n6095), .C2(n6066), .A(n4821), .B(n4820), .ZN(U3012)
         );
  NOR2_X1 U5972 ( .A1(n4823), .A2(n4822), .ZN(n6420) );
  OAI22_X1 U5973 ( .A1(n4824), .A2(n6318), .B1(n5322), .B2(n5609), .ZN(n4825)
         );
  OAI21_X1 U5974 ( .B1(n6420), .B2(n4825), .A(n6181), .ZN(n4826) );
  OAI21_X1 U5975 ( .B1(n6181), .B2(n6188), .A(n4826), .ZN(U3465) );
  INV_X1 U5976 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6009) );
  INV_X1 U5977 ( .A(DATAI_0_), .ZN(n4827) );
  OAI222_X1 U5978 ( .A1(n5669), .A2(n5329), .B1(n5392), .B2(n6009), .C1(n5083), 
        .C2(n4827), .ZN(U2891) );
  INV_X1 U5979 ( .A(DATAI_6_), .ZN(n5981) );
  OAI222_X1 U5980 ( .A1(n5981), .A2(n5083), .B1(n5669), .B2(n6064), .C1(n4828), 
        .C2(n5392), .ZN(U2885) );
  NOR2_X1 U5981 ( .A1(n6313), .A2(n4829), .ZN(n4836) );
  NOR2_X1 U5982 ( .A1(n4947), .A2(n4830), .ZN(n6310) );
  AOI22_X1 U5983 ( .A1(n4836), .A2(n6272), .B1(n6325), .B2(n6310), .ZN(n4866)
         );
  NOR3_X1 U5984 ( .A1(n4837), .A2(n6262), .A3(n6318), .ZN(n4831) );
  NOR2_X1 U5985 ( .A1(n4831), .A2(n6322), .ZN(n4835) );
  NOR2_X1 U5986 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4832), .ZN(n4863)
         );
  INV_X1 U5987 ( .A(n4863), .ZN(n4833) );
  OAI21_X1 U5988 ( .B1(n6310), .B2(n4986), .A(n4946), .ZN(n6324) );
  AOI211_X1 U5989 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4833), .A(n6309), .B(
        n6324), .ZN(n4834) );
  NAND2_X1 U5990 ( .A1(n4859), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4840) );
  OAI22_X1 U5991 ( .A1(n4861), .A2(n6294), .B1(n6355), .B2(n4860), .ZN(n4838)
         );
  AOI21_X1 U5992 ( .B1(n6350), .B2(n4863), .A(n4838), .ZN(n4839) );
  OAI211_X1 U5993 ( .C1(n4866), .C2(n6251), .A(n4840), .B(n4839), .ZN(U3088)
         );
  NAND2_X1 U5994 ( .A1(n4859), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4843) );
  OAI22_X1 U5995 ( .A1(n4861), .A2(n6201), .B1(n6337), .B2(n4860), .ZN(n4841)
         );
  AOI21_X1 U5996 ( .B1(n6332), .B2(n4863), .A(n4841), .ZN(n4842) );
  OAI211_X1 U5997 ( .C1(n4866), .C2(n6240), .A(n4843), .B(n4842), .ZN(U3085)
         );
  NAND2_X1 U5998 ( .A1(n4859), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4846) );
  OAI22_X1 U5999 ( .A1(n4861), .A2(n6301), .B1(n6367), .B2(n4860), .ZN(n4844)
         );
  AOI21_X1 U6000 ( .B1(n6362), .B2(n4863), .A(n4844), .ZN(n4845) );
  OAI211_X1 U6001 ( .C1(n4866), .C2(n6258), .A(n4846), .B(n4845), .ZN(U3090)
         );
  NAND2_X1 U6002 ( .A1(n4859), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4849) );
  OAI22_X1 U6003 ( .A1(n4861), .A2(n6198), .B1(n6331), .B2(n4860), .ZN(n4847)
         );
  AOI21_X1 U6004 ( .B1(n6316), .B2(n4863), .A(n4847), .ZN(n4848) );
  OAI211_X1 U6005 ( .C1(n4866), .C2(n6236), .A(n4849), .B(n4848), .ZN(U3084)
         );
  NAND2_X1 U6006 ( .A1(n4859), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4852) );
  OAI22_X1 U6007 ( .A1(n4861), .A2(n6212), .B1(n6361), .B2(n4860), .ZN(n4850)
         );
  AOI21_X1 U6008 ( .B1(n6356), .B2(n4863), .A(n4850), .ZN(n4851) );
  OAI211_X1 U6009 ( .C1(n4866), .C2(n6255), .A(n4852), .B(n4851), .ZN(U3089)
         );
  NAND2_X1 U6010 ( .A1(n4859), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4855) );
  OAI22_X1 U6011 ( .A1(n4861), .A2(n6222), .B1(n6378), .B2(n4860), .ZN(n4853)
         );
  AOI21_X1 U6012 ( .B1(n6369), .B2(n4863), .A(n4853), .ZN(n4854) );
  OAI211_X1 U6013 ( .C1(n4866), .C2(n6266), .A(n4855), .B(n4854), .ZN(U3091)
         );
  NAND2_X1 U6014 ( .A1(n4859), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4858) );
  OAI22_X1 U6015 ( .A1(n4861), .A2(n6204), .B1(n6343), .B2(n4860), .ZN(n4856)
         );
  AOI21_X1 U6016 ( .B1(n6338), .B2(n4863), .A(n4856), .ZN(n4857) );
  OAI211_X1 U6017 ( .C1(n4866), .C2(n6244), .A(n4858), .B(n4857), .ZN(U3086)
         );
  NAND2_X1 U6018 ( .A1(n4859), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4865) );
  OAI22_X1 U6019 ( .A1(n4861), .A2(n6207), .B1(n6349), .B2(n4860), .ZN(n4862)
         );
  AOI21_X1 U6020 ( .B1(n6344), .B2(n4863), .A(n4862), .ZN(n4864) );
  OAI211_X1 U6021 ( .C1(n4866), .C2(n6248), .A(n4865), .B(n4864), .ZN(U3087)
         );
  OR2_X1 U6022 ( .A1(n4470), .A2(n2979), .ZN(n6191) );
  INV_X1 U6023 ( .A(n6191), .ZN(n6226) );
  INV_X1 U6024 ( .A(n4932), .ZN(n4867) );
  AOI21_X1 U6025 ( .B1(n4868), .B2(n6226), .A(n4867), .ZN(n4871) );
  INV_X1 U6026 ( .A(n4871), .ZN(n4869) );
  AOI22_X1 U6027 ( .A1(n4869), .A2(n6272), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4874), .ZN(n4938) );
  AOI21_X1 U6028 ( .B1(n4870), .B2(n2978), .A(n6063), .ZN(n4872) );
  OAI21_X1 U6029 ( .B1(n4872), .B2(n6322), .A(n4871), .ZN(n4873) );
  OAI211_X1 U6030 ( .C1(n6272), .C2(n4874), .A(n4873), .B(n6231), .ZN(n4936)
         );
  INV_X1 U6031 ( .A(n6183), .ZN(n4875) );
  NOR2_X1 U6032 ( .A1(n4876), .A2(n4875), .ZN(n5152) );
  OAI22_X1 U6033 ( .A1(n6378), .A2(n5179), .B1(n4931), .B2(n6222), .ZN(n4879)
         );
  NOR2_X1 U6034 ( .A1(n4877), .A2(n4932), .ZN(n4878) );
  AOI211_X1 U6035 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4936), .A(n4879), 
        .B(n4878), .ZN(n4880) );
  OAI21_X1 U6036 ( .B1(n4938), .B2(n6266), .A(n4880), .ZN(U3147) );
  OAI22_X1 U6037 ( .A1(n6349), .A2(n5179), .B1(n4931), .B2(n6207), .ZN(n4883)
         );
  NOR2_X1 U6038 ( .A1(n4881), .A2(n4932), .ZN(n4882) );
  AOI211_X1 U6039 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n4936), .A(n4883), 
        .B(n4882), .ZN(n4884) );
  OAI21_X1 U6040 ( .B1(n4938), .B2(n6248), .A(n4884), .ZN(U3143) );
  OAI22_X1 U6041 ( .A1(n6343), .A2(n5179), .B1(n4931), .B2(n6204), .ZN(n4887)
         );
  NOR2_X1 U6042 ( .A1(n4885), .A2(n4932), .ZN(n4886) );
  AOI211_X1 U6043 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n4936), .A(n4887), 
        .B(n4886), .ZN(n4888) );
  OAI21_X1 U6044 ( .B1(n4938), .B2(n6244), .A(n4888), .ZN(U3142) );
  OAI22_X1 U6045 ( .A1(n6367), .A2(n5179), .B1(n4931), .B2(n6301), .ZN(n4891)
         );
  NOR2_X1 U6046 ( .A1(n4889), .A2(n4932), .ZN(n4890) );
  AOI211_X1 U6047 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n4936), .A(n4891), 
        .B(n4890), .ZN(n4892) );
  OAI21_X1 U6048 ( .B1(n4938), .B2(n6258), .A(n4892), .ZN(U3146) );
  OAI21_X1 U6049 ( .B1(n4895), .B2(n4894), .A(n4893), .ZN(n6129) );
  NAND2_X1 U6050 ( .A1(n6059), .A2(n5303), .ZN(n4896) );
  NAND2_X1 U6051 ( .A1(n6171), .A2(REIP_REG_7__SCAN_IN), .ZN(n6126) );
  OAI211_X1 U6052 ( .C1(n5483), .C2(n4897), .A(n4896), .B(n6126), .ZN(n4898)
         );
  AOI21_X1 U6053 ( .B1(n4899), .B2(n6075), .A(n4898), .ZN(n4900) );
  OAI21_X1 U6054 ( .B1(n6129), .B2(n6065), .A(n4900), .ZN(U2979) );
  NAND2_X1 U6055 ( .A1(n4361), .A2(n4903), .ZN(n4904) );
  NAND2_X1 U6056 ( .A1(n4902), .A2(n4904), .ZN(n5926) );
  AOI22_X1 U6057 ( .A1(n5134), .A2(DATAI_9_), .B1(n5944), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4905) );
  OAI21_X1 U6058 ( .B1(n5926), .B2(n5669), .A(n4905), .ZN(U2882) );
  NAND2_X1 U6059 ( .A1(n5028), .A2(n4256), .ZN(n4906) );
  INV_X1 U6060 ( .A(n4907), .ZN(n4912) );
  INV_X1 U6061 ( .A(n4908), .ZN(n6142) );
  AOI22_X1 U6062 ( .A1(n5906), .A2(n6142), .B1(n5903), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4909) );
  OAI211_X1 U6063 ( .C1(n5889), .C2(n4910), .A(n4909), .B(n5301), .ZN(n4911)
         );
  AOI21_X1 U6064 ( .B1(n5912), .B2(n4912), .A(n4911), .ZN(n4917) );
  OR2_X1 U6065 ( .A1(n5826), .A2(n4913), .ZN(n5307) );
  INV_X1 U6066 ( .A(n5307), .ZN(n4915) );
  OAI21_X1 U6067 ( .B1(n5826), .B2(n4914), .A(n5064), .ZN(n5878) );
  OAI21_X1 U6068 ( .B1(n4915), .B2(REIP_REG_5__SCAN_IN), .A(n5878), .ZN(n4916)
         );
  OAI211_X1 U6069 ( .C1(n4918), .C2(n5910), .A(n4917), .B(n4916), .ZN(U2822)
         );
  OAI22_X1 U6070 ( .A1(n6361), .A2(n5179), .B1(n4931), .B2(n6212), .ZN(n4921)
         );
  NOR2_X1 U6071 ( .A1(n4919), .A2(n4932), .ZN(n4920) );
  AOI211_X1 U6072 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n4936), .A(n4921), 
        .B(n4920), .ZN(n4922) );
  OAI21_X1 U6073 ( .B1(n4938), .B2(n6255), .A(n4922), .ZN(U3145) );
  OAI22_X1 U6074 ( .A1(n6337), .A2(n5179), .B1(n4931), .B2(n6201), .ZN(n4925)
         );
  NOR2_X1 U6075 ( .A1(n4923), .A2(n4932), .ZN(n4924) );
  AOI211_X1 U6076 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n4936), .A(n4925), 
        .B(n4924), .ZN(n4926) );
  OAI21_X1 U6077 ( .B1(n4938), .B2(n6240), .A(n4926), .ZN(U3141) );
  OAI22_X1 U6078 ( .A1(n6331), .A2(n5179), .B1(n4931), .B2(n6198), .ZN(n4929)
         );
  NOR2_X1 U6079 ( .A1(n4927), .A2(n4932), .ZN(n4928) );
  AOI211_X1 U6080 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n4936), .A(n4929), 
        .B(n4928), .ZN(n4930) );
  OAI21_X1 U6081 ( .B1(n4938), .B2(n6236), .A(n4930), .ZN(U3140) );
  OAI22_X1 U6082 ( .A1(n6355), .A2(n5179), .B1(n4931), .B2(n6294), .ZN(n4935)
         );
  NOR2_X1 U6083 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  AOI211_X1 U6084 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n4936), .A(n4935), 
        .B(n4934), .ZN(n4937) );
  OAI21_X1 U6085 ( .B1(n4938), .B2(n6251), .A(n4937), .ZN(U3144) );
  INV_X1 U6086 ( .A(n4947), .ZN(n4980) );
  NOR2_X1 U6087 ( .A1(n4980), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6185)
         );
  AOI22_X1 U6088 ( .A1(n4943), .A2(n6272), .B1(n6325), .B2(n6185), .ZN(n4977)
         );
  NOR2_X1 U6089 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4939), .ZN(n4974)
         );
  INV_X1 U6090 ( .A(n4971), .ZN(n4941) );
  OAI21_X1 U6091 ( .B1(n4942), .B2(n4941), .A(n4940), .ZN(n4945) );
  INV_X1 U6092 ( .A(n4943), .ZN(n4944) );
  NAND2_X1 U6093 ( .A1(n4945), .A2(n4944), .ZN(n4948) );
  OAI21_X1 U6094 ( .B1(n4947), .B2(n4986), .A(n4946), .ZN(n5149) );
  NOR2_X1 U6095 ( .A1(n6309), .A2(n5149), .ZN(n4985) );
  NAND2_X1 U6096 ( .A1(n4970), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4951) );
  OAI22_X1 U6097 ( .A1(n6349), .A2(n4972), .B1(n4971), .B2(n6207), .ZN(n4949)
         );
  AOI21_X1 U6098 ( .B1(n6344), .B2(n4974), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6099 ( .C1(n4977), .C2(n6248), .A(n4951), .B(n4950), .ZN(U3039)
         );
  NAND2_X1 U6100 ( .A1(n4970), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4954) );
  OAI22_X1 U6101 ( .A1(n6343), .A2(n4972), .B1(n4971), .B2(n6204), .ZN(n4952)
         );
  AOI21_X1 U6102 ( .B1(n6338), .B2(n4974), .A(n4952), .ZN(n4953) );
  OAI211_X1 U6103 ( .C1(n4977), .C2(n6244), .A(n4954), .B(n4953), .ZN(U3038)
         );
  NAND2_X1 U6104 ( .A1(n4970), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4957) );
  OAI22_X1 U6105 ( .A1(n6355), .A2(n4972), .B1(n4971), .B2(n6294), .ZN(n4955)
         );
  AOI21_X1 U6106 ( .B1(n6350), .B2(n4974), .A(n4955), .ZN(n4956) );
  OAI211_X1 U6107 ( .C1(n4977), .C2(n6251), .A(n4957), .B(n4956), .ZN(U3040)
         );
  NAND2_X1 U6108 ( .A1(n4970), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4960) );
  OAI22_X1 U6109 ( .A1(n6361), .A2(n4972), .B1(n4971), .B2(n6212), .ZN(n4958)
         );
  AOI21_X1 U6110 ( .B1(n6356), .B2(n4974), .A(n4958), .ZN(n4959) );
  OAI211_X1 U6111 ( .C1(n4977), .C2(n6255), .A(n4960), .B(n4959), .ZN(U3041)
         );
  NAND2_X1 U6112 ( .A1(n4970), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4963) );
  OAI22_X1 U6113 ( .A1(n6378), .A2(n4972), .B1(n4971), .B2(n6222), .ZN(n4961)
         );
  AOI21_X1 U6114 ( .B1(n6369), .B2(n4974), .A(n4961), .ZN(n4962) );
  OAI211_X1 U6115 ( .C1(n4977), .C2(n6266), .A(n4963), .B(n4962), .ZN(U3043)
         );
  NAND2_X1 U6116 ( .A1(n4970), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4966) );
  OAI22_X1 U6117 ( .A1(n6367), .A2(n4972), .B1(n4971), .B2(n6301), .ZN(n4964)
         );
  AOI21_X1 U6118 ( .B1(n6362), .B2(n4974), .A(n4964), .ZN(n4965) );
  OAI211_X1 U6119 ( .C1(n4977), .C2(n6258), .A(n4966), .B(n4965), .ZN(U3042)
         );
  NAND2_X1 U6120 ( .A1(n4970), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4969) );
  OAI22_X1 U6121 ( .A1(n6331), .A2(n4972), .B1(n4971), .B2(n6198), .ZN(n4967)
         );
  AOI21_X1 U6122 ( .B1(n6316), .B2(n4974), .A(n4967), .ZN(n4968) );
  OAI211_X1 U6123 ( .C1(n4977), .C2(n6236), .A(n4969), .B(n4968), .ZN(U3036)
         );
  NAND2_X1 U6124 ( .A1(n4970), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4976) );
  OAI22_X1 U6125 ( .A1(n6337), .A2(n4972), .B1(n4971), .B2(n6201), .ZN(n4973)
         );
  AOI21_X1 U6126 ( .B1(n6332), .B2(n4974), .A(n4973), .ZN(n4975) );
  OAI211_X1 U6127 ( .C1(n4977), .C2(n6240), .A(n4976), .B(n4975), .ZN(U3037)
         );
  NAND2_X1 U6128 ( .A1(n5009), .A2(n6307), .ZN(n4978) );
  AOI21_X1 U6129 ( .B1(n4978), .B2(STATEBS16_REG_SCAN_IN), .A(n6318), .ZN(
        n4983) );
  AND2_X1 U6130 ( .A1(n4979), .A2(n4437), .ZN(n6275) );
  NOR2_X1 U6131 ( .A1(n4980), .A2(n6390), .ZN(n5148) );
  AOI22_X1 U6132 ( .A1(n4983), .A2(n6275), .B1(n6325), .B2(n5148), .ZN(n5014)
         );
  INV_X1 U6133 ( .A(n6275), .ZN(n4982) );
  NAND3_X1 U6134 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6665), .ZN(n6280) );
  NOR2_X1 U6135 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6280), .ZN(n5011)
         );
  INV_X1 U6136 ( .A(n5011), .ZN(n4981) );
  AOI22_X1 U6137 ( .A1(n4983), .A2(n4982), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4981), .ZN(n4984) );
  NAND2_X1 U6138 ( .A1(n5008), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4989)
         );
  OAI22_X1 U6139 ( .A1(n5009), .A2(n6331), .B1(n6307), .B2(n6198), .ZN(n4987)
         );
  AOI21_X1 U6140 ( .B1(n6316), .B2(n5011), .A(n4987), .ZN(n4988) );
  OAI211_X1 U6141 ( .C1(n5014), .C2(n6236), .A(n4989), .B(n4988), .ZN(U3100)
         );
  NAND2_X1 U6142 ( .A1(n5008), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4992)
         );
  OAI22_X1 U6143 ( .A1(n5009), .A2(n6349), .B1(n6307), .B2(n6207), .ZN(n4990)
         );
  AOI21_X1 U6144 ( .B1(n6344), .B2(n5011), .A(n4990), .ZN(n4991) );
  OAI211_X1 U6145 ( .C1(n5014), .C2(n6248), .A(n4992), .B(n4991), .ZN(U3103)
         );
  NAND2_X1 U6146 ( .A1(n5008), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4995)
         );
  OAI22_X1 U6147 ( .A1(n5009), .A2(n6355), .B1(n6307), .B2(n6294), .ZN(n4993)
         );
  AOI21_X1 U6148 ( .B1(n6350), .B2(n5011), .A(n4993), .ZN(n4994) );
  OAI211_X1 U6149 ( .C1(n5014), .C2(n6251), .A(n4995), .B(n4994), .ZN(U3104)
         );
  NAND2_X1 U6150 ( .A1(n5008), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4998)
         );
  OAI22_X1 U6151 ( .A1(n5009), .A2(n6367), .B1(n6307), .B2(n6301), .ZN(n4996)
         );
  AOI21_X1 U6152 ( .B1(n6362), .B2(n5011), .A(n4996), .ZN(n4997) );
  OAI211_X1 U6153 ( .C1(n5014), .C2(n6258), .A(n4998), .B(n4997), .ZN(U3106)
         );
  NAND2_X1 U6154 ( .A1(n5008), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5001)
         );
  OAI22_X1 U6155 ( .A1(n5009), .A2(n6361), .B1(n6307), .B2(n6212), .ZN(n4999)
         );
  AOI21_X1 U6156 ( .B1(n6356), .B2(n5011), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6157 ( .C1(n5014), .C2(n6255), .A(n5001), .B(n5000), .ZN(U3105)
         );
  NAND2_X1 U6158 ( .A1(n5008), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5004)
         );
  OAI22_X1 U6159 ( .A1(n5009), .A2(n6378), .B1(n6307), .B2(n6222), .ZN(n5002)
         );
  AOI21_X1 U6160 ( .B1(n6369), .B2(n5011), .A(n5002), .ZN(n5003) );
  OAI211_X1 U6161 ( .C1(n5014), .C2(n6266), .A(n5004), .B(n5003), .ZN(U3107)
         );
  NAND2_X1 U6162 ( .A1(n5008), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5007)
         );
  OAI22_X1 U6163 ( .A1(n5009), .A2(n6337), .B1(n6307), .B2(n6201), .ZN(n5005)
         );
  AOI21_X1 U6164 ( .B1(n6332), .B2(n5011), .A(n5005), .ZN(n5006) );
  OAI211_X1 U6165 ( .C1(n5014), .C2(n6240), .A(n5007), .B(n5006), .ZN(U3101)
         );
  NAND2_X1 U6166 ( .A1(n5008), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5013)
         );
  OAI22_X1 U6167 ( .A1(n5009), .A2(n6343), .B1(n6307), .B2(n6204), .ZN(n5010)
         );
  AOI21_X1 U6168 ( .B1(n6338), .B2(n5011), .A(n5010), .ZN(n5012) );
  OAI211_X1 U6169 ( .C1(n5014), .C2(n6244), .A(n5013), .B(n5012), .ZN(U3102)
         );
  OAI21_X1 U6170 ( .B1(n5017), .B2(n5016), .A(n5015), .ZN(n6118) );
  INV_X1 U6171 ( .A(n5018), .ZN(n5022) );
  AOI22_X1 U6172 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6171), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5019) );
  OAI21_X1 U6173 ( .B1(n5020), .B2(n6090), .A(n5019), .ZN(n5021) );
  AOI21_X1 U6174 ( .B1(n5022), .B2(n6075), .A(n5021), .ZN(n5023) );
  OAI21_X1 U6175 ( .B1(n6118), .B2(n6065), .A(n5023), .ZN(U2978) );
  OAI21_X1 U6176 ( .B1(n5826), .B2(REIP_REG_1__SCAN_IN), .A(n5064), .ZN(n5902)
         );
  NAND2_X1 U6177 ( .A1(n6459), .A2(REIP_REG_1__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U6178 ( .A1(n5906), .A2(n6170), .B1(n5903), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5026) );
  INV_X1 U6179 ( .A(n6089), .ZN(n5024) );
  AOI22_X1 U6180 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n5905), .B1(n5912), 
        .B2(n5024), .ZN(n5025) );
  OAI211_X1 U6181 ( .C1(n5826), .C2(n5027), .A(n5026), .B(n5025), .ZN(n5032)
         );
  INV_X1 U6182 ( .A(n5028), .ZN(n5030) );
  NOR2_X1 U6183 ( .A1(n5030), .A2(n5029), .ZN(n5904) );
  INV_X1 U6184 ( .A(n5904), .ZN(n5323) );
  OAI22_X1 U6185 ( .A1(n5323), .A2(n4470), .B1(n5910), .B2(n6081), .ZN(n5031)
         );
  AOI211_X1 U6186 ( .C1(REIP_REG_2__SCAN_IN), .C2(n5902), .A(n5032), .B(n5031), 
        .ZN(n5033) );
  INV_X1 U6187 ( .A(n5033), .ZN(U2825) );
  OAI21_X1 U6188 ( .B1(n3541), .B2(n3540), .A(n5035), .ZN(n5849) );
  AOI22_X1 U6189 ( .A1(n5134), .A2(DATAI_10_), .B1(n5944), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5036) );
  OAI21_X1 U6190 ( .B1(n5849), .B2(n5669), .A(n5036), .ZN(U2881) );
  XNOR2_X1 U6191 ( .A(n5861), .B(n5832), .ZN(n5846) );
  OAI222_X1 U6192 ( .A1(n5390), .A2(n5849), .B1(n5037), .B2(n5934), .C1(n5925), 
        .C2(n5846), .ZN(U2849) );
  INV_X1 U6193 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6006) );
  AOI22_X1 U6194 ( .A1(n5966), .A2(UWORD_REG_14__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5038) );
  OAI21_X1 U6195 ( .B1(n6006), .B2(n5050), .A(n5038), .ZN(U2893) );
  INV_X1 U6196 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5989) );
  AOI22_X1 U6197 ( .A1(n5966), .A2(UWORD_REG_8__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5039) );
  OAI21_X1 U6198 ( .B1(n5989), .B2(n5050), .A(n5039), .ZN(U2899) );
  AOI22_X1 U6199 ( .A1(n5966), .A2(UWORD_REG_0__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5040) );
  OAI21_X1 U6200 ( .B1(n3635), .B2(n5050), .A(n5040), .ZN(U2907) );
  INV_X1 U6201 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5980) );
  AOI22_X1 U6202 ( .A1(n5966), .A2(UWORD_REG_5__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5041) );
  OAI21_X1 U6203 ( .B1(n5980), .B2(n5050), .A(n5041), .ZN(U2902) );
  AOI22_X1 U6204 ( .A1(n5966), .A2(UWORD_REG_4__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5042) );
  OAI21_X1 U6205 ( .B1(n3709), .B2(n5050), .A(n5042), .ZN(U2903) );
  INV_X1 U6206 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6567) );
  AOI22_X1 U6207 ( .A1(n5966), .A2(UWORD_REG_12__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5043) );
  OAI21_X1 U6208 ( .B1(n6567), .B2(n5050), .A(n5043), .ZN(U2895) );
  AOI22_X1 U6209 ( .A1(n5966), .A2(UWORD_REG_10__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5044) );
  OAI21_X1 U6210 ( .B1(n3832), .B2(n5050), .A(n5044), .ZN(U2897) );
  INV_X1 U6211 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5986) );
  AOI22_X1 U6212 ( .A1(n5966), .A2(UWORD_REG_7__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5045) );
  OAI21_X1 U6213 ( .B1(n5986), .B2(n5050), .A(n5045), .ZN(U2900) );
  INV_X1 U6214 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5983) );
  AOI22_X1 U6215 ( .A1(n5966), .A2(UWORD_REG_6__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5046) );
  OAI21_X1 U6216 ( .B1(n5983), .B2(n5050), .A(n5046), .ZN(U2901) );
  INV_X1 U6217 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5975) );
  AOI22_X1 U6218 ( .A1(n5956), .A2(UWORD_REG_2__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5047) );
  OAI21_X1 U6219 ( .B1(n5975), .B2(n5050), .A(n5047), .ZN(U2905) );
  AOI22_X1 U6220 ( .A1(n5956), .A2(UWORD_REG_1__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5048) );
  OAI21_X1 U6221 ( .B1(n3655), .B2(n5050), .A(n5048), .ZN(U2906) );
  INV_X1 U6222 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5977) );
  AOI22_X1 U6223 ( .A1(n5956), .A2(UWORD_REG_3__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5049) );
  OAI21_X1 U6224 ( .B1(n5977), .B2(n5050), .A(n5049), .ZN(U2904) );
  AOI21_X1 U6225 ( .B1(n5052), .B2(n5035), .A(n5051), .ZN(n6060) );
  INV_X1 U6226 ( .A(n6060), .ZN(n5054) );
  AOI22_X1 U6227 ( .A1(n5134), .A2(DATAI_11_), .B1(n5944), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5053) );
  OAI21_X1 U6228 ( .B1(n5054), .B2(n5669), .A(n5053), .ZN(U2880) );
  XNOR2_X1 U6229 ( .A(n2967), .B(n6103), .ZN(n5056) );
  XNOR2_X1 U6230 ( .A(n5055), .B(n5056), .ZN(n6114) );
  NAND2_X1 U6231 ( .A1(n6114), .A2(n6085), .ZN(n5060) );
  INV_X1 U6232 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U6233 ( .A1(n6092), .A2(n5057), .ZN(n6111) );
  AND2_X1 U6234 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5058)
         );
  AOI211_X1 U6235 ( .C1(n5867), .C2(n6059), .A(n6111), .B(n5058), .ZN(n5059)
         );
  OAI211_X1 U6236 ( .C1(n6063), .C2(n5926), .A(n5060), .B(n5059), .ZN(U2977)
         );
  XOR2_X1 U6237 ( .A(n5061), .B(n5051), .Z(n5117) );
  INV_X1 U6238 ( .A(n5117), .ZN(n5082) );
  AOI21_X1 U6239 ( .B1(n5062), .B2(n5833), .A(n2999), .ZN(n5111) );
  AOI22_X1 U6240 ( .A1(n5930), .A2(n5111), .B1(EBX_REG_12__SCAN_IN), .B2(n5386), .ZN(n5063) );
  OAI21_X1 U6241 ( .B1(n5082), .B2(n5390), .A(n5063), .ZN(U2847) );
  OAI21_X1 U6242 ( .B1(n5826), .B2(n5836), .A(n5064), .ZN(n5842) );
  INV_X1 U6243 ( .A(n5842), .ZN(n5825) );
  INV_X1 U6244 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6245 ( .A1(n5117), .A2(n5879), .ZN(n5073) );
  INV_X1 U6246 ( .A(n5115), .ZN(n5065) );
  NAND2_X1 U6247 ( .A1(n5912), .A2(n5065), .ZN(n5067) );
  NAND2_X1 U6248 ( .A1(n5905), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5066)
         );
  NAND3_X1 U6249 ( .A1(n5067), .A2(n5066), .A3(n5301), .ZN(n5071) );
  NAND2_X1 U6250 ( .A1(n5836), .A2(n5095), .ZN(n5069) );
  INV_X1 U6251 ( .A(n5111), .ZN(n5068) );
  OAI22_X1 U6252 ( .A1(n5826), .A2(n5069), .B1(n5874), .B2(n5068), .ZN(n5070)
         );
  AOI211_X1 U6253 ( .C1(n5903), .C2(EBX_REG_12__SCAN_IN), .A(n5071), .B(n5070), 
        .ZN(n5072) );
  OAI211_X1 U6254 ( .C1(n5825), .C2(n5095), .A(n5073), .B(n5072), .ZN(U2815)
         );
  NAND2_X1 U6255 ( .A1(n6054), .A2(n5075), .ZN(n5076) );
  XNOR2_X1 U6256 ( .A(n5074), .B(n5076), .ZN(n6107) );
  NAND2_X1 U6257 ( .A1(n6107), .A2(n6085), .ZN(n5080) );
  INV_X1 U6258 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U6259 ( .A1(n6092), .A2(n5077), .ZN(n6104) );
  NOR2_X1 U6260 ( .A1(n6090), .A2(n5850), .ZN(n5078) );
  AOI211_X1 U6261 ( .C1(n6080), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6104), 
        .B(n5078), .ZN(n5079) );
  OAI211_X1 U6262 ( .C1(n6063), .C2(n5849), .A(n5080), .B(n5079), .ZN(U2976)
         );
  INV_X1 U6263 ( .A(DATAI_12_), .ZN(n5998) );
  OAI222_X1 U6264 ( .A1(n5083), .A2(n5998), .B1(n5669), .B2(n5082), .C1(n5081), 
        .C2(n5392), .ZN(U2879) );
  INV_X1 U6265 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6266 ( .A1(n2991), .A2(n5085), .ZN(n5087) );
  INV_X1 U6267 ( .A(n5919), .ZN(n5089) );
  AOI22_X1 U6268 ( .A1(n5134), .A2(DATAI_13_), .B1(n5944), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5088) );
  OAI21_X1 U6269 ( .B1(n5089), .B2(n5669), .A(n5088), .ZN(U2878) );
  INV_X1 U6270 ( .A(n5091), .ZN(n5092) );
  NOR2_X1 U6271 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  XNOR2_X1 U6272 ( .A(n5090), .B(n5094), .ZN(n5119) );
  NOR2_X1 U6273 ( .A1(n6092), .A2(n5095), .ZN(n5113) );
  AOI22_X1 U6274 ( .A1(n5099), .A2(n5097), .B1(n6172), .B2(n5096), .ZN(n5098)
         );
  INV_X1 U6275 ( .A(n5098), .ZN(n5595) );
  AOI21_X1 U6276 ( .B1(n5100), .B2(n5099), .A(n5595), .ZN(n6091) );
  OAI21_X1 U6277 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5592), .ZN(n5109) );
  AOI21_X1 U6278 ( .B1(n5103), .B2(n5102), .A(n5101), .ZN(n5104) );
  INV_X1 U6279 ( .A(n5104), .ZN(n5105) );
  AOI21_X1 U6280 ( .B1(n6102), .B2(n6172), .A(n5105), .ZN(n6135) );
  INV_X1 U6281 ( .A(n6135), .ZN(n5106) );
  OAI22_X1 U6282 ( .A1(n5107), .A2(n5106), .B1(n5586), .B2(n5105), .ZN(n6101)
         );
  OAI22_X1 U6283 ( .A1(n6091), .A2(n5109), .B1(n5108), .B2(n6101), .ZN(n5110)
         );
  AOI211_X1 U6284 ( .C1(n6169), .C2(n5111), .A(n5113), .B(n5110), .ZN(n5112)
         );
  OAI21_X1 U6285 ( .B1(n5119), .B2(n6095), .A(n5112), .ZN(U3006) );
  AOI21_X1 U6286 ( .B1(n6080), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5113), 
        .ZN(n5114) );
  OAI21_X1 U6287 ( .B1(n5115), .B2(n6090), .A(n5114), .ZN(n5116) );
  AOI21_X1 U6288 ( .B1(n5117), .B2(n6075), .A(n5116), .ZN(n5118) );
  OAI21_X1 U6289 ( .B1(n5119), .B2(n6065), .A(n5118), .ZN(U2974) );
  OAI21_X1 U6290 ( .B1(n5121), .B2(n5123), .A(n5122), .ZN(n5814) );
  AOI22_X1 U6291 ( .A1(n5134), .A2(DATAI_14_), .B1(n5944), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5124) );
  OAI21_X1 U6292 ( .B1(n5814), .B2(n5669), .A(n5124), .ZN(U2877) );
  OR2_X1 U6293 ( .A1(n5763), .A2(n5125), .ZN(n5126) );
  NAND2_X1 U6294 ( .A1(n5131), .A2(n5126), .ZN(n5811) );
  OAI222_X1 U6295 ( .A1(n5811), .A2(n5925), .B1(n5934), .B2(n4077), .C1(n5814), 
        .C2(n5390), .ZN(U2845) );
  NAND2_X1 U6296 ( .A1(n5122), .A2(n5128), .ZN(n5129) );
  NAND2_X1 U6297 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  AND2_X1 U6298 ( .A1(n5283), .A2(n5132), .ZN(n5752) );
  AOI22_X1 U6299 ( .A1(n5930), .A2(n5752), .B1(EBX_REG_15__SCAN_IN), .B2(n5386), .ZN(n5133) );
  OAI21_X1 U6300 ( .B1(n5300), .B2(n5390), .A(n5133), .ZN(U2844) );
  AOI22_X1 U6301 ( .A1(n5134), .A2(DATAI_15_), .B1(n5944), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5135) );
  OAI21_X1 U6302 ( .B1(n5300), .B2(n5669), .A(n5135), .ZN(U2876) );
  INV_X1 U6303 ( .A(n5136), .ZN(n5147) );
  INV_X1 U6304 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5138) );
  AOI22_X1 U6305 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5138), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5137), .ZN(n5188) );
  NOR2_X1 U6306 ( .A1(n6418), .A2(n5189), .ZN(n5144) );
  NOR3_X1 U6307 ( .A1(n5139), .A2(n4799), .A3(n4436), .ZN(n5140) );
  AOI21_X1 U6308 ( .B1(n5141), .B2(n3112), .A(n5140), .ZN(n5142) );
  OAI21_X1 U6309 ( .B1(n2979), .B2(n5143), .A(n5142), .ZN(n6381) );
  AOI222_X1 U6310 ( .A1(n5186), .A2(n5145), .B1(n5188), .B2(n5144), .C1(n6381), 
        .C2(n5194), .ZN(n5146) );
  INV_X1 U6311 ( .A(n5775), .ZN(n5196) );
  OAI22_X1 U6312 ( .A1(n5147), .A2(n3112), .B1(n5146), .B2(n5196), .ZN(U3460)
         );
  NOR2_X1 U6313 ( .A1(n6191), .A2(n6318), .ZN(n6186) );
  AOI22_X1 U6314 ( .A1(n6186), .A2(n4437), .B1(n6309), .B2(n5148), .ZN(n5185)
         );
  NOR2_X1 U6315 ( .A1(n6325), .A2(n5149), .ZN(n6195) );
  NOR2_X1 U6316 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5150), .ZN(n5182)
         );
  INV_X1 U6317 ( .A(n5182), .ZN(n5151) );
  AOI21_X1 U6318 ( .B1(n5151), .B2(STATE2_REG_3__SCAN_IN), .A(n6390), .ZN(
        n5156) );
  NOR3_X1 U6319 ( .A1(n5153), .A2(n5152), .A3(n6318), .ZN(n5154) );
  OAI21_X1 U6320 ( .B1(n5154), .B2(n6322), .A(n6191), .ZN(n5155) );
  NAND3_X1 U6321 ( .A1(n6195), .A2(n5156), .A3(n5155), .ZN(n5178) );
  NAND2_X1 U6322 ( .A1(n5178), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5159)
         );
  OAI22_X1 U6323 ( .A1(n5180), .A2(n6378), .B1(n6222), .B2(n5179), .ZN(n5157)
         );
  AOI21_X1 U6324 ( .B1(n6369), .B2(n5182), .A(n5157), .ZN(n5158) );
  OAI211_X1 U6325 ( .C1(n5185), .C2(n6266), .A(n5159), .B(n5158), .ZN(U3139)
         );
  NAND2_X1 U6326 ( .A1(n5178), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5162)
         );
  OAI22_X1 U6327 ( .A1(n5180), .A2(n6367), .B1(n6301), .B2(n5179), .ZN(n5160)
         );
  AOI21_X1 U6328 ( .B1(n6362), .B2(n5182), .A(n5160), .ZN(n5161) );
  OAI211_X1 U6329 ( .C1(n5185), .C2(n6258), .A(n5162), .B(n5161), .ZN(U3138)
         );
  NAND2_X1 U6330 ( .A1(n5178), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5165)
         );
  OAI22_X1 U6331 ( .A1(n5180), .A2(n6361), .B1(n6212), .B2(n5179), .ZN(n5163)
         );
  AOI21_X1 U6332 ( .B1(n6356), .B2(n5182), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6333 ( .C1(n5185), .C2(n6255), .A(n5165), .B(n5164), .ZN(U3137)
         );
  NAND2_X1 U6334 ( .A1(n5178), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5168)
         );
  OAI22_X1 U6335 ( .A1(n5180), .A2(n6355), .B1(n6294), .B2(n5179), .ZN(n5166)
         );
  AOI21_X1 U6336 ( .B1(n6350), .B2(n5182), .A(n5166), .ZN(n5167) );
  OAI211_X1 U6337 ( .C1(n5185), .C2(n6251), .A(n5168), .B(n5167), .ZN(U3136)
         );
  NAND2_X1 U6338 ( .A1(n5178), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5171)
         );
  OAI22_X1 U6339 ( .A1(n5180), .A2(n6349), .B1(n6207), .B2(n5179), .ZN(n5169)
         );
  AOI21_X1 U6340 ( .B1(n6344), .B2(n5182), .A(n5169), .ZN(n5170) );
  OAI211_X1 U6341 ( .C1(n5185), .C2(n6248), .A(n5171), .B(n5170), .ZN(U3135)
         );
  NAND2_X1 U6342 ( .A1(n5178), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5174)
         );
  OAI22_X1 U6343 ( .A1(n5180), .A2(n6343), .B1(n6204), .B2(n5179), .ZN(n5172)
         );
  AOI21_X1 U6344 ( .B1(n6338), .B2(n5182), .A(n5172), .ZN(n5173) );
  OAI211_X1 U6345 ( .C1(n5185), .C2(n6244), .A(n5174), .B(n5173), .ZN(U3134)
         );
  NAND2_X1 U6346 ( .A1(n5178), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5177)
         );
  OAI22_X1 U6347 ( .A1(n5180), .A2(n6337), .B1(n6201), .B2(n5179), .ZN(n5175)
         );
  AOI21_X1 U6348 ( .B1(n6332), .B2(n5182), .A(n5175), .ZN(n5176) );
  OAI211_X1 U6349 ( .C1(n5185), .C2(n6240), .A(n5177), .B(n5176), .ZN(U3133)
         );
  NAND2_X1 U6350 ( .A1(n5178), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5184)
         );
  OAI22_X1 U6351 ( .A1(n5180), .A2(n6331), .B1(n6198), .B2(n5179), .ZN(n5181)
         );
  AOI21_X1 U6352 ( .B1(n6316), .B2(n5182), .A(n5181), .ZN(n5183) );
  OAI211_X1 U6353 ( .C1(n5185), .C2(n6236), .A(n5184), .B(n5183), .ZN(U3132)
         );
  AOI21_X1 U6354 ( .B1(n5191), .B2(n5186), .A(n5196), .ZN(n5198) );
  INV_X1 U6355 ( .A(n5187), .ZN(n5195) );
  NOR3_X1 U6356 ( .A1(n6418), .A2(n5189), .A3(n5188), .ZN(n5193) );
  NOR3_X1 U6357 ( .A1(n5191), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5190), 
        .ZN(n5192) );
  AOI211_X1 U6358 ( .C1(n5195), .C2(n5194), .A(n5193), .B(n5192), .ZN(n5197)
         );
  OAI22_X1 U6359 ( .A1(n5198), .A2(n3110), .B1(n5197), .B2(n5196), .ZN(U3459)
         );
  AND2_X1 U6360 ( .A1(n5242), .A2(n5200), .ZN(n5201) );
  NOR2_X1 U6361 ( .A1(n5202), .A2(n5201), .ZN(n5215) );
  AOI22_X1 U6362 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5903), .B1(n5203), .B2(n5912), .ZN(n5204) );
  OAI21_X1 U6363 ( .B1(n5205), .B2(n5889), .A(n5204), .ZN(n5206) );
  AOI21_X1 U6364 ( .B1(n5215), .B2(n5906), .A(n5206), .ZN(n5207) );
  OAI21_X1 U6365 ( .B1(n5219), .B2(REIP_REG_29__SCAN_IN), .A(n5207), .ZN(n5208) );
  AOI21_X1 U6366 ( .B1(n5248), .B2(REIP_REG_29__SCAN_IN), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6367 ( .B1(n5199), .B2(n5659), .A(n5209), .ZN(U2798) );
  AOI22_X1 U6368 ( .A1(n5941), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5944), .ZN(n5214) );
  AND2_X1 U6369 ( .A1(n3222), .A2(n5211), .ZN(n5212) );
  NAND2_X1 U6370 ( .A1(n5945), .A2(DATAI_13_), .ZN(n5213) );
  OAI211_X1 U6371 ( .C1(n5199), .C2(n5669), .A(n5214), .B(n5213), .ZN(U2862)
         );
  INV_X1 U6372 ( .A(n5215), .ZN(n5513) );
  OAI222_X1 U6373 ( .A1(n5390), .A2(n5199), .B1(n5216), .B2(n5934), .C1(n5513), 
        .C2(n5925), .ZN(U2830) );
  INV_X1 U6374 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6504) );
  INV_X1 U6375 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5218) );
  OAI21_X1 U6376 ( .B1(n5219), .B2(n6504), .A(n5218), .ZN(n5231) );
  INV_X1 U6377 ( .A(n5221), .ZN(n5220) );
  OAI21_X1 U6378 ( .B1(n5224), .B2(n5242), .A(n5220), .ZN(n5225) );
  INV_X1 U6379 ( .A(n5242), .ZN(n5222) );
  OAI21_X1 U6380 ( .B1(n5222), .B2(n4080), .A(n5221), .ZN(n5223) );
  OAI22_X1 U6381 ( .A1(n5226), .A2(n5225), .B1(n5224), .B2(n5223), .ZN(n5502)
         );
  AOI22_X1 U6382 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5905), .B1(n5912), 
        .B2(n5227), .ZN(n5229) );
  NAND2_X1 U6383 ( .A1(n5903), .A2(EBX_REG_30__SCAN_IN), .ZN(n5228) );
  OAI211_X1 U6384 ( .C1(n5502), .C2(n5874), .A(n5229), .B(n5228), .ZN(n5230)
         );
  AOI21_X1 U6385 ( .B1(n5232), .B2(n5231), .A(n5230), .ZN(n5233) );
  OAI21_X1 U6386 ( .B1(n5217), .B2(n5659), .A(n5233), .ZN(U2797) );
  AOI22_X1 U6387 ( .A1(n5941), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5944), .ZN(n5235) );
  NAND2_X1 U6388 ( .A1(n5945), .A2(DATAI_14_), .ZN(n5234) );
  OAI211_X1 U6389 ( .C1(n5217), .C2(n5669), .A(n5235), .B(n5234), .ZN(U2861)
         );
  INV_X1 U6390 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5236) );
  OAI222_X1 U6391 ( .A1(n5390), .A2(n5217), .B1(n5236), .B2(n5934), .C1(n5502), 
        .C2(n5925), .ZN(U2829) );
  AOI21_X1 U6392 ( .B1(n5239), .B2(n5237), .A(n5238), .ZN(n5417) );
  INV_X1 U6393 ( .A(n5417), .ZN(n5399) );
  NAND2_X1 U6394 ( .A1(n5254), .A2(n5240), .ZN(n5241) );
  NAND2_X1 U6395 ( .A1(n5242), .A2(n5241), .ZN(n5521) );
  INV_X1 U6396 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6588) );
  NAND3_X1 U6397 ( .A1(n5259), .A2(REIP_REG_27__SCAN_IN), .A3(n6588), .ZN(
        n5246) );
  INV_X1 U6398 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5243) );
  OAI22_X1 U6399 ( .A1(n5243), .A2(n5889), .B1(n5883), .B2(n5415), .ZN(n5244)
         );
  AOI21_X1 U6400 ( .B1(n5903), .B2(EBX_REG_28__SCAN_IN), .A(n5244), .ZN(n5245)
         );
  OAI211_X1 U6401 ( .C1(n5874), .C2(n5521), .A(n5246), .B(n5245), .ZN(n5247)
         );
  AOI21_X1 U6402 ( .B1(n5248), .B2(REIP_REG_28__SCAN_IN), .A(n5247), .ZN(n5249) );
  OAI21_X1 U6403 ( .B1(n5399), .B2(n5659), .A(n5249), .ZN(U2799) );
  INV_X1 U6404 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6498) );
  OR2_X1 U6405 ( .A1(n5339), .A2(n5252), .ZN(n5253) );
  NAND2_X1 U6406 ( .A1(n5254), .A2(n5253), .ZN(n5531) );
  INV_X1 U6407 ( .A(n5425), .ZN(n5255) );
  OAI22_X1 U6408 ( .A1(n5531), .A2(n5874), .B1(n5255), .B2(n5883), .ZN(n5258)
         );
  AOI22_X1 U6409 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5903), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5905), .ZN(n5256) );
  OAI21_X1 U6410 ( .B1(n5615), .B2(n6498), .A(n5256), .ZN(n5257) );
  AOI211_X1 U6411 ( .C1(n5259), .C2(n6498), .A(n5258), .B(n5257), .ZN(n5260)
         );
  OAI21_X1 U6412 ( .B1(n5423), .B2(n5659), .A(n5260), .ZN(U2800) );
  INV_X1 U6413 ( .A(n2988), .ZN(n5264) );
  OAI21_X1 U6414 ( .B1(n5261), .B2(n5467), .A(n5262), .ZN(n5263) );
  NAND2_X1 U6415 ( .A1(n5264), .A2(n5263), .ZN(n5676) );
  INV_X1 U6416 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6488) );
  NOR2_X1 U6417 ( .A1(n6488), .A2(n5641), .ZN(n5630) );
  INV_X1 U6418 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6492) );
  OAI21_X1 U6419 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5641), .A(n5640), .ZN(n5267) );
  AOI22_X1 U6420 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5903), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5905), .ZN(n5265) );
  OAI21_X1 U6421 ( .B1(n5461), .B2(n5883), .A(n5265), .ZN(n5266) );
  AOI221_X1 U6422 ( .B1(n5630), .B2(n6492), .C1(n5267), .C2(
        REIP_REG_22__SCAN_IN), .A(n5266), .ZN(n5272) );
  INV_X1 U6423 ( .A(n5268), .ZN(n5270) );
  INV_X1 U6424 ( .A(n5575), .ZN(n5269) );
  AOI21_X1 U6425 ( .B1(n5270), .B2(n5269), .A(n5354), .ZN(n5567) );
  NAND2_X1 U6426 ( .A1(n5567), .A2(n5906), .ZN(n5271) );
  OAI211_X1 U6427 ( .C1(n5676), .C2(n5659), .A(n5272), .B(n5271), .ZN(U2805)
         );
  XOR2_X1 U6428 ( .A(n5273), .B(n2980), .Z(n5938) );
  INV_X1 U6429 ( .A(n5938), .ZN(n5388) );
  NAND2_X1 U6430 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5287) );
  INV_X1 U6431 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U6432 ( .B1(n5287), .B2(n5296), .A(n6667), .ZN(n5276) );
  OAI22_X1 U6433 ( .A1(n5274), .A2(n5864), .B1(n6631), .B2(n5889), .ZN(n5275)
         );
  AOI211_X1 U6434 ( .C1(n5277), .C2(n5276), .A(n5892), .B(n5275), .ZN(n5280)
         );
  AOI21_X1 U6435 ( .B1(n5278), .B2(n5285), .A(n5382), .ZN(n5737) );
  AOI22_X1 U6436 ( .A1(n5906), .A2(n5737), .B1(n5703), .B2(n5912), .ZN(n5279)
         );
  OAI211_X1 U6437 ( .C1(n5388), .C2(n5659), .A(n5280), .B(n5279), .ZN(U2810)
         );
  AOI21_X1 U6438 ( .B1(n5281), .B2(n5127), .A(n2980), .ZN(n5943) );
  INV_X1 U6439 ( .A(n5943), .ZN(n5391) );
  NAND2_X1 U6440 ( .A1(n5283), .A2(n5282), .ZN(n5284) );
  NAND2_X1 U6441 ( .A1(n5285), .A2(n5284), .ZN(n5744) );
  INV_X1 U6442 ( .A(n5744), .ZN(n5292) );
  NAND2_X1 U6443 ( .A1(n5912), .A2(n5485), .ZN(n5286) );
  OAI211_X1 U6444 ( .C1(n5889), .C2(n6637), .A(n5286), .B(n5301), .ZN(n5291)
         );
  INV_X1 U6445 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5751) );
  INV_X1 U6446 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6481) );
  AOI21_X1 U6447 ( .B1(n5751), .B2(n6481), .A(n5296), .ZN(n5288) );
  AOI22_X1 U6448 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5903), .B1(n5288), .B2(n5287), .ZN(n5289) );
  OAI21_X1 U6449 ( .B1(n5819), .B2(n5751), .A(n5289), .ZN(n5290) );
  AOI211_X1 U6450 ( .C1(n5292), .C2(n5906), .A(n5291), .B(n5290), .ZN(n5293)
         );
  OAI21_X1 U6451 ( .B1(n5391), .B2(n5659), .A(n5293), .ZN(U2811) );
  INV_X1 U6452 ( .A(n5752), .ZN(n5294) );
  OAI22_X1 U6453 ( .A1(n5491), .A2(n5883), .B1(n5874), .B2(n5294), .ZN(n5298)
         );
  AOI21_X1 U6454 ( .B1(n5905), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5892), 
        .ZN(n5295) );
  OAI221_X1 U6455 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5296), .C1(n6481), .C2(
        n5819), .A(n5295), .ZN(n5297) );
  AOI211_X1 U6456 ( .C1(EBX_REG_15__SCAN_IN), .C2(n5903), .A(n5298), .B(n5297), 
        .ZN(n5299) );
  OAI21_X1 U6457 ( .B1(n5300), .B2(n5659), .A(n5299), .ZN(U2812) );
  AOI22_X1 U6458 ( .A1(n5906), .A2(n6128), .B1(n5903), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5302) );
  OAI211_X1 U6459 ( .C1(n5889), .C2(n4897), .A(n5302), .B(n5301), .ZN(n5306)
         );
  INV_X1 U6460 ( .A(n5303), .ZN(n5304) );
  NOR2_X1 U6461 ( .A1(n5883), .A2(n5304), .ZN(n5305) );
  AOI211_X1 U6462 ( .C1(REIP_REG_7__SCAN_IN), .C2(n5878), .A(n5306), .B(n5305), 
        .ZN(n5310) );
  NOR2_X1 U6463 ( .A1(n5307), .A2(n6465), .ZN(n5877) );
  INV_X1 U6464 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6467) );
  INV_X1 U6465 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6469) );
  AOI22_X1 U6466 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .B1(
        n6467), .B2(n6469), .ZN(n5308) );
  NAND2_X1 U6467 ( .A1(n5877), .A2(n5308), .ZN(n5309) );
  OAI211_X1 U6468 ( .C1(n5311), .C2(n5659), .A(n5310), .B(n5309), .ZN(U2820)
         );
  NOR2_X1 U6469 ( .A1(n5889), .A2(n5312), .ZN(n5315) );
  AOI22_X1 U6470 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5903), .B1(n5888), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5313) );
  OAI21_X1 U6471 ( .B1(n5883), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5313), 
        .ZN(n5314) );
  AOI211_X1 U6472 ( .C1(n5904), .C2(n5316), .A(n5315), .B(n5314), .ZN(n5319)
         );
  INV_X1 U6473 ( .A(n5826), .ZN(n5897) );
  AOI22_X1 U6474 ( .A1(n5897), .A2(n6584), .B1(n5906), .B2(n5317), .ZN(n5318)
         );
  OAI211_X1 U6475 ( .C1(n5910), .C2(n5320), .A(n5319), .B(n5318), .ZN(U2826)
         );
  OAI22_X1 U6476 ( .A1(n5323), .A2(n5322), .B1(n5321), .B2(n5864), .ZN(n5324)
         );
  AOI21_X1 U6477 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5886), .A(n5324), .ZN(n5328)
         );
  NAND2_X1 U6478 ( .A1(n5889), .A2(n5883), .ZN(n5326) );
  AOI22_X1 U6479 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5326), .B1(n5906), 
        .B2(n5325), .ZN(n5327) );
  OAI211_X1 U6480 ( .C1(n5910), .C2(n5329), .A(n5328), .B(n5327), .ZN(U2827)
         );
  INV_X1 U6481 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5330) );
  OAI22_X1 U6482 ( .A1(n5331), .A2(n5925), .B1(n5934), .B2(n5330), .ZN(U2828)
         );
  OAI222_X1 U6483 ( .A1(n5390), .A2(n5399), .B1(n5332), .B2(n5934), .C1(n5521), 
        .C2(n5925), .ZN(U2831) );
  INV_X1 U6484 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5333) );
  OAI222_X1 U6485 ( .A1(n5390), .A2(n5423), .B1(n5333), .B2(n5934), .C1(n5531), 
        .C2(n5925), .ZN(U2832) );
  AND2_X1 U6486 ( .A1(n5334), .A2(n5335), .ZN(n5336) );
  NOR2_X1 U6487 ( .A1(n5346), .A2(n5337), .ZN(n5338) );
  OR2_X1 U6488 ( .A1(n5339), .A2(n5338), .ZN(n5613) );
  OAI222_X1 U6489 ( .A1(n5390), .A2(n5427), .B1(n5340), .B2(n5934), .C1(n5613), 
        .C2(n5925), .ZN(U2833) );
  NAND2_X1 U6490 ( .A1(n4318), .A2(n5341), .ZN(n5342) );
  AND2_X1 U6491 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NOR2_X1 U6492 ( .A1(n5346), .A2(n5345), .ZN(n5712) );
  INV_X1 U6493 ( .A(n5712), .ZN(n5347) );
  OAI222_X1 U6494 ( .A1(n5435), .A2(n5390), .B1(n5348), .B2(n5934), .C1(n5925), 
        .C2(n5347), .ZN(U2834) );
  NOR2_X1 U6495 ( .A1(n5934), .A2(n6647), .ZN(n5349) );
  AOI21_X1 U6496 ( .B1(n5553), .B2(n5930), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6497 ( .B1(n5404), .B2(n5390), .A(n5350), .ZN(U2835) );
  NOR2_X1 U6498 ( .A1(n2988), .A2(n5351), .ZN(n5352) );
  OR2_X1 U6499 ( .A1(n4319), .A2(n5352), .ZN(n5629) );
  INV_X1 U6500 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5357) );
  OR2_X1 U6501 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6502 ( .A1(n5356), .A2(n5355), .ZN(n5631) );
  OAI222_X1 U6503 ( .A1(n5390), .A2(n5629), .B1(n5357), .B2(n5934), .C1(n5631), 
        .C2(n5925), .ZN(U2836) );
  AOI22_X1 U6504 ( .A1(n5567), .A2(n5930), .B1(EBX_REG_22__SCAN_IN), .B2(n5386), .ZN(n5358) );
  OAI21_X1 U6505 ( .B1(n5676), .B2(n5390), .A(n5358), .ZN(U2837) );
  NAND2_X1 U6506 ( .A1(n5359), .A2(n5360), .ZN(n5361) );
  AND2_X1 U6507 ( .A1(n5261), .A2(n5361), .ZN(n5689) );
  INV_X1 U6508 ( .A(n5689), .ZN(n5647) );
  INV_X1 U6509 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5364) );
  MUX2_X1 U6510 ( .A(n5367), .B(n4121), .S(n5370), .Z(n5363) );
  XNOR2_X1 U6511 ( .A(n5363), .B(n5362), .ZN(n5722) );
  INV_X1 U6512 ( .A(n5722), .ZN(n5646) );
  OAI222_X1 U6513 ( .A1(n5647), .A2(n5390), .B1(n5364), .B2(n5934), .C1(n5925), 
        .C2(n5646), .ZN(U2839) );
  OAI21_X1 U6514 ( .B1(n5365), .B2(n5366), .A(n5359), .ZN(n5660) );
  MUX2_X1 U6515 ( .A(n5368), .B(n5367), .S(n4080), .Z(n5381) );
  INV_X1 U6516 ( .A(n5381), .ZN(n5369) );
  OR2_X1 U6517 ( .A1(n5370), .A2(n5369), .ZN(n5373) );
  NAND2_X1 U6518 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  NAND2_X1 U6519 ( .A1(n5383), .A2(n3048), .ZN(n5372) );
  NOR2_X1 U6520 ( .A1(n5934), .A2(n5374), .ZN(n5375) );
  AOI21_X1 U6521 ( .B1(n5657), .B2(n5930), .A(n5375), .ZN(n5376) );
  OAI21_X1 U6522 ( .B1(n5660), .B2(n5390), .A(n5376), .ZN(U2840) );
  INV_X1 U6523 ( .A(n5377), .ZN(n5378) );
  NOR2_X1 U6524 ( .A1(n5378), .A2(n5379), .ZN(n5380) );
  OR2_X1 U6525 ( .A1(n5365), .A2(n5380), .ZN(n5696) );
  OR2_X1 U6526 ( .A1(n5382), .A2(n5381), .ZN(n5384) );
  AOI22_X1 U6527 ( .A1(n5806), .A2(n5930), .B1(EBX_REG_18__SCAN_IN), .B2(n5386), .ZN(n5385) );
  OAI21_X1 U6528 ( .B1(n5696), .B2(n5390), .A(n5385), .ZN(U2841) );
  AOI22_X1 U6529 ( .A1(n5737), .A2(n5930), .B1(EBX_REG_17__SCAN_IN), .B2(n5386), .ZN(n5387) );
  OAI21_X1 U6530 ( .B1(n5388), .B2(n5390), .A(n5387), .ZN(U2842) );
  OAI222_X1 U6531 ( .A1(n5391), .A2(n5390), .B1(n5389), .B2(n5934), .C1(n5925), 
        .C2(n5744), .ZN(U2843) );
  AOI22_X1 U6532 ( .A1(n5941), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5944), .ZN(n5395) );
  NAND2_X1 U6533 ( .A1(n5396), .A2(n5395), .ZN(U2860) );
  AOI22_X1 U6534 ( .A1(n5941), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5944), .ZN(n5398) );
  NAND2_X1 U6535 ( .A1(n5945), .A2(DATAI_12_), .ZN(n5397) );
  OAI211_X1 U6536 ( .C1(n5399), .C2(n5669), .A(n5398), .B(n5397), .ZN(U2863)
         );
  AOI22_X1 U6537 ( .A1(n5941), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5944), .ZN(n5401) );
  NAND2_X1 U6538 ( .A1(n5945), .A2(DATAI_11_), .ZN(n5400) );
  OAI211_X1 U6539 ( .C1(n5423), .C2(n5669), .A(n5401), .B(n5400), .ZN(U2864)
         );
  AOI22_X1 U6540 ( .A1(n5945), .A2(DATAI_8_), .B1(n5944), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6541 ( .A1(n5941), .A2(DATAI_24_), .ZN(n5402) );
  OAI211_X1 U6542 ( .C1(n5404), .C2(n5669), .A(n5403), .B(n5402), .ZN(U2867)
         );
  AOI22_X1 U6543 ( .A1(n5945), .A2(DATAI_7_), .B1(n5944), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6544 ( .A1(n5941), .A2(DATAI_23_), .ZN(n5405) );
  OAI211_X1 U6545 ( .C1(n5629), .C2(n5669), .A(n5406), .B(n5405), .ZN(U2868)
         );
  AOI22_X1 U6546 ( .A1(n5945), .A2(DATAI_3_), .B1(n5944), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6547 ( .A1(n5941), .A2(DATAI_19_), .ZN(n5407) );
  OAI211_X1 U6548 ( .C1(n5660), .C2(n5669), .A(n5408), .B(n5407), .ZN(U2872)
         );
  NAND3_X1 U6549 ( .A1(n5409), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n2967), .ZN(n5412) );
  NAND2_X1 U6550 ( .A1(n5716), .A2(n6613), .ZN(n5539) );
  OR2_X1 U6551 ( .A1(n2967), .A2(n5539), .ZN(n5411) );
  OR2_X1 U6552 ( .A1(n5410), .A2(n5411), .ZN(n5419) );
  AOI22_X1 U6553 ( .A1(n5412), .A2(n5419), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6613), .ZN(n5413) );
  XNOR2_X1 U6554 ( .A(n5413), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5528)
         );
  OR2_X1 U6555 ( .A1(n6092), .A2(n6588), .ZN(n5523) );
  NAND2_X1 U6556 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5414)
         );
  OAI211_X1 U6557 ( .C1(n6090), .C2(n5415), .A(n5523), .B(n5414), .ZN(n5416)
         );
  AOI21_X1 U6558 ( .B1(n5417), .B2(n6075), .A(n5416), .ZN(n5418) );
  OAI21_X1 U6559 ( .B1(n6065), .B2(n5528), .A(n5418), .ZN(U2958) );
  NAND2_X1 U6560 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  XNOR2_X1 U6561 ( .A(n5421), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5538)
         );
  NAND2_X1 U6562 ( .A1(n6171), .A2(REIP_REG_27__SCAN_IN), .ZN(n5530) );
  OAI21_X1 U6563 ( .B1(n5483), .B2(n5422), .A(n5530), .ZN(n5424) );
  XNOR2_X1 U6564 ( .A(n2967), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5426)
         );
  XNOR2_X1 U6565 ( .A(n5409), .B(n5426), .ZN(n5546) );
  NAND2_X1 U6566 ( .A1(n6171), .A2(REIP_REG_26__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U6567 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5428)
         );
  OAI211_X1 U6568 ( .C1(n6090), .C2(n5619), .A(n5541), .B(n5428), .ZN(n5429)
         );
  AOI21_X1 U6569 ( .B1(n5670), .B2(n6075), .A(n5429), .ZN(n5430) );
  OAI21_X1 U6570 ( .B1(n6065), .B2(n5546), .A(n5430), .ZN(U2960) );
  AOI21_X1 U6571 ( .B1(n5432), .B2(n5410), .A(n5431), .ZN(n5711) );
  INV_X1 U6572 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5433) );
  OAI22_X1 U6573 ( .A1(n5483), .A2(n5434), .B1(n6092), .B2(n5433), .ZN(n5437)
         );
  NOR2_X1 U6574 ( .A1(n5435), .A2(n6063), .ZN(n5436) );
  OAI21_X1 U6575 ( .B1(n5711), .B2(n6065), .A(n5438), .ZN(U2961) );
  NOR2_X1 U6576 ( .A1(n2967), .A2(n5474), .ZN(n5439) );
  OAI22_X1 U6577 ( .A1(n5472), .A2(n5439), .B1(n4219), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5688) );
  INV_X1 U6578 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5726) );
  AND2_X1 U6579 ( .A1(n2967), .A2(n5726), .ZN(n5686) );
  OR2_X1 U6580 ( .A1(n2967), .A2(n5726), .ZN(n5685) );
  XNOR2_X1 U6581 ( .A(n2967), .B(n6670), .ZN(n5466) );
  NAND4_X1 U6582 ( .A1(n5460), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n2967), .ZN(n5442) );
  NOR2_X1 U6583 ( .A1(n2967), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5458)
         );
  NAND2_X1 U6584 ( .A1(n5440), .A2(n5559), .ZN(n5441) );
  NAND2_X1 U6585 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  XNOR2_X1 U6586 ( .A(n5443), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5555)
         );
  NAND2_X1 U6587 ( .A1(n6171), .A2(REIP_REG_24__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6588 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5444)
         );
  OAI211_X1 U6589 ( .C1(n6090), .C2(n5445), .A(n5547), .B(n5444), .ZN(n5446)
         );
  AOI21_X1 U6590 ( .B1(n5447), .B2(n6075), .A(n5446), .ZN(n5448) );
  OAI21_X1 U6591 ( .B1(n5555), .B2(n6065), .A(n5448), .ZN(U2962) );
  NOR3_X1 U6592 ( .A1(n5449), .A2(n4219), .A3(n5693), .ZN(n5699) );
  NAND4_X1 U6593 ( .A1(n5699), .A2(n5583), .A3(n5451), .A4(n5450), .ZN(n5452)
         );
  NAND2_X1 U6594 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  XNOR2_X1 U6595 ( .A(n5454), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5562)
         );
  NAND2_X1 U6596 ( .A1(n6171), .A2(REIP_REG_23__SCAN_IN), .ZN(n5556) );
  OAI21_X1 U6597 ( .B1(n5483), .B2(n5638), .A(n5556), .ZN(n5456) );
  NOR2_X1 U6598 ( .A1(n5629), .A2(n6063), .ZN(n5455) );
  AOI211_X1 U6599 ( .C1(n6059), .C2(n5628), .A(n5456), .B(n5455), .ZN(n5457)
         );
  OAI21_X1 U6600 ( .B1(n5562), .B2(n6065), .A(n5457), .ZN(U2963) );
  AOI21_X1 U6601 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2967), .A(n5458), 
        .ZN(n5459) );
  XNOR2_X1 U6602 ( .A(n5460), .B(n5459), .ZN(n5563) );
  NAND2_X1 U6603 ( .A1(n5563), .A2(n6085), .ZN(n5464) );
  NOR2_X1 U6604 ( .A1(n6092), .A2(n6492), .ZN(n5566) );
  NOR2_X1 U6605 ( .A1(n6090), .A2(n5461), .ZN(n5462) );
  AOI211_X1 U6606 ( .C1(n6080), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5566), 
        .B(n5462), .ZN(n5463) );
  OAI211_X1 U6607 ( .C1(n6063), .C2(n5676), .A(n5464), .B(n5463), .ZN(U2964)
         );
  AOI21_X1 U6608 ( .B1(n5466), .B2(n5465), .A(n2983), .ZN(n5582) );
  XOR2_X1 U6609 ( .A(n5467), .B(n5261), .Z(n5680) );
  INV_X1 U6610 ( .A(n5639), .ZN(n5469) );
  NOR2_X1 U6611 ( .A1(n6092), .A2(n6488), .ZN(n5576) );
  AOI21_X1 U6612 ( .B1(n6080), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5576), 
        .ZN(n5468) );
  OAI21_X1 U6613 ( .B1(n5469), .B2(n6090), .A(n5468), .ZN(n5470) );
  AOI21_X1 U6614 ( .B1(n5680), .B2(n6075), .A(n5470), .ZN(n5471) );
  OAI21_X1 U6615 ( .B1(n5582), .B2(n6065), .A(n5471), .ZN(U2965) );
  INV_X1 U6616 ( .A(n5472), .ZN(n5473) );
  AOI22_X1 U6617 ( .A1(n4219), .A2(n5473), .B1(n5699), .B2(n5583), .ZN(n5475)
         );
  XNOR2_X1 U6618 ( .A(n5475), .B(n5474), .ZN(n5590) );
  INV_X1 U6619 ( .A(n5660), .ZN(n5479) );
  INV_X1 U6620 ( .A(n5663), .ZN(n5477) );
  AOI22_X1 U6621 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6171), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5476) );
  OAI21_X1 U6622 ( .B1(n5477), .B2(n6090), .A(n5476), .ZN(n5478) );
  AOI21_X1 U6623 ( .B1(n5479), .B2(n6075), .A(n5478), .ZN(n5480) );
  OAI21_X1 U6624 ( .B1(n5590), .B2(n6065), .A(n5480), .ZN(U2967) );
  OAI21_X1 U6625 ( .B1(n4219), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5481), 
        .ZN(n5482) );
  XNOR2_X1 U6626 ( .A(n5449), .B(n5482), .ZN(n5745) );
  OAI22_X1 U6627 ( .A1(n5483), .A2(n6637), .B1(n6092), .B2(n5751), .ZN(n5484)
         );
  AOI21_X1 U6628 ( .B1(n6059), .B2(n5485), .A(n5484), .ZN(n5487) );
  NAND2_X1 U6629 ( .A1(n5943), .A2(n6075), .ZN(n5486) );
  OAI211_X1 U6630 ( .C1(n5745), .C2(n6065), .A(n5487), .B(n5486), .ZN(U2970)
         );
  XNOR2_X1 U6631 ( .A(n2967), .B(n5756), .ZN(n5489) );
  XNOR2_X1 U6632 ( .A(n5488), .B(n5489), .ZN(n5753) );
  INV_X1 U6633 ( .A(n5753), .ZN(n5495) );
  AOI22_X1 U6634 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6171), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5490) );
  OAI21_X1 U6635 ( .B1(n5491), .B2(n6090), .A(n5490), .ZN(n5492) );
  AOI21_X1 U6636 ( .B1(n5493), .B2(n6075), .A(n5492), .ZN(n5494) );
  OAI21_X1 U6637 ( .B1(n5495), .B2(n6065), .A(n5494), .ZN(U2971) );
  XNOR2_X1 U6638 ( .A(n2967), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5497)
         );
  XNOR2_X1 U6639 ( .A(n5496), .B(n5497), .ZN(n5604) );
  NAND2_X1 U6640 ( .A1(n5604), .A2(n6085), .ZN(n5501) );
  INV_X1 U6641 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U6642 ( .A1(n6092), .A2(n5498), .ZN(n5597) );
  AND2_X1 U6643 ( .A1(n6080), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5499)
         );
  AOI211_X1 U6644 ( .C1(n5815), .C2(n6059), .A(n5597), .B(n5499), .ZN(n5500)
         );
  OAI211_X1 U6645 ( .C1(n6063), .C2(n5814), .A(n5501), .B(n5500), .ZN(U2972)
         );
  INV_X1 U6646 ( .A(n5502), .ZN(n5506) );
  NOR4_X1 U6647 ( .A1(n5529), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5519), 
        .A4(n5511), .ZN(n5505) );
  INV_X1 U6648 ( .A(n5503), .ZN(n5504) );
  AOI211_X1 U6649 ( .C1(n5506), .C2(n6169), .A(n5505), .B(n5504), .ZN(n5509)
         );
  INV_X1 U6650 ( .A(n5717), .ZN(n5544) );
  INV_X1 U6651 ( .A(n5519), .ZN(n5507) );
  OAI211_X1 U6652 ( .C1(n5507), .C2(n6106), .A(n5532), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U6653 ( .C1(n5586), .C2(n5544), .A(n5516), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5508) );
  OAI211_X1 U6654 ( .C1(n5510), .C2(n6095), .A(n5509), .B(n5508), .ZN(U2988)
         );
  OAI21_X1 U6655 ( .B1(n5529), .B2(n5519), .A(n5511), .ZN(n5515) );
  OAI21_X1 U6656 ( .B1(n5513), .B2(n6094), .A(n5512), .ZN(n5514) );
  AOI21_X1 U6657 ( .B1(n5516), .B2(n5515), .A(n5514), .ZN(n5517) );
  OAI21_X1 U6658 ( .B1(n5518), .B2(n6095), .A(n5517), .ZN(U2989) );
  INV_X1 U6659 ( .A(n5532), .ZN(n5526) );
  NAND2_X1 U6660 ( .A1(n5520), .A2(n5519), .ZN(n5524) );
  OR2_X1 U6661 ( .A1(n5521), .A2(n6094), .ZN(n5522) );
  OAI211_X1 U6662 ( .C1(n5529), .C2(n5524), .A(n5523), .B(n5522), .ZN(n5525)
         );
  AOI21_X1 U6663 ( .B1(n5526), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5525), 
        .ZN(n5527) );
  OAI21_X1 U6664 ( .B1(n5528), .B2(n6095), .A(n5527), .ZN(U2990) );
  INV_X1 U6665 ( .A(n5529), .ZN(n5536) );
  OAI21_X1 U6666 ( .B1(n5531), .B2(n6094), .A(n5530), .ZN(n5534) );
  NOR2_X1 U6667 ( .A1(n5532), .A2(n5535), .ZN(n5533) );
  AOI211_X1 U6668 ( .C1(n5536), .C2(n5535), .A(n5534), .B(n5533), .ZN(n5537)
         );
  OAI21_X1 U6669 ( .B1(n5538), .B2(n6095), .A(n5537), .ZN(U2991) );
  NAND3_X1 U6670 ( .A1(n5710), .A2(n5540), .A3(n5539), .ZN(n5542) );
  OAI211_X1 U6671 ( .C1(n6094), .C2(n5613), .A(n5542), .B(n5541), .ZN(n5543)
         );
  AOI21_X1 U6672 ( .B1(n5544), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5543), 
        .ZN(n5545) );
  OAI21_X1 U6673 ( .B1(n5546), .B2(n6095), .A(n5545), .ZN(U2992) );
  INV_X1 U6674 ( .A(n5547), .ZN(n5552) );
  INV_X1 U6675 ( .A(n5560), .ZN(n5549) );
  AOI211_X1 U6676 ( .C1(n5550), .C2(n5549), .A(n5548), .B(n5717), .ZN(n5551)
         );
  AOI211_X1 U6677 ( .C1(n6169), .C2(n5553), .A(n5552), .B(n5551), .ZN(n5554)
         );
  OAI21_X1 U6678 ( .B1(n5555), .B2(n6095), .A(n5554), .ZN(U2994) );
  OAI21_X1 U6679 ( .B1(n5631), .B2(n6094), .A(n5556), .ZN(n5558) );
  NOR2_X1 U6680 ( .A1(n5571), .A2(n5559), .ZN(n5557) );
  AOI211_X1 U6681 ( .C1(n5560), .C2(n5559), .A(n5558), .B(n5557), .ZN(n5561)
         );
  OAI21_X1 U6682 ( .B1(n5562), .B2(n6095), .A(n5561), .ZN(U2995) );
  NAND2_X1 U6683 ( .A1(n5563), .A2(n6175), .ZN(n5569) );
  NOR2_X1 U6684 ( .A1(n5564), .A2(n6670), .ZN(n5565) );
  AOI211_X1 U6685 ( .C1(n6169), .C2(n5567), .A(n5566), .B(n5565), .ZN(n5568)
         );
  OAI211_X1 U6686 ( .C1(n5571), .C2(n5570), .A(n5569), .B(n5568), .ZN(U2996)
         );
  AND2_X1 U6687 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  NOR2_X1 U6688 ( .A1(n5575), .A2(n5574), .ZN(n5666) );
  AOI21_X1 U6689 ( .B1(n5666), .B2(n6169), .A(n5576), .ZN(n5577) );
  OAI21_X1 U6690 ( .B1(n5578), .B2(n6670), .A(n5577), .ZN(n5579) );
  AOI21_X1 U6691 ( .B1(n5580), .B2(n6670), .A(n5579), .ZN(n5581) );
  OAI21_X1 U6692 ( .B1(n5582), .B2(n6095), .A(n5581), .ZN(U2997) );
  NAND2_X1 U6693 ( .A1(n5583), .A2(n5739), .ZN(n5718) );
  OAI221_X1 U6694 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5585), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5584), .A(n5735), .ZN(n5729) );
  AOI21_X1 U6695 ( .B1(n5730), .B2(n5586), .A(n5729), .ZN(n5727) );
  NAND2_X1 U6696 ( .A1(n6171), .A2(REIP_REG_19__SCAN_IN), .ZN(n5587) );
  OAI221_X1 U6697 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5718), .C1(
        n5474), .C2(n5727), .A(n5587), .ZN(n5588) );
  AOI21_X1 U6698 ( .B1(n5657), .B2(n6169), .A(n5588), .ZN(n5589) );
  OAI21_X1 U6699 ( .B1(n5590), .B2(n6095), .A(n5589), .ZN(U2999) );
  NOR2_X1 U6700 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5592), .ZN(n5760)
         );
  NAND2_X1 U6701 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  OAI211_X1 U6702 ( .C1(n5599), .C2(n5594), .A(n6101), .B(n5593), .ZN(n5764)
         );
  AOI21_X1 U6703 ( .B1(n5760), .B2(n5595), .A(n5764), .ZN(n5596) );
  NOR2_X1 U6704 ( .A1(n5596), .A2(n4226), .ZN(n5603) );
  INV_X1 U6705 ( .A(n5597), .ZN(n5601) );
  NOR2_X1 U6706 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6091), .ZN(n5598)
         );
  NAND2_X1 U6707 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  OAI211_X1 U6708 ( .C1(n6094), .C2(n5811), .A(n5601), .B(n5600), .ZN(n5602)
         );
  AOI211_X1 U6709 ( .C1(n5604), .C2(n6175), .A(n5603), .B(n5602), .ZN(n5605)
         );
  INV_X1 U6710 ( .A(n5605), .ZN(U3004) );
  OAI21_X1 U6711 ( .B1(n2978), .B2(STATEBS16_REG_SCAN_IN), .A(n6272), .ZN(
        n5606) );
  OAI22_X1 U6712 ( .A1(n5606), .A2(n6271), .B1(n2979), .B2(n5609), .ZN(n5607)
         );
  MUX2_X1 U6713 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5607), .S(n6181), 
        .Z(U3464) );
  XNOR2_X1 U6714 ( .A(n5608), .B(n6271), .ZN(n5610) );
  OAI22_X1 U6715 ( .A1(n5610), .A2(n6318), .B1(n4470), .B2(n5609), .ZN(n5611)
         );
  MUX2_X1 U6716 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5611), .S(n6181), 
        .Z(U3463) );
  AND2_X1 U6717 ( .A1(n5960), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6718 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5903), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5905), .ZN(n5618) );
  NOR2_X1 U6719 ( .A1(n6494), .A2(n5612), .ZN(n5620) );
  AOI21_X1 U6720 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5620), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5614) );
  OAI22_X1 U6721 ( .A1(n5615), .A2(n5614), .B1(n5613), .B2(n5874), .ZN(n5616)
         );
  AOI21_X1 U6722 ( .B1(n5670), .B2(n5879), .A(n5616), .ZN(n5617) );
  OAI211_X1 U6723 ( .C1(n5619), .C2(n5883), .A(n5618), .B(n5617), .ZN(U2801)
         );
  AOI22_X1 U6724 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5903), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5905), .ZN(n5627) );
  AOI22_X1 U6725 ( .A1(n5621), .A2(n5912), .B1(n5620), .B2(n5433), .ZN(n5626)
         );
  AOI22_X1 U6726 ( .A1(n5673), .A2(n5879), .B1(n5906), .B2(n5712), .ZN(n5625)
         );
  OAI21_X1 U6727 ( .B1(n5623), .B2(n5622), .A(REIP_REG_25__SCAN_IN), .ZN(n5624) );
  NAND4_X1 U6728 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(U2802)
         );
  AOI22_X1 U6729 ( .A1(EBX_REG_23__SCAN_IN), .A2(n5903), .B1(n5628), .B2(n5912), .ZN(n5637) );
  INV_X1 U6730 ( .A(n5629), .ZN(n5635) );
  AOI21_X1 U6731 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5630), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5632) );
  OAI22_X1 U6732 ( .A1(n5633), .A2(n5632), .B1(n5631), .B2(n5874), .ZN(n5634)
         );
  AOI21_X1 U6733 ( .B1(n5635), .B2(n5879), .A(n5634), .ZN(n5636) );
  OAI211_X1 U6734 ( .C1(n5638), .C2(n5889), .A(n5637), .B(n5636), .ZN(U2804)
         );
  AOI22_X1 U6735 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5905), .B1(n5639), 
        .B2(n5912), .ZN(n5645) );
  INV_X1 U6736 ( .A(n5640), .ZN(n5650) );
  AOI22_X1 U6737 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5903), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5650), .ZN(n5644) );
  AOI22_X1 U6738 ( .A1(n5680), .A2(n5879), .B1(n5906), .B2(n5666), .ZN(n5643)
         );
  OR2_X1 U6739 ( .A1(n5641), .A2(REIP_REG_21__SCAN_IN), .ZN(n5642) );
  NAND4_X1 U6740 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(U2806)
         );
  AOI22_X1 U6741 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5903), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5905), .ZN(n5652) );
  OAI22_X1 U6742 ( .A1(n5647), .A2(n5659), .B1(n5874), .B2(n5646), .ZN(n5648)
         );
  AOI221_X1 U6743 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5650), .C1(n5649), .C2(
        n5650), .A(n5648), .ZN(n5651) );
  OAI211_X1 U6744 ( .C1(n5692), .C2(n5883), .A(n5652), .B(n5651), .ZN(U2807)
         );
  OAI22_X1 U6745 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5654), .B1(n5653), .B2(
        n5889), .ZN(n5655) );
  AOI211_X1 U6746 ( .C1(n5903), .C2(EBX_REG_19__SCAN_IN), .A(n5892), .B(n5655), 
        .ZN(n5665) );
  INV_X1 U6747 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U6748 ( .A1(n5656), .A2(n6485), .ZN(n5802) );
  AOI21_X1 U6749 ( .B1(n5804), .B2(n5802), .A(n6487), .ZN(n5662) );
  INV_X1 U6750 ( .A(n5657), .ZN(n5658) );
  OAI22_X1 U6751 ( .A1(n5660), .A2(n5659), .B1(n5874), .B2(n5658), .ZN(n5661)
         );
  AOI211_X1 U6752 ( .C1(n5912), .C2(n5663), .A(n5662), .B(n5661), .ZN(n5664)
         );
  NAND2_X1 U6753 ( .A1(n5665), .A2(n5664), .ZN(U2808) );
  AOI22_X1 U6754 ( .A1(n5680), .A2(n5931), .B1(n5930), .B2(n5666), .ZN(n5667)
         );
  OAI21_X1 U6755 ( .B1(n5934), .B2(n5668), .A(n5667), .ZN(U2838) );
  AOI22_X1 U6756 ( .A1(n5670), .A2(n5942), .B1(n5941), .B2(DATAI_26_), .ZN(
        n5672) );
  AOI22_X1 U6757 ( .A1(n5945), .A2(DATAI_10_), .B1(n5944), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6758 ( .A1(n5672), .A2(n5671), .ZN(U2865) );
  AOI22_X1 U6759 ( .A1(n5673), .A2(n5942), .B1(n5941), .B2(DATAI_25_), .ZN(
        n5675) );
  AOI22_X1 U6760 ( .A1(n5945), .A2(DATAI_9_), .B1(n5944), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6761 ( .A1(n5675), .A2(n5674), .ZN(U2866) );
  INV_X1 U6762 ( .A(n5676), .ZN(n5677) );
  AOI22_X1 U6763 ( .A1(n5677), .A2(n5942), .B1(n5941), .B2(DATAI_22_), .ZN(
        n5679) );
  AOI22_X1 U6764 ( .A1(n5945), .A2(DATAI_6_), .B1(n5944), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6765 ( .A1(n5679), .A2(n5678), .ZN(U2869) );
  AOI22_X1 U6766 ( .A1(n5680), .A2(n5942), .B1(n5941), .B2(DATAI_21_), .ZN(
        n5682) );
  AOI22_X1 U6767 ( .A1(n5945), .A2(DATAI_5_), .B1(n5944), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U6768 ( .A1(n5682), .A2(n5681), .ZN(U2870) );
  AOI22_X1 U6769 ( .A1(n5689), .A2(n5942), .B1(n5941), .B2(DATAI_20_), .ZN(
        n5684) );
  AOI22_X1 U6770 ( .A1(n5945), .A2(DATAI_4_), .B1(n5944), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6771 ( .A1(n5684), .A2(n5683), .ZN(U2871) );
  AOI22_X1 U6772 ( .A1(n6171), .A2(REIP_REG_20__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5691) );
  NOR2_X1 U6773 ( .A1(n3018), .A2(n5686), .ZN(n5687) );
  XNOR2_X1 U6774 ( .A(n5688), .B(n5687), .ZN(n5723) );
  AOI22_X1 U6775 ( .A1(n5723), .A2(n6085), .B1(n6075), .B2(n5689), .ZN(n5690)
         );
  OAI211_X1 U6776 ( .C1(n6090), .C2(n5692), .A(n5691), .B(n5690), .ZN(U2966)
         );
  AOI22_X1 U6777 ( .A1(n6171), .A2(REIP_REG_18__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5698) );
  NAND3_X1 U6778 ( .A1(n5449), .A2(n4219), .A3(n5693), .ZN(n5700) );
  NOR2_X1 U6779 ( .A1(n5700), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5694)
         );
  AOI21_X1 U6780 ( .B1(n5699), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5694), 
        .ZN(n5695) );
  XNOR2_X1 U6781 ( .A(n5695), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5728)
         );
  AOI22_X1 U6782 ( .A1(n5728), .A2(n6085), .B1(n6075), .B2(n5935), .ZN(n5697)
         );
  OAI211_X1 U6783 ( .C1(n6090), .C2(n5809), .A(n5698), .B(n5697), .ZN(U2968)
         );
  INV_X1 U6784 ( .A(n5699), .ZN(n5701) );
  NAND2_X1 U6785 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  XNOR2_X1 U6786 ( .A(n5702), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5742)
         );
  AOI22_X1 U6787 ( .A1(n6171), .A2(REIP_REG_17__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5705) );
  AOI22_X1 U6788 ( .A1(n5938), .A2(n6075), .B1(n5703), .B2(n6059), .ZN(n5704)
         );
  OAI211_X1 U6789 ( .C1(n5742), .C2(n6065), .A(n5705), .B(n5704), .ZN(U2969)
         );
  AOI22_X1 U6790 ( .A1(n6171), .A2(REIP_REG_13__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5709) );
  XNOR2_X1 U6791 ( .A(n5706), .B(n5707), .ZN(n5765) );
  AOI22_X1 U6792 ( .A1(n5765), .A2(n6085), .B1(n6075), .B2(n5919), .ZN(n5708)
         );
  OAI211_X1 U6793 ( .C1(n6090), .C2(n5830), .A(n5709), .B(n5708), .ZN(U2973)
         );
  AOI22_X1 U6794 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6171), .B1(n5710), .B2(
        n5716), .ZN(n5715) );
  INV_X1 U6795 ( .A(n5711), .ZN(n5713) );
  AOI22_X1 U6796 ( .A1(n5713), .A2(n6175), .B1(n6169), .B2(n5712), .ZN(n5714)
         );
  OAI211_X1 U6797 ( .C1(n5717), .C2(n5716), .A(n5715), .B(n5714), .ZN(U2993)
         );
  NOR2_X1 U6798 ( .A1(n5719), .A2(n5718), .ZN(n5721) );
  AOI22_X1 U6799 ( .A1(n6171), .A2(REIP_REG_20__SCAN_IN), .B1(n5721), .B2(
        n5720), .ZN(n5725) );
  AOI22_X1 U6800 ( .A1(n5723), .A2(n6175), .B1(n6169), .B2(n5722), .ZN(n5724)
         );
  OAI211_X1 U6801 ( .C1(n5727), .C2(n5726), .A(n5725), .B(n5724), .ZN(U2998)
         );
  AOI22_X1 U6802 ( .A1(n5728), .A2(n6175), .B1(n6169), .B2(n5806), .ZN(n5734)
         );
  NAND2_X1 U6803 ( .A1(n6171), .A2(REIP_REG_18__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U6804 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5729), .ZN(n5732) );
  NAND3_X1 U6805 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5730), .A3(n5739), .ZN(n5731) );
  NAND4_X1 U6806 ( .A1(n5734), .A2(n5733), .A3(n5732), .A4(n5731), .ZN(U3000)
         );
  INV_X1 U6807 ( .A(n5735), .ZN(n5736) );
  AOI22_X1 U6808 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5736), .B1(n6171), .B2(REIP_REG_17__SCAN_IN), .ZN(n5741) );
  AOI22_X1 U6809 ( .A1(n5739), .A2(n5738), .B1(n5737), .B2(n6169), .ZN(n5740)
         );
  OAI211_X1 U6810 ( .C1(n5742), .C2(n6095), .A(n5741), .B(n5740), .ZN(U3001)
         );
  INV_X1 U6811 ( .A(n5747), .ZN(n5743) );
  OAI21_X1 U6812 ( .B1(n5743), .B2(n6106), .A(n6101), .ZN(n5755) );
  OAI22_X1 U6813 ( .A1(n5745), .A2(n6095), .B1(n6094), .B2(n5744), .ZN(n5746)
         );
  AOI21_X1 U6814 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5755), .A(n5746), 
        .ZN(n5750) );
  NOR2_X1 U6815 ( .A1(n6091), .A2(n5747), .ZN(n5757) );
  OAI211_X1 U6816 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5757), .B(n5748), .ZN(n5749) );
  OAI211_X1 U6817 ( .C1(n5751), .C2(n6092), .A(n5750), .B(n5749), .ZN(U3002)
         );
  AOI22_X1 U6818 ( .A1(n5753), .A2(n6175), .B1(n6169), .B2(n5752), .ZN(n5759)
         );
  NOR2_X1 U6819 ( .A1(n6092), .A2(n6481), .ZN(n5754) );
  AOI221_X1 U6820 ( .B1(n5757), .B2(n5756), .C1(n5755), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5754), .ZN(n5758) );
  NAND2_X1 U6821 ( .A1(n5759), .A2(n5758), .ZN(U3003) );
  INV_X1 U6822 ( .A(n5760), .ZN(n5768) );
  NOR2_X1 U6823 ( .A1(n2999), .A2(n5761), .ZN(n5762) );
  OR2_X1 U6824 ( .A1(n5763), .A2(n5762), .ZN(n5917) );
  INV_X1 U6825 ( .A(n5917), .ZN(n5821) );
  AOI22_X1 U6826 ( .A1(n6169), .A2(n5821), .B1(n6171), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5767) );
  AOI22_X1 U6827 ( .A1(n5765), .A2(n6175), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5764), .ZN(n5766) );
  OAI211_X1 U6828 ( .C1(n6091), .C2(n5768), .A(n5767), .B(n5766), .ZN(U3005)
         );
  OR4_X1 U6829 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n5773) );
  OAI21_X1 U6830 ( .B1(n5775), .B2(n5774), .A(n5773), .ZN(U3455) );
  INV_X1 U6831 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6590) );
  INV_X1 U6832 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6448) );
  AOI21_X1 U6833 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6590), .A(n6448), .ZN(n5782) );
  INV_X1 U6834 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5776) );
  AOI21_X1 U6835 ( .B1(n5782), .B2(n5776), .A(n6537), .ZN(U2789) );
  OAI21_X1 U6836 ( .B1(n6398), .B2(n5777), .A(n2962), .ZN(n5778) );
  OAI21_X1 U6837 ( .B1(n6414), .B2(n4256), .A(n5778), .ZN(n5786) );
  INV_X1 U6838 ( .A(n6429), .ZN(n6425) );
  OAI21_X1 U6839 ( .B1(n5786), .B2(n6425), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5779) );
  OAI21_X1 U6840 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5780), .A(n5779), .ZN(
        U2790) );
  INV_X2 U6841 ( .A(n6537), .ZN(n6505) );
  NOR2_X1 U6842 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5783) );
  OAI21_X1 U6843 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5783), .A(n6505), .ZN(n5781)
         );
  OAI21_X1 U6844 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6505), .A(n5781), .ZN(
        U2791) );
  NOR2_X1 U6845 ( .A1(n6537), .A2(n5782), .ZN(n6701) );
  OAI21_X1 U6846 ( .B1(BS16_N), .B2(n5783), .A(n6701), .ZN(n6699) );
  OAI21_X1 U6847 ( .B1(n6701), .B2(n5784), .A(n6699), .ZN(U2792) );
  AOI21_X1 U6848 ( .B1(n5785), .B2(n6445), .A(READY_N), .ZN(n6530) );
  NOR2_X1 U6849 ( .A1(n5786), .A2(n6530), .ZN(n6404) );
  NOR2_X1 U6850 ( .A1(n6404), .A2(n6425), .ZN(n6524) );
  OAI21_X1 U6851 ( .B1(n6524), .B2(n6572), .A(n6065), .ZN(U2793) );
  NOR4_X1 U6852 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5790) );
  NOR4_X1 U6853 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5789) );
  NOR4_X1 U6854 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5788) );
  NOR4_X1 U6855 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5787) );
  NAND4_X1 U6856 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n5796)
         );
  NOR4_X1 U6857 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n5794) );
  AOI211_X1 U6858 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_24__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5793) );
  NOR4_X1 U6859 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5792) );
  NOR4_X1 U6860 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5791) );
  NAND4_X1 U6861 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n5795)
         );
  NOR2_X1 U6862 ( .A1(n5796), .A2(n5795), .ZN(n6521) );
  INV_X1 U6863 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5798) );
  NOR3_X1 U6864 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5799) );
  OAI21_X1 U6865 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5799), .A(n6521), .ZN(n5797)
         );
  OAI21_X1 U6866 ( .B1(n6521), .B2(n5798), .A(n5797), .ZN(U2794) );
  INV_X1 U6867 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6700) );
  AOI21_X1 U6868 ( .B1(n6584), .B2(n6700), .A(n5799), .ZN(n5801) );
  INV_X1 U6869 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5800) );
  INV_X1 U6870 ( .A(n6521), .ZN(n6518) );
  AOI22_X1 U6871 ( .A1(n6521), .A2(n5801), .B1(n5800), .B2(n6518), .ZN(U2795)
         );
  AOI21_X1 U6872 ( .B1(n5905), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5892), 
        .ZN(n5803) );
  OAI211_X1 U6873 ( .C1(n5804), .C2(n6485), .A(n5803), .B(n5802), .ZN(n5805)
         );
  AOI21_X1 U6874 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5903), .A(n5805), .ZN(n5808)
         );
  AOI22_X1 U6875 ( .A1(n5935), .A2(n5879), .B1(n5906), .B2(n5806), .ZN(n5807)
         );
  OAI211_X1 U6876 ( .C1(n5809), .C2(n5883), .A(n5808), .B(n5807), .ZN(U2809)
         );
  NOR2_X1 U6877 ( .A1(n5826), .A2(n5810), .ZN(n5822) );
  AOI21_X1 U6878 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5822), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5820) );
  OAI22_X1 U6879 ( .A1(n5812), .A2(n5889), .B1(n5874), .B2(n5811), .ZN(n5813)
         );
  AOI211_X1 U6880 ( .C1(n5903), .C2(EBX_REG_14__SCAN_IN), .A(n5892), .B(n5813), 
        .ZN(n5818) );
  INV_X1 U6881 ( .A(n5814), .ZN(n5816) );
  AOI22_X1 U6882 ( .A1(n5816), .A2(n5879), .B1(n5912), .B2(n5815), .ZN(n5817)
         );
  OAI211_X1 U6883 ( .C1(n5820), .C2(n5819), .A(n5818), .B(n5817), .ZN(U2813)
         );
  INV_X1 U6884 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6478) );
  AOI22_X1 U6885 ( .A1(n5822), .A2(n6478), .B1(n5906), .B2(n5821), .ZN(n5823)
         );
  OAI21_X1 U6886 ( .B1(n5921), .B2(n5864), .A(n5823), .ZN(n5824) );
  AOI211_X1 U6887 ( .C1(n5905), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5892), 
        .B(n5824), .ZN(n5829) );
  OAI21_X1 U6888 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5826), .A(n5825), .ZN(n5827) );
  AOI22_X1 U6889 ( .A1(n5919), .A2(n5879), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5827), .ZN(n5828) );
  OAI211_X1 U6890 ( .C1(n5830), .C2(n5883), .A(n5829), .B(n5828), .ZN(U2814)
         );
  OAI21_X1 U6891 ( .B1(n5861), .B2(n5832), .A(n5831), .ZN(n5834) );
  NAND2_X1 U6892 ( .A1(n5834), .A2(n5833), .ZN(n6093) );
  INV_X1 U6893 ( .A(n6093), .ZN(n5922) );
  INV_X1 U6894 ( .A(n5835), .ZN(n5838) );
  INV_X1 U6895 ( .A(n5836), .ZN(n5837) );
  AND3_X1 U6896 ( .A1(n5897), .A2(n5838), .A3(n5837), .ZN(n5839) );
  AOI21_X1 U6897 ( .B1(n5922), .B2(n5906), .A(n5839), .ZN(n5845) );
  OAI22_X1 U6898 ( .A1(n6662), .A2(n5864), .B1(n5840), .B2(n5889), .ZN(n5841)
         );
  AOI211_X1 U6899 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5842), .A(n5892), .B(n5841), .ZN(n5844) );
  AOI22_X1 U6900 ( .A1(n6060), .A2(n5879), .B1(n5912), .B2(n6058), .ZN(n5843)
         );
  NAND3_X1 U6901 ( .A1(n5845), .A2(n5844), .A3(n5843), .ZN(U2816) );
  INV_X1 U6902 ( .A(n5846), .ZN(n6105) );
  AOI22_X1 U6903 ( .A1(n5906), .A2(n6105), .B1(n5903), .B2(EBX_REG_10__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6904 ( .A1(n5897), .A2(n5847), .ZN(n5853) );
  NOR3_X1 U6905 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5057), .A3(n5853), .ZN(n5848) );
  AOI211_X1 U6906 ( .C1(n5905), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5892), 
        .B(n5848), .ZN(n5856) );
  INV_X1 U6907 ( .A(n5849), .ZN(n5852) );
  INV_X1 U6908 ( .A(n5850), .ZN(n5851) );
  AOI22_X1 U6909 ( .A1(n5852), .A2(n5879), .B1(n5851), .B2(n5912), .ZN(n5855)
         );
  NOR2_X1 U6910 ( .A1(n5853), .A2(REIP_REG_9__SCAN_IN), .ZN(n5862) );
  OAI21_X1 U6911 ( .B1(n5862), .B2(n5866), .A(REIP_REG_10__SCAN_IN), .ZN(n5854) );
  NAND4_X1 U6912 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(U2817)
         );
  OR2_X1 U6913 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  NAND2_X1 U6914 ( .A1(n5861), .A2(n5860), .ZN(n5924) );
  INV_X1 U6915 ( .A(n5924), .ZN(n6112) );
  AOI21_X1 U6916 ( .B1(n6112), .B2(n5906), .A(n5862), .ZN(n5871) );
  OAI22_X1 U6917 ( .A1(n5929), .A2(n5864), .B1(n5863), .B2(n5889), .ZN(n5865)
         );
  AOI211_X1 U6918 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5866), .A(n5892), .B(n5865), 
        .ZN(n5870) );
  INV_X1 U6919 ( .A(n5926), .ZN(n5868) );
  AOI22_X1 U6920 ( .A1(n5868), .A2(n5879), .B1(n5912), .B2(n5867), .ZN(n5869)
         );
  NAND3_X1 U6921 ( .A1(n5871), .A2(n5870), .A3(n5869), .ZN(U2818) );
  AOI21_X1 U6922 ( .B1(n5905), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5892), 
        .ZN(n5873) );
  NAND2_X1 U6923 ( .A1(n5903), .A2(EBX_REG_6__SCAN_IN), .ZN(n5872) );
  OAI211_X1 U6924 ( .C1(n5875), .C2(n5874), .A(n5873), .B(n5872), .ZN(n5876)
         );
  AOI221_X1 U6925 ( .B1(n5878), .B2(REIP_REG_6__SCAN_IN), .C1(n5877), .C2(
        n6467), .A(n5876), .ZN(n5882) );
  INV_X1 U6926 ( .A(n6064), .ZN(n5880) );
  NAND2_X1 U6927 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  OAI211_X1 U6928 ( .C1(n5883), .C2(n6070), .A(n5882), .B(n5881), .ZN(U2821)
         );
  XNOR2_X1 U6929 ( .A(n5885), .B(n5884), .ZN(n6149) );
  AOI22_X1 U6930 ( .A1(n5906), .A2(n6149), .B1(n5903), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n5901) );
  INV_X1 U6931 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6463) );
  INV_X1 U6932 ( .A(n5896), .ZN(n5887) );
  OAI21_X1 U6933 ( .B1(n5888), .B2(n5887), .A(n5886), .ZN(n5916) );
  OAI22_X1 U6934 ( .A1(n5890), .A2(n5889), .B1(n6463), .B2(n5916), .ZN(n5891)
         );
  AOI211_X1 U6935 ( .C1(n5893), .C2(n5904), .A(n5892), .B(n5891), .ZN(n5900)
         );
  INV_X1 U6936 ( .A(n5910), .ZN(n5895) );
  INV_X1 U6937 ( .A(n6079), .ZN(n5894) );
  AOI22_X1 U6938 ( .A1(n5895), .A2(n6076), .B1(n5894), .B2(n5912), .ZN(n5899)
         );
  NAND3_X1 U6939 ( .A1(n5897), .A2(n5896), .A3(n6463), .ZN(n5898) );
  NAND4_X1 U6940 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(U2823)
         );
  OR2_X1 U6941 ( .A1(n5902), .A2(n6459), .ZN(n5915) );
  AOI22_X1 U6942 ( .A1(n5904), .A2(n4437), .B1(EBX_REG_3__SCAN_IN), .B2(n5903), 
        .ZN(n5908) );
  AOI22_X1 U6943 ( .A1(n5906), .A2(n6157), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n5905), .ZN(n5907) );
  OAI211_X1 U6944 ( .C1(n5910), .C2(n5909), .A(n5908), .B(n5907), .ZN(n5911)
         );
  AOI21_X1 U6945 ( .B1(n5913), .B2(n5912), .A(n5911), .ZN(n5914) );
  OAI221_X1 U6946 ( .B1(n5916), .B2(n6461), .C1(n5916), .C2(n5915), .A(n5914), 
        .ZN(U2824) );
  NOR2_X1 U6947 ( .A1(n5925), .A2(n5917), .ZN(n5918) );
  AOI21_X1 U6948 ( .B1(n5919), .B2(n5931), .A(n5918), .ZN(n5920) );
  OAI21_X1 U6949 ( .B1(n5934), .B2(n5921), .A(n5920), .ZN(U2846) );
  AOI22_X1 U6950 ( .A1(n6060), .A2(n5931), .B1(n5930), .B2(n5922), .ZN(n5923)
         );
  OAI21_X1 U6951 ( .B1(n5934), .B2(n6662), .A(n5923), .ZN(U2848) );
  OAI22_X1 U6952 ( .A1(n5926), .A2(n5390), .B1(n5925), .B2(n5924), .ZN(n5927)
         );
  INV_X1 U6953 ( .A(n5927), .ZN(n5928) );
  OAI21_X1 U6954 ( .B1(n5934), .B2(n5929), .A(n5928), .ZN(U2850) );
  AOI22_X1 U6955 ( .A1(n6076), .A2(n5931), .B1(n5930), .B2(n6149), .ZN(n5932)
         );
  OAI21_X1 U6956 ( .B1(n5934), .B2(n5933), .A(n5932), .ZN(U2855) );
  AOI22_X1 U6957 ( .A1(n5935), .A2(n5942), .B1(n5941), .B2(DATAI_18_), .ZN(
        n5937) );
  AOI22_X1 U6958 ( .A1(n5945), .A2(DATAI_2_), .B1(n5944), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U6959 ( .A1(n5937), .A2(n5936), .ZN(U2873) );
  AOI22_X1 U6960 ( .A1(n5938), .A2(n5942), .B1(n5941), .B2(DATAI_17_), .ZN(
        n5940) );
  AOI22_X1 U6961 ( .A1(n5945), .A2(DATAI_1_), .B1(n5944), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U6962 ( .A1(n5940), .A2(n5939), .ZN(U2874) );
  AOI22_X1 U6963 ( .A1(n5943), .A2(n5942), .B1(n5941), .B2(DATAI_16_), .ZN(
        n5947) );
  AOI22_X1 U6964 ( .A1(n5945), .A2(DATAI_0_), .B1(n5944), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U6965 ( .A1(n5947), .A2(n5946), .ZN(U2875) );
  INV_X1 U6966 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6053) );
  AOI22_X1 U6967 ( .A1(n5966), .A2(LWORD_REG_15__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U6968 ( .B1(n6053), .B2(n5968), .A(n5949), .ZN(U2908) );
  INV_X1 U6969 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U6970 ( .A1(n5956), .A2(LWORD_REG_14__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5950) );
  OAI21_X1 U6971 ( .B1(n6048), .B2(n5968), .A(n5950), .ZN(U2909) );
  INV_X1 U6972 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6045) );
  AOI22_X1 U6973 ( .A1(n5956), .A2(LWORD_REG_13__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5951) );
  OAI21_X1 U6974 ( .B1(n6045), .B2(n5968), .A(n5951), .ZN(U2910) );
  AOI22_X1 U6975 ( .A1(n5956), .A2(LWORD_REG_12__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5952) );
  OAI21_X1 U6976 ( .B1(n5081), .B2(n5968), .A(n5952), .ZN(U2911) );
  INV_X1 U6977 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6039) );
  AOI22_X1 U6978 ( .A1(n5956), .A2(LWORD_REG_11__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U6979 ( .B1(n6039), .B2(n5968), .A(n5953), .ZN(U2912) );
  INV_X1 U6980 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6036) );
  AOI22_X1 U6981 ( .A1(n5956), .A2(LWORD_REG_10__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U6982 ( .B1(n6036), .B2(n5968), .A(n5954), .ZN(U2913) );
  INV_X1 U6983 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6033) );
  AOI22_X1 U6984 ( .A1(n5956), .A2(LWORD_REG_9__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5955) );
  OAI21_X1 U6985 ( .B1(n6033), .B2(n5968), .A(n5955), .ZN(U2914) );
  INV_X1 U6986 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6030) );
  AOI22_X1 U6987 ( .A1(n5956), .A2(LWORD_REG_8__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5957) );
  OAI21_X1 U6988 ( .B1(n6030), .B2(n5968), .A(n5957), .ZN(U2915) );
  INV_X1 U6989 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6027) );
  AOI22_X1 U6990 ( .A1(n5966), .A2(LWORD_REG_7__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5958) );
  OAI21_X1 U6991 ( .B1(n6027), .B2(n5968), .A(n5958), .ZN(U2916) );
  AOI22_X1 U6992 ( .A1(n5966), .A2(LWORD_REG_6__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5959) );
  OAI21_X1 U6993 ( .B1(n4828), .B2(n5968), .A(n5959), .ZN(U2917) );
  AOI22_X1 U6994 ( .A1(n5966), .A2(LWORD_REG_5__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U6995 ( .B1(n3483), .B2(n5968), .A(n5961), .ZN(U2918) );
  AOI22_X1 U6996 ( .A1(n5966), .A2(LWORD_REG_4__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5962) );
  OAI21_X1 U6997 ( .B1(n6020), .B2(n5968), .A(n5962), .ZN(U2919) );
  AOI22_X1 U6998 ( .A1(n5966), .A2(LWORD_REG_3__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U6999 ( .B1(n6017), .B2(n5968), .A(n5963), .ZN(U2920) );
  AOI22_X1 U7000 ( .A1(n5966), .A2(LWORD_REG_2__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5964) );
  OAI21_X1 U7001 ( .B1(n6014), .B2(n5968), .A(n5964), .ZN(U2921) );
  INV_X1 U7002 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7003 ( .A1(n5966), .A2(LWORD_REG_1__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U7004 ( .B1(n6601), .B2(n5968), .A(n5965), .ZN(U2922) );
  AOI22_X1 U7005 ( .A1(n5966), .A2(LWORD_REG_0__SCAN_IN), .B1(n5960), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U7006 ( .B1(n6009), .B2(n5968), .A(n5967), .ZN(U2923) );
  INV_X1 U7007 ( .A(n5969), .ZN(n5970) );
  INV_X1 U7008 ( .A(n6004), .ZN(n6049) );
  AND2_X1 U7009 ( .A1(n6049), .A2(DATAI_0_), .ZN(n6007) );
  AOI21_X1 U7010 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6050), .A(n6007), .ZN(n5971) );
  OAI21_X1 U7011 ( .B1(n3635), .B2(n6052), .A(n5971), .ZN(U2924) );
  INV_X1 U7012 ( .A(DATAI_1_), .ZN(n5972) );
  NOR2_X1 U7013 ( .A1(n6004), .A2(n5972), .ZN(n6010) );
  AOI21_X1 U7014 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6050), .A(n6010), .ZN(n5973) );
  OAI21_X1 U7015 ( .B1(n3655), .B2(n6052), .A(n5973), .ZN(U2925) );
  AND2_X1 U7016 ( .A1(n6049), .A2(DATAI_2_), .ZN(n6012) );
  AOI21_X1 U7017 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6050), .A(n6012), .ZN(n5974) );
  OAI21_X1 U7018 ( .B1(n5975), .B2(n6052), .A(n5974), .ZN(U2926) );
  AND2_X1 U7019 ( .A1(n6049), .A2(DATAI_3_), .ZN(n6015) );
  AOI21_X1 U7020 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6050), .A(n6015), .ZN(n5976) );
  OAI21_X1 U7021 ( .B1(n5977), .B2(n6052), .A(n5976), .ZN(U2927) );
  AND2_X1 U7022 ( .A1(n6049), .A2(DATAI_4_), .ZN(n6018) );
  AOI21_X1 U7023 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6050), .A(n6018), .ZN(n5978) );
  OAI21_X1 U7024 ( .B1(n3709), .B2(n6052), .A(n5978), .ZN(U2928) );
  AND2_X1 U7025 ( .A1(n6049), .A2(DATAI_5_), .ZN(n6021) );
  AOI21_X1 U7026 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6050), .A(n6021), .ZN(n5979) );
  OAI21_X1 U7027 ( .B1(n5980), .B2(n6052), .A(n5979), .ZN(U2929) );
  NOR2_X1 U7028 ( .A1(n6004), .A2(n5981), .ZN(n6023) );
  AOI21_X1 U7029 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6050), .A(n6023), .ZN(n5982) );
  OAI21_X1 U7030 ( .B1(n5983), .B2(n6052), .A(n5982), .ZN(U2930) );
  INV_X1 U7031 ( .A(DATAI_7_), .ZN(n5984) );
  NOR2_X1 U7032 ( .A1(n6004), .A2(n5984), .ZN(n6025) );
  AOI21_X1 U7033 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6050), .A(n6025), .ZN(n5985) );
  OAI21_X1 U7034 ( .B1(n5986), .B2(n6052), .A(n5985), .ZN(U2931) );
  INV_X1 U7035 ( .A(DATAI_8_), .ZN(n5987) );
  NOR2_X1 U7036 ( .A1(n6004), .A2(n5987), .ZN(n6028) );
  AOI21_X1 U7037 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6050), .A(n6028), .ZN(n5988) );
  OAI21_X1 U7038 ( .B1(n5989), .B2(n6052), .A(n5988), .ZN(U2932) );
  INV_X1 U7039 ( .A(DATAI_9_), .ZN(n5990) );
  NOR2_X1 U7040 ( .A1(n6004), .A2(n5990), .ZN(n6031) );
  AOI21_X1 U7041 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6050), .A(n6031), .ZN(n5991) );
  OAI21_X1 U7042 ( .B1(n5992), .B2(n6052), .A(n5991), .ZN(U2933) );
  INV_X1 U7043 ( .A(DATAI_10_), .ZN(n5993) );
  NOR2_X1 U7044 ( .A1(n6004), .A2(n5993), .ZN(n6034) );
  AOI21_X1 U7045 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6050), .A(n6034), .ZN(
        n5994) );
  OAI21_X1 U7046 ( .B1(n3832), .B2(n6052), .A(n5994), .ZN(U2934) );
  INV_X1 U7047 ( .A(DATAI_11_), .ZN(n5995) );
  NOR2_X1 U7048 ( .A1(n6004), .A2(n5995), .ZN(n6037) );
  AOI21_X1 U7049 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6050), .A(n6037), .ZN(
        n5996) );
  OAI21_X1 U7050 ( .B1(n5997), .B2(n6052), .A(n5996), .ZN(U2935) );
  NOR2_X1 U7051 ( .A1(n6004), .A2(n5998), .ZN(n6040) );
  AOI21_X1 U7052 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6050), .A(n6040), .ZN(
        n5999) );
  OAI21_X1 U7053 ( .B1(n6567), .B2(n6052), .A(n5999), .ZN(U2936) );
  INV_X1 U7054 ( .A(DATAI_13_), .ZN(n6000) );
  NOR2_X1 U7055 ( .A1(n6004), .A2(n6000), .ZN(n6042) );
  AOI21_X1 U7056 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6050), .A(n6042), .ZN(
        n6001) );
  OAI21_X1 U7057 ( .B1(n6002), .B2(n6052), .A(n6001), .ZN(U2937) );
  INV_X1 U7058 ( .A(DATAI_14_), .ZN(n6003) );
  NOR2_X1 U7059 ( .A1(n6004), .A2(n6003), .ZN(n6046) );
  AOI21_X1 U7060 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6043), .A(n6046), .ZN(
        n6005) );
  OAI21_X1 U7061 ( .B1(n6006), .B2(n6052), .A(n6005), .ZN(U2938) );
  AOI21_X1 U7062 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6050), .A(n6007), .ZN(n6008) );
  OAI21_X1 U7063 ( .B1(n6009), .B2(n6052), .A(n6008), .ZN(U2939) );
  AOI21_X1 U7064 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6043), .A(n6010), .ZN(n6011) );
  OAI21_X1 U7065 ( .B1(n6601), .B2(n6052), .A(n6011), .ZN(U2940) );
  AOI21_X1 U7066 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6050), .A(n6012), .ZN(n6013) );
  OAI21_X1 U7067 ( .B1(n6014), .B2(n6052), .A(n6013), .ZN(U2941) );
  AOI21_X1 U7068 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6050), .A(n6015), .ZN(n6016) );
  OAI21_X1 U7069 ( .B1(n6017), .B2(n6052), .A(n6016), .ZN(U2942) );
  AOI21_X1 U7070 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6050), .A(n6018), .ZN(n6019) );
  OAI21_X1 U7071 ( .B1(n6020), .B2(n6052), .A(n6019), .ZN(U2943) );
  AOI21_X1 U7072 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6050), .A(n6021), .ZN(n6022) );
  OAI21_X1 U7073 ( .B1(n3483), .B2(n6052), .A(n6022), .ZN(U2944) );
  AOI21_X1 U7074 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6043), .A(n6023), .ZN(n6024) );
  OAI21_X1 U7075 ( .B1(n4828), .B2(n6052), .A(n6024), .ZN(U2945) );
  AOI21_X1 U7076 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6043), .A(n6025), .ZN(n6026) );
  OAI21_X1 U7077 ( .B1(n6027), .B2(n6052), .A(n6026), .ZN(U2946) );
  AOI21_X1 U7078 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6043), .A(n6028), .ZN(n6029) );
  OAI21_X1 U7079 ( .B1(n6030), .B2(n6052), .A(n6029), .ZN(U2947) );
  AOI21_X1 U7080 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6043), .A(n6031), .ZN(n6032) );
  OAI21_X1 U7081 ( .B1(n6033), .B2(n6052), .A(n6032), .ZN(U2948) );
  AOI21_X1 U7082 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6043), .A(n6034), .ZN(
        n6035) );
  OAI21_X1 U7083 ( .B1(n6036), .B2(n6052), .A(n6035), .ZN(U2949) );
  AOI21_X1 U7084 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6043), .A(n6037), .ZN(
        n6038) );
  OAI21_X1 U7085 ( .B1(n6039), .B2(n6052), .A(n6038), .ZN(U2950) );
  AOI21_X1 U7086 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6043), .A(n6040), .ZN(
        n6041) );
  OAI21_X1 U7087 ( .B1(n5081), .B2(n6052), .A(n6041), .ZN(U2951) );
  AOI21_X1 U7088 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6043), .A(n6042), .ZN(
        n6044) );
  OAI21_X1 U7089 ( .B1(n6045), .B2(n6052), .A(n6044), .ZN(U2952) );
  AOI21_X1 U7090 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6043), .A(n6046), .ZN(
        n6047) );
  OAI21_X1 U7091 ( .B1(n6048), .B2(n6052), .A(n6047), .ZN(U2953) );
  AOI22_X1 U7092 ( .A1(n6050), .A2(LWORD_REG_15__SCAN_IN), .B1(n6049), .B2(
        DATAI_15_), .ZN(n6051) );
  OAI21_X1 U7093 ( .B1(n6053), .B2(n6052), .A(n6051), .ZN(U2954) );
  NAND2_X1 U7094 ( .A1(n6055), .A2(n6054), .ZN(n6057) );
  XNOR2_X1 U7095 ( .A(n2967), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6056)
         );
  XNOR2_X1 U7096 ( .A(n6057), .B(n6056), .ZN(n6096) );
  AOI22_X1 U7097 ( .A1(n6171), .A2(REIP_REG_11__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6062) );
  AOI22_X1 U7098 ( .A1(n6060), .A2(n6075), .B1(n6059), .B2(n6058), .ZN(n6061)
         );
  OAI211_X1 U7099 ( .C1(n6096), .C2(n6065), .A(n6062), .B(n6061), .ZN(U2975)
         );
  AOI22_X1 U7100 ( .A1(n6171), .A2(REIP_REG_6__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6069) );
  OAI22_X1 U7101 ( .A1(n6066), .A2(n6065), .B1(n6064), .B2(n6063), .ZN(n6067)
         );
  INV_X1 U7102 ( .A(n6067), .ZN(n6068) );
  OAI211_X1 U7103 ( .C1(n6090), .C2(n6070), .A(n6069), .B(n6068), .ZN(U2980)
         );
  AOI22_X1 U7104 ( .A1(n6171), .A2(REIP_REG_4__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7105 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  AND2_X1 U7106 ( .A1(n6074), .A2(n6073), .ZN(n6150) );
  AOI22_X1 U7107 ( .A1(n6076), .A2(n6075), .B1(n6150), .B2(n6085), .ZN(n6077)
         );
  OAI211_X1 U7108 ( .C1(n6090), .C2(n6079), .A(n6078), .B(n6077), .ZN(U2982)
         );
  AOI22_X1 U7109 ( .A1(n6171), .A2(REIP_REG_2__SCAN_IN), .B1(n6080), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6088) );
  INV_X1 U7110 ( .A(n6081), .ZN(n6086) );
  XNOR2_X1 U7111 ( .A(n6082), .B(n6179), .ZN(n6084) );
  XNOR2_X1 U7112 ( .A(n6084), .B(n6083), .ZN(n6174) );
  AOI22_X1 U7113 ( .A1(n6075), .A2(n6086), .B1(n6174), .B2(n6085), .ZN(n6087)
         );
  OAI211_X1 U7114 ( .C1(n6090), .C2(n6089), .A(n6088), .B(n6087), .ZN(U2984)
         );
  INV_X1 U7115 ( .A(n6091), .ZN(n6099) );
  OAI22_X1 U7116 ( .A1(n6094), .A2(n6093), .B1(n6475), .B2(n6092), .ZN(n6098)
         );
  NOR2_X1 U7117 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  AOI211_X1 U7118 ( .C1(n6685), .C2(n6099), .A(n6098), .B(n6097), .ZN(n6100)
         );
  OAI21_X1 U7119 ( .B1(n6685), .B2(n6101), .A(n6100), .ZN(U3007) );
  NOR2_X1 U7120 ( .A1(n6158), .A2(n6102), .ZN(n6131) );
  NAND2_X1 U7121 ( .A1(n6121), .A2(n6131), .ZN(n6117) );
  AOI22_X1 U7122 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n4218), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6103), .ZN(n6110) );
  AOI21_X1 U7123 ( .B1(n6169), .B2(n6105), .A(n6104), .ZN(n6109) );
  OAI21_X1 U7124 ( .B1(n6106), .B2(n6121), .A(n6135), .ZN(n6113) );
  AOI22_X1 U7125 ( .A1(n6107), .A2(n6175), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6113), .ZN(n6108) );
  OAI211_X1 U7126 ( .C1(n6117), .C2(n6110), .A(n6109), .B(n6108), .ZN(U3008)
         );
  AOI21_X1 U7127 ( .B1(n6169), .B2(n6112), .A(n6111), .ZN(n6116) );
  AOI22_X1 U7128 ( .A1(n6114), .A2(n6175), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6113), .ZN(n6115) );
  OAI211_X1 U7129 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6117), .A(n6116), 
        .B(n6115), .ZN(U3009) );
  INV_X1 U7130 ( .A(n6118), .ZN(n6119) );
  AOI222_X1 U7131 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6171), .B1(n6169), .B2(
        n6120), .C1(n6175), .C2(n6119), .ZN(n6124) );
  INV_X1 U7132 ( .A(n6121), .ZN(n6122) );
  OAI211_X1 U7133 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6131), .B(n6122), .ZN(n6123) );
  OAI211_X1 U7134 ( .C1(n6135), .C2(n6125), .A(n6124), .B(n6123), .ZN(U3010)
         );
  INV_X1 U7135 ( .A(n6126), .ZN(n6127) );
  AOI21_X1 U7136 ( .B1(n6169), .B2(n6128), .A(n6127), .ZN(n6133) );
  INV_X1 U7137 ( .A(n6129), .ZN(n6130) );
  AOI22_X1 U7138 ( .A1(n6131), .A2(n6134), .B1(n6130), .B2(n6175), .ZN(n6132)
         );
  OAI211_X1 U7139 ( .C1(n6135), .C2(n6134), .A(n6133), .B(n6132), .ZN(U3011)
         );
  OAI21_X1 U7140 ( .B1(n6138), .B2(n6137), .A(n6136), .ZN(n6139) );
  AOI21_X1 U7141 ( .B1(n6172), .B2(n6140), .A(n6139), .ZN(n6146) );
  INV_X1 U7142 ( .A(n6141), .ZN(n6143) );
  AOI22_X1 U7143 ( .A1(n6143), .A2(n6175), .B1(n6169), .B2(n6142), .ZN(n6145)
         );
  NAND2_X1 U7144 ( .A1(n6171), .A2(REIP_REG_5__SCAN_IN), .ZN(n6144) );
  OAI211_X1 U7145 ( .C1(n6147), .C2(n6146), .A(n6145), .B(n6144), .ZN(U3013)
         );
  AOI21_X1 U7146 ( .B1(n6172), .B2(n6166), .A(n6148), .ZN(n6165) );
  AOI22_X1 U7147 ( .A1(n6169), .A2(n6149), .B1(n6171), .B2(REIP_REG_4__SCAN_IN), .ZN(n6154) );
  AOI211_X1 U7148 ( .C1(n6164), .C2(n6155), .A(n6158), .B(n6166), .ZN(n6152)
         );
  AOI22_X1 U7149 ( .A1(n6152), .A2(n6151), .B1(n6175), .B2(n6150), .ZN(n6153)
         );
  OAI211_X1 U7150 ( .C1(n6165), .C2(n6155), .A(n6154), .B(n6153), .ZN(U3014)
         );
  AOI21_X1 U7151 ( .B1(n6169), .B2(n6157), .A(n6156), .ZN(n6163) );
  NOR2_X1 U7152 ( .A1(n6166), .A2(n6158), .ZN(n6161) );
  INV_X1 U7153 ( .A(n6159), .ZN(n6160) );
  AOI22_X1 U7154 ( .A1(n6161), .A2(n6164), .B1(n6175), .B2(n6160), .ZN(n6162)
         );
  OAI211_X1 U7155 ( .C1(n6165), .C2(n6164), .A(n6163), .B(n6162), .ZN(U3015)
         );
  NAND2_X1 U7156 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6168) );
  INV_X1 U7157 ( .A(n6166), .ZN(n6167) );
  OAI21_X1 U7158 ( .B1(n6168), .B2(n6179), .A(n6167), .ZN(n6173) );
  AOI222_X1 U7159 ( .A1(n6173), .A2(n6172), .B1(REIP_REG_2__SCAN_IN), .B2(
        n6171), .C1(n6170), .C2(n6169), .ZN(n6178) );
  AOI22_X1 U7160 ( .A1(n6176), .A2(n6179), .B1(n6175), .B2(n6174), .ZN(n6177)
         );
  OAI211_X1 U7161 ( .C1(n6180), .C2(n6179), .A(n6178), .B(n6177), .ZN(U3016)
         );
  NOR2_X1 U7162 ( .A1(n6182), .A2(n6181), .ZN(U3019) );
  AOI22_X1 U7163 ( .A1(n6186), .A2(n6313), .B1(n6185), .B2(n6309), .ZN(n6187)
         );
  NAND2_X1 U7164 ( .A1(n6188), .A2(n6233), .ZN(n6189) );
  INV_X1 U7165 ( .A(n6189), .ZN(n6215) );
  AOI22_X1 U7166 ( .A1(n6317), .A2(n6216), .B1(n6316), .B2(n6215), .ZN(n6197)
         );
  AOI21_X1 U7167 ( .B1(n6189), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6194) );
  NOR3_X1 U7168 ( .A1(n6217), .A2(n6259), .A3(n6318), .ZN(n6192) );
  OAI21_X1 U7169 ( .B1(n6192), .B2(n6322), .A(n6191), .ZN(n6193) );
  NAND3_X1 U7170 ( .A1(n6195), .A2(n6194), .A3(n6193), .ZN(n6218) );
  AOI22_X1 U7171 ( .A1(n6218), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6228), 
        .B2(n6217), .ZN(n6196) );
  OAI211_X1 U7172 ( .C1(n6198), .C2(n6221), .A(n6197), .B(n6196), .ZN(U3068)
         );
  AOI22_X1 U7173 ( .A1(n6333), .A2(n6216), .B1(n6332), .B2(n6215), .ZN(n6200)
         );
  AOI22_X1 U7174 ( .A1(n6218), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6237), 
        .B2(n6217), .ZN(n6199) );
  OAI211_X1 U7175 ( .C1(n6201), .C2(n6221), .A(n6200), .B(n6199), .ZN(U3069)
         );
  AOI22_X1 U7176 ( .A1(n6339), .A2(n6216), .B1(n6338), .B2(n6215), .ZN(n6203)
         );
  AOI22_X1 U7177 ( .A1(n6218), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6241), 
        .B2(n6217), .ZN(n6202) );
  OAI211_X1 U7178 ( .C1(n6204), .C2(n6221), .A(n6203), .B(n6202), .ZN(U3070)
         );
  AOI22_X1 U7179 ( .A1(n6345), .A2(n6216), .B1(n6344), .B2(n6215), .ZN(n6206)
         );
  AOI22_X1 U7180 ( .A1(n6218), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6245), 
        .B2(n6217), .ZN(n6205) );
  OAI211_X1 U7181 ( .C1(n6207), .C2(n6221), .A(n6206), .B(n6205), .ZN(U3071)
         );
  AOI22_X1 U7182 ( .A1(n6351), .A2(n6216), .B1(n6350), .B2(n6215), .ZN(n6209)
         );
  AOI22_X1 U7183 ( .A1(n6218), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6291), 
        .B2(n6217), .ZN(n6208) );
  OAI211_X1 U7184 ( .C1(n6294), .C2(n6221), .A(n6209), .B(n6208), .ZN(U3072)
         );
  AOI22_X1 U7185 ( .A1(n6357), .A2(n6216), .B1(n6356), .B2(n6215), .ZN(n6211)
         );
  AOI22_X1 U7186 ( .A1(n6218), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6252), 
        .B2(n6217), .ZN(n6210) );
  OAI211_X1 U7187 ( .C1(n6212), .C2(n6221), .A(n6211), .B(n6210), .ZN(U3073)
         );
  AOI22_X1 U7188 ( .A1(n6363), .A2(n6216), .B1(n6362), .B2(n6215), .ZN(n6214)
         );
  AOI22_X1 U7189 ( .A1(n6218), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6297), 
        .B2(n6217), .ZN(n6213) );
  OAI211_X1 U7190 ( .C1(n6301), .C2(n6221), .A(n6214), .B(n6213), .ZN(U3074)
         );
  AOI22_X1 U7191 ( .A1(n6371), .A2(n6216), .B1(n6369), .B2(n6215), .ZN(n6220)
         );
  AOI22_X1 U7192 ( .A1(n6218), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6260), 
        .B2(n6217), .ZN(n6219) );
  OAI211_X1 U7193 ( .C1(n6222), .C2(n6221), .A(n6220), .B(n6219), .ZN(U3075)
         );
  INV_X1 U7194 ( .A(n6223), .ZN(n6225) );
  INV_X1 U7195 ( .A(n6224), .ZN(n6261) );
  AOI21_X1 U7196 ( .B1(n6226), .B2(n6225), .A(n6261), .ZN(n6229) );
  NOR2_X1 U7197 ( .A1(n6229), .A2(n6318), .ZN(n6227) );
  AOI21_X1 U7198 ( .B1(n6233), .B2(STATE2_REG_2__SCAN_IN), .A(n6227), .ZN(
        n6267) );
  AOI22_X1 U7199 ( .A1(n6316), .A2(n6261), .B1(n6228), .B2(n6259), .ZN(n6235)
         );
  NAND3_X1 U7200 ( .A1(n6230), .A2(n6272), .A3(n6229), .ZN(n6232) );
  OAI211_X1 U7201 ( .C1(n6233), .C2(n6272), .A(n6232), .B(n6231), .ZN(n6263)
         );
  AOI22_X1 U7202 ( .A1(n6263), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n6328), 
        .B2(n6262), .ZN(n6234) );
  OAI211_X1 U7203 ( .C1(n6267), .C2(n6236), .A(n6235), .B(n6234), .ZN(U3076)
         );
  AOI22_X1 U7204 ( .A1(n6332), .A2(n6261), .B1(n6237), .B2(n6259), .ZN(n6239)
         );
  AOI22_X1 U7205 ( .A1(n6263), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6334), 
        .B2(n6262), .ZN(n6238) );
  OAI211_X1 U7206 ( .C1(n6267), .C2(n6240), .A(n6239), .B(n6238), .ZN(U3077)
         );
  AOI22_X1 U7207 ( .A1(n6338), .A2(n6261), .B1(n6340), .B2(n6262), .ZN(n6243)
         );
  AOI22_X1 U7208 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6263), .B1(n6241), 
        .B2(n6259), .ZN(n6242) );
  OAI211_X1 U7209 ( .C1(n6267), .C2(n6244), .A(n6243), .B(n6242), .ZN(U3078)
         );
  AOI22_X1 U7210 ( .A1(n6344), .A2(n6261), .B1(n6245), .B2(n6259), .ZN(n6247)
         );
  AOI22_X1 U7211 ( .A1(n6263), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6346), 
        .B2(n6262), .ZN(n6246) );
  OAI211_X1 U7212 ( .C1(n6267), .C2(n6248), .A(n6247), .B(n6246), .ZN(U3079)
         );
  AOI22_X1 U7213 ( .A1(n6350), .A2(n6261), .B1(n6352), .B2(n6262), .ZN(n6250)
         );
  AOI22_X1 U7214 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6263), .B1(n6291), 
        .B2(n6259), .ZN(n6249) );
  OAI211_X1 U7215 ( .C1(n6267), .C2(n6251), .A(n6250), .B(n6249), .ZN(U3080)
         );
  AOI22_X1 U7216 ( .A1(n6356), .A2(n6261), .B1(n6252), .B2(n6259), .ZN(n6254)
         );
  AOI22_X1 U7217 ( .A1(n6263), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6358), 
        .B2(n6262), .ZN(n6253) );
  OAI211_X1 U7218 ( .C1(n6267), .C2(n6255), .A(n6254), .B(n6253), .ZN(U3081)
         );
  AOI22_X1 U7219 ( .A1(n6362), .A2(n6261), .B1(n6364), .B2(n6262), .ZN(n6257)
         );
  AOI22_X1 U7220 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6263), .B1(n6297), 
        .B2(n6259), .ZN(n6256) );
  OAI211_X1 U7221 ( .C1(n6267), .C2(n6258), .A(n6257), .B(n6256), .ZN(U3082)
         );
  AOI22_X1 U7222 ( .A1(n6369), .A2(n6261), .B1(n6260), .B2(n6259), .ZN(n6265)
         );
  AOI22_X1 U7223 ( .A1(n6263), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6373), 
        .B2(n6262), .ZN(n6264) );
  OAI211_X1 U7224 ( .C1(n6267), .C2(n6266), .A(n6265), .B(n6264), .ZN(U3083)
         );
  NOR2_X1 U7225 ( .A1(n6268), .A2(n6390), .ZN(n6302) );
  AOI22_X1 U7226 ( .A1(n6316), .A2(n6302), .B1(n6328), .B2(n6319), .ZN(n6284)
         );
  INV_X1 U7227 ( .A(n6271), .ZN(n6273) );
  OAI21_X1 U7228 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(n6282) );
  AOI21_X1 U7229 ( .B1(n6275), .B2(n3446), .A(n6302), .ZN(n6281) );
  INV_X1 U7230 ( .A(n6281), .ZN(n6278) );
  AOI21_X1 U7231 ( .B1(n6318), .B2(n6280), .A(n6276), .ZN(n6277) );
  OAI21_X1 U7232 ( .B1(n6282), .B2(n6278), .A(n6277), .ZN(n6304) );
  OAI22_X1 U7233 ( .A1(n6282), .A2(n6281), .B1(n6280), .B2(n6279), .ZN(n6303)
         );
  AOI22_X1 U7234 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6304), .B1(n6317), 
        .B2(n6303), .ZN(n6283) );
  OAI211_X1 U7235 ( .C1(n6331), .C2(n6307), .A(n6284), .B(n6283), .ZN(U3108)
         );
  AOI22_X1 U7236 ( .A1(n6332), .A2(n6302), .B1(n6334), .B2(n6319), .ZN(n6286)
         );
  AOI22_X1 U7237 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6304), .B1(n6333), 
        .B2(n6303), .ZN(n6285) );
  OAI211_X1 U7238 ( .C1(n6337), .C2(n6307), .A(n6286), .B(n6285), .ZN(U3109)
         );
  AOI22_X1 U7239 ( .A1(n6338), .A2(n6302), .B1(n6340), .B2(n6319), .ZN(n6288)
         );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6304), .B1(n6339), 
        .B2(n6303), .ZN(n6287) );
  OAI211_X1 U7241 ( .C1(n6343), .C2(n6307), .A(n6288), .B(n6287), .ZN(U3110)
         );
  AOI22_X1 U7242 ( .A1(n6344), .A2(n6302), .B1(n6346), .B2(n6319), .ZN(n6290)
         );
  AOI22_X1 U7243 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6304), .B1(n6345), 
        .B2(n6303), .ZN(n6289) );
  OAI211_X1 U7244 ( .C1(n6349), .C2(n6307), .A(n6290), .B(n6289), .ZN(U3111)
         );
  INV_X1 U7245 ( .A(n6307), .ZN(n6298) );
  AOI22_X1 U7246 ( .A1(n6350), .A2(n6302), .B1(n6298), .B2(n6291), .ZN(n6293)
         );
  AOI22_X1 U7247 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6304), .B1(n6351), 
        .B2(n6303), .ZN(n6292) );
  OAI211_X1 U7248 ( .C1(n6294), .C2(n6377), .A(n6293), .B(n6292), .ZN(U3112)
         );
  AOI22_X1 U7249 ( .A1(n6356), .A2(n6302), .B1(n6358), .B2(n6319), .ZN(n6296)
         );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6304), .B1(n6357), 
        .B2(n6303), .ZN(n6295) );
  OAI211_X1 U7251 ( .C1(n6361), .C2(n6307), .A(n6296), .B(n6295), .ZN(U3113)
         );
  AOI22_X1 U7252 ( .A1(n6362), .A2(n6302), .B1(n6298), .B2(n6297), .ZN(n6300)
         );
  AOI22_X1 U7253 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6304), .B1(n6363), 
        .B2(n6303), .ZN(n6299) );
  OAI211_X1 U7254 ( .C1(n6301), .C2(n6377), .A(n6300), .B(n6299), .ZN(U3114)
         );
  AOI22_X1 U7255 ( .A1(n6369), .A2(n6302), .B1(n6373), .B2(n6319), .ZN(n6306)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6304), .B1(n6371), 
        .B2(n6303), .ZN(n6305) );
  OAI211_X1 U7257 ( .C1(n6378), .C2(n6307), .A(n6306), .B(n6305), .ZN(U3115)
         );
  INV_X1 U7258 ( .A(n6308), .ZN(n6314) );
  INV_X1 U7259 ( .A(n6309), .ZN(n6312) );
  INV_X1 U7260 ( .A(n6310), .ZN(n6311) );
  OAI22_X1 U7261 ( .A1(n6314), .A2(n6313), .B1(n6312), .B2(n6311), .ZN(n6370)
         );
  NOR2_X1 U7262 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6315), .ZN(n6368)
         );
  AOI22_X1 U7263 ( .A1(n6317), .A2(n6370), .B1(n6316), .B2(n6368), .ZN(n6330)
         );
  NOR3_X1 U7264 ( .A1(n6319), .A2(n6372), .A3(n6318), .ZN(n6323) );
  OAI22_X1 U7265 ( .A1(n6323), .A2(n6322), .B1(n6321), .B2(n6320), .ZN(n6327)
         );
  NOR2_X1 U7266 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  AOI22_X1 U7267 ( .A1(n6374), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6328), 
        .B2(n6372), .ZN(n6329) );
  OAI211_X1 U7268 ( .C1(n6331), .C2(n6377), .A(n6330), .B(n6329), .ZN(U3116)
         );
  AOI22_X1 U7269 ( .A1(n6333), .A2(n6370), .B1(n6332), .B2(n6368), .ZN(n6336)
         );
  AOI22_X1 U7270 ( .A1(n6374), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6334), 
        .B2(n6372), .ZN(n6335) );
  OAI211_X1 U7271 ( .C1(n6337), .C2(n6377), .A(n6336), .B(n6335), .ZN(U3117)
         );
  AOI22_X1 U7272 ( .A1(n6339), .A2(n6370), .B1(n6338), .B2(n6368), .ZN(n6342)
         );
  AOI22_X1 U7273 ( .A1(n6374), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6340), 
        .B2(n6372), .ZN(n6341) );
  OAI211_X1 U7274 ( .C1(n6343), .C2(n6377), .A(n6342), .B(n6341), .ZN(U3118)
         );
  AOI22_X1 U7275 ( .A1(n6345), .A2(n6370), .B1(n6344), .B2(n6368), .ZN(n6348)
         );
  AOI22_X1 U7276 ( .A1(n6374), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6346), 
        .B2(n6372), .ZN(n6347) );
  OAI211_X1 U7277 ( .C1(n6349), .C2(n6377), .A(n6348), .B(n6347), .ZN(U3119)
         );
  AOI22_X1 U7278 ( .A1(n6351), .A2(n6370), .B1(n6350), .B2(n6368), .ZN(n6354)
         );
  AOI22_X1 U7279 ( .A1(n6374), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6352), 
        .B2(n6372), .ZN(n6353) );
  OAI211_X1 U7280 ( .C1(n6355), .C2(n6377), .A(n6354), .B(n6353), .ZN(U3120)
         );
  AOI22_X1 U7281 ( .A1(n6357), .A2(n6370), .B1(n6356), .B2(n6368), .ZN(n6360)
         );
  AOI22_X1 U7282 ( .A1(n6374), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6358), 
        .B2(n6372), .ZN(n6359) );
  OAI211_X1 U7283 ( .C1(n6361), .C2(n6377), .A(n6360), .B(n6359), .ZN(U3121)
         );
  AOI22_X1 U7284 ( .A1(n6363), .A2(n6370), .B1(n6362), .B2(n6368), .ZN(n6366)
         );
  AOI22_X1 U7285 ( .A1(n6374), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6364), 
        .B2(n6372), .ZN(n6365) );
  OAI211_X1 U7286 ( .C1(n6367), .C2(n6377), .A(n6366), .B(n6365), .ZN(U3122)
         );
  AOI22_X1 U7287 ( .A1(n6371), .A2(n6370), .B1(n6369), .B2(n6368), .ZN(n6376)
         );
  AOI22_X1 U7288 ( .A1(n6374), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6373), 
        .B2(n6372), .ZN(n6375) );
  OAI211_X1 U7289 ( .C1(n6378), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3123)
         );
  INV_X1 U7290 ( .A(n6391), .ZN(n6393) );
  AND3_X1 U7291 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6380), .A3(n6379), 
        .ZN(n6384) );
  NAND2_X1 U7292 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  AOI222_X1 U7293 ( .A1(n6384), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6384), .B2(n6383), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6383), 
        .ZN(n6385) );
  NAND2_X1 U7294 ( .A1(n6665), .A2(n6385), .ZN(n6387) );
  INV_X1 U7295 ( .A(n6385), .ZN(n6386) );
  AOI22_X1 U7296 ( .A1(n6388), .A2(n6387), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6386), .ZN(n6389) );
  AOI21_X1 U7297 ( .B1(n6391), .B2(n6390), .A(n6389), .ZN(n6392) );
  AOI211_X1 U7298 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6393), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6392), .ZN(n6410) );
  INV_X1 U7299 ( .A(n6394), .ZN(n6409) );
  AND3_X1 U7300 ( .A1(n2962), .A2(n6395), .A3(n6406), .ZN(n6402) );
  NAND2_X1 U7301 ( .A1(n6398), .A2(n6397), .ZN(n6401) );
  NAND2_X1 U7302 ( .A1(n6414), .A2(n6399), .ZN(n6400) );
  OAI211_X1 U7303 ( .C1(n6414), .C2(n6402), .A(n6401), .B(n6400), .ZN(n6403)
         );
  INV_X1 U7304 ( .A(n6403), .ZN(n6523) );
  OAI21_X1 U7305 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6404), 
        .ZN(n6405) );
  NAND4_X1 U7306 ( .A1(n6407), .A2(n6523), .A3(n6406), .A4(n6405), .ZN(n6408)
         );
  NOR3_X1 U7307 ( .A1(n6410), .A2(n6409), .A3(n6408), .ZN(n6426) );
  NOR2_X1 U7308 ( .A1(n6514), .A2(n6434), .ZN(n6415) );
  OAI21_X1 U7309 ( .B1(n6412), .B2(n6411), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6413) );
  AOI221_X1 U7310 ( .B1(n6418), .B2(n6419), .C1(n4249), .C2(n6419), .A(n6413), 
        .ZN(n6417) );
  AOI21_X1 U7311 ( .B1(n6415), .B2(n6414), .A(n6417), .ZN(n6416) );
  INV_X1 U7312 ( .A(n6416), .ZN(n6422) );
  OAI221_X1 U7313 ( .B1(n6419), .B2(n6426), .C1(n6419), .C2(n6418), .A(n6417), 
        .ZN(n6513) );
  OAI21_X1 U7314 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4249), .A(n6513), .ZN(
        n6427) );
  NOR2_X1 U7315 ( .A1(n6420), .A2(n6427), .ZN(n6421) );
  MUX2_X1 U7316 ( .A(n6422), .B(n6421), .S(STATE2_REG_0__SCAN_IN), .Z(n6424)
         );
  OAI211_X1 U7317 ( .C1(n6426), .C2(n6425), .A(n6424), .B(n6423), .ZN(U3148)
         );
  NOR2_X1 U7318 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6437) );
  NAND2_X1 U7319 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6427), .ZN(n6432) );
  OAI221_X1 U7320 ( .B1(n6429), .B2(n6428), .C1(n6429), .C2(n4249), .A(n6513), 
        .ZN(n6431) );
  OAI211_X1 U7321 ( .C1(n6437), .C2(n6432), .A(n6431), .B(n6430), .ZN(U3149)
         );
  INV_X1 U7322 ( .A(n6433), .ZN(n6511) );
  OAI211_X1 U7323 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4249), .A(n6511), .B(
        n6434), .ZN(n6436) );
  OAI21_X1 U7324 ( .B1(n6437), .B2(n6436), .A(n6435), .ZN(U3150) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6438), .ZN(U3151) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6438), .ZN(U3152) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6438), .ZN(U3153) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6438), .ZN(U3154) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6438), .ZN(U3155) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6438), .ZN(U3156) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6438), .ZN(U3157) );
  AND2_X1 U7332 ( .A1(n6438), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7333 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6438), .ZN(U3159) );
  AND2_X1 U7334 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6438), .ZN(U3160) );
  AND2_X1 U7335 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6438), .ZN(U3161) );
  AND2_X1 U7336 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6438), .ZN(U3162) );
  AND2_X1 U7337 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6438), .ZN(U3163) );
  AND2_X1 U7338 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6438), .ZN(U3164) );
  AND2_X1 U7339 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6438), .ZN(U3165) );
  AND2_X1 U7340 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6438), .ZN(U3166) );
  AND2_X1 U7341 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6438), .ZN(U3167) );
  AND2_X1 U7342 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6438), .ZN(U3168) );
  AND2_X1 U7343 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6438), .ZN(U3169) );
  AND2_X1 U7344 ( .A1(n6438), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6438), .ZN(U3171) );
  AND2_X1 U7346 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6438), .ZN(U3172) );
  AND2_X1 U7347 ( .A1(n6438), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6438), .ZN(U3174) );
  AND2_X1 U7349 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6438), .ZN(U3175) );
  AND2_X1 U7350 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6438), .ZN(U3176) );
  AND2_X1 U7351 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6438), .ZN(U3177) );
  AND2_X1 U7352 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6438), .ZN(U3178) );
  AND2_X1 U7353 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6438), .ZN(U3179) );
  AND2_X1 U7354 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6438), .ZN(U3180) );
  NAND2_X1 U7355 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6443) );
  NAND2_X1 U7356 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6442) );
  NAND2_X1 U7357 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7358 ( .A1(n6442), .A2(n6450), .ZN(n6439) );
  INV_X1 U7359 ( .A(NA_N), .ZN(n6451) );
  AOI221_X1 U7360 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6451), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6455) );
  AOI21_X1 U7361 ( .B1(n6440), .B2(n6439), .A(n6455), .ZN(n6441) );
  OAI221_X1 U7362 ( .B1(n6537), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6537), 
        .C2(n6443), .A(n6441), .ZN(U3181) );
  INV_X1 U7363 ( .A(n6442), .ZN(n6447) );
  INV_X1 U7364 ( .A(n6443), .ZN(n6444) );
  AOI21_X1 U7365 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6444), .ZN(n6446) );
  OAI211_X1 U7366 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n6450), .ZN(U3182)
         );
  AOI221_X1 U7367 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4249), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6449) );
  AOI221_X1 U7368 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6449), .C2(HOLD), .A(n6448), .ZN(n6456) );
  INV_X1 U7369 ( .A(n6450), .ZN(n6452) );
  NAND4_X1 U7370 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6452), .A4(n6451), .ZN(n6454) );
  NAND3_X1 U7371 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .A3(
        STATE_REG_2__SCAN_IN), .ZN(n6453) );
  OAI211_X1 U7372 ( .C1(n6456), .C2(n6455), .A(n6454), .B(n6453), .ZN(U3183)
         );
  NAND2_X1 U7373 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6537), .ZN(n6503) );
  NOR2_X2 U7374 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6505), .ZN(n6501) );
  AOI22_X1 U7375 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6505), .ZN(n6457) );
  OAI21_X1 U7376 ( .B1(n6584), .B2(n6503), .A(n6457), .ZN(U3184) );
  AOI22_X1 U7377 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6505), .ZN(n6458) );
  OAI21_X1 U7378 ( .B1(n6459), .B2(n6503), .A(n6458), .ZN(U3185) );
  AOI22_X1 U7379 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6505), .ZN(n6460) );
  OAI21_X1 U7380 ( .B1(n6461), .B2(n6503), .A(n6460), .ZN(U3186) );
  AOI22_X1 U7381 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6505), .ZN(n6462) );
  OAI21_X1 U7382 ( .B1(n6463), .B2(n6503), .A(n6462), .ZN(U3187) );
  AOI22_X1 U7383 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6505), .ZN(n6464) );
  OAI21_X1 U7384 ( .B1(n6465), .B2(n6503), .A(n6464), .ZN(U3188) );
  AOI22_X1 U7385 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6505), .ZN(n6466) );
  OAI21_X1 U7386 ( .B1(n6467), .B2(n6503), .A(n6466), .ZN(U3189) );
  AOI22_X1 U7387 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6505), .ZN(n6468) );
  OAI21_X1 U7388 ( .B1(n6469), .B2(n6503), .A(n6468), .ZN(U3190) );
  AOI22_X1 U7389 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6505), .ZN(n6470) );
  OAI21_X1 U7390 ( .B1(n6471), .B2(n6503), .A(n6470), .ZN(U3191) );
  AOI22_X1 U7391 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6505), .ZN(n6472) );
  OAI21_X1 U7392 ( .B1(n5057), .B2(n6503), .A(n6472), .ZN(U3192) );
  INV_X1 U7393 ( .A(n6503), .ZN(n6506) );
  AOI22_X1 U7394 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6505), .ZN(n6473) );
  OAI21_X1 U7395 ( .B1(n6475), .B2(n6508), .A(n6473), .ZN(U3193) );
  AOI22_X1 U7396 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6505), .ZN(n6474) );
  OAI21_X1 U7397 ( .B1(n6475), .B2(n6503), .A(n6474), .ZN(U3194) );
  AOI22_X1 U7398 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6505), .ZN(n6476) );
  OAI21_X1 U7399 ( .B1(n6478), .B2(n6508), .A(n6476), .ZN(U3195) );
  AOI22_X1 U7400 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6505), .ZN(n6477) );
  OAI21_X1 U7401 ( .B1(n6478), .B2(n6503), .A(n6477), .ZN(U3196) );
  AOI222_X1 U7402 ( .A1(n6501), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6505), .C1(REIP_REG_14__SCAN_IN), .C2(
        n6506), .ZN(n6479) );
  INV_X1 U7403 ( .A(n6479), .ZN(U3197) );
  AOI22_X1 U7404 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6505), .ZN(n6480) );
  OAI21_X1 U7405 ( .B1(n6481), .B2(n6503), .A(n6480), .ZN(U3198) );
  AOI22_X1 U7406 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6505), .ZN(n6482) );
  OAI21_X1 U7407 ( .B1(n6667), .B2(n6508), .A(n6482), .ZN(U3199) );
  AOI22_X1 U7408 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6505), .ZN(n6483) );
  OAI21_X1 U7409 ( .B1(n6485), .B2(n6508), .A(n6483), .ZN(U3200) );
  AOI22_X1 U7410 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6505), .ZN(n6484) );
  OAI21_X1 U7411 ( .B1(n6485), .B2(n6503), .A(n6484), .ZN(U3201) );
  AOI22_X1 U7412 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6505), .ZN(n6486) );
  OAI21_X1 U7413 ( .B1(n6487), .B2(n6503), .A(n6486), .ZN(U3202) );
  INV_X1 U7414 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6640) );
  INV_X1 U7415 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6489) );
  OAI222_X1 U7416 ( .A1(n6503), .A2(n6640), .B1(n6489), .B2(n6537), .C1(n6488), 
        .C2(n6508), .ZN(U3203) );
  AOI22_X1 U7417 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6505), .ZN(n6490) );
  OAI21_X1 U7418 ( .B1(n6492), .B2(n6508), .A(n6490), .ZN(U3204) );
  AOI22_X1 U7419 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6505), .ZN(n6491) );
  OAI21_X1 U7420 ( .B1(n6492), .B2(n6503), .A(n6491), .ZN(U3205) );
  AOI22_X1 U7421 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6505), .ZN(n6493) );
  OAI21_X1 U7422 ( .B1(n6494), .B2(n6508), .A(n6493), .ZN(U3206) );
  AOI22_X1 U7423 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6505), .ZN(n6495) );
  OAI21_X1 U7424 ( .B1(n5433), .B2(n6508), .A(n6495), .ZN(U3207) );
  AOI22_X1 U7425 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6505), .ZN(n6496) );
  OAI21_X1 U7426 ( .B1(n5433), .B2(n6503), .A(n6496), .ZN(U3208) );
  AOI22_X1 U7427 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6505), .ZN(n6497) );
  OAI21_X1 U7428 ( .B1(n6498), .B2(n6508), .A(n6497), .ZN(U3209) );
  AOI22_X1 U7429 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6505), .ZN(n6499) );
  OAI21_X1 U7430 ( .B1(n6588), .B2(n6508), .A(n6499), .ZN(U3210) );
  AOI22_X1 U7431 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6505), .ZN(n6500) );
  OAI21_X1 U7432 ( .B1(n6504), .B2(n6508), .A(n6500), .ZN(U3211) );
  AOI22_X1 U7433 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6501), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6505), .ZN(n6502) );
  OAI21_X1 U7434 ( .B1(n6504), .B2(n6503), .A(n6502), .ZN(U3212) );
  AOI22_X1 U7435 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6505), .ZN(n6507) );
  OAI21_X1 U7436 ( .B1(n6509), .B2(n6508), .A(n6507), .ZN(U3213) );
  MUX2_X1 U7437 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6537), .Z(U3445) );
  MUX2_X1 U7438 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6537), .Z(U3446) );
  MUX2_X1 U7439 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6537), .Z(U3447) );
  MUX2_X1 U7440 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6537), .Z(U3448) );
  OAI21_X1 U7441 ( .B1(n6701), .B2(DATAWIDTH_REG_0__SCAN_IN), .A(n6699), .ZN(
        n6510) );
  INV_X1 U7442 ( .A(n6510), .ZN(U3451) );
  OAI211_X1 U7443 ( .C1(n6514), .C2(n6513), .A(n6512), .B(n6511), .ZN(U3453)
         );
  AOI21_X1 U7444 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6515) );
  OAI22_X1 U7445 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6584), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6515), .ZN(n6517) );
  INV_X1 U7446 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6516) );
  AOI22_X1 U7447 ( .A1(n6521), .A2(n6517), .B1(n6516), .B2(n6518), .ZN(U3468)
         );
  NOR2_X1 U7448 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6520) );
  INV_X1 U7449 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6519) );
  AOI22_X1 U7450 ( .A1(n6521), .A2(n6520), .B1(n6519), .B2(n6518), .ZN(U3469)
         );
  INV_X1 U7451 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6582) );
  MUX2_X1 U7452 ( .A(W_R_N_REG_SCAN_IN), .B(n6582), .S(n6537), .Z(U3470) );
  INV_X1 U7453 ( .A(MORE_REG_SCAN_IN), .ZN(n6682) );
  INV_X1 U7454 ( .A(n6524), .ZN(n6522) );
  AOI22_X1 U7455 ( .A1(n6524), .A2(n6523), .B1(n6682), .B2(n6522), .ZN(U3471)
         );
  INV_X1 U7456 ( .A(n6525), .ZN(n6529) );
  OAI211_X1 U7457 ( .C1(READY_N), .C2(n6527), .A(n6526), .B(n6318), .ZN(n6528)
         );
  NOR2_X1 U7458 ( .A1(n6529), .A2(n6528), .ZN(n6536) );
  OAI211_X1 U7459 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6531), .A(n6530), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6533) );
  AOI21_X1 U7460 ( .B1(n6533), .B2(STATE2_REG_0__SCAN_IN), .A(n6532), .ZN(
        n6535) );
  NAND2_X1 U7461 ( .A1(n6536), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6534) );
  OAI21_X1 U7462 ( .B1(n6536), .B2(n6535), .A(n6534), .ZN(U3472) );
  MUX2_X1 U7463 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6537), .Z(U3473) );
  NOR2_X1 U7464 ( .A1(keyinput0), .A2(keyinput45), .ZN(n6538) );
  NAND3_X1 U7465 ( .A1(keyinput14), .A2(keyinput1), .A3(n6538), .ZN(n6543) );
  NAND3_X1 U7466 ( .A1(keyinput40), .A2(keyinput39), .A3(keyinput17), .ZN(
        n6542) );
  NOR3_X1 U7467 ( .A1(keyinput2), .A2(keyinput21), .A3(keyinput44), .ZN(n6540)
         );
  NOR3_X1 U7468 ( .A1(keyinput22), .A2(keyinput20), .A3(keyinput42), .ZN(n6539) );
  NAND4_X1 U7469 ( .A1(keyinput18), .A2(n6540), .A3(keyinput32), .A4(n6539), 
        .ZN(n6541) );
  NOR4_X1 U7470 ( .A1(keyinput29), .A2(n6543), .A3(n6542), .A4(n6541), .ZN(
        n6698) );
  NAND2_X1 U7471 ( .A1(keyinput4), .A2(keyinput61), .ZN(n6544) );
  NOR3_X1 U7472 ( .A1(keyinput26), .A2(keyinput8), .A3(n6544), .ZN(n6549) );
  NOR3_X1 U7473 ( .A1(keyinput52), .A2(keyinput33), .A3(keyinput16), .ZN(n6548) );
  NAND4_X1 U7474 ( .A1(keyinput37), .A2(keyinput9), .A3(keyinput6), .A4(
        keyinput48), .ZN(n6546) );
  NAND2_X1 U7475 ( .A1(keyinput41), .A2(keyinput27), .ZN(n6545) );
  NOR4_X1 U7476 ( .A1(keyinput10), .A2(keyinput47), .A3(n6546), .A4(n6545), 
        .ZN(n6547) );
  NAND4_X1 U7477 ( .A1(n6549), .A2(keyinput46), .A3(n6548), .A4(n6547), .ZN(
        n6564) );
  NAND4_X1 U7478 ( .A1(keyinput23), .A2(keyinput24), .A3(keyinput49), .A4(
        keyinput53), .ZN(n6563) );
  NOR2_X1 U7479 ( .A1(keyinput62), .A2(keyinput50), .ZN(n6554) );
  NAND2_X1 U7480 ( .A1(keyinput63), .A2(keyinput13), .ZN(n6552) );
  INV_X1 U7481 ( .A(keyinput5), .ZN(n6550) );
  NAND4_X1 U7482 ( .A1(keyinput19), .A2(keyinput55), .A3(keyinput31), .A4(
        n6550), .ZN(n6551) );
  NOR4_X1 U7483 ( .A1(keyinput15), .A2(keyinput35), .A3(n6552), .A4(n6551), 
        .ZN(n6553) );
  NAND4_X1 U7484 ( .A1(keyinput28), .A2(keyinput38), .A3(n6554), .A4(n6553), 
        .ZN(n6562) );
  NOR2_X1 U7485 ( .A1(keyinput56), .A2(keyinput11), .ZN(n6560) );
  NAND2_X1 U7486 ( .A1(keyinput54), .A2(keyinput59), .ZN(n6558) );
  NOR3_X1 U7487 ( .A1(keyinput51), .A2(keyinput57), .A3(keyinput3), .ZN(n6556)
         );
  NOR3_X1 U7488 ( .A1(keyinput58), .A2(keyinput36), .A3(keyinput30), .ZN(n6555) );
  NAND4_X1 U7489 ( .A1(keyinput7), .A2(n6556), .A3(keyinput43), .A4(n6555), 
        .ZN(n6557) );
  NOR4_X1 U7490 ( .A1(keyinput12), .A2(keyinput34), .A3(n6558), .A4(n6557), 
        .ZN(n6559) );
  NAND4_X1 U7491 ( .A1(keyinput25), .A2(keyinput60), .A3(n6560), .A4(n6559), 
        .ZN(n6561) );
  NOR4_X1 U7492 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n6697)
         );
  INV_X1 U7493 ( .A(keyinput37), .ZN(n6566) );
  AOI22_X1 U7494 ( .A1(n6567), .A2(keyinput9), .B1(DATAO_REG_26__SCAN_IN), 
        .B2(n6566), .ZN(n6565) );
  OAI221_X1 U7495 ( .B1(n6567), .B2(keyinput9), .C1(n6566), .C2(
        DATAO_REG_26__SCAN_IN), .A(n6565), .ZN(n6579) );
  INV_X1 U7496 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U7497 ( .A1(n6570), .A2(keyinput6), .B1(n6569), .B2(keyinput48), 
        .ZN(n6568) );
  OAI221_X1 U7498 ( .B1(n6570), .B2(keyinput6), .C1(n6569), .C2(keyinput48), 
        .A(n6568), .ZN(n6578) );
  INV_X1 U7499 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6573) );
  AOI22_X1 U7500 ( .A1(n6573), .A2(keyinput61), .B1(keyinput8), .B2(n6572), 
        .ZN(n6571) );
  OAI221_X1 U7501 ( .B1(n6573), .B2(keyinput61), .C1(n6572), .C2(keyinput8), 
        .A(n6571), .ZN(n6577) );
  INV_X1 U7502 ( .A(keyinput4), .ZN(n6575) );
  AOI22_X1 U7503 ( .A1(n5216), .A2(keyinput26), .B1(ADDRESS_REG_19__SCAN_IN), 
        .B2(n6575), .ZN(n6574) );
  OAI221_X1 U7504 ( .B1(n5216), .B2(keyinput26), .C1(n6575), .C2(
        ADDRESS_REG_19__SCAN_IN), .A(n6574), .ZN(n6576) );
  NOR4_X1 U7505 ( .A1(n6579), .A2(n6578), .A3(n6577), .A4(n6576), .ZN(n6628)
         );
  INV_X1 U7506 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6581) );
  AOI22_X1 U7507 ( .A1(n6582), .A2(keyinput41), .B1(n6581), .B2(keyinput47), 
        .ZN(n6580) );
  OAI221_X1 U7508 ( .B1(n6582), .B2(keyinput41), .C1(n6581), .C2(keyinput47), 
        .A(n6580), .ZN(n6595) );
  INV_X1 U7509 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6585) );
  AOI22_X1 U7510 ( .A1(n6585), .A2(keyinput27), .B1(keyinput10), .B2(n6584), 
        .ZN(n6583) );
  OAI221_X1 U7511 ( .B1(n6585), .B2(keyinput27), .C1(n6584), .C2(keyinput10), 
        .A(n6583), .ZN(n6594) );
  INV_X1 U7512 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7513 ( .A1(n6588), .A2(keyinput52), .B1(n6587), .B2(keyinput33), 
        .ZN(n6586) );
  OAI221_X1 U7514 ( .B1(n6588), .B2(keyinput52), .C1(n6587), .C2(keyinput33), 
        .A(n6586), .ZN(n6593) );
  AOI22_X1 U7515 ( .A1(n6591), .A2(keyinput46), .B1(n6590), .B2(keyinput16), 
        .ZN(n6589) );
  OAI221_X1 U7516 ( .B1(n6591), .B2(keyinput46), .C1(n6590), .C2(keyinput16), 
        .A(n6589), .ZN(n6592) );
  NOR4_X1 U7517 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6627)
         );
  INV_X1 U7518 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6598) );
  INV_X1 U7519 ( .A(keyinput62), .ZN(n6597) );
  AOI22_X1 U7520 ( .A1(n6598), .A2(keyinput28), .B1(ADDRESS_REG_22__SCAN_IN), 
        .B2(n6597), .ZN(n6596) );
  OAI221_X1 U7521 ( .B1(n6598), .B2(keyinput28), .C1(n6597), .C2(
        ADDRESS_REG_22__SCAN_IN), .A(n6596), .ZN(n6610) );
  INV_X1 U7522 ( .A(DATAI_17_), .ZN(n6600) );
  AOI22_X1 U7523 ( .A1(n6601), .A2(keyinput50), .B1(keyinput38), .B2(n6600), 
        .ZN(n6599) );
  OAI221_X1 U7524 ( .B1(n6601), .B2(keyinput50), .C1(n6600), .C2(keyinput38), 
        .A(n6599), .ZN(n6609) );
  INV_X1 U7525 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6603) );
  AOI22_X1 U7526 ( .A1(n6000), .A2(keyinput23), .B1(n6603), .B2(keyinput24), 
        .ZN(n6602) );
  OAI221_X1 U7527 ( .B1(n6000), .B2(keyinput23), .C1(n6603), .C2(keyinput24), 
        .A(n6602), .ZN(n6608) );
  INV_X1 U7528 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6606) );
  INV_X1 U7529 ( .A(keyinput53), .ZN(n6605) );
  AOI22_X1 U7530 ( .A1(n6606), .A2(keyinput49), .B1(HOLD), .B2(n6605), .ZN(
        n6604) );
  OAI221_X1 U7531 ( .B1(n6606), .B2(keyinput49), .C1(n6605), .C2(HOLD), .A(
        n6604), .ZN(n6607) );
  NOR4_X1 U7532 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n6626)
         );
  INV_X1 U7533 ( .A(keyinput55), .ZN(n6612) );
  AOI22_X1 U7534 ( .A1(n6613), .A2(keyinput31), .B1(DATAWIDTH_REG_12__SCAN_IN), 
        .B2(n6612), .ZN(n6611) );
  OAI221_X1 U7535 ( .B1(n6613), .B2(keyinput31), .C1(n6612), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6611), .ZN(n6624) );
  INV_X1 U7536 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U7537 ( .A1(n6615), .A2(keyinput63), .B1(keyinput15), .B2(n4226), 
        .ZN(n6614) );
  OAI221_X1 U7538 ( .B1(n6615), .B2(keyinput63), .C1(n4226), .C2(keyinput15), 
        .A(n6614), .ZN(n6623) );
  INV_X1 U7539 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6617) );
  AOI22_X1 U7540 ( .A1(n6618), .A2(keyinput5), .B1(n6617), .B2(keyinput19), 
        .ZN(n6616) );
  OAI221_X1 U7541 ( .B1(n6618), .B2(keyinput5), .C1(n6617), .C2(keyinput19), 
        .A(n6616), .ZN(n6622) );
  XOR2_X1 U7542 ( .A(n4077), .B(keyinput35), .Z(n6620) );
  XNOR2_X1 U7543 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput13), .ZN(
        n6619) );
  NAND2_X1 U7544 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NOR4_X1 U7545 ( .A1(n6624), .A2(n6623), .A3(n6622), .A4(n6621), .ZN(n6625)
         );
  NAND4_X1 U7546 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(n6696)
         );
  INV_X1 U7547 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6630) );
  INV_X1 U7548 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6634) );
  INV_X1 U7549 ( .A(keyinput21), .ZN(n6633) );
  AOI22_X1 U7550 ( .A1(n6634), .A2(keyinput2), .B1(ADDRESS_REG_24__SCAN_IN), 
        .B2(n6633), .ZN(n6632) );
  OAI221_X1 U7551 ( .B1(n6634), .B2(keyinput2), .C1(n6633), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n6632), .ZN(n6643) );
  INV_X1 U7552 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6636) );
  AOI22_X1 U7553 ( .A1(n6637), .A2(keyinput20), .B1(n6636), .B2(keyinput42), 
        .ZN(n6635) );
  OAI221_X1 U7554 ( .B1(n6637), .B2(keyinput20), .C1(n6636), .C2(keyinput42), 
        .A(n6635), .ZN(n6642) );
  AOI22_X1 U7555 ( .A1(n6640), .A2(keyinput32), .B1(n6639), .B2(keyinput22), 
        .ZN(n6638) );
  OAI221_X1 U7556 ( .B1(n6640), .B2(keyinput32), .C1(n6639), .C2(keyinput22), 
        .A(n6638), .ZN(n6641) );
  NOR4_X1 U7557 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6694)
         );
  INV_X1 U7558 ( .A(keyinput0), .ZN(n6646) );
  AOI22_X1 U7559 ( .A1(n6647), .A2(keyinput45), .B1(NA_N), .B2(n6646), .ZN(
        n6645) );
  OAI221_X1 U7560 ( .B1(n6647), .B2(keyinput45), .C1(n6646), .C2(NA_N), .A(
        n6645), .ZN(n6659) );
  INV_X1 U7561 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7562 ( .A1(n6650), .A2(keyinput1), .B1(n6649), .B2(keyinput14), 
        .ZN(n6648) );
  OAI221_X1 U7563 ( .B1(n6650), .B2(keyinput1), .C1(n6649), .C2(keyinput14), 
        .A(n6648), .ZN(n6658) );
  AOI22_X1 U7564 ( .A1(n5998), .A2(keyinput39), .B1(n6652), .B2(keyinput17), 
        .ZN(n6651) );
  OAI221_X1 U7565 ( .B1(n5998), .B2(keyinput39), .C1(n6652), .C2(keyinput17), 
        .A(n6651), .ZN(n6657) );
  INV_X1 U7566 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6655) );
  INV_X1 U7567 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7568 ( .A1(n6655), .A2(keyinput29), .B1(n6654), .B2(keyinput40), 
        .ZN(n6653) );
  OAI221_X1 U7569 ( .B1(n6655), .B2(keyinput29), .C1(n6654), .C2(keyinput40), 
        .A(n6653), .ZN(n6656) );
  NOR4_X1 U7570 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6693)
         );
  INV_X1 U7571 ( .A(keyinput43), .ZN(n6661) );
  AOI22_X1 U7572 ( .A1(n6662), .A2(keyinput30), .B1(DATAWIDTH_REG_9__SCAN_IN), 
        .B2(n6661), .ZN(n6660) );
  OAI221_X1 U7573 ( .B1(n6662), .B2(keyinput30), .C1(n6661), .C2(
        DATAWIDTH_REG_9__SCAN_IN), .A(n6660), .ZN(n6675) );
  INV_X1 U7574 ( .A(keyinput58), .ZN(n6664) );
  AOI22_X1 U7575 ( .A1(n6665), .A2(keyinput36), .B1(ADDRESS_REG_13__SCAN_IN), 
        .B2(n6664), .ZN(n6663) );
  OAI221_X1 U7576 ( .B1(n6665), .B2(keyinput36), .C1(n6664), .C2(
        ADDRESS_REG_13__SCAN_IN), .A(n6663), .ZN(n6674) );
  INV_X1 U7577 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6668) );
  AOI22_X1 U7578 ( .A1(n6668), .A2(keyinput12), .B1(keyinput34), .B2(n6667), 
        .ZN(n6666) );
  OAI221_X1 U7579 ( .B1(n6668), .B2(keyinput12), .C1(n6667), .C2(keyinput34), 
        .A(n6666), .ZN(n6673) );
  INV_X1 U7580 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7581 ( .A1(n6671), .A2(keyinput54), .B1(keyinput59), .B2(n6670), 
        .ZN(n6669) );
  OAI221_X1 U7582 ( .B1(n6671), .B2(keyinput54), .C1(n6670), .C2(keyinput59), 
        .A(n6669), .ZN(n6672) );
  NOR4_X1 U7583 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6692)
         );
  INV_X1 U7584 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6678) );
  INV_X1 U7585 ( .A(keyinput3), .ZN(n6677) );
  AOI22_X1 U7586 ( .A1(n6678), .A2(keyinput7), .B1(DATAWIDTH_REG_24__SCAN_IN), 
        .B2(n6677), .ZN(n6676) );
  OAI221_X1 U7587 ( .B1(n6678), .B2(keyinput7), .C1(n6677), .C2(
        DATAWIDTH_REG_24__SCAN_IN), .A(n6676), .ZN(n6690) );
  INV_X1 U7588 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6680) );
  AOI22_X1 U7589 ( .A1(n3832), .A2(keyinput51), .B1(n6680), .B2(keyinput57), 
        .ZN(n6679) );
  OAI221_X1 U7590 ( .B1(n3832), .B2(keyinput51), .C1(n6680), .C2(keyinput57), 
        .A(n6679), .ZN(n6689) );
  INV_X1 U7591 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7592 ( .A1(n6683), .A2(keyinput11), .B1(keyinput60), .B2(n6682), 
        .ZN(n6681) );
  OAI221_X1 U7593 ( .B1(n6683), .B2(keyinput11), .C1(n6682), .C2(keyinput60), 
        .A(n6681), .ZN(n6688) );
  INV_X1 U7594 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6686) );
  AOI22_X1 U7595 ( .A1(n6686), .A2(keyinput56), .B1(n6685), .B2(keyinput25), 
        .ZN(n6684) );
  OAI221_X1 U7596 ( .B1(n6686), .B2(keyinput56), .C1(n6685), .C2(keyinput25), 
        .A(n6684), .ZN(n6687) );
  NOR4_X1 U7597 ( .A1(n6690), .A2(n6689), .A3(n6688), .A4(n6687), .ZN(n6691)
         );
  NAND4_X1 U7598 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .ZN(n6695)
         );
  AOI211_X1 U7599 ( .C1(n6698), .C2(n6697), .A(n6696), .B(n6695), .ZN(n6703)
         );
  OAI21_X1 U7600 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6702) );
  XOR2_X1 U7601 ( .A(n6703), .B(n6702), .Z(U3452) );
  AND2_X2 U3896 ( .A1(n5145), .A2(n3118), .ZN(n3329) );
  BUF_X2 U3430 ( .A(n3904), .Z(n2975) );
  CLKBUF_X1 U3424 ( .A(n3879), .Z(n3819) );
endmodule

