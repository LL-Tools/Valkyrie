

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9715, n9716, n9717, n9719, n9720, n9721, n9722, n9723, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760;

  NAND2_X1 U11160 ( .A1(n13151), .A2(n13727), .ZN(n15969) );
  OR2_X1 U11161 ( .A1(n12851), .A2(n12985), .ZN(n12972) );
  NOR2_X1 U11162 ( .A1(n13040), .A2(n13119), .ZN(n13120) );
  INV_X2 U11163 ( .A(n12822), .ZN(n12994) );
  CLKBUF_X2 U11164 ( .A(n11740), .Z(n9723) );
  INV_X1 U11165 ( .A(n17550), .ZN(n18410) );
  NAND2_X1 U11166 ( .A1(n12144), .A2(n12143), .ZN(n12146) );
  INV_X1 U11167 ( .A(n12624), .ZN(n12793) );
  NAND2_X2 U11168 ( .A1(n10987), .A2(n10991), .ZN(n11133) );
  NAND2_X1 U11169 ( .A1(n12612), .A2(n12991), .ZN(n12620) );
  AND2_X2 U11170 ( .A1(n9747), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12273) );
  BUF_X1 U11171 ( .A(n11769), .Z(n18517) );
  AND2_X2 U11172 ( .A1(n9748), .A2(n11984), .ZN(n12278) );
  CLKBUF_X1 U11173 ( .A(n10931), .Z(n11670) );
  CLKBUF_X2 U11174 ( .A(n10818), .Z(n11700) );
  INV_X2 U11175 ( .A(n18505), .ZN(n18611) );
  CLKBUF_X2 U11176 ( .A(n12125), .Z(n14904) );
  INV_X2 U11177 ( .A(n11836), .ZN(n18505) );
  AND2_X2 U11178 ( .A1(n14788), .A2(n11984), .ZN(n14803) );
  INV_X1 U11179 ( .A(n18261), .ZN(n17549) );
  CLKBUF_X1 U11180 ( .A(n12080), .Z(n14609) );
  BUF_X1 U11181 ( .A(n12090), .Z(n20400) );
  AND4_X1 U11182 ( .A1(n10707), .A2(n10706), .A3(n10705), .A4(n10704), .ZN(
        n10708) );
  INV_X1 U11183 ( .A(n18261), .ZN(n18612) );
  AND2_X1 U11184 ( .A1(n10524), .A2(n14113), .ZN(n11836) );
  INV_X2 U11185 ( .A(n10540), .ZN(n11843) );
  AND2_X1 U11187 ( .A1(n10702), .A2(n16091), .ZN(n10960) );
  AND3_X1 U11188 ( .A1(n14997), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n15095), .ZN(n11258) );
  AND2_X1 U11189 ( .A1(n16091), .A2(n10701), .ZN(n10961) );
  AND2_X2 U11190 ( .A1(n10346), .A2(n10703), .ZN(n10837) );
  INV_X4 U11191 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11984) );
  INV_X1 U11192 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14209) );
  CLKBUF_X1 U11193 ( .A(n14021), .Z(n9715) );
  NOR2_X1 U11194 ( .A1(n15585), .A2(n17666), .ZN(n14021) );
  CLKBUF_X1 U11195 ( .A(n14023), .Z(n9716) );
  NOR2_X1 U11196 ( .A1(n17666), .A2(n14022), .ZN(n14023) );
  CLKBUF_X3 U11198 ( .A(n10834), .Z(n11650) );
  AND2_X1 U11199 ( .A1(n12997), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12116) );
  AND2_X1 U11200 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12187) );
  INV_X1 U11201 ( .A(n11711), .ZN(n13406) );
  BUF_X1 U11202 ( .A(n12419), .Z(n9725) );
  AND2_X1 U11203 ( .A1(n10521), .A2(n10524), .ZN(n11769) );
  OR2_X1 U11204 ( .A1(n14045), .A2(n13032), .ZN(n13124) );
  AND4_X2 U11205 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n13032) );
  NAND2_X1 U11206 ( .A1(n15001), .A2(n16091), .ZN(n10723) );
  NAND2_X1 U11207 ( .A1(n12968), .A2(n12972), .ZN(n12992) );
  NAND2_X1 U11208 ( .A1(n12901), .A2(n12972), .ZN(n12910) );
  INV_X1 U11209 ( .A(n12547), .ZN(n12557) );
  AND2_X1 U11210 ( .A1(n12176), .A2(n12175), .ZN(n20709) );
  AND2_X1 U11213 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14113) );
  AOI21_X1 U11214 ( .B1(n13869), .B2(n13868), .A(n11105), .ZN(n14372) );
  OR3_X1 U11215 ( .A1(n21069), .A2(n12388), .A3(n15163), .ZN(n20260) );
  NOR2_X1 U11216 ( .A1(n16727), .A2(n16726), .ZN(n16725) );
  NAND2_X1 U11217 ( .A1(n13769), .A2(n12089), .ZN(n12609) );
  INV_X2 U11218 ( .A(n12091), .ZN(n9874) );
  INV_X1 U11219 ( .A(n19390), .ZN(n19406) );
  INV_X1 U11220 ( .A(n21137), .ZN(n21130) );
  INV_X1 U11221 ( .A(n15644), .ZN(n15637) );
  XNOR2_X1 U11222 ( .A(n10095), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13469) );
  NOR2_X2 U11224 ( .A1(n14075), .A2(n14074), .ZN(n16155) );
  XNOR2_X1 U11225 ( .A(n10413), .B(n12158), .ZN(n13834) );
  NOR2_X1 U11226 ( .A1(n17731), .A2(n17732), .ZN(n20364) );
  AND2_X1 U11227 ( .A1(n14707), .A2(n14709), .ZN(n17397) );
  NAND2_X1 U11228 ( .A1(n21030), .A2(n20368), .ZN(n20813) );
  NOR2_X1 U11229 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17942), .ZN(n17913) );
  CLKBUF_X2 U11230 ( .A(n10512), .Z(n18132) );
  INV_X1 U11231 ( .A(n19178), .ZN(n19128) );
  INV_X2 U11232 ( .A(n21185), .ZN(n21170) );
  OR2_X1 U11233 ( .A1(n17602), .A2(n21089), .ZN(n21094) );
  OAI21_X1 U11234 ( .B1(n13841), .B2(n13842), .A(n13948), .ZN(n21036) );
  OR2_X1 U11235 ( .A1(n19959), .A2(n19976), .ZN(n17853) );
  AND2_X1 U11236 ( .A1(n10338), .A2(n10337), .ZN(n13499) );
  OR2_X1 U11237 ( .A1(n17853), .A2(n20089), .ZN(n19210) );
  AND2_X2 U11238 ( .A1(n12455), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9747) );
  AND2_X2 U11239 ( .A1(n12455), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9748) );
  NAND2_X4 U11240 ( .A1(n11987), .A2(n11986), .ZN(n12602) );
  AND2_X1 U11241 ( .A1(n9890), .A2(n12859), .ZN(n9717) );
  OR3_X4 U11242 ( .A1(n19095), .A2(n19055), .A3(n10325), .ZN(n18954) );
  NOR2_X2 U11243 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18001), .ZN(n17989) );
  NAND2_X2 U11244 ( .A1(n12374), .A2(n12373), .ZN(n17067) );
  XNOR2_X1 U11245 ( .A(n9886), .B(n17368), .ZN(n17365) );
  NOR2_X4 U11246 ( .A1(n10503), .A2(n10481), .ZN(n10507) );
  NAND2_X2 U11247 ( .A1(n11964), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10503) );
  XNOR2_X2 U11248 ( .A(n11878), .B(n11876), .ZN(n19188) );
  NAND4_X2 U11249 ( .A1(n10162), .A2(n10160), .A3(n10161), .A4(n9923), .ZN(
        n10941) );
  OAI21_X2 U11250 ( .B1(n13354), .B2(n13355), .A(n10012), .ZN(n9885) );
  NAND2_X2 U11251 ( .A1(n10329), .A2(n10327), .ZN(n11878) );
  XNOR2_X2 U11252 ( .A(n12371), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17084) );
  AND2_X1 U11253 ( .A1(n15011), .A2(n10702), .ZN(n10818) );
  AND3_X1 U11254 ( .A1(n10009), .A2(n10316), .A3(n10317), .ZN(n12318) );
  NAND3_X2 U11255 ( .A1(n10112), .A2(n14111), .A3(n13924), .ZN(n18440) );
  AND2_X2 U11256 ( .A1(n10693), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10703) );
  BUF_X4 U11257 ( .A(n18230), .Z(n11841) );
  NOR3_X2 U11258 ( .A1(n17151), .A2(n17152), .A3(n13259), .ZN(n17137) );
  NOR2_X2 U11259 ( .A1(n14045), .A2(n10861), .ZN(n10878) );
  BUF_X4 U11261 ( .A(n11623), .Z(n9719) );
  INV_X1 U11262 ( .A(n10834), .ZN(n11623) );
  BUF_X4 U11263 ( .A(n11842), .Z(n18439) );
  NAND2_X1 U11264 ( .A1(n12090), .A2(n12089), .ZN(n12095) );
  INV_X1 U11265 ( .A(n12090), .ZN(n13769) );
  AND2_X1 U11266 ( .A1(n10346), .A2(n16091), .ZN(n11004) );
  XNOR2_X1 U11267 ( .A(n11077), .B(n11076), .ZN(n13782) );
  AND2_X2 U11268 ( .A1(n17366), .A2(n17365), .ZN(n13491) );
  BUF_X1 U11269 ( .A(n11258), .Z(n9721) );
  CLKBUF_X1 U11271 ( .A(n10846), .Z(n9722) );
  NOR2_X1 U11272 ( .A1(n21077), .A2(n12605), .ZN(n12122) );
  AOI22_X2 U11273 ( .A1(n20638), .A2(n20637), .B1(n20636), .B2(n20864), .ZN(
        n20666) );
  INV_X4 U11274 ( .A(n18258), .ZN(n18251) );
  AOI21_X2 U11275 ( .B1(n10494), .B2(n10201), .A(n10199), .ZN(n17969) );
  OAI21_X2 U11276 ( .B1(n10068), .B2(n10065), .A(n10064), .ZN(n14740) );
  NAND2_X2 U11278 ( .A1(n9733), .A2(n19061), .ZN(n10482) );
  NOR2_X4 U11279 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10702) );
  NAND2_X1 U11280 ( .A1(n11086), .A2(n14045), .ZN(n13144) );
  NOR2_X2 U11281 ( .A1(n19120), .A2(n19110), .ZN(n19102) );
  OR2_X1 U11283 ( .A1(n14719), .A2(n14718), .ZN(n10154) );
  AND2_X1 U11284 ( .A1(n13251), .A2(n9742), .ZN(n16901) );
  AND2_X1 U11285 ( .A1(n17244), .A2(n10174), .ZN(n14719) );
  AND2_X1 U11286 ( .A1(n14711), .A2(n14710), .ZN(n17244) );
  NAND2_X1 U11287 ( .A1(n10169), .A2(n9786), .ZN(n9947) );
  NAND2_X1 U11288 ( .A1(n14900), .A2(n14899), .ZN(n14905) );
  AND2_X1 U11289 ( .A1(n19039), .A2(n13233), .ZN(n18965) );
  NAND2_X1 U11290 ( .A1(n10086), .A2(n12318), .ZN(n12347) );
  AND2_X2 U11291 ( .A1(n15203), .A2(n15202), .ZN(n21185) );
  NAND2_X1 U11292 ( .A1(n11884), .A2(n19174), .ZN(n18963) );
  INV_X1 U11293 ( .A(n12318), .ZN(n9895) );
  INV_X1 U11294 ( .A(n14127), .ZN(n12507) );
  NAND2_X1 U11295 ( .A1(n11042), .A2(n11043), .ZN(n11126) );
  INV_X2 U11296 ( .A(n15664), .ZN(n15831) );
  XNOR2_X1 U11297 ( .A(n11104), .B(n13041), .ZN(n13869) );
  CLKBUF_X2 U11298 ( .A(n15664), .Z(n15840) );
  CLKBUF_X1 U11299 ( .A(n13430), .Z(n15618) );
  OR2_X1 U11300 ( .A1(n9905), .A2(n9737), .ZN(n12208) );
  NAND2_X1 U11301 ( .A1(n13841), .A2(n13842), .ZN(n13948) );
  OR2_X1 U11302 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  OR2_X1 U11303 ( .A1(n11882), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11883) );
  AND2_X1 U11304 ( .A1(n13024), .A2(n14679), .ZN(n13151) );
  NAND2_X1 U11305 ( .A1(n12178), .A2(n12174), .ZN(n14594) );
  AND2_X1 U11306 ( .A1(n12178), .A2(n12175), .ZN(n9880) );
  AND2_X1 U11307 ( .A1(n12178), .A2(n12171), .ZN(n14396) );
  INV_X1 U11308 ( .A(n19177), .ZN(n18981) );
  CLKBUF_X2 U11309 ( .A(n13834), .Z(n16661) );
  AND2_X1 U11310 ( .A1(n9964), .A2(n9963), .ZN(n12998) );
  AND2_X1 U11311 ( .A1(n10090), .A2(n9835), .ZN(n13997) );
  NAND3_X1 U11312 ( .A1(n17536), .A2(n20087), .A3(n17535), .ZN(n18644) );
  OR2_X1 U11313 ( .A1(n11865), .A2(n11927), .ZN(n11870) );
  BUF_X2 U11314 ( .A(n18178), .Z(n9750) );
  NOR2_X1 U11315 ( .A1(n10507), .A2(n10509), .ZN(n10510) );
  NAND2_X1 U11316 ( .A1(n19493), .A2(n20089), .ZN(n11919) );
  NAND3_X1 U11317 ( .A1(n19500), .A2(n19508), .A3(n19515), .ZN(n10649) );
  INV_X4 U11318 ( .A(n19521), .ZN(n18697) );
  INV_X4 U11319 ( .A(n14904), .ZN(n21078) );
  AND2_X1 U11320 ( .A1(n10878), .A2(n10881), .ZN(n10426) );
  AND2_X1 U11321 ( .A1(n10546), .A2(n10545), .ZN(n19521) );
  CLKBUF_X2 U11322 ( .A(n10868), .Z(n14051) );
  AND2_X1 U11323 ( .A1(n13409), .A2(n15557), .ZN(n13134) );
  INV_X1 U11324 ( .A(n13032), .ZN(n10883) );
  NAND2_X2 U11326 ( .A1(n10479), .A2(n9776), .ZN(n14057) );
  AND4_X1 U11327 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10709) );
  BUF_X2 U11328 ( .A(n10923), .Z(n11701) );
  CLKBUF_X2 U11329 ( .A(n11012), .Z(n11628) );
  AND2_X2 U11330 ( .A1(n18058), .A2(n19106), .ZN(n19061) );
  INV_X1 U11331 ( .A(n10833), .ZN(n10923) );
  INV_X2 U11332 ( .A(n18498), .ZN(n9726) );
  CLKBUF_X2 U11333 ( .A(n11004), .Z(n11655) );
  CLKBUF_X2 U11334 ( .A(n10808), .Z(n11606) );
  INV_X2 U11336 ( .A(n18606), .ZN(n18592) );
  CLKBUF_X2 U11337 ( .A(n18230), .Z(n17545) );
  BUF_X4 U11338 ( .A(n18317), .Z(n18614) );
  CLKBUF_X2 U11339 ( .A(n10960), .Z(n11521) );
  CLKBUF_X2 U11340 ( .A(n10961), .Z(n11629) );
  AND2_X2 U11341 ( .A1(n10346), .A2(n15011), .ZN(n10808) );
  AND2_X2 U11342 ( .A1(n12043), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12353) );
  CLKBUF_X1 U11343 ( .A(n12043), .Z(n9727) );
  AND2_X1 U11344 ( .A1(n10093), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10346) );
  INV_X4 U11345 ( .A(n18440), .ZN(n9728) );
  AOI21_X1 U11347 ( .B1(n10151), .B2(n14718), .A(n10149), .ZN(n10148) );
  AND2_X1 U11348 ( .A1(n9962), .A2(n9961), .ZN(n17162) );
  AOI21_X1 U11349 ( .B1(n14674), .B2(n17719), .A(n10197), .ZN(n14676) );
  NAND2_X1 U11350 ( .A1(n9904), .A2(n17168), .ZN(n17174) );
  AOI21_X1 U11351 ( .B1(n13286), .B2(n13442), .A(n13285), .ZN(n16943) );
  AOI21_X1 U11352 ( .B1(n17146), .B2(n17719), .A(n16880), .ZN(n16881) );
  XNOR2_X1 U11353 ( .A(n13359), .B(n13358), .ZN(n14674) );
  AOI21_X1 U11354 ( .B1(n10037), .B2(n10356), .A(n10036), .ZN(n16958) );
  AND2_X1 U11355 ( .A1(n10354), .A2(n10351), .ZN(n13283) );
  NAND2_X1 U11356 ( .A1(n10446), .A2(n16879), .ZN(n16880) );
  OAI21_X1 U11357 ( .B1(n16907), .B2(n16871), .A(n16905), .ZN(n10087) );
  NOR2_X1 U11358 ( .A1(n13268), .A2(n13267), .ZN(n13269) );
  AND2_X1 U11359 ( .A1(n13362), .A2(n13363), .ZN(n9949) );
  OAI21_X1 U11360 ( .B1(n9947), .B2(n9946), .A(n9944), .ZN(n9943) );
  NAND2_X1 U11361 ( .A1(n17067), .A2(n17068), .ZN(n10080) );
  OAI21_X1 U11362 ( .B1(n15182), .B2(n17098), .A(n14675), .ZN(n10197) );
  AND2_X1 U11363 ( .A1(n9909), .A2(n9908), .ZN(n16690) );
  OR2_X1 U11364 ( .A1(n16447), .A2(n16464), .ZN(n17159) );
  NAND2_X1 U11365 ( .A1(n10034), .A2(n15840), .ZN(n10035) );
  NAND2_X1 U11366 ( .A1(n9974), .A2(n19174), .ZN(n17426) );
  XNOR2_X1 U11367 ( .A(n13361), .B(n13360), .ZN(n15182) );
  NAND2_X1 U11368 ( .A1(n9992), .A2(n9991), .ZN(n15674) );
  AND2_X1 U11369 ( .A1(n15695), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15704) );
  AND2_X1 U11370 ( .A1(n11169), .A2(n9937), .ZN(n15696) );
  AND2_X2 U11371 ( .A1(n16484), .A2(n9828), .ZN(n13361) );
  NAND2_X1 U11372 ( .A1(n12846), .A2(n17069), .ZN(n10070) );
  NAND2_X1 U11373 ( .A1(n13491), .A2(n10072), .ZN(n10071) );
  INV_X1 U11374 ( .A(n15373), .ZN(n10442) );
  XNOR2_X1 U11375 ( .A(n12375), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17068) );
  NAND2_X1 U11376 ( .A1(n10406), .A2(n10410), .ZN(n17105) );
  NOR3_X1 U11377 ( .A1(n10051), .A2(n10050), .A3(n10047), .ZN(n15222) );
  NAND2_X1 U11378 ( .A1(n12288), .A2(n20363), .ZN(n10079) );
  NAND2_X1 U11379 ( .A1(n9950), .A2(n17114), .ZN(n9897) );
  OR2_X1 U11380 ( .A1(n12376), .A2(n12994), .ZN(n12375) );
  NAND2_X1 U11381 ( .A1(n12845), .A2(n16620), .ZN(n17069) );
  NAND2_X1 U11382 ( .A1(n10392), .A2(n9830), .ZN(n16707) );
  OR2_X1 U11383 ( .A1(n16725), .A2(n10394), .ZN(n10392) );
  AOI211_X1 U11384 ( .C1(n17583), .C2(n17501), .A(n17500), .B(n17499), .ZN(
        n17502) );
  NAND2_X1 U11385 ( .A1(n17131), .A2(n12994), .ZN(n12826) );
  NAND2_X1 U11386 ( .A1(n17890), .A2(n10506), .ZN(n17891) );
  AND2_X1 U11387 ( .A1(n10096), .A2(n9784), .ZN(n15769) );
  NAND2_X1 U11388 ( .A1(n9895), .A2(n10176), .ZN(n10013) );
  OR2_X2 U11389 ( .A1(n15203), .A2(n15201), .ZN(n21137) );
  XNOR2_X1 U11390 ( .A(n10267), .B(n13195), .ZN(n15212) );
  NOR2_X2 U11391 ( .A1(n20671), .A2(n20539), .ZN(n20857) );
  INV_X1 U11392 ( .A(n13130), .ZN(n10267) );
  AND2_X1 U11393 ( .A1(n12340), .A2(n12339), .ZN(n12348) );
  NAND2_X1 U11394 ( .A1(n12775), .A2(n10301), .ZN(n16512) );
  NOR2_X2 U11395 ( .A1(n20569), .A2(n20869), .ZN(n20622) );
  NAND2_X1 U11396 ( .A1(n21030), .A2(n20421), .ZN(n20671) );
  AND2_X1 U11397 ( .A1(n16733), .A2(n9821), .ZN(n14817) );
  NOR2_X1 U11398 ( .A1(n10099), .A2(n9935), .ZN(n10098) );
  NAND2_X1 U11399 ( .A1(n10326), .A2(n19174), .ZN(n11885) );
  INV_X1 U11400 ( .A(n20422), .ZN(n21030) );
  OR2_X1 U11401 ( .A1(n15216), .A2(n15215), .ZN(n15870) );
  NOR2_X1 U11402 ( .A1(n13464), .A2(n13463), .ZN(n13465) );
  NAND2_X2 U11403 ( .A1(n14012), .A2(n13951), .ZN(n20422) );
  NAND2_X1 U11404 ( .A1(n11126), .A2(n11125), .ZN(n11226) );
  NOR2_X1 U11405 ( .A1(n11153), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9935) );
  OR2_X1 U11406 ( .A1(n15729), .A2(n16040), .ZN(n15823) );
  NOR2_X1 U11407 ( .A1(n12215), .A2(n12214), .ZN(n12225) );
  AOI21_X1 U11408 ( .B1(n19339), .B2(n19948), .A(n10275), .ZN(n19322) );
  NAND2_X1 U11409 ( .A1(n12992), .A2(n12966), .ZN(n12979) );
  NAND2_X1 U11410 ( .A1(n10342), .A2(n10341), .ZN(n19092) );
  INV_X4 U11411 ( .A(n15664), .ZN(n15729) );
  AND2_X1 U11412 ( .A1(n11061), .A2(n11060), .ZN(n11214) );
  AND2_X1 U11413 ( .A1(n13946), .A2(n14574), .ZN(n13949) );
  CLKBUF_X1 U11414 ( .A(n15559), .Z(n15620) );
  AOI22_X1 U11415 ( .A1(n20862), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20599), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12179) );
  NAND2_X1 U11416 ( .A1(n10032), .A2(n10116), .ZN(n11061) );
  NAND2_X1 U11417 ( .A1(n9990), .A2(n11093), .ZN(n11104) );
  INV_X1 U11418 ( .A(n14594), .ZN(n14601) );
  NAND2_X1 U11419 ( .A1(n12947), .A2(n10378), .ZN(n16489) );
  NAND2_X1 U11420 ( .A1(n9984), .A2(n11879), .ZN(n11882) );
  AND2_X1 U11421 ( .A1(n11094), .A2(n11026), .ZN(n10348) );
  OAI22_X1 U11422 ( .A1(n16771), .A2(n20393), .B1(n20392), .B2(n20391), .ZN(
        n20906) );
  NAND2_X1 U11423 ( .A1(n10227), .A2(n11011), .ZN(n11094) );
  AND2_X1 U11424 ( .A1(n12882), .A2(n12885), .ZN(n20174) );
  NOR2_X2 U11425 ( .A1(n14506), .A2(n14505), .ZN(n14507) );
  NAND2_X1 U11426 ( .A1(n11083), .A2(n11082), .ZN(n13788) );
  NAND2_X1 U11427 ( .A1(n18735), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18731) );
  AND2_X1 U11428 ( .A1(n10002), .A2(n9782), .ZN(n11956) );
  AND2_X1 U11429 ( .A1(n16674), .A2(n16684), .ZN(n12174) );
  OR2_X1 U11430 ( .A1(n12915), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12885) );
  NAND2_X2 U11431 ( .A1(n17853), .A2(n9845), .ZN(n19202) );
  OAI21_X1 U11432 ( .B1(n16684), .B2(n13833), .A(n13639), .ZN(n13771) );
  INV_X2 U11433 ( .A(n18777), .ZN(n18784) );
  NAND2_X1 U11434 ( .A1(n14029), .A2(n10940), .ZN(n14337) );
  NAND2_X1 U11435 ( .A1(n10941), .A2(n10909), .ZN(n10995) );
  NAND2_X1 U11436 ( .A1(n12166), .A2(n12165), .ZN(n16684) );
  OAI221_X1 U11437 ( .B1(n13997), .B2(n13996), .C1(n13997), .C2(n17535), .A(
        n20087), .ZN(n18655) );
  NAND2_X1 U11438 ( .A1(n19346), .A2(n19253), .ZN(n19440) );
  OAI21_X1 U11439 ( .B1(n17458), .B2(n10004), .A(n10003), .ZN(n13815) );
  NOR2_X1 U11440 ( .A1(n15144), .A2(n20933), .ZN(n16678) );
  NOR2_X1 U11441 ( .A1(n10332), .A2(n10333), .ZN(n10330) );
  NOR2_X1 U11442 ( .A1(n13487), .A2(n14015), .ZN(n10415) );
  AND2_X1 U11443 ( .A1(n9971), .A2(n17462), .ZN(n9970) );
  NOR2_X1 U11444 ( .A1(n12851), .A2(n10370), .ZN(n12905) );
  AND2_X1 U11445 ( .A1(n10092), .A2(n11906), .ZN(n17565) );
  AND2_X1 U11446 ( .A1(n11069), .A2(n10165), .ZN(n10160) );
  INV_X1 U11447 ( .A(n12559), .ZN(n12552) );
  NAND2_X1 U11448 ( .A1(n10388), .A2(n10387), .ZN(n12160) );
  INV_X1 U11449 ( .A(n10891), .ZN(n10907) );
  AOI21_X1 U11450 ( .B1(n18132), .B2(n19036), .A(n19024), .ZN(n10201) );
  NAND2_X1 U11451 ( .A1(n11855), .A2(n11854), .ZN(n11858) );
  NOR2_X1 U11453 ( .A1(n17852), .A2(n11919), .ZN(n13927) );
  AND2_X1 U11454 ( .A1(n11903), .A2(n20089), .ZN(n9936) );
  OR2_X1 U11455 ( .A1(n10654), .A2(n19500), .ZN(n17852) );
  OAI211_X1 U11456 ( .C1(n12620), .C2(n12604), .A(n12622), .B(n12603), .ZN(
        n13746) );
  NAND2_X1 U11457 ( .A1(n11369), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11368) );
  CLKBUF_X1 U11458 ( .A(n12425), .Z(n9741) );
  AND2_X1 U11459 ( .A1(n10831), .A2(n14057), .ZN(n13013) );
  CLKBUF_X2 U11460 ( .A(n12625), .Z(n12794) );
  INV_X1 U11461 ( .A(n18798), .ZN(n19493) );
  INV_X2 U11462 ( .A(n13800), .ZN(n13040) );
  INV_X2 U11463 ( .A(n13119), .ZN(n13196) );
  OR2_X1 U11464 ( .A1(n11269), .A2(n15460), .ZN(n11274) );
  AND2_X1 U11466 ( .A1(n14057), .A2(n10868), .ZN(n10827) );
  OR2_X1 U11467 ( .A1(n12194), .A2(n12193), .ZN(n12635) );
  INV_X2 U11468 ( .A(n17803), .ZN(n17800) );
  NAND2_X1 U11469 ( .A1(n14287), .A2(n10883), .ZN(n14283) );
  NOR2_X2 U11470 ( .A1(n14287), .A2(n13032), .ZN(n13800) );
  CLKBUF_X2 U11471 ( .A(n10830), .Z(n10879) );
  CLKBUF_X1 U11472 ( .A(n12103), .Z(n14604) );
  NAND3_X1 U11473 ( .A1(n10461), .A2(n9778), .A3(n12239), .ZN(n13563) );
  OR2_X1 U11474 ( .A1(n10967), .A2(n10966), .ZN(n11150) );
  INV_X1 U11475 ( .A(n10777), .ZN(n13409) );
  OR2_X1 U11476 ( .A1(n12251), .A2(n12250), .ZN(n12611) );
  NAND4_X2 U11477 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n20089) );
  OR2_X2 U11478 ( .A1(n10859), .A2(n10858), .ZN(n14045) );
  NAND4_X1 U11479 ( .A1(n10760), .A2(n10759), .A3(n10758), .A4(n10757), .ZN(
        n10777) );
  NAND2_X1 U11480 ( .A1(n11999), .A2(n11998), .ZN(n12080) );
  NAND2_X1 U11481 ( .A1(n12050), .A2(n12049), .ZN(n12090) );
  NAND2_X1 U11482 ( .A1(n10478), .A2(n10477), .ZN(n10861) );
  NAND4_X1 U11483 ( .A1(n10817), .A2(n10476), .A3(n10816), .A4(n10815), .ZN(
        n10830) );
  INV_X2 U11484 ( .A(U214), .ZN(n17798) );
  AND4_X1 U11485 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n10758) );
  AND4_X1 U11486 ( .A1(n10756), .A2(n10755), .A3(n10754), .A4(n10753), .ZN(
        n10757) );
  AND4_X1 U11487 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10478) );
  AND4_X1 U11488 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n10731) );
  AND4_X1 U11489 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11753) );
  AND2_X1 U11490 ( .A1(n12000), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12005) );
  INV_X1 U11491 ( .A(n18498), .ZN(n9745) );
  AND2_X1 U11492 ( .A1(n11217), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11227) );
  INV_X1 U11493 ( .A(n18498), .ZN(n9744) );
  AND4_X1 U11494 ( .A1(n10812), .A2(n10811), .A3(n10810), .A4(n10809), .ZN(
        n10817) );
  AND3_X1 U11495 ( .A1(n12007), .A2(n12006), .A3(n11984), .ZN(n12011) );
  BUF_X2 U11496 ( .A(n10973), .Z(n11699) );
  NOR2_X2 U11497 ( .A1(n17446), .A2(n19134), .ZN(n18058) );
  INV_X2 U11498 ( .A(n18189), .ZN(n13366) );
  BUF_X2 U11499 ( .A(n10968), .Z(n11533) );
  BUF_X2 U11500 ( .A(n12180), .Z(n14952) );
  INV_X2 U11501 ( .A(n21085), .ZN(n20999) );
  INV_X2 U11502 ( .A(n17841), .ZN(n17843) );
  NAND2_X1 U11503 ( .A1(n15011), .A2(n10701), .ZN(n10834) );
  AND2_X1 U11504 ( .A1(n10694), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10425) );
  AND2_X1 U11505 ( .A1(n11909), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10522) );
  NOR2_X1 U11506 ( .A1(n21563), .A2(n18951), .ZN(n18936) );
  AND2_X1 U11507 ( .A1(n19926), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13935) );
  AND2_X2 U11508 ( .A1(n14784), .A2(n12188), .ZN(n12234) );
  AND2_X2 U11509 ( .A1(n14784), .A2(n12187), .ZN(n12233) );
  AND2_X1 U11510 ( .A1(n9942), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10521) );
  NOR2_X1 U11511 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10696) );
  AND2_X1 U11512 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14997) );
  AND2_X2 U11513 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16091) );
  AND2_X1 U11514 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10701) );
  NOR2_X2 U11515 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14114) );
  AND2_X1 U11516 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14667) );
  INV_X2 U11517 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11909) );
  NOR2_X2 U11518 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10524) );
  INV_X1 U11519 ( .A(n17459), .ZN(n9730) );
  INV_X1 U11520 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19110) );
  NOR3_X1 U11521 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18194) );
  NAND2_X1 U11522 ( .A1(n17575), .A2(n17483), .ZN(n17425) );
  OR2_X2 U11523 ( .A1(n12447), .A2(n9736), .ZN(n12066) );
  NOR2_X1 U11524 ( .A1(n19173), .A2(n9983), .ZN(n9731) );
  AND2_X1 U11525 ( .A1(n10464), .A2(n9732), .ZN(n9733) );
  INV_X1 U11526 ( .A(n19063), .ZN(n9732) );
  AND2_X1 U11527 ( .A1(n19061), .A2(n9732), .ZN(n10487) );
  INV_X1 U11528 ( .A(n13528), .ZN(n9734) );
  CLKBUF_X1 U11529 ( .A(n12109), .Z(n13634) );
  OR2_X1 U11530 ( .A1(n21077), .A2(n12605), .ZN(n9735) );
  NOR2_X4 U11531 ( .A1(n14630), .A2(n13318), .ZN(n16744) );
  NOR2_X2 U11532 ( .A1(n11484), .A2(n15743), .ZN(n11485) );
  NOR2_X2 U11533 ( .A1(n11274), .A2(n15849), .ZN(n11293) );
  NAND2_X2 U11534 ( .A1(n15722), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11169) );
  OAI21_X4 U11535 ( .B1(n17653), .B2(n9998), .A(n9995), .ZN(n15765) );
  OR2_X1 U11536 ( .A1(n12125), .A2(n14609), .ZN(n9736) );
  INV_X1 U11537 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9737) );
  NOR2_X2 U11538 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18049), .ZN(n18031) );
  NOR2_X2 U11539 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18148), .ZN(n18133) );
  OAI22_X1 U11540 ( .A1(n17105), .A2(n17104), .B1(n20261), .B2(n20363), .ZN(
        n9738) );
  OAI22_X1 U11541 ( .A1(n17105), .A2(n17104), .B1(n20261), .B2(n20363), .ZN(
        n17366) );
  AND2_X2 U11542 ( .A1(n12455), .A2(n14248), .ZN(n9749) );
  AND3_X1 U11543 ( .A1(n12131), .A2(n12130), .A3(n12129), .ZN(n9739) );
  CLKBUF_X1 U11544 ( .A(n12562), .Z(n9740) );
  XNOR2_X1 U11545 ( .A(n13201), .B(n13200), .ZN(n15497) );
  NOR2_X2 U11546 ( .A1(n15336), .A2(n10276), .ZN(n10279) );
  OR2_X2 U11547 ( .A1(n15266), .A2(n10260), .ZN(n9773) );
  NOR2_X2 U11548 ( .A1(n15350), .A2(n15352), .ZN(n15335) );
  AND2_X2 U11549 ( .A1(n12605), .A2(n20821), .ZN(n12632) );
  AND2_X2 U11550 ( .A1(n11896), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10177) );
  AND2_X1 U11551 ( .A1(n13767), .A2(n16684), .ZN(n12175) );
  XNOR2_X1 U11552 ( .A(n12159), .B(n12160), .ZN(n12167) );
  AOI21_X1 U11553 ( .B1(n12156), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12157), .ZN(n12482) );
  NAND2_X1 U11554 ( .A1(n17175), .A2(n13253), .ZN(n9742) );
  INV_X1 U11555 ( .A(n21077), .ZN(n12419) );
  INV_X1 U11556 ( .A(n12605), .ZN(n12125) );
  AND2_X1 U11557 ( .A1(n9886), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13490) );
  AND2_X1 U11558 ( .A1(n13252), .A2(n9860), .ZN(n13344) );
  NAND2_X1 U11559 ( .A1(n9900), .A2(n13301), .ZN(n17026) );
  INV_X1 U11560 ( .A(n11733), .ZN(n9743) );
  NAND2_X1 U11561 ( .A1(n13935), .A2(n14114), .ZN(n11733) );
  AND2_X1 U11562 ( .A1(n12186), .A2(n14209), .ZN(n9746) );
  AND3_X4 U11563 ( .A1(n10290), .A2(n10289), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12180) );
  AND2_X4 U11564 ( .A1(n12187), .A2(n14209), .ZN(n12043) );
  NOR2_X2 U11565 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17903), .ZN(n17902) );
  INV_X1 U11566 ( .A(n17056), .ZN(n9900) );
  NAND2_X1 U11567 ( .A1(n17057), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17056) );
  AND3_X4 U11568 ( .A1(n10289), .A2(n11974), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12001) );
  NOR2_X2 U11569 ( .A1(n10482), .A2(n10202), .ZN(n11964) );
  INV_X2 U11570 ( .A(n12161), .ZN(n9877) );
  OAI21_X1 U11571 ( .B1(n13379), .B2(n17136), .A(n13187), .ZN(n10107) );
  XNOR2_X1 U11572 ( .A(n10108), .B(n9783), .ZN(n13379) );
  NAND2_X1 U11573 ( .A1(n16929), .A2(n12954), .ZN(n16923) );
  NOR2_X2 U11574 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18022), .ZN(n18014) );
  NOR2_X2 U11575 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17897), .ZN(n17881) );
  AND2_X2 U11576 ( .A1(n10507), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10490) );
  INV_X1 U11577 ( .A(n10512), .ZN(n18178) );
  INV_X1 U11578 ( .A(n11095), .ZN(n10116) );
  MUX2_X1 U11579 ( .A(n12635), .B(n12408), .S(n12388), .Z(n12811) );
  OR2_X1 U11580 ( .A1(n12263), .A2(n12262), .ZN(n12443) );
  INV_X1 U11581 ( .A(n14503), .ZN(n12763) );
  INV_X1 U11582 ( .A(n13297), .ZN(n12775) );
  AND4_X1 U11583 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12369) );
  AND4_X1 U11584 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12368) );
  NOR2_X1 U11585 ( .A1(n10654), .A2(n11904), .ZN(n11906) );
  OR2_X1 U11586 ( .A1(n17628), .A2(n14687), .ZN(n15476) );
  NAND3_X1 U11587 ( .A1(n10018), .A2(n10017), .A3(n11052), .ZN(n11181) );
  AND2_X1 U11588 ( .A1(n10994), .A2(n10955), .ZN(n10017) );
  AND2_X1 U11589 ( .A1(n13175), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10368) );
  AND2_X1 U11590 ( .A1(n9965), .A2(n20929), .ZN(n9964) );
  NAND2_X1 U11591 ( .A1(n14287), .A2(n10884), .ZN(n10885) );
  NOR2_X1 U11592 ( .A1(n10232), .A2(n11125), .ZN(n10231) );
  AND2_X1 U11593 ( .A1(n10348), .A2(n11054), .ZN(n10032) );
  AND2_X1 U11594 ( .A1(n10897), .A2(n10896), .ZN(n13137) );
  AND2_X1 U11595 ( .A1(n11595), .A2(n15264), .ZN(n11596) );
  NOR2_X1 U11596 ( .A1(n10117), .A2(n14329), .ZN(n15387) );
  NOR2_X1 U11597 ( .A1(n9848), .A2(n15538), .ZN(n10121) );
  OR2_X1 U11598 ( .A1(n14057), .A2(n14687), .ZN(n11711) );
  NAND2_X1 U11599 ( .A1(n15782), .A2(n15768), .ZN(n10096) );
  AND2_X1 U11600 ( .A1(n10879), .A2(n14057), .ZN(n13417) );
  NAND3_X1 U11601 ( .A1(n14337), .A2(n21654), .A3(n10941), .ZN(n10018) );
  NOR2_X1 U11602 ( .A1(n12849), .A2(n12848), .ZN(n12854) );
  NAND2_X1 U11603 ( .A1(n12123), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U11604 ( .A1(n12813), .A2(n12812), .ZN(n12815) );
  NAND2_X1 U11605 ( .A1(n12388), .A2(n12441), .ZN(n12442) );
  NOR2_X1 U11606 ( .A1(n9794), .A2(n10391), .ZN(n10068) );
  INV_X1 U11607 ( .A(n14011), .ZN(n10391) );
  NOR2_X1 U11608 ( .A1(n16691), .A2(n10384), .ZN(n10383) );
  INV_X1 U11609 ( .A(n16697), .ZN(n10384) );
  NAND2_X1 U11610 ( .A1(n16733), .A2(n9824), .ZN(n10395) );
  AND2_X1 U11611 ( .A1(n21078), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13770) );
  INV_X1 U11612 ( .A(n13296), .ZN(n12774) );
  AND2_X1 U11613 ( .A1(n14751), .A2(n16750), .ZN(n10399) );
  NAND3_X1 U11614 ( .A1(n9897), .A2(n10079), .A3(n17362), .ZN(n10001) );
  NOR2_X1 U11615 ( .A1(n10021), .A2(n10024), .ZN(n10320) );
  AND2_X1 U11616 ( .A1(n12179), .A2(n12173), .ZN(n10319) );
  NAND2_X1 U11617 ( .A1(n12160), .A2(n12159), .ZN(n9893) );
  AND2_X1 U11618 ( .A1(n16743), .A2(n10419), .ZN(n10418) );
  INV_X1 U11619 ( .A(n13294), .ZN(n10419) );
  NAND2_X1 U11620 ( .A1(n9988), .A2(n10030), .ZN(n9987) );
  AND2_X1 U11621 ( .A1(n10029), .A2(n10078), .ZN(n9988) );
  INV_X1 U11622 ( .A(n14714), .ZN(n10300) );
  INV_X1 U11623 ( .A(n14278), .ZN(n12764) );
  NAND3_X1 U11624 ( .A1(n10071), .A2(n10031), .A3(n9717), .ZN(n10030) );
  AND2_X1 U11625 ( .A1(n10070), .A2(n10362), .ZN(n10031) );
  INV_X1 U11626 ( .A(n9914), .ZN(n10362) );
  NAND2_X1 U11627 ( .A1(n10294), .A2(n13859), .ZN(n10293) );
  INV_X1 U11628 ( .A(n10295), .ZN(n10294) );
  NAND2_X1 U11629 ( .A1(n12645), .A2(n12644), .ZN(n14561) );
  INV_X1 U11630 ( .A(n14569), .ZN(n12644) );
  INV_X1 U11631 ( .A(n14565), .ZN(n12645) );
  NAND2_X1 U11632 ( .A1(n9985), .A2(n16631), .ZN(n9886) );
  NOR2_X1 U11633 ( .A1(n12463), .A2(n13178), .ZN(n12465) );
  AND3_X1 U11634 ( .A1(n12639), .A2(n12638), .A3(n12637), .ZN(n14566) );
  AND2_X2 U11635 ( .A1(n12083), .A2(n12081), .ZN(n12576) );
  NAND2_X1 U11636 ( .A1(n13834), .A2(n13766), .ZN(n13836) );
  NOR2_X1 U11637 ( .A1(n14897), .A2(n13944), .ZN(n13945) );
  INV_X1 U11638 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13944) );
  NOR2_X1 U11639 ( .A1(n21494), .A2(n21692), .ZN(n20863) );
  AOI21_X1 U11640 ( .B1(n10673), .B2(n10672), .A(n10671), .ZN(n11917) );
  AND2_X1 U11641 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19943), .ZN(
        n10671) );
  OR2_X1 U11642 ( .A1(n11916), .A2(n10668), .ZN(n11924) );
  AND2_X1 U11643 ( .A1(n10521), .A2(n13935), .ZN(n18230) );
  NAND2_X1 U11644 ( .A1(n18697), .A2(n10639), .ZN(n11903) );
  NOR2_X1 U11645 ( .A1(n13927), .A2(n18856), .ZN(n11902) );
  NAND2_X1 U11646 ( .A1(n10521), .A2(n14667), .ZN(n10611) );
  AND4_X1 U11647 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10729) );
  AND4_X1 U11648 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10730) );
  OR2_X1 U11649 ( .A1(n17628), .A2(n21335), .ZN(n15201) );
  OR2_X1 U11650 ( .A1(n15216), .A2(n13119), .ZN(n13197) );
  OR2_X1 U11651 ( .A1(n13168), .A2(n13203), .ZN(n10215) );
  NAND2_X1 U11652 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15687), .ZN(
        n9991) );
  OAI22_X1 U11653 ( .A1(n15758), .A2(n9856), .B1(n15840), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9937) );
  OR2_X1 U11654 ( .A1(n13023), .A2(n13022), .ZN(n13024) );
  NAND2_X1 U11655 ( .A1(n10217), .A2(n10216), .ZN(n13023) );
  INV_X1 U11656 ( .A(n10992), .ZN(n10019) );
  NAND2_X1 U11657 ( .A1(n10230), .A2(n10229), .ZN(n10228) );
  INV_X1 U11658 ( .A(n10996), .ZN(n10229) );
  INV_X1 U11659 ( .A(n10995), .ZN(n10230) );
  CLKBUF_X1 U11660 ( .A(n14028), .Z(n15024) );
  OAI21_X1 U11661 ( .B1(n16486), .B2(n10238), .A(n16909), .ZN(n16474) );
  INV_X1 U11662 ( .A(n12812), .ZN(n12985) );
  AND2_X1 U11663 ( .A1(n10381), .A2(n14940), .ZN(n10054) );
  NAND2_X1 U11664 ( .A1(n13347), .A2(n13346), .ZN(n14964) );
  NAND2_X1 U11665 ( .A1(n10183), .A2(n10186), .ZN(n13354) );
  AOI21_X1 U11666 ( .B1(n10188), .B2(n10189), .A(n10187), .ZN(n10186) );
  INV_X1 U11667 ( .A(n13185), .ZN(n10187) );
  NOR2_X1 U11668 ( .A1(n17194), .A2(n17181), .ZN(n10133) );
  INV_X1 U11669 ( .A(n13252), .ZN(n9904) );
  INV_X1 U11670 ( .A(n16512), .ZN(n12782) );
  AND2_X1 U11671 ( .A1(n9771), .A2(n12594), .ZN(n10132) );
  NAND2_X1 U11672 ( .A1(n12416), .A2(n12415), .ZN(n14314) );
  NAND2_X1 U11673 ( .A1(n9888), .A2(n21057), .ZN(n12415) );
  XNOR2_X1 U11674 ( .A(n13771), .B(n13829), .ZN(n13772) );
  NAND2_X1 U11675 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20475) );
  NAND2_X1 U11676 ( .A1(n20422), .A2(n20368), .ZN(n20569) );
  NAND2_X1 U11677 ( .A1(n10136), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n10135) );
  INV_X1 U11678 ( .A(n10137), .ZN(n10136) );
  AND4_X1 U11679 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10638) );
  AND4_X1 U11680 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10635) );
  AND4_X1 U11681 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10637) );
  AOI211_X1 U11682 ( .C1(n19949), .C2(n19303), .A(n19256), .B(n19300), .ZN(
        n19271) );
  NAND2_X1 U11683 ( .A1(n10219), .A2(n10052), .ZN(n15196) );
  NOR2_X1 U11684 ( .A1(n13408), .A2(n21089), .ZN(n10052) );
  NAND2_X1 U11685 ( .A1(n17620), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21089) );
  NAND2_X1 U11686 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  AOI21_X1 U11687 ( .B1(n15229), .B2(P1_REIP_REG_29__SCAN_IN), .A(n15220), 
        .ZN(n10048) );
  NAND2_X1 U11688 ( .A1(n15221), .A2(n21176), .ZN(n10049) );
  AOI21_X1 U11689 ( .B1(n13207), .B2(n13206), .A(n10211), .ZN(n13208) );
  OR2_X1 U11690 ( .A1(n13205), .A2(n13466), .ZN(n10211) );
  NAND2_X1 U11691 ( .A1(n16448), .A2(n13179), .ZN(n9908) );
  INV_X1 U11692 ( .A(n13361), .ZN(n9909) );
  CLKBUF_X1 U11693 ( .A(n12161), .Z(n12166) );
  INV_X1 U11694 ( .A(n16976), .ZN(n16963) );
  INV_X1 U11695 ( .A(n14717), .ZN(n10150) );
  INV_X1 U11696 ( .A(n20355), .ZN(n17372) );
  NAND2_X1 U11697 ( .A1(n20709), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n9879) );
  INV_X1 U11698 ( .A(n11058), .ZN(n11026) );
  AND2_X1 U11699 ( .A1(n10795), .A2(n10794), .ZN(n10797) );
  OR2_X1 U11700 ( .A1(n10954), .A2(n10953), .ZN(n11084) );
  OR2_X1 U11701 ( .A1(n14051), .A2(n21654), .ZN(n10991) );
  NAND2_X1 U11702 ( .A1(n13134), .A2(n14090), .ZN(n10867) );
  CLKBUF_X1 U11703 ( .A(n10910), .Z(n10911) );
  AOI21_X1 U11704 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n17600), .A(
        n10797), .ZN(n10800) );
  INV_X1 U11705 ( .A(n13004), .ZN(n10801) );
  AND2_X1 U11706 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12055) );
  INV_X1 U11707 ( .A(n14642), .ZN(n10067) );
  OAI21_X1 U11708 ( .B1(n9915), .B2(n13275), .A(n13277), .ZN(n9914) );
  AND2_X1 U11709 ( .A1(n9838), .A2(n10318), .ZN(n10316) );
  AOI22_X1 U11710 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11996) );
  AOI21_X1 U11711 ( .B1(n10660), .B2(n19926), .A(n10662), .ZN(n10673) );
  INV_X1 U11712 ( .A(n13822), .ZN(n10332) );
  INV_X1 U11713 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10626) );
  AND2_X1 U11714 ( .A1(n11901), .A2(n11900), .ZN(n11921) );
  AND2_X1 U11715 ( .A1(n11594), .A2(n15275), .ZN(n15264) );
  AND2_X1 U11716 ( .A1(n15334), .A2(n10127), .ZN(n10126) );
  AND2_X1 U11717 ( .A1(n14514), .A2(n10466), .ZN(n10443) );
  INV_X1 U11718 ( .A(n11061), .ZN(n11042) );
  AND2_X1 U11719 ( .A1(n11044), .A2(n11383), .ZN(n10129) );
  NAND2_X1 U11720 ( .A1(n10263), .A2(n15241), .ZN(n10262) );
  INV_X1 U11721 ( .A(n15267), .ZN(n10263) );
  NAND2_X1 U11722 ( .A1(n15695), .A2(n15674), .ZN(n10033) );
  AND2_X1 U11723 ( .A1(n10349), .A2(n11160), .ZN(n10167) );
  NAND2_X1 U11724 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  INV_X1 U11725 ( .A(n15409), .ZN(n10269) );
  INV_X1 U11726 ( .A(n10271), .ZN(n10270) );
  OR2_X1 U11727 ( .A1(n15729), .A2(n16069), .ZN(n15766) );
  NAND2_X1 U11728 ( .A1(n11143), .A2(n11142), .ZN(n11144) );
  AND2_X1 U11729 ( .A1(n10280), .A2(n13052), .ZN(n10281) );
  INV_X1 U11730 ( .A(n14334), .ZN(n10280) );
  INV_X1 U11731 ( .A(n13047), .ZN(n13127) );
  NAND2_X1 U11732 ( .A1(n13852), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9990) );
  AND4_X1 U11733 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n10760) );
  AND4_X1 U11734 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n10759) );
  OR2_X1 U11735 ( .A1(n10979), .A2(n10978), .ZN(n11085) );
  NAND2_X1 U11736 ( .A1(n10163), .A2(n10907), .ZN(n10162) );
  NOR2_X1 U11737 ( .A1(n10907), .A2(n10889), .ZN(n10164) );
  NAND2_X1 U11738 ( .A1(n15197), .A2(n10899), .ZN(n10101) );
  OR2_X1 U11739 ( .A1(n11010), .A2(n11009), .ZN(n11045) );
  AND2_X1 U11740 ( .A1(n10042), .A2(n14697), .ZN(n11132) );
  INV_X1 U11741 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15029) );
  OAI21_X1 U11742 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n10913), .ZN(n16164) );
  INV_X1 U11743 ( .A(n11054), .ZN(n15022) );
  NAND2_X1 U11744 ( .A1(n12394), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12412) );
  NAND2_X1 U11745 ( .A1(n16502), .A2(n15144), .ZN(n10237) );
  NOR2_X1 U11746 ( .A1(n12878), .A2(n12874), .ZN(n10377) );
  NAND2_X1 U11747 ( .A1(n10374), .A2(n10375), .ZN(n10373) );
  INV_X1 U11748 ( .A(n12852), .ZN(n10374) );
  OR2_X1 U11749 ( .A1(n12851), .A2(n10373), .ZN(n12892) );
  AND2_X1 U11750 ( .A1(n13257), .A2(n16463), .ZN(n10424) );
  NOR2_X1 U11751 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14784) );
  CLKBUF_X1 U11752 ( .A(n14783), .Z(n14948) );
  NOR2_X1 U11753 ( .A1(n10308), .A2(n10307), .ZN(n10306) );
  INV_X1 U11754 ( .A(n13265), .ZN(n10307) );
  NAND2_X1 U11755 ( .A1(n9820), .A2(n16719), .ZN(n10393) );
  NAND2_X1 U11756 ( .A1(n10309), .A2(n16483), .ZN(n10308) );
  INV_X1 U11757 ( .A(n16497), .ZN(n10309) );
  INV_X1 U11758 ( .A(n10394), .ZN(n10061) );
  NOR2_X1 U11759 ( .A1(n10393), .A2(n14874), .ZN(n10063) );
  NAND2_X1 U11760 ( .A1(n10395), .A2(n9820), .ZN(n10394) );
  NOR2_X1 U11761 ( .A1(n10246), .A2(n15175), .ZN(n10244) );
  INV_X1 U11762 ( .A(n10247), .ZN(n10245) );
  NOR2_X1 U11763 ( .A1(n15121), .A2(n20187), .ZN(n15123) );
  NOR2_X1 U11764 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  INV_X1 U11765 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U11766 ( .A1(n14409), .A2(n14415), .ZN(n10421) );
  NAND2_X1 U11767 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10252) );
  AND2_X1 U11768 ( .A1(n10424), .A2(n16449), .ZN(n10423) );
  NAND2_X1 U11769 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  INV_X1 U11770 ( .A(n13282), .ZN(n10358) );
  NAND2_X1 U11771 ( .A1(n9779), .A2(n10360), .ZN(n10359) );
  NAND2_X1 U11772 ( .A1(n12764), .A2(n9829), .ZN(n13332) );
  OAI21_X1 U11773 ( .B1(n9915), .B2(n9913), .A(n9912), .ZN(n10029) );
  NAND2_X1 U11774 ( .A1(n13274), .A2(n16984), .ZN(n9913) );
  NAND2_X1 U11775 ( .A1(n9914), .A2(n16984), .ZN(n9912) );
  NAND2_X1 U11776 ( .A1(n10313), .A2(n14002), .ZN(n10312) );
  INV_X1 U11777 ( .A(n10314), .ZN(n10313) );
  OR2_X1 U11778 ( .A1(n20217), .A2(n12994), .ZN(n12933) );
  INV_X1 U11779 ( .A(n13757), .ZN(n12666) );
  NOR2_X1 U11780 ( .A1(n17122), .A2(n17732), .ZN(n10411) );
  INV_X1 U11781 ( .A(n16641), .ZN(n10408) );
  NOR2_X1 U11782 ( .A1(n9874), .A2(n12089), .ZN(n9873) );
  INV_X1 U11783 ( .A(n12138), .ZN(n10388) );
  NAND2_X1 U11784 ( .A1(n12562), .A2(n9832), .ZN(n10387) );
  NOR2_X1 U11785 ( .A1(n12605), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12612) );
  AND2_X1 U11786 ( .A1(n12631), .A2(n12640), .ZN(n10292) );
  CLKBUF_X1 U11787 ( .A(n12186), .Z(n14242) );
  AND2_X2 U11788 ( .A1(n9901), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14241) );
  INV_X1 U11789 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13837) );
  NAND2_X1 U11790 ( .A1(n13839), .A2(n13838), .ZN(n13947) );
  INV_X1 U11791 ( .A(n12213), .ZN(n12298) );
  AND4_X1 U11792 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12566), .ZN(
        n14225) );
  NAND2_X1 U11793 ( .A1(n12123), .A2(n13769), .ZN(n12096) );
  AND2_X1 U11794 ( .A1(n18659), .A2(n11922), .ZN(n10648) );
  INV_X1 U11795 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11796 ( .A1(n10524), .A2(n14114), .ZN(n10540) );
  NAND2_X1 U11797 ( .A1(n10205), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10204) );
  INV_X1 U11798 ( .A(n10206), .ZN(n10205) );
  NOR2_X1 U11799 ( .A1(n19113), .A2(n10181), .ZN(n10179) );
  NAND2_X1 U11800 ( .A1(n19176), .A2(n9754), .ZN(n10182) );
  NAND2_X1 U11801 ( .A1(n19188), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9984) );
  OAI21_X1 U11802 ( .B1(n13885), .B2(n9973), .A(n9970), .ZN(n11864) );
  AND2_X1 U11803 ( .A1(n13227), .A2(n11922), .ZN(n13222) );
  INV_X1 U11804 ( .A(n19950), .ZN(n13994) );
  INV_X1 U11805 ( .A(n10436), .ZN(n10435) );
  NAND2_X1 U11806 ( .A1(n10438), .A2(n10437), .ZN(n10436) );
  INV_X1 U11807 ( .A(n10439), .ZN(n10437) );
  INV_X1 U11808 ( .A(n13407), .ZN(n10433) );
  AND2_X1 U11809 ( .A1(n15422), .A2(n15405), .ZN(n15406) );
  AND3_X1 U11810 ( .A1(n11273), .A2(n11272), .A3(n11271), .ZN(n15538) );
  NAND2_X1 U11811 ( .A1(n11184), .A2(n11183), .ZN(n13794) );
  INV_X1 U11812 ( .A(n15675), .ZN(n9941) );
  NAND2_X1 U11813 ( .A1(n9994), .A2(n9993), .ZN(n15650) );
  NAND2_X1 U11814 ( .A1(n10034), .A2(n9759), .ZN(n9994) );
  NAND2_X1 U11815 ( .A1(n10033), .A2(n10035), .ZN(n15675) );
  NAND2_X1 U11816 ( .A1(n15313), .A2(n10277), .ZN(n10276) );
  NOR2_X1 U11817 ( .A1(n15310), .A2(n15325), .ZN(n10277) );
  NAND2_X1 U11818 ( .A1(n9996), .A2(n9792), .ZN(n9938) );
  AOI22_X1 U11819 ( .A1(n17653), .A2(n9999), .B1(n9998), .B2(n9997), .ZN(n9996) );
  NAND2_X1 U11820 ( .A1(n15664), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15801) );
  XNOR2_X1 U11821 ( .A(n11144), .B(n17690), .ZN(n17652) );
  NAND2_X1 U11822 ( .A1(n17653), .A2(n17652), .ZN(n17651) );
  AND2_X1 U11823 ( .A1(n11068), .A2(n11067), .ZN(n11108) );
  OAI21_X1 U11824 ( .B1(n17660), .B2(n17658), .A(n17695), .ZN(n11112) );
  NAND2_X1 U11825 ( .A1(n10018), .A2(n10955), .ZN(n11179) );
  AND2_X1 U11826 ( .A1(n11181), .A2(n11052), .ZN(n11053) );
  OR2_X1 U11827 ( .A1(n15024), .A2(n14070), .ZN(n16159) );
  INV_X1 U11828 ( .A(n14075), .ZN(n14541) );
  NOR2_X1 U11829 ( .A1(n14443), .A2(n14687), .ZN(n16203) );
  AND2_X1 U11830 ( .A1(n15024), .A2(n16291), .ZN(n15053) );
  INV_X1 U11831 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17600) );
  NAND2_X1 U11832 ( .A1(n21654), .A2(n14032), .ZN(n16202) );
  NOR2_X1 U11833 ( .A1(n11176), .A2(n15022), .ZN(n21280) );
  INV_X1 U11834 ( .A(n13523), .ZN(n14260) );
  NAND2_X1 U11835 ( .A1(n12413), .A2(n12412), .ZN(n12449) );
  OR2_X1 U11836 ( .A1(n12411), .A2(n21553), .ZN(n12413) );
  INV_X1 U11837 ( .A(n9956), .ZN(n12445) );
  OAI21_X1 U11838 ( .B1(n16433), .B2(n10238), .A(n16434), .ZN(n16435) );
  NAND2_X1 U11839 ( .A1(n12910), .A2(n9790), .ZN(n12888) );
  INV_X1 U11840 ( .A(n12889), .ZN(n12862) );
  NAND2_X1 U11841 ( .A1(n12823), .A2(n9916), .ZN(n12849) );
  NOR2_X1 U11842 ( .A1(n9917), .A2(n9918), .ZN(n9916) );
  AND2_X1 U11843 ( .A1(n14876), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14572) );
  NAND3_X1 U11844 ( .A1(n14901), .A2(n14905), .A3(n9827), .ZN(n10381) );
  OR2_X1 U11845 ( .A1(n14900), .A2(n14899), .ZN(n14901) );
  INV_X1 U11846 ( .A(n10395), .ZN(n14818) );
  AND2_X1 U11847 ( .A1(n10399), .A2(n10398), .ZN(n10397) );
  INV_X1 U11848 ( .A(n16740), .ZN(n10398) );
  NAND2_X1 U11849 ( .A1(n14314), .A2(n21078), .ZN(n14219) );
  AND2_X1 U11850 ( .A1(n15133), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15135) );
  NAND2_X1 U11851 ( .A1(n9987), .A2(n13278), .ZN(n14712) );
  NOR2_X1 U11852 ( .A1(n14014), .A2(n10414), .ZN(n14129) );
  INV_X1 U11853 ( .A(n10415), .ZN(n10414) );
  AND2_X1 U11854 ( .A1(n10318), .A2(n12264), .ZN(n10175) );
  AND2_X1 U11855 ( .A1(n9896), .A2(n12286), .ZN(n17131) );
  AND2_X1 U11856 ( .A1(n13353), .A2(n13356), .ZN(n10012) );
  NOR2_X1 U11857 ( .A1(n16454), .A2(n12994), .ZN(n16874) );
  OAI21_X1 U11858 ( .B1(n16872), .B2(n16873), .A(n16905), .ZN(n9945) );
  NOR2_X1 U11859 ( .A1(n16885), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9946) );
  AND2_X1 U11860 ( .A1(n17212), .A2(n12594), .ZN(n12585) );
  AND2_X1 U11861 ( .A1(n13454), .A2(n12380), .ZN(n13451) );
  AND2_X1 U11862 ( .A1(n10418), .A2(n10417), .ZN(n10416) );
  INV_X1 U11863 ( .A(n13448), .ZN(n10417) );
  AND2_X1 U11864 ( .A1(n9826), .A2(n16529), .ZN(n10301) );
  OR2_X1 U11865 ( .A1(n10460), .A2(n10011), .ZN(n10010) );
  INV_X1 U11866 ( .A(n10357), .ZN(n10351) );
  NAND2_X1 U11867 ( .A1(n9987), .A2(n9986), .ZN(n10354) );
  AND2_X1 U11868 ( .A1(n9810), .A2(n13278), .ZN(n9986) );
  NAND2_X1 U11869 ( .A1(n10354), .A2(n10352), .ZN(n13443) );
  NOR2_X1 U11870 ( .A1(n10357), .A2(n10353), .ZN(n10352) );
  INV_X1 U11871 ( .A(n13284), .ZN(n10353) );
  NAND2_X1 U11872 ( .A1(n10360), .A2(n13328), .ZN(n10355) );
  INV_X1 U11873 ( .A(n14712), .ZN(n10037) );
  AND2_X1 U11874 ( .A1(n10361), .A2(n13328), .ZN(n10356) );
  CLKBUF_X1 U11875 ( .A(n13332), .Z(n16841) );
  NAND2_X1 U11876 ( .A1(n12721), .A2(n9846), .ZN(n10314) );
  AOI21_X1 U11877 ( .B1(n13275), .B2(n17006), .A(n10367), .ZN(n10366) );
  INV_X1 U11878 ( .A(n17008), .ZN(n10367) );
  NAND2_X1 U11879 ( .A1(n17005), .A2(n13275), .ZN(n10365) );
  CLKBUF_X1 U11880 ( .A(n13857), .Z(n13858) );
  OR3_X1 U11881 ( .A1(n12376), .A2(n12994), .A3(n17341), .ZN(n12377) );
  NAND2_X1 U11882 ( .A1(n17113), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U11883 ( .A(n10412), .ZN(n10409) );
  NAND2_X1 U11884 ( .A1(n13637), .A2(n20821), .ZN(n13941) );
  OR2_X1 U11885 ( .A1(n13771), .A2(n13830), .ZN(n13831) );
  OR2_X1 U11886 ( .A1(n14013), .A2(n13945), .ZN(n13946) );
  INV_X1 U11887 ( .A(n12289), .ZN(n20374) );
  AND2_X1 U11889 ( .A1(n21028), .A2(n20818), .ZN(n20706) );
  AND3_X1 U11890 ( .A1(n21028), .A2(n13940), .A3(n20871), .ZN(n14600) );
  NAND2_X1 U11891 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21050), .ZN(
        n20672) );
  NAND2_X1 U11892 ( .A1(n14390), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20820) );
  NAND2_X1 U11893 ( .A1(n14395), .A2(n14394), .ZN(n20874) );
  NAND2_X1 U11894 ( .A1(n14393), .A2(n21072), .ZN(n14394) );
  NAND2_X1 U11895 ( .A1(n17418), .A2(n21075), .ZN(n14395) );
  INV_X1 U11896 ( .A(n20874), .ZN(n20823) );
  NAND2_X1 U11897 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17409), .ZN(n14316) );
  NOR2_X1 U11898 ( .A1(n17565), .A2(n10655), .ZN(n19952) );
  NOR2_X1 U11899 ( .A1(n18010), .A2(n18178), .ZN(n18004) );
  NAND2_X1 U11900 ( .A1(n10512), .A2(n10210), .ZN(n10209) );
  NAND2_X1 U11901 ( .A1(n10492), .A2(n18221), .ZN(n10210) );
  NAND2_X1 U11902 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10532) );
  NOR2_X1 U11903 ( .A1(n19496), .A2(n19493), .ZN(n17536) );
  OR2_X1 U11904 ( .A1(n17565), .A2(n10091), .ZN(n10090) );
  OAI21_X1 U11905 ( .B1(n17452), .B2(n18177), .A(n19507), .ZN(n19062) );
  NAND2_X1 U11906 ( .A1(n11894), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10109) );
  NOR2_X1 U11907 ( .A1(n19154), .A2(n9768), .ZN(n19069) );
  NOR2_X1 U11908 ( .A1(n9768), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U11909 ( .A1(n11902), .A2(n10641), .ZN(n11905) );
  AND2_X1 U11910 ( .A1(n13917), .A2(n19926), .ZN(n11740) );
  INV_X1 U11911 ( .A(n11922), .ZN(n19515) );
  INV_X1 U11912 ( .A(n21173), .ZN(n17640) );
  NOR2_X1 U11913 ( .A1(n21432), .A2(n14686), .ZN(n17628) );
  NAND2_X1 U11914 ( .A1(n13198), .A2(n13197), .ZN(n13201) );
  NAND2_X1 U11915 ( .A1(n13440), .A2(n13439), .ZN(n15544) );
  INV_X1 U11916 ( .A(n15611), .ZN(n15617) );
  NAND2_X1 U11917 ( .A1(n13415), .A2(n13414), .ZN(n15644) );
  XNOR2_X1 U11918 ( .A(n13465), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15203) );
  NAND2_X1 U11919 ( .A1(n15865), .A2(n10212), .ZN(n13207) );
  AND2_X1 U11920 ( .A1(n10213), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10212) );
  AND2_X1 U11921 ( .A1(n13151), .A2(n13131), .ZN(n21250) );
  NAND2_X1 U11922 ( .A1(n14687), .A2(n17711), .ZN(n16385) );
  INV_X1 U11923 ( .A(n16385), .ZN(n21274) );
  OR3_X1 U11924 ( .A1(n14260), .A2(n13519), .A3(n13521), .ZN(n13532) );
  INV_X1 U11925 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20814) );
  INV_X1 U11926 ( .A(n15182), .ZN(n10256) );
  NAND2_X1 U11927 ( .A1(n10255), .A2(n15180), .ZN(n10254) );
  NAND2_X1 U11928 ( .A1(n15181), .A2(n20235), .ZN(n10255) );
  OAI21_X1 U11929 ( .B1(n15178), .B2(n20260), .A(n15177), .ZN(n15179) );
  AOI21_X1 U11930 ( .B1(n16474), .B2(n15144), .A(n16897), .ZN(n16465) );
  NAND2_X1 U11931 ( .A1(n9866), .A2(n9864), .ZN(n9863) );
  INV_X1 U11932 ( .A(n9865), .ZN(n9864) );
  OR2_X1 U11933 ( .A1(n16793), .A2(n20267), .ZN(n9866) );
  OAI21_X1 U11934 ( .B1(n16479), .B2(n20260), .A(n16478), .ZN(n9865) );
  OR2_X1 U11935 ( .A1(n16476), .A2(n16678), .ZN(n9868) );
  NAND2_X1 U11936 ( .A1(n14498), .A2(n14572), .ZN(n14578) );
  OR2_X1 U11937 ( .A1(n13771), .A2(n13641), .ZN(n20368) );
  AND2_X1 U11938 ( .A1(n13742), .A2(n20929), .ZN(n14282) );
  NAND2_X1 U11939 ( .A1(n10185), .A2(n10189), .ZN(n10108) );
  NAND2_X1 U11940 ( .A1(n16923), .A2(n10192), .ZN(n10185) );
  INV_X1 U11941 ( .A(n17201), .ZN(n9883) );
  XNOR2_X1 U11942 ( .A(n14712), .B(n14713), .ZN(n16970) );
  NAND2_X1 U11943 ( .A1(n17723), .A2(n21041), .ZN(n17098) );
  AND2_X1 U11944 ( .A1(n17723), .A2(n13564), .ZN(n17714) );
  INV_X1 U11945 ( .A(n17098), .ZN(n17716) );
  AND2_X1 U11946 ( .A1(n13186), .A2(n21078), .ZN(n17719) );
  AOI21_X1 U11947 ( .B1(n9968), .B2(n13349), .A(n13350), .ZN(n13351) );
  OAI21_X1 U11948 ( .B1(n13348), .B2(n13384), .A(n12582), .ZN(n9968) );
  XNOR2_X1 U11949 ( .A(n13344), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14677) );
  AOI21_X1 U11950 ( .B1(n16690), .B2(n20356), .A(n13388), .ZN(n10298) );
  OR2_X1 U11951 ( .A1(n16772), .A2(n17372), .ZN(n10299) );
  NAND2_X1 U11952 ( .A1(n13251), .A2(n17152), .ZN(n9961) );
  XNOR2_X1 U11953 ( .A(n10087), .B(n9760), .ZN(n16903) );
  NOR2_X1 U11954 ( .A1(n13317), .A2(n13316), .ZN(n13340) );
  NAND2_X1 U11955 ( .A1(n16970), .A2(n17383), .ZN(n9922) );
  NAND2_X1 U11956 ( .A1(n17380), .A2(n17243), .ZN(n10174) );
  NAND2_X1 U11957 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  NAND2_X1 U11958 ( .A1(n17251), .A2(n14716), .ZN(n10152) );
  NAND2_X1 U11959 ( .A1(n16963), .A2(n17726), .ZN(n10153) );
  AND2_X1 U11960 ( .A1(n12998), .A2(n12804), .ZN(n20355) );
  INV_X1 U11961 ( .A(n17352), .ZN(n20356) );
  INV_X1 U11962 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21050) );
  INV_X1 U11963 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21692) );
  INV_X1 U11964 ( .A(n21065), .ZN(n21028) );
  NOR2_X1 U11965 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20546), .ZN(
        n20533) );
  NOR2_X1 U11966 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14595), .ZN(
        n20785) );
  NOR2_X1 U11967 ( .A1(n19980), .A2(n20102), .ZN(n20087) );
  NAND2_X1 U11968 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18417), .ZN(n18399) );
  AND2_X1 U11969 ( .A1(n18464), .A2(n10139), .ZN(n18417) );
  NOR2_X1 U11970 ( .A1(n18697), .A2(n10140), .ZN(n10139) );
  INV_X1 U11971 ( .A(n10141), .ZN(n10140) );
  NAND2_X1 U11972 ( .A1(n10138), .A2(n9769), .ZN(n10137) );
  NOR2_X1 U11973 ( .A1(n18644), .A2(n10135), .ZN(n18635) );
  AND2_X1 U11974 ( .A1(n18677), .A2(n9858), .ZN(n18661) );
  INV_X1 U11975 ( .A(n13245), .ZN(n18769) );
  NOR2_X1 U11976 ( .A1(n19521), .A2(n18655), .ZN(n18777) );
  NOR2_X1 U11977 ( .A1(n14115), .A2(n18655), .ZN(n18786) );
  NAND2_X1 U11978 ( .A1(n10340), .A2(n10339), .ZN(n10338) );
  NAND2_X1 U11979 ( .A1(n18910), .A2(n19113), .ZN(n10339) );
  INV_X1 U11980 ( .A(n13500), .ZN(n10337) );
  NOR2_X1 U11981 ( .A1(n19258), .A2(n10286), .ZN(n10285) );
  NAND2_X1 U11982 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  NAND2_X1 U11983 ( .A1(n19949), .A2(n19259), .ZN(n10287) );
  AOI21_X1 U11984 ( .B1(n10283), .B2(n19261), .A(n19459), .ZN(n10282) );
  OR2_X1 U11985 ( .A1(n19262), .A2(n19260), .ZN(n10283) );
  AND2_X1 U11986 ( .A1(n19443), .A2(n13245), .ZN(n19377) );
  INV_X1 U11987 ( .A(n19466), .ZN(n19468) );
  AND2_X1 U11988 ( .A1(n9879), .A2(n9878), .ZN(n12293) );
  AND2_X1 U11989 ( .A1(n14975), .A2(n15466), .ZN(n10901) );
  NAND2_X1 U11990 ( .A1(n10832), .A2(n13013), .ZN(n10895) );
  INV_X1 U11991 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U11992 ( .A1(n20709), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12207) );
  AND2_X1 U11993 ( .A1(n9921), .A2(n9920), .ZN(n12184) );
  NAND2_X1 U11994 ( .A1(n14952), .A2(n9793), .ZN(n9920) );
  NAND2_X1 U11995 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9921) );
  AOI22_X1 U11996 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U11997 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U11998 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12045) );
  AOI21_X1 U11999 ( .B1(n10667), .B2(n10665), .A(n10658), .ZN(n10660) );
  AND2_X1 U12000 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19938), .ZN(
        n10658) );
  OR2_X1 U12001 ( .A1(n10771), .A2(n10774), .ZN(n10773) );
  AND2_X1 U12002 ( .A1(n10773), .A2(n10762), .ZN(n10764) );
  OR2_X1 U12003 ( .A1(n10846), .A2(n10710), .ZN(n10714) );
  OR2_X1 U12004 ( .A1(n11124), .A2(n11123), .ZN(n11139) );
  AOI22_X1 U12005 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U12006 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10923), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U12007 ( .A1(n20446), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10025) );
  NAND2_X1 U12008 ( .A1(n14396), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U12009 ( .A1(n20446), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n9898) );
  NAND2_X1 U12010 ( .A1(n20599), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n9903) );
  NOR2_X1 U12011 ( .A1(n16479), .A2(n12994), .ZN(n12974) );
  NAND2_X1 U12012 ( .A1(n12609), .A2(n14604), .ZN(n12105) );
  NAND2_X1 U12013 ( .A1(n9957), .A2(n9955), .ZN(n9954) );
  NAND2_X1 U12014 ( .A1(n9956), .A2(n12388), .ZN(n9955) );
  NAND2_X1 U12015 ( .A1(n12410), .A2(n12453), .ZN(n9957) );
  INV_X1 U12016 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10290) );
  NAND2_X1 U12017 ( .A1(n9747), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U12018 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12007) );
  NAND2_X1 U12019 ( .A1(n12097), .A2(n12091), .ZN(n12424) );
  INV_X1 U12020 ( .A(n12432), .ZN(n12097) );
  OR2_X1 U12021 ( .A1(n10797), .A2(n10796), .ZN(n13004) );
  NAND2_X1 U12022 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10793), .ZN(
        n13005) );
  INV_X1 U12023 ( .A(n16094), .ZN(n13146) );
  INV_X1 U12024 ( .A(n15557), .ZN(n10881) );
  NAND2_X1 U12025 ( .A1(n15213), .A2(n10440), .ZN(n10439) );
  INV_X1 U12026 ( .A(n15225), .ZN(n10440) );
  AND2_X1 U12027 ( .A1(n11425), .A2(n11403), .ZN(n10441) );
  NAND2_X1 U12028 ( .A1(n13146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11685) );
  XNOR2_X1 U12029 ( .A(n11148), .B(n11137), .ZN(n11233) );
  AND2_X1 U12030 ( .A1(n9784), .A2(n11160), .ZN(n10097) );
  INV_X1 U12031 ( .A(n9818), .ZN(n9997) );
  NOR2_X1 U12032 ( .A1(n11161), .A2(n15793), .ZN(n15768) );
  NAND2_X1 U12033 ( .A1(n10272), .A2(n13080), .ZN(n10271) );
  INV_X1 U12034 ( .A(n10273), .ZN(n10272) );
  NAND2_X1 U12035 ( .A1(n15527), .A2(n10274), .ZN(n10273) );
  INV_X1 U12036 ( .A(n15533), .ZN(n10274) );
  INV_X1 U12037 ( .A(n11145), .ZN(n10099) );
  INV_X1 U12038 ( .A(n17652), .ZN(n10000) );
  OR2_X1 U12039 ( .A1(n14374), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11068) );
  OR2_X1 U12040 ( .A1(n11025), .A2(n11024), .ZN(n11062) );
  AND2_X1 U12041 ( .A1(n13906), .A2(n13166), .ZN(n13155) );
  OAI211_X1 U12042 ( .C1(n13040), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13034), .B(
        n13196), .ZN(n13035) );
  OR2_X1 U12043 ( .A1(n11179), .A2(n14287), .ZN(n11090) );
  NAND2_X1 U12044 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  NOR2_X1 U12045 ( .A1(n13011), .A2(n14090), .ZN(n10218) );
  NAND2_X1 U12046 ( .A1(n13012), .A2(n14090), .ZN(n10216) );
  INV_X1 U12047 ( .A(n10991), .ZN(n10984) );
  INV_X1 U12048 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14983) );
  NAND2_X1 U12049 ( .A1(n13134), .A2(n13119), .ZN(n14975) );
  NOR2_X1 U12050 ( .A1(n10882), .A2(n13144), .ZN(n14976) );
  NAND2_X1 U12051 ( .A1(n10867), .A2(n10866), .ZN(n10872) );
  NAND2_X1 U12052 ( .A1(n10922), .A2(n10921), .ZN(n14152) );
  OAI21_X1 U12053 ( .B1(n17708), .B2(n16074), .A(n16112), .ZN(n14032) );
  NAND2_X1 U12054 ( .A1(n10040), .A2(n10042), .ZN(n10805) );
  AND2_X1 U12055 ( .A1(n14697), .A2(n11146), .ZN(n10040) );
  NOR2_X1 U12056 ( .A1(n9755), .A2(n9833), .ZN(n10220) );
  NAND2_X1 U12057 ( .A1(n12811), .A2(n12816), .ZN(n9956) );
  OAI21_X1 U12058 ( .B1(n10238), .B2(n10241), .A(n16888), .ZN(n10240) );
  NOR2_X1 U12059 ( .A1(n16914), .A2(n10236), .ZN(n10235) );
  INV_X1 U12060 ( .A(n16909), .ZN(n10236) );
  NAND2_X1 U12061 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12064) );
  CLKBUF_X1 U12062 ( .A(n12001), .Z(n14953) );
  AND2_X1 U12063 ( .A1(n14801), .A2(n14800), .ZN(n14836) );
  INV_X1 U12064 ( .A(n16730), .ZN(n10069) );
  INV_X1 U12065 ( .A(n10066), .ZN(n10065) );
  AND2_X1 U12066 ( .A1(n14497), .A2(n10067), .ZN(n10066) );
  INV_X1 U12067 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U12068 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10247) );
  AND2_X1 U12069 ( .A1(n12977), .A2(n16882), .ZN(n10194) );
  NAND2_X1 U12070 ( .A1(n16919), .A2(n16920), .ZN(n10191) );
  NOR2_X1 U12071 ( .A1(n9813), .A2(n10247), .ZN(n15152) );
  NAND2_X1 U12072 ( .A1(n15135), .A2(n9767), .ZN(n15142) );
  NOR2_X1 U12073 ( .A1(n15136), .A2(n10259), .ZN(n10258) );
  INV_X1 U12074 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U12075 ( .A1(n15106), .A2(n10249), .ZN(n15113) );
  NAND2_X1 U12076 ( .A1(n10250), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10249) );
  AND2_X1 U12077 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U12078 ( .A1(n14904), .A2(n12195), .ZN(n10318) );
  NOR2_X1 U12079 ( .A1(n10190), .A2(n10173), .ZN(n10184) );
  INV_X1 U12080 ( .A(n10192), .ZN(n10188) );
  NAND2_X1 U12081 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  INV_X1 U12082 ( .A(n16460), .ZN(n10305) );
  OR2_X1 U12083 ( .A1(n12974), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13255) );
  AOI21_X1 U12084 ( .B1(n10171), .B2(n10172), .A(n10193), .ZN(n10170) );
  INV_X1 U12085 ( .A(n10402), .ZN(n10171) );
  AND2_X1 U12086 ( .A1(n16930), .A2(n10403), .ZN(n10402) );
  NAND2_X1 U12087 ( .A1(n10404), .A2(n16934), .ZN(n10403) );
  INV_X1 U12088 ( .A(n16933), .ZN(n10404) );
  INV_X1 U12089 ( .A(n13459), .ZN(n10302) );
  INV_X1 U12090 ( .A(n13490), .ZN(n12847) );
  NAND2_X1 U12091 ( .A1(n12845), .A2(n9823), .ZN(n10072) );
  NAND2_X1 U12092 ( .A1(n13490), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9890) );
  INV_X1 U12093 ( .A(n13278), .ZN(n10077) );
  AND2_X1 U12094 ( .A1(n9757), .A2(n14619), .ZN(n10420) );
  INV_X1 U12095 ( .A(n10366), .ZN(n10364) );
  NOR2_X1 U12096 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  INV_X1 U12097 ( .A(n14280), .ZN(n10311) );
  NAND2_X1 U12098 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  INV_X1 U12099 ( .A(n13807), .ZN(n10296) );
  INV_X1 U12100 ( .A(n13777), .ZN(n10297) );
  INV_X1 U12101 ( .A(n12347), .ZN(n10130) );
  AND3_X1 U12102 ( .A1(n12643), .A2(n12642), .A3(n12641), .ZN(n14569) );
  NOR2_X1 U12103 ( .A1(n10459), .A2(n12153), .ZN(n12154) );
  NAND2_X1 U12104 ( .A1(n12466), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12155) );
  OAI21_X1 U12105 ( .B1(n12499), .B2(n12152), .A(n12151), .ZN(n12153) );
  NAND2_X1 U12106 ( .A1(n9894), .A2(n12149), .ZN(n12480) );
  NAND2_X1 U12107 ( .A1(n9952), .A2(n9951), .ZN(n12416) );
  NAND2_X1 U12108 ( .A1(n21075), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9951) );
  NAND2_X1 U12109 ( .A1(n9953), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U12110 ( .A1(n9954), .A2(n12449), .ZN(n9953) );
  NAND2_X1 U12111 ( .A1(n12576), .A2(n12122), .ZN(n12568) );
  NAND2_X1 U12112 ( .A1(n14876), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13829) );
  NAND2_X1 U12113 ( .A1(n21045), .A2(n20874), .ZN(n14398) );
  AND2_X1 U12114 ( .A1(n21076), .A2(n21073), .ZN(n14204) );
  NOR3_X1 U12115 ( .A1(n18993), .A2(n18987), .A3(n10486), .ZN(n18937) );
  INV_X1 U12116 ( .A(n10328), .ZN(n10327) );
  OAI21_X1 U12117 ( .B1(n11869), .B2(n10332), .A(n11873), .ZN(n10328) );
  AND4_X1 U12118 ( .A1(n10630), .A2(n10629), .A3(n10628), .A4(n10627), .ZN(
        n10636) );
  NAND2_X1 U12119 ( .A1(n10182), .A2(n10114), .ZN(n10113) );
  INV_X1 U12120 ( .A(n10326), .ZN(n10114) );
  NAND2_X1 U12121 ( .A1(n10182), .A2(n19113), .ZN(n10115) );
  AND2_X1 U12122 ( .A1(n9852), .A2(n10345), .ZN(n10344) );
  OAI21_X1 U12123 ( .B1(n11924), .B2(n10674), .A(n11917), .ZN(n17850) );
  AND2_X1 U12124 ( .A1(n10652), .A2(n10468), .ZN(n13218) );
  OR2_X1 U12125 ( .A1(n10643), .A2(n10648), .ZN(n10652) );
  OR2_X1 U12126 ( .A1(n19414), .A2(n19174), .ZN(n19176) );
  NAND2_X1 U12127 ( .A1(n11930), .A2(n13998), .ZN(n11857) );
  OR2_X1 U12128 ( .A1(n10588), .A2(n10587), .ZN(n11898) );
  OR2_X1 U12129 ( .A1(n10560), .A2(n10559), .ZN(n10639) );
  OR2_X1 U12130 ( .A1(n10602), .A2(n10601), .ZN(n11899) );
  OR2_X1 U12131 ( .A1(n10616), .A2(n10617), .ZN(n11922) );
  OAI221_X1 U12132 ( .B1(n20102), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n19481), .A(n14124), .ZN(n19491) );
  NAND2_X1 U12133 ( .A1(n11921), .A2(n13918), .ZN(n13995) );
  NOR3_X1 U12134 ( .A1(n15432), .A2(n10045), .A3(n14694), .ZN(n15293) );
  INV_X1 U12135 ( .A(n14693), .ZN(n10046) );
  INV_X1 U12136 ( .A(n14057), .ZN(n15558) );
  NAND2_X1 U12137 ( .A1(n13970), .A2(n11194), .ZN(n13963) );
  NAND2_X1 U12138 ( .A1(n11642), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11668) );
  INV_X1 U12139 ( .A(n11644), .ZN(n11642) );
  NAND2_X1 U12140 ( .A1(n11618), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11619) );
  INV_X1 U12141 ( .A(n11617), .ZN(n11618) );
  NOR2_X1 U12142 ( .A1(n10427), .A2(n10125), .ZN(n10124) );
  INV_X1 U12143 ( .A(n10126), .ZN(n10125) );
  NAND2_X1 U12144 ( .A1(n11596), .A2(n10430), .ZN(n10427) );
  OR2_X1 U12145 ( .A1(n11574), .A2(n11503), .ZN(n11566) );
  NAND2_X1 U12146 ( .A1(n11485), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11574) );
  INV_X1 U12147 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U12148 ( .A1(n15349), .A2(n10128), .ZN(n10127) );
  INV_X1 U12149 ( .A(n10441), .ZN(n10128) );
  NAND2_X1 U12150 ( .A1(n11405), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11426) );
  INV_X1 U12151 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15364) );
  INV_X1 U12152 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15397) );
  AND3_X1 U12153 ( .A1(n15391), .A2(n15421), .A3(n15438), .ZN(n15422) );
  AND2_X1 U12154 ( .A1(n11293), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11369) );
  CLKBUF_X1 U12155 ( .A(n15387), .Z(n15388) );
  INV_X1 U12156 ( .A(n15538), .ZN(n10119) );
  AND2_X1 U12157 ( .A1(n10443), .A2(n15546), .ZN(n10123) );
  INV_X1 U12158 ( .A(n11234), .ZN(n11235) );
  NAND2_X1 U12159 ( .A1(n10129), .A2(n11126), .ZN(n11225) );
  OAI21_X1 U12160 ( .B1(n11176), .B2(n11364), .A(n11175), .ZN(n11177) );
  OR2_X1 U12161 ( .A1(n17587), .A2(n13026), .ZN(n17602) );
  OR2_X1 U12162 ( .A1(n13780), .A2(n11189), .ZN(n13796) );
  AND2_X1 U12163 ( .A1(n10449), .A2(n15653), .ZN(n10168) );
  OR3_X1 U12164 ( .A1(n15252), .A2(n10262), .A3(n10261), .ZN(n10260) );
  INV_X1 U12165 ( .A(n15227), .ZN(n10261) );
  NOR3_X1 U12166 ( .A1(n15266), .A2(n15252), .A3(n15267), .ZN(n15239) );
  NAND2_X1 U12167 ( .A1(n9940), .A2(n9939), .ZN(n15722) );
  INV_X1 U12168 ( .A(n10166), .ZN(n9940) );
  OAI21_X1 U12169 ( .B1(n11167), .B2(n10350), .A(n15729), .ZN(n10166) );
  AND2_X1 U12170 ( .A1(n13109), .A2(n13108), .ZN(n15310) );
  OR2_X1 U12171 ( .A1(n15958), .A2(n13158), .ZN(n15933) );
  AND2_X1 U12172 ( .A1(n13102), .A2(n13101), .ZN(n15325) );
  NAND2_X1 U12173 ( .A1(n15335), .A2(n13099), .ZN(n15336) );
  INV_X1 U12174 ( .A(n15338), .ZN(n13099) );
  NOR2_X1 U12175 ( .A1(n11157), .A2(n15816), .ZN(n10016) );
  NAND2_X1 U12176 ( .A1(n15729), .A2(n16040), .ZN(n15822) );
  CLKBUF_X1 U12177 ( .A(n15456), .Z(n15457) );
  INV_X1 U12178 ( .A(n15540), .ZN(n13069) );
  AND2_X1 U12179 ( .A1(n13053), .A2(n9839), .ZN(n15551) );
  NAND2_X1 U12180 ( .A1(n13053), .A2(n10281), .ZN(n14430) );
  INV_X1 U12181 ( .A(n13155), .ZN(n15965) );
  CLKBUF_X1 U12182 ( .A(n13028), .Z(n13559) );
  NAND2_X1 U12183 ( .A1(n15092), .A2(n21654), .ZN(n11720) );
  NAND2_X1 U12184 ( .A1(n13782), .A2(n11080), .ZN(n11083) );
  NAND2_X1 U12185 ( .A1(n10228), .A2(n9924), .ZN(n10227) );
  AND2_X1 U12186 ( .A1(n9925), .A2(n21654), .ZN(n9924) );
  NAND2_X1 U12187 ( .A1(n11181), .A2(n11052), .ZN(n11095) );
  CLKBUF_X1 U12188 ( .A(n10870), .Z(n16094) );
  AND2_X1 U12189 ( .A1(n14680), .A2(n14691), .ZN(n16090) );
  OR2_X1 U12190 ( .A1(n14024), .A2(n14069), .ZN(n14075) );
  INV_X1 U12191 ( .A(n14160), .ZN(n14340) );
  NAND2_X1 U12192 ( .A1(n14069), .A2(n15022), .ZN(n14160) );
  AND2_X1 U12193 ( .A1(n16248), .A2(n15019), .ZN(n16166) );
  AND3_X1 U12194 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21654), .A3(n14032), 
        .ZN(n14091) );
  INV_X1 U12195 ( .A(n9720), .ZN(n14156) );
  NOR2_X1 U12196 ( .A1(n16291), .A2(n16290), .ZN(n21272) );
  NOR2_X1 U12197 ( .A1(n14687), .A2(n21335), .ZN(n16074) );
  NAND2_X1 U12198 ( .A1(n12462), .A2(n12461), .ZN(n13178) );
  NOR2_X1 U12199 ( .A1(n12979), .A2(n9844), .ZN(n12984) );
  NAND2_X1 U12200 ( .A1(n10471), .A2(n13381), .ZN(n13383) );
  OAI211_X1 U12201 ( .C1(n10238), .C2(n10237), .A(n10234), .B(n10239), .ZN(
        n16450) );
  OR2_X1 U12202 ( .A1(n10238), .A2(n10235), .ZN(n10234) );
  INV_X1 U12204 ( .A(n10240), .ZN(n10239) );
  NOR2_X1 U12205 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  OR2_X1 U12206 ( .A1(n12956), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10380) );
  AND2_X1 U12207 ( .A1(n10237), .A2(n10242), .ZN(n16486) );
  INV_X1 U12208 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U12209 ( .A1(n12868), .A2(n10377), .ZN(n12876) );
  NAND2_X1 U12210 ( .A1(n20166), .A2(n16967), .ZN(n20146) );
  INV_X1 U12211 ( .A(n17012), .ZN(n9869) );
  NAND2_X1 U12212 ( .A1(n12910), .A2(n12899), .ZN(n12903) );
  NAND2_X1 U12214 ( .A1(n10372), .A2(n10371), .ZN(n10370) );
  INV_X1 U12215 ( .A(n10373), .ZN(n10372) );
  OAI211_X1 U12216 ( .C1(n12892), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12972), .B(
        n9919), .ZN(n20217) );
  NAND2_X1 U12217 ( .A1(n12892), .A2(n9825), .ZN(n9919) );
  OR2_X1 U12218 ( .A1(n16613), .A2(n17096), .ZN(n20241) );
  NAND2_X1 U12219 ( .A1(n20274), .A2(n17712), .ZN(n16613) );
  NAND2_X1 U12220 ( .A1(n12823), .A2(n12840), .ZN(n12820) );
  MUX2_X1 U12221 ( .A(n12807), .B(n12806), .S(n12123), .Z(n12827) );
  INV_X1 U12222 ( .A(n20255), .ZN(n20258) );
  NAND2_X1 U12223 ( .A1(n15170), .A2(n15169), .ZN(n20245) );
  NAND2_X2 U12224 ( .A1(n12605), .A2(n21077), .ZN(n12388) );
  OAI21_X1 U12225 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_0__SCAN_IN), .A(n9871), .ZN(n16665) );
  NAND2_X1 U12226 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9871) );
  NAND2_X1 U12227 ( .A1(n21069), .A2(n15173), .ZN(n20249) );
  INV_X1 U12228 ( .A(n16496), .ZN(n10303) );
  INV_X1 U12229 ( .A(n14874), .ZN(n10396) );
  AOI21_X1 U12230 ( .B1(n10394), .B2(n9837), .A(n10063), .ZN(n10058) );
  NAND2_X1 U12231 ( .A1(n16733), .A2(n16735), .ZN(n16734) );
  AND2_X1 U12232 ( .A1(n12773), .A2(n12772), .ZN(n13296) );
  NAND2_X1 U12233 ( .A1(n12775), .A2(n12774), .ZN(n13295) );
  OR2_X1 U12234 ( .A1(n14739), .A2(n14738), .ZN(n16750) );
  AND2_X1 U12235 ( .A1(n12766), .A2(n12765), .ZN(n14714) );
  AND2_X1 U12236 ( .A1(n12762), .A2(n12761), .ZN(n14503) );
  CLKBUF_X1 U12237 ( .A(n14561), .Z(n14562) );
  INV_X1 U12238 ( .A(n14506), .ZN(n14504) );
  INV_X1 U12239 ( .A(n12602), .ZN(n13751) );
  NOR2_X1 U12240 ( .A1(n9813), .A2(n10243), .ZN(n13393) );
  NAND2_X1 U12241 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  NOR2_X1 U12242 ( .A1(n12978), .A2(n10193), .ZN(n10192) );
  INV_X1 U12243 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16895) );
  NOR2_X1 U12244 ( .A1(n15142), .A2(n16916), .ZN(n15146) );
  NAND2_X1 U12245 ( .A1(n15135), .A2(n10258), .ZN(n15139) );
  AND2_X1 U12246 ( .A1(n10324), .A2(n9861), .ZN(n10323) );
  AND2_X1 U12247 ( .A1(n15125), .A2(n9841), .ZN(n15133) );
  NAND2_X1 U12248 ( .A1(n15125), .A2(n9766), .ZN(n15131) );
  NAND2_X1 U12249 ( .A1(n9911), .A2(n9910), .ZN(n14630) );
  AND2_X1 U12250 ( .A1(n15125), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15129) );
  NOR2_X1 U12251 ( .A1(n13288), .A2(n17268), .ZN(n10324) );
  NOR2_X1 U12252 ( .A1(n13287), .A2(n17329), .ZN(n10156) );
  OR2_X1 U12253 ( .A1(n17305), .A2(n13302), .ZN(n13287) );
  INV_X1 U12254 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20202) );
  INV_X1 U12255 ( .A(n15106), .ZN(n10248) );
  NOR2_X1 U12256 ( .A1(n15106), .A2(n10252), .ZN(n15111) );
  NOR2_X1 U12257 ( .A1(n15106), .A2(n17089), .ZN(n15107) );
  AND2_X1 U12258 ( .A1(n12344), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9966) );
  NAND2_X1 U12259 ( .A1(n10001), .A2(n12342), .ZN(n12343) );
  NAND2_X1 U12260 ( .A1(n10233), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15100) );
  NOR2_X1 U12261 ( .A1(n15100), .A2(n20259), .ZN(n15101) );
  NAND2_X1 U12262 ( .A1(n9891), .A2(n9892), .ZN(n10413) );
  NAND2_X1 U12263 ( .A1(n12161), .A2(n9893), .ZN(n9891) );
  AND2_X1 U12264 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15099) );
  INV_X1 U12265 ( .A(n13179), .ZN(n10422) );
  AND2_X1 U12266 ( .A1(n13254), .A2(n16905), .ZN(n16882) );
  NAND2_X1 U12267 ( .A1(n13252), .A2(n17153), .ZN(n13251) );
  NAND2_X1 U12268 ( .A1(n10169), .A2(n10170), .ZN(n16907) );
  AND2_X1 U12269 ( .A1(n12784), .A2(n12783), .ZN(n16497) );
  NOR2_X1 U12270 ( .A1(n17333), .A2(n12581), .ZN(n17212) );
  INV_X1 U12271 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17214) );
  AND2_X1 U12272 ( .A1(n12769), .A2(n12768), .ZN(n16840) );
  NAND2_X1 U12273 ( .A1(n16994), .A2(n10323), .ZN(n16953) );
  NOR3_X1 U12274 ( .A1(n14713), .A2(n10077), .A3(n10078), .ZN(n10074) );
  OR3_X1 U12275 ( .A1(n17278), .A2(n17268), .A3(n13302), .ZN(n17238) );
  CLKBUF_X1 U12276 ( .A(n14278), .Z(n14279) );
  AND2_X1 U12277 ( .A1(n17017), .A2(n17018), .ZN(n17007) );
  AND3_X1 U12278 ( .A1(n12720), .A2(n12719), .A3(n12718), .ZN(n13896) );
  NOR2_X1 U12279 ( .A1(n17030), .A2(n17032), .ZN(n17017) );
  OR2_X1 U12280 ( .A1(n13754), .A2(n13777), .ZN(n13806) );
  AND3_X1 U12281 ( .A1(n12665), .A2(n12664), .A3(n12663), .ZN(n13757) );
  CLKBUF_X1 U12282 ( .A(n13754), .Z(n13755) );
  INV_X1 U12283 ( .A(n17369), .ZN(n17259) );
  NAND2_X1 U12284 ( .A1(n9967), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17363) );
  AND2_X1 U12285 ( .A1(n17397), .A2(n17396), .ZN(n17369) );
  NAND2_X1 U12286 ( .A1(n17122), .A2(n17732), .ZN(n10410) );
  NOR2_X1 U12287 ( .A1(n10411), .A2(n10408), .ZN(n10407) );
  NAND2_X1 U12288 ( .A1(n9895), .A2(n12287), .ZN(n17114) );
  INV_X1 U12289 ( .A(n17106), .ZN(n12490) );
  INV_X1 U12290 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U12291 ( .A1(n14193), .A2(n14192), .ZN(n14195) );
  NAND2_X1 U12292 ( .A1(n14191), .A2(n12631), .ZN(n14567) );
  AOI21_X1 U12293 ( .B1(n13767), .B2(n13766), .A(n10400), .ZN(n13773) );
  INV_X1 U12294 ( .A(n13768), .ZN(n10400) );
  CLKBUF_X1 U12295 ( .A(n12455), .Z(n14229) );
  INV_X1 U12296 ( .A(n13840), .ZN(n13842) );
  INV_X1 U12297 ( .A(n20599), .ZN(n20604) );
  INV_X1 U12298 ( .A(n12218), .ZN(n20635) );
  NOR3_X1 U12299 ( .A1(n14396), .A2(n20806), .A3(n20864), .ZN(n14401) );
  OR2_X1 U12300 ( .A1(n21036), .A2(n21043), .ZN(n20539) );
  INV_X1 U12301 ( .A(n20405), .ZN(n20393) );
  INV_X1 U12302 ( .A(n20406), .ZN(n20391) );
  AND2_X1 U12303 ( .A1(n20874), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20407) );
  OR2_X1 U12304 ( .A1(n21036), .A2(n20369), .ZN(n20869) );
  NOR2_X2 U12305 ( .A1(n14399), .A2(n14398), .ZN(n20405) );
  NOR2_X2 U12306 ( .A1(n14505), .A2(n14398), .ZN(n20406) );
  AND2_X1 U12307 ( .A1(n12431), .A2(n12449), .ZN(n13523) );
  OR2_X1 U12308 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  INV_X1 U12309 ( .A(n12096), .ZN(n10390) );
  INV_X1 U12310 ( .A(n19992), .ZN(n20088) );
  AND2_X1 U12311 ( .A1(n11918), .A2(n11917), .ZN(n19950) );
  INV_X1 U12312 ( .A(n13243), .ZN(n19955) );
  INV_X1 U12313 ( .A(n10200), .ZN(n10199) );
  AOI21_X1 U12314 ( .B1(n10201), .B2(n9750), .A(n9750), .ZN(n10200) );
  NAND2_X1 U12315 ( .A1(n10494), .A2(n10493), .ZN(n17991) );
  NOR2_X1 U12316 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18074), .ZN(n18061) );
  NAND2_X1 U12317 ( .A1(n14113), .A2(n14667), .ZN(n18258) );
  NAND2_X1 U12318 ( .A1(n20105), .A2(n18798), .ZN(n10677) );
  OR2_X1 U12319 ( .A1(n10147), .A2(n21576), .ZN(n10146) );
  NAND2_X1 U12320 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .ZN(n10147) );
  AND2_X1 U12321 ( .A1(n9772), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U12322 ( .A1(n18464), .A2(n10141), .ZN(n18400) );
  NOR2_X1 U12323 ( .A1(n18531), .A2(n18514), .ZN(n18464) );
  NOR2_X1 U12324 ( .A1(n21456), .A2(n10145), .ZN(n10144) );
  INV_X1 U12325 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n10145) );
  AND2_X1 U12326 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10112) );
  OR2_X1 U12327 ( .A1(n11816), .A2(n11815), .ZN(n11950) );
  AND4_X1 U12328 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11786) );
  AOI22_X1 U12329 ( .A1(n11769), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U12330 ( .A1(n19515), .A2(n18659), .ZN(n14115) );
  OAI21_X1 U12331 ( .B1(n13927), .B2(n19967), .A(n20088), .ZN(n18796) );
  NOR4_X2 U12332 ( .A1(n19493), .A2(n11903), .A3(n18659), .A4(n10649), .ZN(
        n18856) );
  NAND2_X1 U12333 ( .A1(n10203), .A2(n10451), .ZN(n10202) );
  INV_X1 U12334 ( .A(n10204), .ZN(n10203) );
  NOR2_X1 U12335 ( .A1(n10483), .A2(n10488), .ZN(n10498) );
  NAND2_X1 U12336 ( .A1(n19202), .A2(n19059), .ZN(n17452) );
  INV_X1 U12337 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19133) );
  NAND2_X1 U12338 ( .A1(n10002), .A2(n9787), .ZN(n19185) );
  CLKBUF_X1 U12339 ( .A(n17446), .Z(n17447) );
  NOR2_X1 U12340 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20102), .ZN(n19059) );
  AND2_X1 U12341 ( .A1(n17578), .A2(n17741), .ZN(n9975) );
  AND2_X1 U12342 ( .A1(n19080), .A2(n13236), .ZN(n17512) );
  OR2_X1 U12343 ( .A1(n19398), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U12344 ( .A1(n18963), .A2(n11886), .ZN(n19039) );
  AND2_X1 U12345 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19037) );
  NAND2_X1 U12346 ( .A1(n9754), .A2(n10179), .ZN(n10178) );
  NOR2_X1 U12347 ( .A1(n19380), .A2(n19068), .ZN(n19329) );
  NAND2_X1 U12348 ( .A1(n19176), .A2(n11883), .ZN(n19115) );
  NAND2_X1 U12349 ( .A1(n10342), .A2(n10344), .ZN(n19125) );
  NAND2_X1 U12350 ( .A1(n10342), .A2(n10345), .ZN(n19143) );
  INV_X1 U12351 ( .A(n17850), .ZN(n19953) );
  NAND2_X1 U12352 ( .A1(n19174), .A2(n9983), .ZN(n9982) );
  NAND2_X2 U12353 ( .A1(n11883), .A2(n19081), .ZN(n19414) );
  NAND2_X1 U12354 ( .A1(n10005), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10004) );
  NAND2_X1 U12355 ( .A1(n11947), .A2(n10005), .ZN(n10003) );
  INV_X1 U12356 ( .A(n13816), .ZN(n10005) );
  NOR2_X1 U12357 ( .A1(n17458), .A2(n19449), .ZN(n17457) );
  NOR2_X2 U12358 ( .A1(n20106), .A2(n13995), .ZN(n19949) );
  AND2_X1 U12359 ( .A1(n14113), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13917) );
  INV_X1 U12360 ( .A(n11905), .ZN(n10092) );
  INV_X1 U12361 ( .A(n20089), .ZN(n19496) );
  INV_X1 U12362 ( .A(n11898), .ZN(n19500) );
  INV_X1 U12363 ( .A(n10639), .ZN(n19503) );
  INV_X1 U12364 ( .A(n11899), .ZN(n19508) );
  INV_X1 U12365 ( .A(n19565), .ZN(n19783) );
  INV_X1 U12366 ( .A(n19507), .ZN(n19871) );
  NAND2_X1 U12367 ( .A1(n20092), .A2(n19491), .ZN(n19565) );
  AOI21_X1 U12368 ( .B1(n19948), .B2(n19950), .A(n11926), .ZN(n19959) );
  NOR2_X1 U12369 ( .A1(n19955), .A2(n19947), .ZN(n11926) );
  NAND2_X2 U12370 ( .A1(n13484), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n14505)
         );
  NAND2_X1 U12371 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  NAND2_X1 U12372 ( .A1(n15196), .A2(n15194), .ZN(n21432) );
  INV_X1 U12373 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15460) );
  OR2_X1 U12374 ( .A1(n15476), .A2(n14689), .ZN(n21161) );
  NAND2_X1 U12375 ( .A1(n10043), .A2(n9849), .ZN(n21173) );
  INV_X1 U12376 ( .A(n15476), .ZN(n10043) );
  OR2_X1 U12377 ( .A1(n17628), .A2(n17711), .ZN(n21149) );
  OR2_X1 U12378 ( .A1(n15476), .A2(n14701), .ZN(n21122) );
  INV_X1 U12379 ( .A(n21149), .ZN(n21174) );
  INV_X1 U12380 ( .A(n21161), .ZN(n21176) );
  INV_X1 U12381 ( .A(n15545), .ZN(n15554) );
  INV_X1 U12382 ( .A(n15544), .ZN(n15553) );
  INV_X1 U12383 ( .A(n15536), .ZN(n15530) );
  INV_X1 U12384 ( .A(n15639), .ZN(n15646) );
  INV_X1 U12385 ( .A(n21220), .ZN(n21206) );
  INV_X2 U12386 ( .A(n21218), .ZN(n21435) );
  OR3_X1 U12387 ( .A1(n17587), .A2(n13673), .A3(n21089), .ZN(n21220) );
  AOI21_X1 U12388 ( .B1(n16090), .B2(n14690), .A(n17613), .ZN(n13673) );
  AND2_X1 U12389 ( .A1(n14283), .A2(n21340), .ZN(n14284) );
  OAI211_X1 U12390 ( .C1(n15223), .C2(n10434), .A(n10432), .B(n10431), .ZN(
        n14678) );
  NAND2_X1 U12391 ( .A1(n10436), .A2(n10433), .ZN(n10431) );
  NAND2_X1 U12392 ( .A1(n10435), .A2(n13407), .ZN(n10434) );
  INV_X1 U12393 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15743) );
  INV_X1 U12394 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15761) );
  INV_X1 U12395 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15849) );
  INV_X1 U12396 ( .A(n17665), .ZN(n17655) );
  AND2_X1 U12397 ( .A1(n15450), .A2(n15547), .ZN(n21131) );
  INV_X1 U12398 ( .A(n17669), .ZN(n15856) );
  INV_X1 U12399 ( .A(n17671), .ZN(n15857) );
  NAND2_X1 U12400 ( .A1(n21430), .A2(n14159), .ZN(n17666) );
  NAND2_X1 U12401 ( .A1(n15652), .A2(n15651), .ZN(n15654) );
  NAND2_X1 U12402 ( .A1(n9941), .A2(n10449), .ZN(n15652) );
  OR2_X1 U12403 ( .A1(n15933), .A2(n13161), .ZN(n15908) );
  INV_X1 U12404 ( .A(n10035), .ZN(n15689) );
  AND2_X1 U12405 ( .A1(n13162), .A2(n10222), .ZN(n10221) );
  AND2_X1 U12406 ( .A1(n10226), .A2(n13163), .ZN(n10222) );
  INV_X1 U12407 ( .A(n13167), .ZN(n10226) );
  NAND2_X1 U12408 ( .A1(n15937), .A2(n10225), .ZN(n15907) );
  AND2_X1 U12409 ( .A1(n13162), .A2(n13163), .ZN(n10225) );
  NOR2_X1 U12410 ( .A1(n10224), .A2(n10223), .ZN(n15917) );
  INV_X1 U12411 ( .A(n13162), .ZN(n10223) );
  OR2_X1 U12412 ( .A1(n15758), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15739) );
  AND2_X1 U12413 ( .A1(n15844), .A2(n15843), .ZN(n16065) );
  NOR2_X1 U12414 ( .A1(n9818), .A2(n9935), .ZN(n15853) );
  NAND2_X1 U12415 ( .A1(n17651), .A2(n11145), .ZN(n15854) );
  AND2_X1 U12416 ( .A1(n9989), .A2(n11114), .ZN(n14424) );
  AND2_X1 U12417 ( .A1(n13984), .A2(n16025), .ZN(n17692) );
  NAND2_X1 U12418 ( .A1(n11181), .A2(n11180), .ZN(n16079) );
  AOI21_X1 U12419 ( .B1(n15021), .B2(n15020), .A(n15019), .ZN(n21258) );
  NOR2_X1 U12420 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15092) );
  NAND2_X1 U12421 ( .A1(n13734), .A2(n13733), .ZN(n16116) );
  OAI21_X1 U12422 ( .B1(n14073), .B2(n14072), .A(n21281), .ZN(n14095) );
  OAI21_X1 U12423 ( .B1(n16159), .B2(n21276), .A(n14071), .ZN(n14093) );
  NAND2_X1 U12424 ( .A1(n14541), .A2(n16345), .ZN(n16190) );
  OAI22_X1 U12425 ( .A1(n14540), .A2(n14539), .B1(n14687), .B2(n16161), .ZN(
        n14556) );
  INV_X1 U12426 ( .A(n16190), .ZN(n14558) );
  NAND2_X1 U12427 ( .A1(n14340), .A2(n16287), .ZN(n16238) );
  INV_X1 U12428 ( .A(n16238), .ZN(n16197) );
  NAND2_X1 U12429 ( .A1(n14340), .A2(n16346), .ZN(n16280) );
  NAND2_X1 U12430 ( .A1(n14340), .A2(n16345), .ZN(n16281) );
  INV_X1 U12431 ( .A(n15083), .ZN(n14181) );
  OAI22_X1 U12432 ( .A1(n15058), .A2(n16385), .B1(n16298), .B2(n15055), .ZN(
        n15087) );
  OAI21_X1 U12433 ( .B1(n15036), .B2(n15035), .A(n21281), .ZN(n21267) );
  INV_X1 U12434 ( .A(n21266), .ZN(n14467) );
  AND2_X1 U12435 ( .A1(n14034), .A2(n9720), .ZN(n21753) );
  NOR2_X1 U12436 ( .A1(n16202), .A2(n14040), .ZN(n21288) );
  NOR2_X1 U12437 ( .A1(n16202), .A2(n14092), .ZN(n21294) );
  NOR2_X1 U12438 ( .A1(n16202), .A2(n14044), .ZN(n21300) );
  NOR2_X1 U12439 ( .A1(n16202), .A2(n14371), .ZN(n21306) );
  NOR2_X1 U12440 ( .A1(n16202), .A2(n14350), .ZN(n21312) );
  NOR2_X1 U12441 ( .A1(n16202), .A2(n14534), .ZN(n21318) );
  NOR2_X1 U12442 ( .A1(n16202), .A2(n15645), .ZN(n21325) );
  OAI21_X1 U12443 ( .B1(n21283), .B2(n21282), .A(n21281), .ZN(n21330) );
  INV_X1 U12444 ( .A(n21329), .ZN(n16375) );
  INV_X1 U12445 ( .A(n21278), .ZN(n16394) );
  INV_X1 U12446 ( .A(n16295), .ZN(n21279) );
  INV_X1 U12447 ( .A(n21288), .ZN(n16399) );
  INV_X1 U12448 ( .A(n16304), .ZN(n21289) );
  INV_X1 U12449 ( .A(n21748), .ZN(n21295) );
  INV_X1 U12450 ( .A(n21294), .ZN(n21750) );
  INV_X1 U12451 ( .A(n21300), .ZN(n16407) );
  INV_X1 U12452 ( .A(n16312), .ZN(n21301) );
  INV_X1 U12453 ( .A(n21312), .ZN(n16417) );
  INV_X1 U12454 ( .A(n16322), .ZN(n21313) );
  INV_X1 U12455 ( .A(n21318), .ZN(n16422) );
  INV_X1 U12456 ( .A(n16327), .ZN(n21319) );
  INV_X1 U12457 ( .A(n21325), .ZN(n16431) );
  NAND2_X1 U12458 ( .A1(n21280), .A2(n16345), .ZN(n16424) );
  INV_X1 U12459 ( .A(n16333), .ZN(n21327) );
  INV_X1 U12460 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21335) );
  INV_X1 U12461 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n17711) );
  INV_X1 U12462 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21357) );
  NAND2_X1 U12463 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21434) );
  INV_X1 U12464 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21359) );
  NAND2_X1 U12465 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n21073) );
  INV_X1 U12466 ( .A(n16688), .ZN(n16651) );
  INV_X1 U12467 ( .A(n20245), .ZN(n20266) );
  AND2_X1 U12468 ( .A1(n12920), .A2(n12919), .ZN(n20189) );
  NAND2_X1 U12469 ( .A1(n20212), .A2(n20211), .ZN(n20215) );
  INV_X1 U12470 ( .A(n20933), .ZN(n20276) );
  INV_X1 U12471 ( .A(n20249), .ZN(n20264) );
  AND2_X1 U12472 ( .A1(n20249), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20255) );
  OR2_X1 U12473 ( .A1(n13450), .A2(n13449), .ZN(n16738) );
  OR2_X1 U12474 ( .A1(n12677), .A2(n12676), .ZN(n14616) );
  NOR2_X1 U12475 ( .A1(n14416), .A2(n14407), .ZN(n14617) );
  OR2_X1 U12476 ( .A1(n12662), .A2(n12661), .ZN(n14474) );
  INV_X2 U12477 ( .A(n20291), .ZN(n16764) );
  INV_X1 U12478 ( .A(n20283), .ZN(n20288) );
  INV_X1 U12479 ( .A(n21043), .ZN(n20369) );
  NAND2_X1 U12480 ( .A1(n12602), .A2(n20291), .ZN(n20283) );
  XNOR2_X1 U12481 ( .A(n10057), .B(n10056), .ZN(n14973) );
  INV_X1 U12482 ( .A(n14963), .ZN(n10056) );
  NAND2_X1 U12483 ( .A1(n10055), .A2(n10054), .ZN(n10057) );
  NAND2_X1 U12484 ( .A1(n10385), .A2(n16697), .ZN(n16692) );
  NAND2_X1 U12485 ( .A1(n14905), .A2(n10386), .ZN(n10385) );
  NOR2_X1 U12486 ( .A1(n16725), .A2(n14818), .ZN(n16720) );
  AND2_X1 U12487 ( .A1(n14282), .A2(n13744), .ZN(n16858) );
  NAND2_X1 U12488 ( .A1(n14504), .A2(n14505), .ZN(n16859) );
  AND2_X1 U12489 ( .A1(n16868), .A2(n20311), .ZN(n14582) );
  NAND2_X1 U12490 ( .A1(n14012), .A2(n14011), .ZN(n14576) );
  OR2_X1 U12491 ( .A1(n14504), .A2(n16858), .ZN(n14579) );
  AND2_X1 U12492 ( .A1(n14282), .A2(n13751), .ZN(n20307) );
  INV_X1 U12493 ( .A(n20311), .ZN(n20295) );
  INV_X1 U12494 ( .A(n14579), .ZN(n20315) );
  AND2_X1 U12495 ( .A1(n13689), .A2(n21076), .ZN(n20321) );
  INV_X1 U12496 ( .A(n13570), .ZN(n20351) );
  AND2_X1 U12497 ( .A1(n16501), .A2(n16500), .ZN(n16918) );
  NAND2_X1 U12498 ( .A1(n16994), .A2(n10322), .ZN(n10321) );
  AND2_X1 U12499 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10322) );
  AND2_X1 U12500 ( .A1(n10156), .A2(n10324), .ZN(n10155) );
  OR2_X1 U12501 ( .A1(n14589), .A2(n14588), .ZN(n17281) );
  INV_X1 U12502 ( .A(n17714), .ZN(n17112) );
  CLKBUF_X1 U12503 ( .A(n13952), .Z(n13953) );
  INV_X1 U12504 ( .A(n13834), .ZN(n13661) );
  NOR2_X1 U12505 ( .A1(n12599), .A2(n12598), .ZN(n12600) );
  XNOR2_X1 U12506 ( .A(n9885), .B(n12996), .ZN(n13399) );
  NOR2_X1 U12507 ( .A1(n15189), .A2(n12994), .ZN(n12995) );
  XNOR2_X1 U12508 ( .A(n12383), .B(n12382), .ZN(n13402) );
  XNOR2_X1 U12509 ( .A(n9943), .B(n16875), .ZN(n17146) );
  INV_X1 U12510 ( .A(n9945), .ZN(n9944) );
  OAI21_X1 U12511 ( .B1(n16913), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n9904), .ZN(n17190) );
  NAND2_X1 U12512 ( .A1(n10401), .A2(n16934), .ZN(n16931) );
  NAND2_X1 U12513 ( .A1(n16935), .A2(n16933), .ZN(n10401) );
  AND2_X1 U12514 ( .A1(n16496), .A2(n16514), .ZN(n17204) );
  NOR2_X1 U12515 ( .A1(n16951), .A2(n20358), .ZN(n13313) );
  AOI21_X1 U12516 ( .B1(n13442), .B2(n13284), .A(n13283), .ZN(n13285) );
  NAND2_X1 U12517 ( .A1(n10355), .A2(n16954), .ZN(n10036) );
  INV_X1 U12518 ( .A(n17238), .ZN(n17251) );
  INV_X1 U12519 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17250) );
  NOR2_X1 U12520 ( .A1(n13858), .A2(n10314), .ZN(n14003) );
  NAND2_X1 U12521 ( .A1(n10365), .A2(n10366), .ZN(n16995) );
  NAND2_X1 U12522 ( .A1(n9899), .A2(n17274), .ZN(n17003) );
  INV_X1 U12523 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17319) );
  OR2_X1 U12524 ( .A1(n17340), .A2(n12591), .ZN(n17333) );
  NAND2_X1 U12525 ( .A1(n20364), .A2(n17367), .ZN(n17340) );
  OR2_X1 U12526 ( .A1(n17397), .A2(n12580), .ZN(n17731) );
  NAND2_X1 U12527 ( .A1(n10412), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17120) );
  NAND2_X1 U12528 ( .A1(n10409), .A2(n17732), .ZN(n17121) );
  NAND2_X1 U12529 ( .A1(n12998), .A2(n12577), .ZN(n14709) );
  INV_X1 U12530 ( .A(n17397), .ZN(n17380) );
  INV_X1 U12531 ( .A(n16684), .ZN(n17393) );
  INV_X1 U12532 ( .A(n20368), .ZN(n20421) );
  NOR2_X1 U12533 ( .A1(n21065), .A2(n20814), .ZN(n21045) );
  INV_X1 U12534 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21494) );
  NOR2_X1 U12535 ( .A1(n20874), .A2(n17405), .ZN(n21051) );
  AOI21_X1 U12536 ( .B1(n13941), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13638), .ZN(n13639) );
  AND2_X1 U12537 ( .A1(n14314), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U12538 ( .B1(n13773), .B2(n13772), .A(n13832), .ZN(n21043) );
  NAND2_X1 U12539 ( .A1(n20376), .A2(n20375), .ZN(n20411) );
  NAND2_X1 U12540 ( .A1(n20447), .A2(n21024), .ZN(n20505) );
  INV_X1 U12541 ( .A(n20492), .ZN(n20508) );
  OAI21_X1 U12542 ( .B1(n20483), .B2(n20482), .A(n20481), .ZN(n20507) );
  OAI21_X1 U12543 ( .B1(n20518), .B2(n20517), .A(n20516), .ZN(n20536) );
  NOR2_X1 U12544 ( .A1(n20514), .A2(n20512), .ZN(n20534) );
  OAI21_X1 U12545 ( .B1(n20547), .B2(n20546), .A(n20545), .ZN(n20565) );
  NOR2_X1 U12546 ( .A1(n20820), .A2(n20570), .ZN(n20592) );
  OAI21_X1 U12547 ( .B1(n20602), .B2(n21065), .A(n20600), .ZN(n20621) );
  OAI21_X1 U12548 ( .B1(n20680), .B2(n20679), .A(n20678), .ZN(n20701) );
  NOR2_X1 U12549 ( .A1(n20671), .A2(n20674), .ZN(n20711) );
  NOR2_X2 U12550 ( .A1(n20813), .A2(n20741), .ZN(n20735) );
  OAI21_X1 U12551 ( .B1(n20740), .B2(n20708), .A(n20707), .ZN(n20730) );
  INV_X1 U12552 ( .A(n20888), .ZN(n20754) );
  INV_X1 U12553 ( .A(n20900), .ZN(n20760) );
  INV_X1 U12554 ( .A(n20906), .ZN(n20763) );
  INV_X1 U12555 ( .A(n20735), .ZN(n20772) );
  OAI21_X1 U12556 ( .B1(n14603), .B2(n20511), .A(n14602), .ZN(n20786) );
  AOI211_X2 U12557 ( .C1(n14595), .C2(n20864), .A(n20571), .B(n14401), .ZN(
        n20807) );
  INV_X1 U12558 ( .A(n20885), .ZN(n20832) );
  INV_X1 U12559 ( .A(n20891), .ZN(n20835) );
  INV_X1 U12560 ( .A(n20903), .ZN(n20843) );
  OAI21_X1 U12561 ( .B1(n20827), .B2(n20826), .A(n20825), .ZN(n20858) );
  AOI211_X2 U12562 ( .C1(n20824), .C2(n20826), .A(n20823), .B(n20822), .ZN(
        n20861) );
  AND2_X1 U12563 ( .A1(n20407), .A2(n21077), .ZN(n20866) );
  AND2_X1 U12564 ( .A1(n20407), .A2(n21078), .ZN(n20880) );
  OAI22_X1 U12565 ( .A1(n17831), .A2(n20393), .B1(n17764), .B2(n20391), .ZN(
        n20888) );
  AND2_X1 U12566 ( .A1(n20407), .A2(n14609), .ZN(n20886) );
  OAI22_X1 U12567 ( .A1(n17762), .A2(n20391), .B1(n17834), .B2(n20393), .ZN(
        n20894) );
  OAI22_X1 U12568 ( .A1(n20387), .A2(n20391), .B1(n16780), .B2(n20393), .ZN(
        n20900) );
  AND2_X1 U12569 ( .A1(n20407), .A2(n9874), .ZN(n20898) );
  AND2_X1 U12570 ( .A1(n20407), .A2(n12812), .ZN(n20904) );
  AND2_X1 U12571 ( .A1(n20407), .A2(n20400), .ZN(n20910) );
  AND2_X1 U12572 ( .A1(n20407), .A2(n12602), .ZN(n20916) );
  AND2_X1 U12573 ( .A1(n20873), .A2(n20865), .ZN(n20919) );
  INV_X1 U12574 ( .A(n14316), .ZN(n12464) );
  INV_X1 U12575 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20864) );
  NOR3_X1 U12576 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20947), .A3(n20949), 
        .ZN(n21076) );
  INV_X1 U12577 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20959) );
  NOR2_X1 U12578 ( .A1(n19952), .A2(n18857), .ZN(n20105) );
  NOR2_X1 U12579 ( .A1(n20050), .A2(n17912), .ZN(n17880) );
  NOR2_X1 U12580 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17979), .ZN(n17970) );
  OAI21_X1 U12581 ( .B1(n10494), .B2(n9750), .A(n10201), .ZN(n17977) );
  INV_X1 U12582 ( .A(n19060), .ZN(n10208) );
  INV_X1 U12583 ( .A(n10209), .ZN(n18011) );
  INV_X1 U12584 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n21456) );
  NOR2_X1 U12585 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18122), .ZN(n18108) );
  INV_X1 U12586 ( .A(n18217), .ZN(n18158) );
  INV_X1 U12587 ( .A(n18171), .ZN(n18226) );
  NAND2_X1 U12588 ( .A1(n18212), .A2(n18205), .ZN(n18156) );
  AND4_X1 U12589 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10545) );
  AND4_X1 U12590 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10546) );
  NAND2_X1 U12591 ( .A1(n18375), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n18367) );
  INV_X1 U12592 ( .A(n18367), .ZN(n18372) );
  NOR3_X1 U12593 ( .A1(n18399), .A2(n17924), .A3(n10146), .ZN(n18375) );
  NOR2_X1 U12594 ( .A1(n18399), .A2(n10146), .ZN(n18380) );
  NAND2_X1 U12595 ( .A1(n18464), .A2(n10467), .ZN(n18465) );
  INV_X1 U12596 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n18514) );
  AND2_X1 U12597 ( .A1(n18601), .A2(n10143), .ZN(n18532) );
  AND2_X1 U12598 ( .A1(n9770), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U12599 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18532), .ZN(n18531) );
  NAND2_X1 U12600 ( .A1(n18601), .A2(n9770), .ZN(n18547) );
  NAND2_X1 U12601 ( .A1(n18601), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n18581) );
  NOR2_X1 U12602 ( .A1(n18097), .A2(n18621), .ZN(n18601) );
  NOR3_X1 U12603 ( .A1(n18626), .A2(n18123), .A3(n18629), .ZN(n18625) );
  OR2_X1 U12604 ( .A1(n18644), .A2(n10134), .ZN(n18626) );
  OR2_X1 U12605 ( .A1(n10135), .A2(n18155), .ZN(n10134) );
  INV_X1 U12606 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18629) );
  INV_X1 U12607 ( .A(n18687), .ZN(n18683) );
  NAND2_X1 U12608 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18683), .ZN(n18682) );
  NOR2_X1 U12609 ( .A1(n18692), .A2(n18697), .ZN(n18688) );
  NAND2_X1 U12610 ( .A1(n18688), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18687) );
  NOR2_X1 U12611 ( .A1(n18731), .A2(n10089), .ZN(n18693) );
  NAND2_X1 U12612 ( .A1(n18693), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18692) );
  NOR3_X1 U12613 ( .A1(n18655), .A2(n18740), .A3(n18654), .ZN(n18656) );
  NOR2_X1 U12614 ( .A1(n18740), .A2(n18739), .ZN(n18771) );
  INV_X1 U12615 ( .A(n11950), .ZN(n18772) );
  OR2_X1 U12616 ( .A1(n11801), .A2(n11800), .ZN(n18775) );
  INV_X1 U12617 ( .A(n18795), .ZN(n18787) );
  NOR2_X1 U12618 ( .A1(n18857), .A2(n18796), .ZN(n18841) );
  CLKBUF_X1 U12619 ( .A(n18898), .Z(n18896) );
  NOR3_X1 U12620 ( .A1(n20089), .A2(n18858), .A3(n18857), .ZN(n18898) );
  NOR2_X1 U12622 ( .A1(n18904), .A2(n19496), .ZN(n18905) );
  OR2_X1 U12623 ( .A1(n18925), .A2(n19225), .ZN(n10008) );
  NOR2_X1 U12624 ( .A1(n19010), .A2(n17578), .ZN(n10007) );
  OR2_X1 U12625 ( .A1(n13515), .A2(n13514), .ZN(n10335) );
  OAI22_X1 U12626 ( .A1(n13216), .A2(n19210), .B1(n17512), .B2(n19177), .ZN(
        n18925) );
  NAND2_X1 U12627 ( .A1(n10207), .A2(n10465), .ZN(n10206) );
  INV_X1 U12628 ( .A(n10483), .ZN(n10207) );
  INV_X1 U12629 ( .A(n19048), .ZN(n19067) );
  OAI22_X1 U12630 ( .A1(n19065), .A2(n19078), .B1(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9934) );
  NOR2_X1 U12631 ( .A1(n19067), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9931) );
  OAI211_X1 U12632 ( .C1(n19066), .C2(n10181), .A(n9929), .B(n9928), .ZN(n9927) );
  OR2_X1 U12633 ( .A1(n19076), .A2(n19065), .ZN(n9929) );
  NAND2_X1 U12634 ( .A1(n19128), .A2(n19325), .ZN(n9928) );
  INV_X1 U12635 ( .A(n19064), .ZN(n9930) );
  NAND2_X1 U12636 ( .A1(n19062), .A2(n19061), .ZN(n19121) );
  INV_X1 U12637 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19481) );
  NAND2_X1 U12638 ( .A1(n18909), .A2(n17578), .ZN(n17576) );
  NAND2_X1 U12639 ( .A1(n13239), .A2(n13238), .ZN(n13241) );
  NOR2_X1 U12640 ( .A1(n18943), .A2(n10110), .ZN(n9980) );
  INV_X1 U12641 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n20102) );
  NOR2_X1 U12642 ( .A1(n19080), .A2(n19381), .ZN(n10275) );
  NAND2_X1 U12643 ( .A1(n10331), .A2(n11869), .ZN(n13823) );
  NAND2_X1 U12644 ( .A1(n13810), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10331) );
  INV_X1 U12645 ( .A(n10002), .ZN(n13820) );
  AND2_X1 U12646 ( .A1(n19948), .A2(n19470), .ZN(n19476) );
  INV_X1 U12647 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10656) );
  INV_X1 U12648 ( .A(n17560), .ZN(n20086) );
  NOR3_X1 U12649 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n17849), .ZN(n19837) );
  INV_X1 U12650 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19938) );
  INV_X1 U12651 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19943) );
  NOR2_X1 U12652 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20070), .ZN(
        n19965) );
  NOR2_X1 U12653 ( .A1(n19492), .A2(n13932), .ZN(n14139) );
  INV_X1 U12654 ( .A(n14139), .ZN(n17569) );
  NOR2_X1 U12655 ( .A1(n19500), .A2(n19520), .ZN(n19885) );
  NOR2_X1 U12656 ( .A1(n19503), .A2(n19520), .ZN(n19891) );
  INV_X1 U12657 ( .A(n20083), .ZN(n20090) );
  NAND2_X1 U12658 ( .A1(n19481), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19980) );
  OAI211_X1 U12659 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n20001), .B(n20062), .ZN(n19992) );
  OR2_X1 U12660 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19988), .ZN(n20099) );
  INV_X1 U12661 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21426) );
  NOR2_X1 U12662 ( .A1(n14505), .A2(n13485), .ZN(n17755) );
  NOR2_X1 U12663 ( .A1(n17798), .A2(n17755), .ZN(n17803) );
  NOR2_X1 U12664 ( .A1(n15219), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U12665 ( .A1(n15648), .A2(n21170), .ZN(n10050) );
  OAI21_X1 U12666 ( .B1(n15212), .B2(n15545), .A(n10265), .ZN(P1_U2842) );
  AOI21_X1 U12667 ( .B1(n15200), .B2(n15536), .A(n10266), .ZN(n10265) );
  NOR2_X1 U12668 ( .A1(n15544), .A2(n13441), .ZN(n10266) );
  INV_X1 U12669 ( .A(n15200), .ZN(n15564) );
  INV_X1 U12670 ( .A(n13208), .ZN(n13209) );
  NAND2_X1 U12671 ( .A1(n10257), .A2(n10253), .ZN(P2_U2825) );
  NAND2_X1 U12672 ( .A1(n15160), .A2(n15161), .ZN(n10257) );
  NAND2_X1 U12673 ( .A1(n9867), .A2(n9862), .ZN(P2_U2829) );
  NAND2_X1 U12674 ( .A1(n16475), .A2(n9868), .ZN(n9867) );
  AOI21_X1 U12675 ( .B1(n16480), .B2(n20269), .A(n9863), .ZN(n9862) );
  INV_X1 U12676 ( .A(n10107), .ZN(n13188) );
  INV_X1 U12677 ( .A(n16893), .ZN(n9959) );
  OAI21_X1 U12678 ( .B1(n17206), .B2(n17116), .A(n9881), .ZN(P2_U2991) );
  AOI21_X1 U12679 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9881) );
  OAI21_X1 U12680 ( .B1(n17199), .B2(n17098), .A(n16932), .ZN(n9882) );
  NOR2_X1 U12681 ( .A1(n17200), .A2(n17136), .ZN(n9884) );
  OR2_X1 U12682 ( .A1(n13341), .A2(n17136), .ZN(n13330) );
  OAI211_X1 U12683 ( .C1(n14677), .C2(n20358), .A(n9949), .B(n9948), .ZN(
        P2_U3016) );
  NAND2_X1 U12684 ( .A1(n14674), .A2(n17383), .ZN(n9948) );
  AND2_X1 U12685 ( .A1(n10299), .A2(n10298), .ZN(n13389) );
  NAND2_X1 U12686 ( .A1(n17162), .A2(n17726), .ZN(n10082) );
  OAI21_X1 U12687 ( .B1(n16903), .B2(n20360), .A(n13269), .ZN(n13270) );
  OR2_X1 U12688 ( .A1(n13341), .A2(n20360), .ZN(n13342) );
  NAND2_X1 U12689 ( .A1(n10154), .A2(n10148), .ZN(P2_U3029) );
  NAND2_X1 U12690 ( .A1(n9922), .A2(n10150), .ZN(n10149) );
  NOR2_X1 U12691 ( .A1(n18399), .A2(n18356), .ZN(n18381) );
  NOR2_X1 U12692 ( .A1(n18644), .A2(n10137), .ZN(n18632) );
  INV_X1 U12693 ( .A(n18661), .ZN(n18665) );
  OAI21_X1 U12694 ( .B1(n10336), .B2(n13499), .A(n10334), .ZN(P3_U2802) );
  OAI21_X1 U12695 ( .B1(n10338), .B2(n10337), .A(n19128), .ZN(n10336) );
  NOR2_X1 U12696 ( .A1(n10335), .A2(n10006), .ZN(n10334) );
  AND2_X1 U12697 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  NAND2_X1 U12698 ( .A1(n9932), .A2(n9926), .ZN(P3_U2814) );
  NAND2_X1 U12699 ( .A1(n19079), .A2(n9933), .ZN(n9932) );
  NOR3_X1 U12700 ( .A1(n9931), .A2(n9930), .A3(n9927), .ZN(n9926) );
  INV_X1 U12701 ( .A(n9934), .ZN(n9933) );
  AOI21_X1 U12702 ( .B1(n10284), .B2(n10282), .A(n9831), .ZN(n19264) );
  CLKBUF_X3 U12703 ( .A(n10603), .Z(n18610) );
  INV_X1 U12704 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20821) );
  INV_X2 U12705 ( .A(n10539), .ZN(n18565) );
  INV_X2 U12706 ( .A(n12089), .ZN(n12123) );
  AND4_X1 U12707 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n9751)
         );
  AND2_X2 U12708 ( .A1(n14242), .A2(n14784), .ZN(n12231) );
  NAND2_X1 U12709 ( .A1(n15758), .A2(n15757), .ZN(n15728) );
  AND4_X1 U12710 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n9752) );
  AND2_X1 U12711 ( .A1(n10442), .A2(n10441), .ZN(n9753) );
  AND2_X1 U12712 ( .A1(n11883), .A2(n19296), .ZN(n9754) );
  INV_X1 U12713 ( .A(n10103), .ZN(n15489) );
  AND2_X1 U12714 ( .A1(n12775), .A2(n9826), .ZN(n13458) );
  NAND2_X1 U12715 ( .A1(n10442), .A2(n10126), .ZN(n15322) );
  NAND2_X1 U12716 ( .A1(n10303), .A2(n10306), .ZN(n13263) );
  INV_X1 U12717 ( .A(n10131), .ZN(n16913) );
  AND2_X1 U12718 ( .A1(n12507), .A2(n10421), .ZN(n14410) );
  NAND2_X1 U12719 ( .A1(n12507), .A2(n12506), .ZN(n14408) );
  AND2_X1 U12720 ( .A1(n13006), .A2(n11133), .ZN(n9755) );
  OR2_X1 U12721 ( .A1(n12851), .A2(n12852), .ZN(n12860) );
  OR3_X1 U12722 ( .A1(n15336), .A2(n10278), .A3(n15325), .ZN(n9756) );
  AND2_X1 U12723 ( .A1(n10421), .A2(n17050), .ZN(n9757) );
  INV_X1 U12724 ( .A(n10428), .ZN(n15314) );
  AND2_X1 U12725 ( .A1(n12764), .A2(n9819), .ZN(n9758) );
  INV_X1 U12726 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9901) );
  INV_X1 U12727 ( .A(n16934), .ZN(n10405) );
  OR2_X1 U12728 ( .A1(n12951), .A2(n17214), .ZN(n16934) );
  AND2_X1 U12729 ( .A1(n19382), .A2(n19296), .ZN(n19080) );
  AND2_X1 U12730 ( .A1(n15840), .A2(n10100), .ZN(n9759) );
  NOR3_X1 U12731 ( .A1(n15266), .A2(n15252), .A3(n10262), .ZN(n15226) );
  AND2_X1 U12732 ( .A1(n13255), .A2(n13254), .ZN(n9760) );
  AND2_X1 U12733 ( .A1(n17007), .A2(n17009), .ZN(n13275) );
  NAND2_X1 U12734 ( .A1(n12868), .A2(n9822), .ZN(n9761) );
  INV_X1 U12735 ( .A(n12954), .ZN(n10173) );
  AND2_X1 U12736 ( .A1(n15191), .A2(n20355), .ZN(n9762) );
  AND2_X1 U12737 ( .A1(n10415), .A2(n14128), .ZN(n9763) );
  AND2_X1 U12738 ( .A1(n9760), .A2(n16904), .ZN(n9764) );
  AND2_X1 U12739 ( .A1(n12507), .A2(n9757), .ZN(n14584) );
  NAND2_X1 U12740 ( .A1(n14740), .A2(n10399), .ZN(n16739) );
  INV_X1 U12741 ( .A(n20358), .ZN(n17726) );
  INV_X1 U12742 ( .A(n10861), .ZN(n11086) );
  INV_X1 U12743 ( .A(n14629), .ZN(n9910) );
  AND2_X1 U12744 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9765) );
  AND2_X1 U12745 ( .A1(n9765), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9766) );
  AND2_X1 U12746 ( .A1(n10258), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9767) );
  NAND2_X1 U12747 ( .A1(n10344), .A2(n10343), .ZN(n9768) );
  AND2_X1 U12748 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_2__SCAN_IN), 
        .ZN(n9769) );
  AND2_X1 U12749 ( .A1(n10144), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9770) );
  AND2_X1 U12750 ( .A1(n13451), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9771) );
  AND2_X1 U12751 ( .A1(n10467), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n9772) );
  INV_X1 U12752 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17152) );
  AND2_X2 U12754 ( .A1(n12181), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12240) );
  AND2_X2 U12755 ( .A1(n14241), .A2(n14784), .ZN(n12232) );
  NOR2_X1 U12756 ( .A1(n15322), .A2(n10429), .ZN(n15263) );
  NOR2_X1 U12757 ( .A1(n15108), .A2(n15107), .ZN(n9774) );
  NAND2_X1 U12758 ( .A1(n12826), .A2(n16641), .ZN(n10412) );
  NAND2_X1 U12759 ( .A1(n13773), .A2(n13772), .ZN(n13832) );
  NAND2_X1 U12760 ( .A1(n13950), .A2(n13949), .ZN(n14012) );
  AND2_X1 U12761 ( .A1(n13800), .A2(n13119), .ZN(n13047) );
  INV_X1 U12762 ( .A(n14713), .ZN(n10361) );
  NAND2_X1 U12763 ( .A1(n10442), .A2(n11403), .ZN(n15360) );
  AND2_X1 U12764 ( .A1(n16744), .A2(n10416), .ZN(n13449) );
  XNOR2_X1 U12765 ( .A(n12561), .B(n12560), .ZN(n15183) );
  NOR2_X1 U12766 ( .A1(n16496), .A2(n16497), .ZN(n16481) );
  AND2_X1 U12767 ( .A1(n10442), .A2(n10124), .ZN(n15250) );
  NAND2_X1 U12768 ( .A1(n16744), .A2(n16743), .ZN(n13291) );
  NAND2_X1 U12769 ( .A1(n17027), .A2(n13274), .ZN(n17005) );
  INV_X2 U12770 ( .A(n14691), .ZN(n14287) );
  NOR2_X1 U12771 ( .A1(n18399), .A2(n10147), .ZN(n9775) );
  INV_X1 U12772 ( .A(n9905), .ZN(n12320) );
  AND4_X1 U12773 ( .A1(n10826), .A2(n10825), .A3(n10824), .A4(n10823), .ZN(
        n9776) );
  AND2_X1 U12774 ( .A1(n10055), .A2(n10381), .ZN(n9777) );
  AND4_X1 U12775 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(
        n9778) );
  AND2_X1 U12776 ( .A1(n10523), .A2(n14114), .ZN(n11725) );
  INV_X1 U12777 ( .A(n11725), .ZN(n10539) );
  OR2_X1 U12778 ( .A1(n15223), .A2(n10439), .ZN(n13404) );
  NOR2_X1 U12779 ( .A1(n14329), .A2(n14330), .ZN(n14331) );
  NOR2_X1 U12780 ( .A1(n16496), .A2(n10308), .ZN(n13264) );
  NAND2_X1 U12781 ( .A1(n16744), .A2(n10418), .ZN(n13292) );
  NAND2_X1 U12782 ( .A1(n14331), .A2(n10123), .ZN(n15451) );
  AND2_X1 U12783 ( .A1(n14331), .A2(n14514), .ZN(n14515) );
  AND2_X1 U12784 ( .A1(n13449), .A2(n16530), .ZN(n16521) );
  AND2_X1 U12785 ( .A1(n16956), .A2(n13328), .ZN(n9779) );
  NAND2_X1 U12786 ( .A1(n15723), .A2(n11169), .ZN(n15658) );
  NAND2_X1 U12787 ( .A1(n10020), .A2(n10019), .ZN(n11052) );
  INV_X1 U12788 ( .A(n12123), .ZN(n12991) );
  INV_X1 U12789 ( .A(n10104), .ZN(n11189) );
  AND2_X1 U12790 ( .A1(n15548), .A2(n15549), .ZN(n9780) );
  AND2_X1 U12791 ( .A1(n9897), .A2(n10079), .ZN(n9781) );
  OR2_X1 U12792 ( .A1(n11952), .A2(n11953), .ZN(n9782) );
  AND2_X1 U12793 ( .A1(n13185), .A2(n13353), .ZN(n9783) );
  AND2_X1 U12794 ( .A1(n13832), .A2(n13831), .ZN(n13841) );
  INV_X1 U12795 ( .A(n16920), .ZN(n10193) );
  INV_X1 U12796 ( .A(n13280), .ZN(n10360) );
  AND2_X1 U12797 ( .A1(n15784), .A2(n15794), .ZN(n9784) );
  NAND2_X1 U12798 ( .A1(n12764), .A2(n12763), .ZN(n14501) );
  NAND2_X1 U12799 ( .A1(n12176), .A2(n12174), .ZN(n12218) );
  XNOR2_X1 U12800 ( .A(n13347), .B(n12801), .ZN(n15191) );
  AND2_X1 U12801 ( .A1(n10442), .A2(n10127), .ZN(n15333) );
  NAND2_X2 U12802 ( .A1(n12079), .A2(n12078), .ZN(n21077) );
  AND2_X1 U12803 ( .A1(n10365), .A2(n10363), .ZN(n9785) );
  AND2_X1 U12804 ( .A1(n10170), .A2(n9764), .ZN(n9786) );
  INV_X1 U12805 ( .A(n13403), .ZN(n10438) );
  INV_X1 U12806 ( .A(n10214), .ZN(n15865) );
  NAND2_X1 U12807 ( .A1(n10053), .A2(n10807), .ZN(n10219) );
  NAND2_X1 U12808 ( .A1(n13160), .A2(n16056), .ZN(n15937) );
  INV_X1 U12809 ( .A(n15937), .ZN(n10224) );
  AND2_X1 U12810 ( .A1(n9782), .A2(n11957), .ZN(n9787) );
  AND2_X1 U12811 ( .A1(n11902), .A2(n9936), .ZN(n9788) );
  INV_X1 U12812 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n21728) );
  NOR2_X1 U12813 ( .A1(n18673), .A2(n18802), .ZN(n9789) );
  AND2_X1 U12814 ( .A1(n12862), .A2(n12899), .ZN(n9790) );
  INV_X1 U12815 ( .A(n10190), .ZN(n10189) );
  OAI21_X1 U12816 ( .B1(n12978), .B2(n10191), .A(n10194), .ZN(n10190) );
  NAND2_X1 U12817 ( .A1(n10109), .A2(n9980), .ZN(n9791) );
  INV_X1 U12819 ( .A(n13134), .ZN(n10864) );
  INV_X1 U12820 ( .A(n10430), .ZN(n10429) );
  NOR2_X1 U12821 ( .A1(n15315), .A2(n15323), .ZN(n10430) );
  NAND2_X1 U12822 ( .A1(n10068), .A2(n14012), .ZN(n14498) );
  NOR2_X1 U12823 ( .A1(n15322), .A2(n15323), .ZN(n10428) );
  INV_X1 U12824 ( .A(n14329), .ZN(n10120) );
  AND2_X1 U12825 ( .A1(n10097), .A2(n10096), .ZN(n9792) );
  INV_X1 U12826 ( .A(n12388), .ZN(n12997) );
  INV_X2 U12827 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19926) );
  AND2_X1 U12828 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n9793) );
  NOR2_X1 U12829 ( .A1(n15266), .A2(n15267), .ZN(n10264) );
  NAND2_X1 U12830 ( .A1(n12782), .A2(n12781), .ZN(n16496) );
  AND2_X1 U12831 ( .A1(n14013), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9794) );
  AND4_X1 U12832 ( .A1(n12293), .A2(n12294), .A3(n12305), .A4(n12306), .ZN(
        n9795) );
  NAND2_X1 U12833 ( .A1(n12025), .A2(n12024), .ZN(n12103) );
  OR2_X1 U12834 ( .A1(n12218), .A2(n10027), .ZN(n9796) );
  INV_X1 U12835 ( .A(n10350), .ZN(n10349) );
  NAND2_X1 U12836 ( .A1(n15757), .A2(n10452), .ZN(n10350) );
  INV_X1 U12837 ( .A(n9915), .ZN(n10363) );
  OR2_X1 U12838 ( .A1(n10364), .A2(n16997), .ZN(n9915) );
  NOR2_X2 U12839 ( .A1(n11897), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18909) );
  INV_X1 U12840 ( .A(n18909), .ZN(n10340) );
  NAND2_X1 U12841 ( .A1(n10030), .A2(n10029), .ZN(n16973) );
  INV_X1 U12842 ( .A(n12139), .ZN(n12150) );
  AND3_X1 U12843 ( .A1(n10443), .A2(n15546), .A3(n10119), .ZN(n9797) );
  AND3_X1 U12844 ( .A1(n10900), .A2(n10905), .A3(n10102), .ZN(n9798) );
  AND3_X1 U12845 ( .A1(n12681), .A2(n12680), .A3(n12679), .ZN(n13777) );
  AND3_X1 U12846 ( .A1(n10281), .A2(n9780), .A3(n15458), .ZN(n9799) );
  AND3_X1 U12847 ( .A1(n10085), .A2(n10084), .A3(n12195), .ZN(n9800) );
  AND2_X1 U12848 ( .A1(n12171), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n9801) );
  AND3_X1 U12849 ( .A1(n12172), .A2(n10083), .A3(n9800), .ZN(n9802) );
  AND2_X1 U12850 ( .A1(n14905), .A2(n10382), .ZN(n9803) );
  INV_X1 U12851 ( .A(n18659), .ZN(n19511) );
  OR2_X1 U12852 ( .A1(n10574), .A2(n10573), .ZN(n18659) );
  NOR2_X1 U12853 ( .A1(n15432), .A2(n10044), .ZN(n9804) );
  NOR2_X1 U12854 ( .A1(n16720), .A2(n16719), .ZN(n9805) );
  NAND2_X1 U12855 ( .A1(n9967), .A2(n9966), .ZN(n12345) );
  NOR2_X1 U12856 ( .A1(n17160), .A2(n17161), .ZN(n9807) );
  AND2_X1 U12857 ( .A1(n15812), .A2(n15823), .ZN(n9808) );
  NOR2_X1 U12858 ( .A1(n16919), .A2(n10173), .ZN(n10172) );
  AND2_X1 U12859 ( .A1(n12174), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9809) );
  AND2_X1 U12860 ( .A1(n9779), .A2(n10361), .ZN(n9810) );
  OR2_X1 U12861 ( .A1(n12957), .A2(n12956), .ZN(n9811) );
  NAND2_X1 U12862 ( .A1(n10172), .A2(n16934), .ZN(n9812) );
  INV_X1 U12863 ( .A(n16974), .ZN(n10078) );
  INV_X1 U12864 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20259) );
  OR2_X1 U12865 ( .A1(n15145), .A2(n16895), .ZN(n9813) );
  NAND2_X1 U12866 ( .A1(n13519), .A2(n9741), .ZN(n12802) );
  INV_X1 U12867 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17409) );
  NOR2_X1 U12868 ( .A1(n15532), .A2(n10273), .ZN(n15424) );
  AND2_X1 U12869 ( .A1(n13118), .A2(n13117), .ZN(n15252) );
  INV_X1 U12870 ( .A(n15556), .ZN(n15536) );
  OAI22_X1 U12871 ( .A1(n14561), .A2(n14563), .B1(n12844), .B2(n12620), .ZN(
        n13489) );
  OR3_X1 U12872 ( .A1(n9813), .A2(n10247), .A3(n10246), .ZN(n9814) );
  NAND2_X1 U12873 ( .A1(n13151), .A2(n13031), .ZN(n16064) );
  INV_X1 U12874 ( .A(n16064), .ZN(n21251) );
  NAND2_X1 U12875 ( .A1(n14498), .A2(n14497), .ZN(n14641) );
  NAND2_X1 U12876 ( .A1(n14740), .A2(n16750), .ZN(n16746) );
  INV_X1 U12877 ( .A(n19174), .ZN(n19113) );
  AND2_X1 U12878 ( .A1(n14740), .A2(n10397), .ZN(n16733) );
  NOR2_X1 U12879 ( .A1(n13754), .A2(n10295), .ZN(n9815) );
  NAND2_X1 U12880 ( .A1(n13053), .A2(n13052), .ZN(n14333) );
  AND2_X1 U12881 ( .A1(n18464), .A2(n9772), .ZN(n9816) );
  NAND2_X1 U12882 ( .A1(n15135), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14720) );
  NAND2_X1 U12883 ( .A1(n10248), .A2(n10250), .ZN(n15110) );
  NAND2_X1 U12884 ( .A1(n15125), .A2(n9765), .ZN(n13320) );
  AND2_X1 U12885 ( .A1(n18601), .A2(n10144), .ZN(n9817) );
  OR2_X1 U12886 ( .A1(n13821), .A2(n19420), .ZN(n10002) );
  AND2_X1 U12887 ( .A1(n11153), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9818) );
  AND2_X1 U12888 ( .A1(n12763), .A2(n10300), .ZN(n9819) );
  NAND2_X1 U12889 ( .A1(n14839), .A2(n14838), .ZN(n9820) );
  NOR2_X1 U12890 ( .A1(n9813), .A2(n16889), .ZN(n15149) );
  NOR2_X1 U12891 ( .A1(n15532), .A2(n15533), .ZN(n15526) );
  NOR2_X1 U12892 ( .A1(n15118), .A2(n20202), .ZN(n15119) );
  NAND2_X1 U12893 ( .A1(n9907), .A2(n12496), .ZN(n13486) );
  NOR2_X1 U12894 ( .A1(n13858), .A2(n10312), .ZN(n14001) );
  AND2_X1 U12895 ( .A1(n15378), .A2(n15379), .ZN(n15362) );
  NAND2_X1 U12896 ( .A1(n10903), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11364) );
  OR2_X1 U12897 ( .A1(n11882), .A2(n9982), .ZN(n19154) );
  BUF_X1 U12898 ( .A(n10861), .Z(n14090) );
  AND2_X1 U12899 ( .A1(n10069), .A2(n16735), .ZN(n9821) );
  AND2_X1 U12900 ( .A1(n10377), .A2(n10376), .ZN(n9822) );
  AND2_X1 U12901 ( .A1(n13875), .A2(n13876), .ZN(n13874) );
  NAND2_X1 U12902 ( .A1(n21077), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n21074) );
  INV_X1 U12903 ( .A(n21074), .ZN(n9888) );
  INV_X1 U12904 ( .A(n12948), .ZN(n10379) );
  OR2_X1 U12905 ( .A1(n19217), .A2(n18769), .ZN(n19178) );
  AND2_X1 U12906 ( .A1(n16620), .A2(n13492), .ZN(n9823) );
  AND2_X1 U12907 ( .A1(n15123), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15125) );
  AND2_X1 U12908 ( .A1(n14839), .A2(n9821), .ZN(n9824) );
  AND2_X1 U12909 ( .A1(n15394), .A2(n13087), .ZN(n15378) );
  AND2_X1 U12910 ( .A1(n12985), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n9825) );
  INV_X1 U12911 ( .A(n11043), .ZN(n10232) );
  INV_X1 U12912 ( .A(n12819), .ZN(n9918) );
  AND2_X1 U12913 ( .A1(n12774), .A2(n10302), .ZN(n9826) );
  OR2_X1 U12914 ( .A1(n14645), .A2(n14644), .ZN(n14647) );
  INV_X1 U12915 ( .A(n14647), .ZN(n9911) );
  AND2_X1 U12916 ( .A1(n10383), .A2(n10382), .ZN(n9827) );
  AND2_X1 U12917 ( .A1(n10423), .A2(n10422), .ZN(n9828) );
  AND2_X1 U12918 ( .A1(n9819), .A2(n13333), .ZN(n9829) );
  INV_X1 U12919 ( .A(n19296), .ZN(n19055) );
  AND2_X1 U12920 ( .A1(n19329), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19296) );
  AND2_X1 U12921 ( .A1(n10393), .A2(n10396), .ZN(n9830) );
  OR2_X1 U12922 ( .A1(n12284), .A2(n12283), .ZN(n12395) );
  AND2_X1 U12923 ( .A1(n19468), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9831) );
  AND2_X1 U12924 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9832) );
  AND2_X1 U12925 ( .A1(n21654), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9833) );
  INV_X1 U12927 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15114) );
  INV_X1 U12928 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13323) );
  INV_X1 U12929 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20137) );
  NAND2_X1 U12930 ( .A1(n12491), .A2(n12490), .ZN(n14014) );
  INV_X1 U12931 ( .A(n14014), .ZN(n9907) );
  INV_X1 U12932 ( .A(n10111), .ZN(n10110) );
  NAND2_X1 U12933 ( .A1(n19113), .A2(n19235), .ZN(n10111) );
  INV_X1 U12934 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17089) );
  AND2_X1 U12935 ( .A1(n11885), .A2(n9978), .ZN(n9834) );
  AND2_X1 U12936 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12464), .ZN(n20929) );
  NOR2_X1 U12937 ( .A1(n17850), .A2(n20090), .ZN(n9835) );
  OR2_X1 U12938 ( .A1(n14709), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9836) );
  AND2_X1 U12939 ( .A1(n10393), .A2(n14874), .ZN(n9837) );
  AND2_X1 U12940 ( .A1(n12264), .A2(n12395), .ZN(n9838) );
  NAND2_X1 U12941 ( .A1(n9907), .A2(n9763), .ZN(n14127) );
  INV_X1 U12942 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19755) );
  AND2_X1 U12943 ( .A1(n14691), .A2(n15557), .ZN(n11146) );
  AND2_X1 U12944 ( .A1(n11225), .A2(n11224), .ZN(n14330) );
  AND2_X1 U12945 ( .A1(n10281), .A2(n9780), .ZN(n9839) );
  OR2_X1 U12946 ( .A1(n15532), .A2(n10271), .ZN(n9840) );
  AND2_X1 U12947 ( .A1(n9766), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9841) );
  AND2_X1 U12948 ( .A1(n9822), .A2(n16544), .ZN(n9842) );
  INV_X1 U12949 ( .A(n16914), .ZN(n10242) );
  AND2_X1 U12950 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9843) );
  INV_X2 U12951 ( .A(n18410), .ZN(n18613) );
  AND2_X1 U12952 ( .A1(n12985), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n9844) );
  INV_X1 U12953 ( .A(n20251), .ZN(n20269) );
  INV_X1 U12954 ( .A(n13767), .ZN(n16674) );
  INV_X1 U12955 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17732) );
  NAND2_X1 U12956 ( .A1(n12998), .A2(n21053), .ZN(n20360) );
  INV_X1 U12957 ( .A(n20360), .ZN(n17383) );
  OR2_X1 U12958 ( .A1(n20086), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n9845) );
  NAND3_X1 U12959 ( .A1(n12735), .A2(n12734), .A3(n12733), .ZN(n9846) );
  AND2_X1 U12960 ( .A1(n17991), .A2(n18132), .ZN(n9847) );
  INV_X1 U12961 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10695) );
  AND2_X1 U12962 ( .A1(n11292), .A2(n11291), .ZN(n9848) );
  NOR2_X1 U12963 ( .A1(n14698), .A2(n13032), .ZN(n9849) );
  NOR2_X1 U12964 ( .A1(n17457), .A2(n11947), .ZN(n9850) );
  INV_X1 U12965 ( .A(n9870), .ZN(n20198) );
  OR2_X1 U12966 ( .A1(n20196), .A2(n10462), .ZN(n9870) );
  INV_X1 U12967 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19380) );
  INV_X1 U12968 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16926) );
  AND2_X1 U12969 ( .A1(n13231), .A2(n20087), .ZN(n19470) );
  INV_X1 U12970 ( .A(n19470), .ZN(n19459) );
  NOR2_X1 U12971 ( .A1(n18644), .A2(n18636), .ZN(n9851) );
  INV_X1 U12972 ( .A(n16897), .ZN(n10241) );
  INV_X1 U12973 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21654) );
  INV_X1 U12974 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16889) );
  AND2_X1 U12975 ( .A1(n19389), .A2(n19142), .ZN(n9852) );
  AND2_X1 U12976 ( .A1(n13502), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17525) );
  INV_X1 U12977 ( .A(n17525), .ZN(n10325) );
  INV_X1 U12978 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10181) );
  INV_X1 U12979 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9983) );
  NOR2_X1 U12980 ( .A1(n10482), .A2(n10204), .ZN(n13505) );
  OR2_X1 U12981 ( .A1(n10482), .A2(n10206), .ZN(n9853) );
  NOR2_X1 U12982 ( .A1(n10482), .A2(n10483), .ZN(n18982) );
  OR2_X1 U12983 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11168), .ZN(
        n9854) );
  AND3_X1 U12984 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17461) );
  INV_X1 U12985 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14111) );
  OR2_X1 U12986 ( .A1(n21028), .A2(n20855), .ZN(n9855) );
  INV_X1 U12987 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17460) );
  OR2_X1 U12988 ( .A1(n9854), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9856) );
  AND2_X1 U12989 ( .A1(n9771), .A2(n10133), .ZN(n9857) );
  INV_X1 U12990 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n18050) );
  INV_X1 U12991 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10345) );
  INV_X1 U12992 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15098) );
  INV_X1 U12993 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10371) );
  INV_X1 U12994 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10375) );
  INV_X1 U12995 ( .A(n18636), .ZN(n10138) );
  INV_X1 U12996 ( .A(n15871), .ZN(n10100) );
  INV_X1 U12997 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10333) );
  INV_X1 U12998 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10142) );
  INV_X1 U12999 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10343) );
  AND3_X1 U13000 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), 
        .A3(P3_EAX_REG_27__SCAN_IN), .ZN(n9858) );
  AND2_X1 U13001 ( .A1(n17153), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9859) );
  AND2_X1 U13002 ( .A1(n10368), .A2(n17153), .ZN(n9860) );
  AND2_X1 U13003 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9861) );
  INV_X1 U13004 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16952) );
  INV_X1 U13005 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13924) );
  INV_X1 U13006 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n20070) );
  AOI22_X2 U13007 ( .A1(DATAI_22_), .A2(n9715), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n9716), .ZN(n16418) );
  AOI22_X2 U13008 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9716), .B1(DATAI_17_), 
        .B2(n9715), .ZN(n16395) );
  AOI22_X2 U13009 ( .A1(DATAI_19_), .A2(n9715), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n9716), .ZN(n16403) );
  AOI22_X2 U13010 ( .A1(DATAI_20_), .A2(n9715), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n9716), .ZN(n16408) );
  AOI22_X2 U13011 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9716), .B1(DATAI_23_), 
        .B2(n9715), .ZN(n16426) );
  AOI22_X2 U13012 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9716), .B1(DATAI_21_), 
        .B2(n9715), .ZN(n16413) );
  NOR3_X2 U13013 ( .A1(n19978), .A2(n19755), .A3(n19610), .ZN(n19583) );
  NOR3_X2 U13014 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19978), .A3(
        n19707), .ZN(n19674) );
  AOI22_X2 U13015 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9716), .B1(DATAI_18_), 
        .B2(n9715), .ZN(n21758) );
  NOR2_X2 U13016 ( .A1(n20132), .A2(n16556), .ZN(n16546) );
  NAND2_X1 U13019 ( .A1(n9872), .A2(n12177), .ZN(n12213) );
  AND2_X2 U13020 ( .A1(n9872), .A2(n12175), .ZN(n20446) );
  AND2_X2 U13021 ( .A1(n9872), .A2(n12171), .ZN(n12297) );
  NAND2_X1 U13022 ( .A1(n9872), .A2(n12174), .ZN(n12289) );
  NAND2_X1 U13023 ( .A1(n9809), .A2(n9872), .ZN(n10085) );
  AND2_X2 U13024 ( .A1(n12170), .A2(n13661), .ZN(n9872) );
  NAND3_X1 U13025 ( .A1(n20400), .A2(n13751), .A3(n9873), .ZN(n12109) );
  NAND2_X2 U13026 ( .A1(n12036), .A2(n12037), .ZN(n12089) );
  NAND3_X1 U13027 ( .A1(n12109), .A2(n12609), .A3(n12125), .ZN(n12127) );
  OAI21_X2 U13028 ( .B1(n16935), .B2(n10405), .A(n10402), .ZN(n16929) );
  AND2_X2 U13029 ( .A1(n9875), .A2(n10010), .ZN(n16935) );
  NAND4_X1 U13030 ( .A1(n10071), .A2(n10070), .A3(n9717), .A4(n12946), .ZN(
        n9875) );
  NAND3_X1 U13031 ( .A1(n12158), .A2(n9876), .A3(n9893), .ZN(n9894) );
  NAND2_X1 U13032 ( .A1(n9892), .A2(n9877), .ZN(n9876) );
  OR2_X2 U13033 ( .A1(n12159), .A2(n12160), .ZN(n9892) );
  NAND2_X1 U13034 ( .A1(n12163), .A2(n12162), .ZN(n12161) );
  NAND2_X1 U13035 ( .A1(n9880), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U13036 ( .A1(n9880), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9902) );
  AOI21_X1 U13037 ( .B1(n9880), .B2(n20821), .A(n9855), .ZN(n20822) );
  OAI21_X1 U13038 ( .B1(n9880), .B2(n20855), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20825) );
  NAND2_X1 U13039 ( .A1(n9880), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n9878) );
  AOI22_X1 U13040 ( .A1(n20635), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9880), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12327) );
  AOI21_X1 U13041 ( .B1(n13399), .B2(n17383), .A(n9762), .ZN(n12999) );
  NAND3_X1 U13042 ( .A1(n12067), .A2(n12066), .A3(n9888), .ZN(n9887) );
  NAND2_X1 U13043 ( .A1(n12067), .A2(n12066), .ZN(n9889) );
  NAND2_X1 U13044 ( .A1(n12094), .A2(n9887), .ZN(n12121) );
  NAND2_X1 U13045 ( .A1(n12563), .A2(n9889), .ZN(n14258) );
  INV_X1 U13046 ( .A(n9947), .ZN(n16884) );
  OR2_X2 U13047 ( .A1(n16935), .A2(n9812), .ZN(n10169) );
  NAND3_X1 U13048 ( .A1(n9896), .A2(n12286), .A3(n12270), .ZN(n17130) );
  NAND2_X1 U13049 ( .A1(n10157), .A2(n10158), .ZN(n9896) );
  OAI21_X1 U13050 ( .B1(n12289), .B2(n12196), .A(n9898), .ZN(n12201) );
  OR2_X2 U13051 ( .A1(n17026), .A2(n17277), .ZN(n9899) );
  AND2_X4 U13052 ( .A1(n14241), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14788) );
  OAI21_X1 U13053 ( .B1(n12343), .B2(n9806), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10315) );
  INV_X1 U13054 ( .A(n12319), .ZN(n9967) );
  NAND2_X1 U13055 ( .A1(n12319), .A2(n17368), .ZN(n17362) );
  NAND2_X1 U13056 ( .A1(n9903), .A2(n9902), .ZN(n12205) );
  AND2_X2 U13057 ( .A1(n16661), .A2(n13952), .ZN(n12178) );
  AND2_X2 U13058 ( .A1(n9906), .A2(n12177), .ZN(n20599) );
  AND2_X2 U13059 ( .A1(n12170), .A2(n16661), .ZN(n9906) );
  NAND3_X1 U13060 ( .A1(n13391), .A2(n13389), .A3(n13390), .ZN(P2_U3017) );
  AND2_X2 U13061 ( .A1(n17057), .A2(n9857), .ZN(n13252) );
  AND2_X2 U13062 ( .A1(n9906), .A2(n12175), .ZN(n12296) );
  AND2_X2 U13063 ( .A1(n9906), .A2(n12174), .ZN(n12291) );
  NAND2_X1 U13064 ( .A1(n9906), .A2(n12171), .ZN(n9905) );
  NAND2_X1 U13065 ( .A1(n9801), .A2(n9906), .ZN(n10084) );
  AND2_X2 U13066 ( .A1(n13252), .A2(n9859), .ZN(n16870) );
  INV_X1 U13067 ( .A(n12840), .ZN(n9917) );
  AND2_X4 U13068 ( .A1(n14952), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14802) );
  AOI22_X1 U13069 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U13070 ( .A1(n9923), .A2(n11071), .ZN(n10983) );
  NAND2_X1 U13071 ( .A1(n9923), .A2(n11069), .ZN(n10940) );
  XNOR2_X1 U13072 ( .A(n11070), .B(n9923), .ZN(n10106) );
  NAND2_X2 U13073 ( .A1(n10893), .A2(n10892), .ZN(n9923) );
  NOR2_X1 U13074 ( .A1(n9925), .A2(n16290), .ZN(n13735) );
  NAND2_X1 U13075 ( .A1(n10228), .A2(n9925), .ZN(n16291) );
  XNOR2_X1 U13076 ( .A(n9925), .B(n14152), .ZN(n14028) );
  NAND2_X2 U13077 ( .A1(n10995), .A2(n10996), .ZN(n9925) );
  NOR2_X2 U13078 ( .A1(n11904), .A2(n9788), .ZN(n13919) );
  NAND3_X1 U13079 ( .A1(n10426), .A2(n13417), .A3(n10898), .ZN(n13027) );
  AND2_X1 U13080 ( .A1(n10426), .A2(n10898), .ZN(n14979) );
  NAND2_X2 U13081 ( .A1(n9938), .A2(n11167), .ZN(n15758) );
  NAND3_X1 U13082 ( .A1(n15765), .A2(n15769), .A3(n10167), .ZN(n9939) );
  NOR2_X4 U13083 ( .A1(n19440), .A2(n20089), .ZN(n19948) );
  NOR2_X4 U13084 ( .A1(n19390), .A2(n19949), .ZN(n19346) );
  NAND4_X1 U13085 ( .A1(n10648), .A2(n10644), .A3(n19508), .A4(n19503), .ZN(
        n10654) );
  AND2_X2 U13086 ( .A1(n11148), .A2(n11147), .ZN(n15664) );
  NAND4_X1 U13087 ( .A1(n10348), .A2(n11054), .A3(n10231), .A4(n10116), .ZN(
        n11148) );
  NAND2_X2 U13088 ( .A1(n17130), .A2(n12272), .ZN(n17113) );
  NAND3_X1 U13089 ( .A1(n9960), .A2(n9959), .A3(n9958), .ZN(P2_U2987) );
  OR2_X1 U13090 ( .A1(n17163), .A2(n17136), .ZN(n9958) );
  NAND2_X1 U13091 ( .A1(n17162), .A2(n17718), .ZN(n9960) );
  INV_X1 U13092 ( .A(n16870), .ZN(n9962) );
  NAND3_X1 U13093 ( .A1(n14219), .A2(n12465), .A3(n12417), .ZN(n9963) );
  NAND4_X1 U13094 ( .A1(n14314), .A2(n21078), .A3(n12465), .A4(n12418), .ZN(
        n9965) );
  NAND2_X1 U13095 ( .A1(n17057), .A2(n9771), .ZN(n13447) );
  NAND2_X1 U13096 ( .A1(n17057), .A2(n10155), .ZN(n16976) );
  NAND2_X1 U13097 ( .A1(n17057), .A2(n13451), .ZN(n13289) );
  AND2_X1 U13098 ( .A1(n17057), .A2(n10156), .ZN(n16994) );
  NAND2_X1 U13099 ( .A1(n17057), .A2(n10132), .ZN(n10131) );
  NAND2_X4 U13100 ( .A1(n10080), .A2(n12377), .ZN(n17057) );
  NAND2_X1 U13101 ( .A1(n9969), .A2(n11859), .ZN(n17464) );
  NAND2_X1 U13102 ( .A1(n13885), .A2(n13884), .ZN(n9969) );
  NAND2_X1 U13103 ( .A1(n11859), .A2(n9972), .ZN(n9971) );
  INV_X1 U13104 ( .A(n13884), .ZN(n9972) );
  INV_X1 U13105 ( .A(n11859), .ZN(n9973) );
  XNOR2_X1 U13106 ( .A(n11858), .B(n11856), .ZN(n13885) );
  NAND2_X1 U13107 ( .A1(n18909), .A2(n9975), .ZN(n9974) );
  NAND2_X1 U13108 ( .A1(n17423), .A2(n17426), .ZN(n9976) );
  XNOR2_X2 U13109 ( .A(n9976), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17491) );
  NAND3_X1 U13110 ( .A1(n9977), .A2(n10180), .A3(n10178), .ZN(n9978) );
  NAND3_X1 U13111 ( .A1(n19414), .A2(n9754), .A3(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9977) );
  NAND3_X1 U13112 ( .A1(n11885), .A2(n19310), .A3(n9978), .ZN(n11884) );
  NAND2_X1 U13113 ( .A1(n11881), .A2(n10455), .ZN(n10326) );
  AND2_X2 U13114 ( .A1(n11896), .A2(n17504), .ZN(n11897) );
  NAND2_X1 U13115 ( .A1(n10109), .A2(n9979), .ZN(n17504) );
  NOR2_X2 U13116 ( .A1(n18943), .A2(n9981), .ZN(n9979) );
  NAND2_X1 U13117 ( .A1(n10111), .A2(n17516), .ZN(n9981) );
  NAND3_X1 U13118 ( .A1(n10013), .A2(n12994), .A3(n12347), .ZN(n9985) );
  NAND3_X1 U13119 ( .A1(n9989), .A2(n11114), .A3(n14423), .ZN(n10159) );
  NAND3_X1 U13120 ( .A1(n11107), .A2(n11108), .A3(n11109), .ZN(n9989) );
  XNOR2_X1 U13121 ( .A(n11091), .B(n13788), .ZN(n13852) );
  NAND2_X1 U13122 ( .A1(n11090), .A2(n11089), .ZN(n11091) );
  NAND2_X1 U13123 ( .A1(n11169), .A2(n15729), .ZN(n15695) );
  NAND3_X1 U13124 ( .A1(n15723), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11169), .ZN(n9992) );
  NAND3_X1 U13125 ( .A1(n15674), .A2(n10100), .A3(n15695), .ZN(n9993) );
  INV_X1 U13126 ( .A(n10098), .ZN(n9998) );
  AOI21_X2 U13127 ( .B1(n10098), .B2(n10000), .A(n9818), .ZN(n9995) );
  NOR2_X1 U13128 ( .A1(n10000), .A2(n9818), .ZN(n9999) );
  NAND2_X1 U13129 ( .A1(n10001), .A2(n17363), .ZN(n12341) );
  XNOR2_X1 U13130 ( .A(n11952), .B(n11953), .ZN(n13821) );
  XNOR2_X2 U13131 ( .A(n11945), .B(n11946), .ZN(n17458) );
  OR2_X1 U13132 ( .A1(n19095), .A2(n19055), .ZN(n19339) );
  INV_X1 U13133 ( .A(n19339), .ZN(n19082) );
  NAND3_X1 U13134 ( .A1(n10009), .A2(n10175), .A3(n10317), .ZN(n12286) );
  NAND4_X1 U13135 ( .A1(n12224), .A2(n12226), .A3(n12227), .A4(n12225), .ZN(
        n10009) );
  NAND2_X1 U13136 ( .A1(n10009), .A2(n12264), .ZN(n10157) );
  NAND3_X1 U13137 ( .A1(n10071), .A2(n9717), .A3(n10070), .ZN(n17027) );
  INV_X1 U13138 ( .A(n12946), .ZN(n10011) );
  AND2_X2 U13139 ( .A1(n17522), .A2(n19174), .ZN(n18943) );
  AOI21_X1 U13140 ( .B1(n10870), .B2(n14045), .A(n10869), .ZN(n10871) );
  NAND2_X1 U13141 ( .A1(n10315), .A2(n12346), .ZN(n17083) );
  NOR3_X2 U13142 ( .A1(n18954), .A2(n18957), .A3(n19235), .ZN(n18941) );
  NOR2_X2 U13143 ( .A1(n17515), .A2(n17476), .ZN(n17739) );
  NAND2_X1 U13144 ( .A1(n12135), .A2(n12134), .ZN(n12159) );
  AOI22_X2 U13145 ( .A1(n11113), .A2(n11112), .B1(n11111), .B2(n11110), .ZN(
        n11114) );
  NAND2_X1 U13146 ( .A1(n15696), .A2(n15661), .ZN(n10034) );
  AND2_X1 U13147 ( .A1(n13028), .A2(n10885), .ZN(n10886) );
  NAND2_X1 U13148 ( .A1(n10013), .A2(n12347), .ZN(n12319) );
  INV_X1 U13149 ( .A(n13144), .ZN(n10015) );
  NOR2_X1 U13150 ( .A1(n10882), .A2(n10014), .ZN(n13028) );
  NAND2_X1 U13151 ( .A1(n10015), .A2(n10883), .ZN(n10014) );
  NAND2_X1 U13152 ( .A1(n10016), .A2(n11158), .ZN(n15782) );
  AOI21_X1 U13153 ( .B1(n15803), .B2(n10016), .A(n15802), .ZN(n15805) );
  NAND2_X1 U13154 ( .A1(n11052), .A2(n10994), .ZN(n11178) );
  NAND2_X1 U13155 ( .A1(n14337), .A2(n10941), .ZN(n14436) );
  INV_X1 U13156 ( .A(n10993), .ZN(n10020) );
  NAND4_X1 U13157 ( .A1(n12169), .A2(n9796), .A3(n10023), .A4(n10022), .ZN(
        n10021) );
  NAND2_X1 U13158 ( .A1(n14601), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U13159 ( .A1(n12296), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10023) );
  NAND3_X1 U13160 ( .A1(n10025), .A2(n10028), .A3(n10026), .ZN(n10024) );
  NAND2_X1 U13161 ( .A1(n20709), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10028) );
  NAND3_X1 U13162 ( .A1(n10033), .A2(n10035), .A3(n10168), .ZN(n13191) );
  NAND2_X1 U13163 ( .A1(n10038), .A2(n13003), .ZN(n10039) );
  INV_X1 U13164 ( .A(n10781), .ZN(n10038) );
  NAND3_X1 U13165 ( .A1(n10041), .A2(n10780), .A3(n10039), .ZN(n10782) );
  NAND2_X1 U13166 ( .A1(n10776), .A2(n10805), .ZN(n10041) );
  AND2_X1 U13167 ( .A1(n14051), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10042) );
  OR2_X1 U13168 ( .A1(n15432), .A2(n10045), .ZN(n15357) );
  NAND3_X1 U13169 ( .A1(n10046), .A2(P1_REIP_REG_15__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .ZN(n10044) );
  NAND4_X1 U13170 ( .A1(n10046), .A2(P1_REIP_REG_15__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_17__SCAN_IN), .ZN(n10045) );
  OR2_X1 U13171 ( .A1(n15432), .A2(n14693), .ZN(n15401) );
  INV_X2 U13172 ( .A(n10219), .ZN(n17587) );
  NAND3_X1 U13173 ( .A1(n10804), .A2(n10220), .A3(n10803), .ZN(n10053) );
  NAND2_X1 U13174 ( .A1(n14920), .A2(n10383), .ZN(n10055) );
  NAND3_X1 U13175 ( .A1(n10059), .A2(n10058), .A3(n10062), .ZN(n16706) );
  NAND2_X1 U13176 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  NOR2_X1 U13177 ( .A1(n16725), .A2(n14874), .ZN(n10060) );
  NAND2_X1 U13178 ( .A1(n16725), .A2(n9837), .ZN(n10062) );
  NAND3_X1 U13179 ( .A1(n13950), .A2(n10066), .A3(n13949), .ZN(n10064) );
  NAND2_X1 U13180 ( .A1(n10075), .A2(n10073), .ZN(n13327) );
  NOR2_X1 U13181 ( .A1(n10074), .A2(n10360), .ZN(n10073) );
  NAND2_X1 U13182 ( .A1(n16973), .A2(n10076), .ZN(n10075) );
  NOR2_X1 U13183 ( .A1(n14713), .A2(n10077), .ZN(n10076) );
  NAND3_X1 U13184 ( .A1(n10082), .A2(n9807), .A3(n10081), .ZN(P2_U3019) );
  OR2_X1 U13185 ( .A1(n17163), .A2(n20360), .ZN(n10081) );
  NAND2_X1 U13186 ( .A1(n12297), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10083) );
  INV_X1 U13187 ( .A(n10176), .ZN(n10086) );
  NAND2_X1 U13188 ( .A1(n18677), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n18673) );
  INV_X1 U13189 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n10088) );
  NAND3_X1 U13190 ( .A1(n9751), .A2(P3_EAX_REG_21__SCAN_IN), .A3(
        P3_EAX_REG_20__SCAN_IN), .ZN(n10089) );
  AND2_X1 U13191 ( .A1(n18856), .A2(n20089), .ZN(n10091) );
  INV_X1 U13192 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10093) );
  AND2_X4 U13193 ( .A1(n14045), .A2(n14691), .ZN(n13119) );
  NAND2_X1 U13194 ( .A1(n10094), .A2(n13470), .ZN(P1_U2968) );
  NAND2_X1 U13195 ( .A1(n13469), .A2(n17668), .ZN(n10094) );
  NAND2_X1 U13196 ( .A1(n13193), .A2(n13194), .ZN(n10095) );
  NAND2_X1 U13197 ( .A1(n15650), .A2(n10454), .ZN(n13192) );
  NAND3_X1 U13198 ( .A1(n13137), .A2(n9798), .A3(n10101), .ZN(n11069) );
  AND2_X1 U13199 ( .A1(n10901), .A2(n13139), .ZN(n10102) );
  CLKBUF_X1 U13200 ( .A(n10106), .Z(n10103) );
  NAND2_X1 U13201 ( .A1(n10106), .A2(n21654), .ZN(n11072) );
  NAND2_X1 U13202 ( .A1(n10103), .A2(n16076), .ZN(n16077) );
  OAI21_X1 U13203 ( .B1(n15489), .B2(n11364), .A(n10105), .ZN(n10104) );
  INV_X1 U13204 ( .A(n11188), .ZN(n10105) );
  AOI21_X1 U13205 ( .B1(n16097), .B2(n10103), .A(n15089), .ZN(n17590) );
  AND2_X2 U13206 ( .A1(n13952), .A2(n13661), .ZN(n12176) );
  NOR2_X2 U13207 ( .A1(n19926), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10523) );
  NAND3_X1 U13208 ( .A1(n10115), .A2(n10113), .A3(n17525), .ZN(n11892) );
  NAND3_X1 U13209 ( .A1(n10116), .A2(n11054), .A3(n11094), .ZN(n11059) );
  INV_X1 U13210 ( .A(n14330), .ZN(n10118) );
  NAND4_X1 U13211 ( .A1(n10118), .A2(n10121), .A3(n15546), .A4(n10443), .ZN(
        n10117) );
  NAND3_X1 U13212 ( .A1(n10120), .A2(n9797), .A3(n10118), .ZN(n10122) );
  INV_X1 U13213 ( .A(n10122), .ZN(n15531) );
  XNOR2_X2 U13214 ( .A(n13404), .B(n10438), .ZN(n15200) );
  XNOR2_X2 U13215 ( .A(n12376), .B(n12994), .ZN(n12371) );
  NAND2_X2 U13216 ( .A1(n10130), .A2(n12348), .ZN(n12376) );
  NAND2_X1 U13217 ( .A1(n10317), .A2(n10318), .ZN(n10158) );
  NAND2_X2 U13218 ( .A1(n10159), .A2(n11131), .ZN(n17653) );
  NAND3_X1 U13219 ( .A1(n10162), .A2(n10165), .A3(n10161), .ZN(n14029) );
  NAND2_X1 U13220 ( .A1(n10890), .A2(n10164), .ZN(n10161) );
  INV_X1 U13221 ( .A(n10890), .ZN(n10163) );
  NAND2_X1 U13222 ( .A1(n10907), .A2(n10889), .ZN(n10165) );
  XNOR2_X2 U13223 ( .A(n11097), .B(n11054), .ZN(n14024) );
  NAND2_X1 U13224 ( .A1(n10195), .A2(n12317), .ZN(n10176) );
  NAND2_X1 U13225 ( .A1(n17504), .A2(n10177), .ZN(n18910) );
  NOR2_X2 U13226 ( .A1(n18910), .A2(n19174), .ZN(n17575) );
  NAND2_X1 U13227 ( .A1(n19174), .A2(n10181), .ZN(n10180) );
  NAND2_X1 U13228 ( .A1(n16929), .A2(n10184), .ZN(n10183) );
  AND2_X1 U13229 ( .A1(n12292), .A2(n12295), .ZN(n10196) );
  NAND4_X1 U13230 ( .A1(n10196), .A2(n9795), .A3(n12304), .A4(n12303), .ZN(
        n10195) );
  NAND2_X1 U13231 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17459) );
  NAND2_X1 U13232 ( .A1(n9730), .A2(n10198), .ZN(n17446) );
  AND2_X1 U13233 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10198) );
  AND2_X1 U13234 ( .A1(n10209), .A2(n10208), .ZN(n18010) );
  INV_X1 U13235 ( .A(n10215), .ZN(n15883) );
  OR2_X1 U13236 ( .A1(n16030), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10213) );
  OAI21_X1 U13237 ( .B1(n13203), .B2(n10100), .A(n10215), .ZN(n10214) );
  NAND2_X1 U13238 ( .A1(n15937), .A2(n10221), .ZN(n15901) );
  NAND3_X1 U13239 ( .A1(n15812), .A2(n15823), .A3(n11163), .ZN(n15780) );
  NAND2_X1 U13240 ( .A1(n15838), .A2(n9808), .ZN(n15803) );
  OAI21_X2 U13241 ( .B1(n15758), .B2(n9854), .A(n15840), .ZN(n15723) );
  NAND4_X1 U13242 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10233), .A3(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15103) );
  AOI21_X1 U13243 ( .B1(n10256), .B2(n20269), .A(n10254), .ZN(n10253) );
  XNOR2_X1 U13244 ( .A(n11931), .B(n19465), .ZN(n19212) );
  XNOR2_X2 U13245 ( .A(n11933), .B(n11930), .ZN(n11931) );
  NAND2_X2 U13246 ( .A1(n14007), .A2(n13998), .ZN(n11933) );
  OR2_X2 U13247 ( .A1(n11849), .A2(n11848), .ZN(n14007) );
  INV_X1 U13248 ( .A(n10264), .ZN(n10469) );
  NOR2_X2 U13249 ( .A1(n11941), .A2(n11942), .ZN(n11945) );
  NOR2_X2 U13250 ( .A1(n15532), .A2(n10268), .ZN(n15394) );
  INV_X2 U13251 ( .A(n10540), .ZN(n11825) );
  NOR2_X2 U13252 ( .A1(n19172), .A2(n11961), .ZN(n19095) );
  NOR2_X1 U13253 ( .A1(n15336), .A2(n15325), .ZN(n15324) );
  INV_X1 U13254 ( .A(n15313), .ZN(n10278) );
  INV_X1 U13255 ( .A(n10279), .ZN(n15289) );
  NAND2_X1 U13256 ( .A1(n9799), .A2(n13053), .ZN(n15456) );
  NAND3_X1 U13257 ( .A1(n19271), .A2(n19272), .A3(n10285), .ZN(n10284) );
  NOR2_X2 U13258 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10291) );
  AND2_X4 U13259 ( .A1(n10291), .A2(n14248), .ZN(n12181) );
  NOR2_X1 U13260 ( .A1(n14229), .A2(n10291), .ZN(n14230) );
  NAND2_X1 U13261 ( .A1(n14191), .A2(n10292), .ZN(n14565) );
  NAND2_X2 U13262 ( .A1(n14189), .A2(n14188), .ZN(n14191) );
  OR2_X2 U13263 ( .A1(n13754), .A2(n10293), .ZN(n13857) );
  NAND2_X1 U13264 ( .A1(n13382), .A2(n13383), .ZN(n16772) );
  INV_X1 U13265 ( .A(n13332), .ZN(n12771) );
  NOR2_X2 U13266 ( .A1(n16496), .A2(n10304), .ZN(n16444) );
  NAND2_X1 U13267 ( .A1(n12722), .A2(n10310), .ZN(n14278) );
  NAND2_X1 U13268 ( .A1(n12722), .A2(n12721), .ZN(n13895) );
  NAND2_X1 U13269 ( .A1(n17083), .A2(n17084), .ZN(n12374) );
  NAND3_X1 U13270 ( .A1(n9802), .A2(n10319), .A3(n10320), .ZN(n10317) );
  NAND2_X1 U13271 ( .A1(n16994), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17239) );
  NAND2_X1 U13272 ( .A1(n10321), .A2(n13307), .ZN(n13290) );
  NAND2_X1 U13273 ( .A1(n12562), .A2(n9843), .ZN(n12144) );
  AND2_X2 U13274 ( .A1(n12562), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U13275 ( .A1(n11885), .A2(n10182), .ZN(n19056) );
  NAND2_X1 U13276 ( .A1(n13810), .A2(n10330), .ZN(n10329) );
  NAND2_X2 U13277 ( .A1(n14114), .A2(n14667), .ZN(n18261) );
  INV_X1 U13278 ( .A(n19154), .ZN(n10342) );
  AND2_X2 U13279 ( .A1(n10346), .A2(n10425), .ZN(n10968) );
  MUX2_X1 U13280 ( .A(n10346), .B(n10695), .S(n16091), .Z(n15000) );
  INV_X1 U13281 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10347) );
  NAND2_X2 U13282 ( .A1(n10939), .A2(n10938), .ZN(n11054) );
  NAND3_X1 U13283 ( .A1(n11126), .A2(n11044), .A3(n11146), .ZN(n11051) );
  NAND2_X1 U13284 ( .A1(n10369), .A2(n12345), .ZN(n13493) );
  NAND2_X1 U13285 ( .A1(n12346), .A2(n12343), .ZN(n10369) );
  INV_X1 U13286 ( .A(n12345), .ZN(n9806) );
  NAND2_X2 U13287 ( .A1(n12116), .A2(n12437), .ZN(n12499) );
  NOR2_X2 U13288 ( .A1(n12096), .A2(n12051), .ZN(n12437) );
  NAND2_X1 U13289 ( .A1(n12868), .A2(n9842), .ZN(n12949) );
  NAND2_X1 U13290 ( .A1(n12868), .A2(n12867), .ZN(n12873) );
  XNOR2_X1 U13291 ( .A(n12979), .B(n9844), .ZN(n16454) );
  INV_X1 U13292 ( .A(n16489), .ZN(n12965) );
  NAND2_X1 U13293 ( .A1(n12947), .A2(n12948), .ZN(n12957) );
  NAND2_X1 U13294 ( .A1(n9803), .A2(n14901), .ZN(n10386) );
  NAND2_X1 U13295 ( .A1(n14901), .A2(n14905), .ZN(n16703) );
  INV_X1 U13296 ( .A(n10386), .ZN(n16701) );
  INV_X1 U13297 ( .A(n16702), .ZN(n10382) );
  NAND2_X2 U13298 ( .A1(n12126), .A2(n14206), .ZN(n12562) );
  NAND2_X1 U13299 ( .A1(n14263), .A2(n9725), .ZN(n12425) );
  NOR2_X2 U13300 ( .A1(n12082), .A2(n12095), .ZN(n14263) );
  INV_X1 U13301 ( .A(n12051), .ZN(n10389) );
  NAND3_X1 U13302 ( .A1(n10390), .A2(n21077), .A3(n10389), .ZN(n13519) );
  OAI211_X2 U13303 ( .C1(n12568), .C2(n12124), .A(n13519), .B(n12425), .ZN(
        n12132) );
  XNOR2_X2 U13304 ( .A(n12167), .B(n9877), .ZN(n13767) );
  XNOR2_X2 U13305 ( .A(n12480), .B(n12479), .ZN(n13952) );
  NAND2_X1 U13306 ( .A1(n12826), .A2(n10407), .ZN(n10406) );
  AND2_X2 U13307 ( .A1(n12507), .A2(n10420), .ZN(n14526) );
  NAND2_X1 U13308 ( .A1(n16484), .A2(n10423), .ZN(n16448) );
  AND2_X1 U13309 ( .A1(n16484), .A2(n10424), .ZN(n16447) );
  AND2_X1 U13310 ( .A1(n16484), .A2(n13257), .ZN(n13256) );
  NAND3_X1 U13312 ( .A1(n13438), .A2(n10426), .A3(n13800), .ZN(n13439) );
  NAND2_X1 U13313 ( .A1(n15223), .A2(n10433), .ZN(n10432) );
  NOR2_X1 U13314 ( .A1(n15223), .A2(n15225), .ZN(n15224) );
  NAND2_X1 U13315 ( .A1(n14515), .A2(n15546), .ZN(n15450) );
  NAND2_X1 U13316 ( .A1(n12771), .A2(n12770), .ZN(n13297) );
  NAND2_X1 U13317 ( .A1(n15159), .A2(n15158), .ZN(n15160) );
  CLKBUF_X1 U13318 ( .A(n14788), .Z(n14949) );
  OAI21_X1 U13319 ( .B1(n13499), .B2(n13214), .A(n13213), .ZN(n13215) );
  NAND2_X1 U13320 ( .A1(n11051), .A2(n11050), .ZN(n11113) );
  NAND2_X1 U13321 ( .A1(n13212), .A2(n13245), .ZN(n13214) );
  NAND2_X1 U13322 ( .A1(n14879), .A2(n14878), .ZN(n14880) );
  INV_X1 U13323 ( .A(n15394), .ZN(n15411) );
  NAND2_X1 U13324 ( .A1(n13181), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15106) );
  AND2_X1 U13325 ( .A1(n16079), .A2(n9720), .ZN(n16345) );
  NOR2_X1 U13326 ( .A1(n16079), .A2(n14156), .ZN(n16287) );
  NOR2_X1 U13327 ( .A1(n16079), .A2(n9720), .ZN(n16346) );
  INV_X1 U13328 ( .A(n15103), .ZN(n13181) );
  INV_X1 U13329 ( .A(n13857), .ZN(n12722) );
  NAND2_X1 U13330 ( .A1(n15650), .A2(n15729), .ZN(n15651) );
  AND3_X1 U13331 ( .A1(n11732), .A2(n11731), .A3(n11730), .ZN(n11737) );
  AND2_X1 U13332 ( .A1(n10656), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11908) );
  AND2_X1 U13333 ( .A1(n12181), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12056) );
  CLKBUF_X1 U13334 ( .A(n12181), .Z(n14947) );
  XNOR2_X1 U13335 ( .A(n13446), .B(n10458), .ZN(n14729) );
  NAND2_X1 U13336 ( .A1(n13634), .A2(n12081), .ZN(n12099) );
  INV_X1 U13337 ( .A(n12843), .ZN(n12342) );
  INV_X1 U13338 ( .A(n12984), .ZN(n12981) );
  AND2_X4 U13339 ( .A1(n10522), .A2(n10524), .ZN(n18317) );
  INV_X1 U13340 ( .A(n12877), .ZN(n12868) );
  AOI22_X1 U13341 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11980) );
  AND2_X1 U13342 ( .A1(n13770), .A2(n13769), .ZN(n14876) );
  INV_X1 U13343 ( .A(n16444), .ZN(n16462) );
  XNOR2_X1 U13344 ( .A(n12347), .B(n12348), .ZN(n12843) );
  INV_X1 U13345 ( .A(n12609), .ZN(n13749) );
  NOR2_X1 U13346 ( .A1(n14584), .A2(n17051), .ZN(n10444) );
  INV_X1 U13347 ( .A(n21246), .ZN(n14349) );
  NAND2_X2 U13348 ( .A1(n15644), .A2(n13899), .ZN(n15643) );
  AND2_X1 U13349 ( .A1(n15497), .A2(n21250), .ZN(n10445) );
  AND2_X1 U13350 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21274), .ZN(n14159) );
  INV_X1 U13351 ( .A(n11190), .ZN(n11715) );
  NAND2_X1 U13352 ( .A1(n21075), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13833) );
  OR2_X1 U13353 ( .A1(n17142), .A2(n17098), .ZN(n10446) );
  INV_X1 U13354 ( .A(n15179), .ZN(n15180) );
  AND2_X1 U13355 ( .A1(n13461), .A2(n13460), .ZN(n10447) );
  AND2_X1 U13356 ( .A1(n13462), .A2(n10447), .ZN(n10448) );
  AND2_X1 U13357 ( .A1(n15840), .A2(n11170), .ZN(n10449) );
  NOR2_X1 U13358 ( .A1(n12651), .A2(n13761), .ZN(n10450) );
  AND2_X1 U13359 ( .A1(n18936), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10451) );
  INV_X1 U13360 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16916) );
  INV_X1 U13361 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16988) );
  AND2_X1 U13362 ( .A1(n15943), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10452) );
  INV_X1 U13363 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17094) );
  AND3_X1 U13364 ( .A1(n11743), .A2(n11742), .A3(n11741), .ZN(n10453) );
  AND2_X1 U13365 ( .A1(n15729), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10454) );
  AND2_X1 U13366 ( .A1(n11880), .A2(n19093), .ZN(n10455) );
  NAND3_X1 U13367 ( .A1(n13229), .A2(n19953), .A3(n17851), .ZN(n10456) );
  INV_X1 U13368 ( .A(n18638), .ZN(n18648) );
  INV_X2 U13369 ( .A(n18648), .ZN(n18642) );
  NAND2_X1 U13370 ( .A1(n18651), .A2(n18697), .ZN(n18638) );
  NOR2_X1 U13371 ( .A1(n14535), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10457) );
  INV_X1 U13372 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12394) );
  NOR2_X1 U13373 ( .A1(n19481), .A2(n19984), .ZN(n18189) );
  AND2_X1 U13374 ( .A1(n13445), .A2(n13444), .ZN(n10458) );
  AND2_X1 U13375 ( .A1(n12139), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10459) );
  INV_X1 U13376 ( .A(n11364), .ZN(n11383) );
  AND3_X1 U13377 ( .A1(n13444), .A2(n13284), .A3(n12924), .ZN(n10460) );
  INV_X1 U13378 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17036) );
  AND3_X1 U13379 ( .A1(n12230), .A2(n12229), .A3(n12228), .ZN(n10461) );
  NOR2_X1 U13380 ( .A1(n15120), .A2(n15119), .ZN(n10462) );
  AND2_X1 U13381 ( .A1(n12128), .A2(n12127), .ZN(n10463) );
  INV_X1 U13382 ( .A(n13845), .ZN(n21221) );
  INV_X1 U13383 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15015) );
  INV_X1 U13384 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13190) );
  AND2_X2 U13385 ( .A1(n13427), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15585)
         );
  INV_X1 U13386 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n21698) );
  AND2_X1 U13387 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10464) );
  AND2_X1 U13388 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10465) );
  NAND2_X1 U13389 ( .A1(n11257), .A2(n11256), .ZN(n10466) );
  INV_X1 U13390 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21584) );
  AND3_X1 U13391 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_17__SCAN_IN), .ZN(n10467) );
  INV_X1 U13393 ( .A(n13785), .ZN(n11078) );
  NOR2_X1 U13394 ( .A1(n10651), .A2(n10650), .ZN(n10468) );
  INV_X1 U13395 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17872) );
  INV_X1 U13396 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n21507) );
  OR2_X1 U13397 ( .A1(n21025), .A2(n15155), .ZN(n12586) );
  INV_X1 U13398 ( .A(n12586), .ZN(n20263) );
  INV_X1 U13399 ( .A(n20263), .ZN(n20169) );
  OR2_X1 U13400 ( .A1(n20321), .A2(n13718), .ZN(n20323) );
  INV_X2 U13401 ( .A(n20323), .ZN(n20344) );
  AND2_X1 U13402 ( .A1(n13295), .A2(n13459), .ZN(n10470) );
  AOI21_X1 U13403 ( .B1(n13799), .B2(n13800), .A(n13039), .ZN(n13875) );
  AND2_X2 U13404 ( .A1(n16444), .A2(n12791), .ZN(n10471) );
  OR2_X1 U13405 ( .A1(n18219), .A2(n17437), .ZN(n10472) );
  INV_X1 U13406 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n14687) );
  INV_X1 U13407 ( .A(n12499), .ZN(n12547) );
  AND2_X1 U13408 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10473) );
  INV_X1 U13409 ( .A(n17575), .ZN(n13212) );
  AND4_X1 U13410 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .ZN(
        n10474) );
  AND4_X1 U13411 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n10475) );
  AND2_X1 U13412 ( .A1(n10814), .A2(n10813), .ZN(n10476) );
  AND4_X1 U13413 ( .A1(n10845), .A2(n10844), .A3(n10843), .A4(n10842), .ZN(
        n10477) );
  AND4_X1 U13414 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10479) );
  AND4_X1 U13415 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10480) );
  INV_X1 U13416 ( .A(n13001), .ZN(n10884) );
  NAND2_X1 U13417 ( .A1(n10645), .A2(n19503), .ZN(n10646) );
  NAND2_X1 U13418 ( .A1(n10865), .A2(n11086), .ZN(n10866) );
  NAND2_X1 U13419 ( .A1(n9874), .A2(n12602), .ZN(n12084) );
  NAND2_X1 U13420 ( .A1(n12208), .A2(n12207), .ZN(n12215) );
  OAI21_X1 U13421 ( .B1(n10647), .B2(n19508), .A(n10646), .ZN(n10651) );
  INV_X1 U13422 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14992) );
  INV_X1 U13423 ( .A(n12123), .ZN(n12812) );
  INV_X1 U13424 ( .A(n10764), .ZN(n10767) );
  INV_X1 U13425 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10710) );
  OR2_X1 U13426 ( .A1(n17620), .A2(n16294), .ZN(n10906) );
  INV_X1 U13427 ( .A(n10779), .ZN(n10788) );
  AND2_X1 U13428 ( .A1(n14390), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12399) );
  AND2_X1 U13429 ( .A1(n16716), .A2(n14875), .ZN(n14873) );
  AOI22_X1 U13430 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12029) );
  INV_X1 U13431 ( .A(n14566), .ZN(n12640) );
  NAND2_X1 U13432 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10481) );
  INV_X1 U13433 ( .A(n14370), .ZN(n11215) );
  INV_X1 U13434 ( .A(n15375), .ZN(n11403) );
  INV_X1 U13435 ( .A(n11715), .ZN(n14683) );
  AND2_X1 U13436 ( .A1(n11146), .A2(n11150), .ZN(n11147) );
  OR2_X1 U13437 ( .A1(n11039), .A2(n11038), .ZN(n11048) );
  AND2_X1 U13438 ( .A1(n14994), .A2(n14993), .ZN(n17596) );
  INV_X1 U13439 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n21722) );
  INV_X1 U13440 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21621) );
  XNOR2_X1 U13441 ( .A(n11984), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12389) );
  AOI22_X1 U13442 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U13443 ( .A1(n12815), .A2(n12814), .ZN(n12824) );
  INV_X1 U13444 ( .A(n16513), .ZN(n12781) );
  NAND2_X1 U13445 ( .A1(n10474), .A2(n10475), .ZN(n12340) );
  INV_X1 U13446 ( .A(n12443), .ZN(n12621) );
  AND2_X1 U13447 ( .A1(n12168), .A2(n17393), .ZN(n12177) );
  AND3_X1 U13448 ( .A1(n10606), .A2(n10605), .A3(n10604), .ZN(n10610) );
  INV_X1 U13449 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15243) );
  INV_X1 U13450 ( .A(n11404), .ZN(n11405) );
  INV_X1 U13451 ( .A(n15395), .ZN(n13087) );
  AND4_X1 U13452 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10728) );
  NAND2_X1 U13453 ( .A1(n11053), .A2(n11094), .ZN(n11097) );
  INV_X1 U13454 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n21554) );
  NOR2_X1 U13455 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12394), .ZN(
        n21553) );
  NAND2_X1 U13456 ( .A1(n12115), .A2(n12114), .ZN(n12163) );
  AND2_X1 U13457 ( .A1(n14872), .A2(n14871), .ZN(n14875) );
  AND2_X1 U13458 ( .A1(n12777), .A2(n12776), .ZN(n13459) );
  INV_X1 U13459 ( .A(n14876), .ZN(n14897) );
  INV_X1 U13460 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15175) );
  INV_X1 U13461 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15136) );
  AND2_X1 U13462 ( .A1(n12928), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13281) );
  OAI211_X1 U13463 ( .C1(n12624), .C2(n20123), .A(n12607), .B(n12606), .ZN(
        n13745) );
  AND2_X1 U13464 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19961), .ZN(
        n10662) );
  INV_X1 U13465 ( .A(n18913), .ZN(n10506) );
  NAND2_X1 U13466 ( .A1(n17738), .A2(n18769), .ZN(n13213) );
  OAI21_X1 U13467 ( .B1(n19503), .B2(n10653), .A(n13218), .ZN(n11904) );
  INV_X1 U13468 ( .A(n11566), .ZN(n11504) );
  AND2_X1 U13469 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11195), .ZN(
        n11208) );
  INV_X1 U13470 ( .A(n14376), .ZN(n13052) );
  AND2_X1 U13471 ( .A1(n14687), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13405) );
  NOR2_X1 U13472 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11190) );
  NAND2_X1 U13473 ( .A1(n11235), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11269) );
  INV_X1 U13474 ( .A(n15969), .ZN(n16027) );
  NAND2_X1 U13475 ( .A1(n14372), .A2(n11106), .ZN(n11107) );
  OR2_X1 U13476 ( .A1(n10937), .A2(n10936), .ZN(n11055) );
  NOR2_X1 U13477 ( .A1(n10894), .A2(n13019), .ZN(n14680) );
  NOR2_X1 U13478 ( .A1(n14160), .A2(n14157), .ZN(n15083) );
  XNOR2_X1 U13479 ( .A(n13393), .B(n13392), .ZN(n15097) );
  OR2_X1 U13480 ( .A1(n12691), .A2(n12690), .ZN(n14477) );
  NOR2_X1 U13481 ( .A1(n14897), .A2(n13837), .ZN(n13838) );
  AND2_X1 U13482 ( .A1(n14855), .A2(n14854), .ZN(n14857) );
  INV_X1 U13483 ( .A(n16840), .ZN(n12770) );
  INV_X1 U13484 ( .A(n13896), .ZN(n12721) );
  NOR2_X1 U13485 ( .A1(n12338), .A2(n12337), .ZN(n12844) );
  INV_X1 U13486 ( .A(n15113), .ZN(n15116) );
  INV_X1 U13487 ( .A(n13281), .ZN(n16956) );
  AND2_X1 U13488 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U13489 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20473) );
  AND2_X1 U13490 ( .A1(n12167), .A2(n17393), .ZN(n12171) );
  INV_X1 U13491 ( .A(n12210), .ZN(n20862) );
  OR2_X1 U13492 ( .A1(n13920), .A2(n11920), .ZN(n13993) );
  OR2_X1 U13493 ( .A1(n9744), .A2(n10626), .ZN(n10630) );
  NAND2_X1 U13494 ( .A1(n11893), .A2(n18963), .ZN(n17521) );
  AND2_X1 U13495 ( .A1(n18997), .A2(n19268), .ZN(n18977) );
  INV_X1 U13496 ( .A(n18775), .ZN(n11927) );
  AND4_X1 U13497 ( .A1(n13481), .A2(n13480), .A3(n13479), .A4(n20960), .ZN(
        n13482) );
  OR2_X1 U13498 ( .A1(n11668), .A2(n15218), .ZN(n13464) );
  NAND2_X1 U13499 ( .A1(n11504), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11557) );
  OR2_X1 U13500 ( .A1(n11446), .A2(n15340), .ZN(n11484) );
  AND2_X1 U13501 ( .A1(n11208), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11217) );
  INV_X1 U13502 ( .A(n15429), .ZN(n21129) );
  INV_X1 U13503 ( .A(n15585), .ZN(n14022) );
  INV_X1 U13504 ( .A(n11640), .ZN(n15238) );
  NAND2_X1 U13505 ( .A1(n17671), .A2(n13789), .ZN(n17665) );
  INV_X1 U13506 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15653) );
  INV_X1 U13507 ( .A(n15335), .ZN(n15351) );
  AND2_X1 U13508 ( .A1(n13095), .A2(n13094), .ZN(n15352) );
  AND2_X1 U13509 ( .A1(n15664), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15793) );
  INV_X1 U13510 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17695) );
  AND2_X1 U13511 ( .A1(n13872), .A2(n13871), .ZN(n16055) );
  INV_X1 U13512 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16099) );
  OR2_X1 U13513 ( .A1(n13730), .A2(n13729), .ZN(n15012) );
  OR2_X1 U13514 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16161), .ZN(
        n16191) );
  INV_X1 U13515 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16294) );
  INV_X1 U13516 ( .A(n14436), .ZN(n16341) );
  AND2_X1 U13517 ( .A1(n14024), .A2(n14025), .ZN(n14034) );
  INV_X1 U13518 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21271) );
  NOR2_X1 U13519 ( .A1(n16203), .A2(n16202), .ZN(n16351) );
  AND2_X1 U13520 ( .A1(n21335), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17620) );
  AND2_X1 U13521 ( .A1(n12788), .A2(n12787), .ZN(n16460) );
  INV_X1 U13522 ( .A(n12947), .ZN(n12871) );
  INV_X1 U13523 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20187) );
  OR2_X1 U13524 ( .A1(n20306), .A2(n13743), .ZN(n14506) );
  AND3_X1 U13525 ( .A1(n12694), .A2(n12693), .A3(n12692), .ZN(n13807) );
  AND2_X1 U13526 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  INV_X1 U13527 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13453) );
  INV_X1 U13528 ( .A(n17723), .ZN(n17109) );
  NAND2_X1 U13529 ( .A1(n16976), .A2(n14708), .ZN(n14711) );
  INV_X1 U13530 ( .A(n13301), .ZN(n17305) );
  AND2_X1 U13531 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17367) );
  AND3_X1 U13532 ( .A1(n12590), .A2(n14662), .A3(n12589), .ZN(n17730) );
  OR3_X1 U13533 ( .A1(n12297), .A2(n20437), .A3(n20864), .ZN(n20419) );
  NOR2_X1 U13534 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21692), .ZN(
        n21552) );
  NAND2_X1 U13535 ( .A1(n21036), .A2(n21043), .ZN(n20741) );
  INV_X1 U13536 ( .A(n14400), .ZN(n20571) );
  NAND2_X1 U13537 ( .A1(n20864), .A2(n20821), .ZN(n21065) );
  OR3_X1 U13538 ( .A1(n20862), .A2(n20917), .A3(n20864), .ZN(n20873) );
  NAND2_X1 U13539 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U13540 ( .A1(n10682), .A2(n10472), .ZN(n10688) );
  INV_X1 U13541 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18967) );
  INV_X1 U13542 ( .A(n18169), .ZN(n18205) );
  INV_X1 U13543 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13510) );
  INV_X1 U13544 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18916) );
  INV_X1 U13545 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21563) );
  INV_X1 U13546 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18993) );
  INV_X1 U13547 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19159) );
  INV_X1 U13548 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19134) );
  INV_X1 U13549 ( .A(n17452), .ZN(n19004) );
  INV_X1 U13550 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19012) );
  AND2_X1 U13551 ( .A1(n13217), .A2(n13222), .ZN(n13243) );
  INV_X1 U13552 ( .A(n19965), .ZN(n14124) );
  INV_X1 U13553 ( .A(n19657), .ZN(n19658) );
  NAND2_X1 U13554 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n20083) );
  INV_X1 U13555 ( .A(n21089), .ZN(n14679) );
  INV_X1 U13556 ( .A(n21147), .ZN(n21163) );
  INV_X1 U13557 ( .A(n21122), .ZN(n21182) );
  AND2_X1 U13558 ( .A1(n15644), .A2(n15558), .ZN(n13416) );
  NOR2_X1 U13559 ( .A1(n15637), .A2(n13899), .ZN(n15639) );
  INV_X2 U13560 ( .A(n14327), .ZN(n21245) );
  NOR2_X2 U13561 ( .A1(n21245), .A2(n14287), .ZN(n21231) );
  INV_X1 U13562 ( .A(n17666), .ZN(n17654) );
  INV_X1 U13563 ( .A(n21094), .ZN(n17668) );
  NOR2_X2 U13564 ( .A1(n15289), .A2(n15290), .ZN(n15291) );
  OAI21_X1 U13565 ( .B1(n13166), .B2(n15090), .A(n13906), .ZN(n16031) );
  INV_X1 U13566 ( .A(n16030), .ZN(n17673) );
  NAND2_X1 U13567 ( .A1(n10219), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16112) );
  INV_X1 U13568 ( .A(n16167), .ZN(n16193) );
  NAND3_X1 U13569 ( .A1(n16166), .A2(n16165), .A3(n16256), .ZN(n16189) );
  AND2_X1 U13570 ( .A1(n16079), .A2(n14156), .ZN(n16118) );
  OAI21_X1 U13571 ( .B1(n16247), .B2(n16208), .A(n16207), .ZN(n16242) );
  INV_X1 U13572 ( .A(n16280), .ZN(n14366) );
  OAI21_X1 U13573 ( .B1(n15025), .B2(n16251), .A(n21281), .ZN(n14184) );
  NOR3_X1 U13574 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15029), .A3(
        n16294), .ZN(n16251) );
  AND2_X1 U13575 ( .A1(n14024), .A2(n14434), .ZN(n21266) );
  OAI211_X1 U13576 ( .C1(n14446), .C2(n14445), .A(n14444), .B(n16166), .ZN(
        n14470) );
  OAI21_X1 U13577 ( .B1(n14037), .B2(n14036), .A(n21281), .ZN(n21754) );
  OAI211_X1 U13578 ( .C1(n16301), .C2(n16300), .A(n16351), .B(n16299), .ZN(
        n16337) );
  AND2_X1 U13579 ( .A1(n14034), .A2(n14156), .ZN(n16336) );
  AND2_X1 U13580 ( .A1(n21280), .A2(n16346), .ZN(n21329) );
  OAI21_X1 U13581 ( .B1(n21277), .B2(n21276), .A(n21275), .ZN(n21324) );
  OAI211_X1 U13582 ( .C1(n16352), .C2(n16377), .A(n16351), .B(n16350), .ZN(
        n16374) );
  NOR2_X1 U13583 ( .A1(n16202), .A2(n14292), .ZN(n21278) );
  INV_X1 U13584 ( .A(n16317), .ZN(n21307) );
  NAND2_X1 U13585 ( .A1(n21281), .A2(n16389), .ZN(n16423) );
  INV_X1 U13586 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21345) );
  INV_X1 U13587 ( .A(n21408), .ZN(n21403) );
  INV_X1 U13588 ( .A(n13718), .ZN(n21070) );
  INV_X1 U13589 ( .A(n20929), .ZN(n13521) );
  OR2_X1 U13590 ( .A1(n10471), .A2(n13381), .ZN(n13382) );
  INV_X1 U13591 ( .A(n20260), .ZN(n20246) );
  AND2_X1 U13592 ( .A1(n20350), .A2(n15164), .ZN(n20235) );
  OR2_X1 U13593 ( .A1(n13950), .A2(n13949), .ZN(n13951) );
  OR2_X1 U13594 ( .A1(n12745), .A2(n12744), .ZN(n14530) );
  OR2_X1 U13595 ( .A1(n12704), .A2(n12703), .ZN(n14618) );
  NOR2_X1 U13596 ( .A1(n14578), .A2(n14476), .ZN(n14406) );
  AND2_X1 U13597 ( .A1(n14919), .A2(n14918), .ZN(n16697) );
  AND3_X1 U13598 ( .A1(n12648), .A2(n12647), .A3(n12646), .ZN(n14563) );
  INV_X1 U13599 ( .A(n14282), .ZN(n20306) );
  INV_X1 U13600 ( .A(n15096), .ZN(n20350) );
  INV_X1 U13601 ( .A(n14505), .ZN(n14399) );
  INV_X1 U13602 ( .A(n17116), .ZN(n17718) );
  AND2_X1 U13603 ( .A1(n12447), .A2(n12448), .ZN(n21056) );
  INV_X1 U13604 ( .A(n16645), .ZN(n21029) );
  NOR2_X1 U13605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20416), .ZN(
        n20394) );
  OR2_X1 U13606 ( .A1(n20452), .A2(n20823), .ZN(n20469) );
  INV_X1 U13607 ( .A(n20505), .ZN(n20498) );
  NOR2_X2 U13608 ( .A1(n20598), .A2(n20741), .ZN(n20535) );
  NOR2_X1 U13609 ( .A1(n20569), .A2(n20539), .ZN(n20564) );
  NOR2_X1 U13610 ( .A1(n20598), .A2(n20539), .ZN(n20588) );
  NAND2_X1 U13611 ( .A1(n20422), .A2(n20421), .ZN(n20598) );
  NAND2_X1 U13612 ( .A1(n21036), .A2(n20369), .ZN(n20674) );
  INV_X1 U13613 ( .A(n20742), .ZN(n20767) );
  NOR2_X2 U13614 ( .A1(n20671), .A2(n20741), .ZN(n20787) );
  NOR2_X2 U13615 ( .A1(n20813), .A2(n20539), .ZN(n20808) );
  INV_X1 U13616 ( .A(n20897), .ZN(n20839) );
  AND2_X1 U13617 ( .A1(n20407), .A2(n14604), .ZN(n20892) );
  NOR2_X2 U13618 ( .A1(n20813), .A2(n20869), .ZN(n20921) );
  AOI21_X1 U13619 ( .B1(n20864), .B2(n17409), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n21072) );
  NOR2_X1 U13620 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20949) );
  INV_X1 U13621 ( .A(n21073), .ZN(n21071) );
  INV_X1 U13622 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20955) );
  NAND2_X1 U13623 ( .A1(n20087), .A2(n19953), .ZN(n18857) );
  OR2_X1 U13624 ( .A1(n10688), .A2(n10687), .ZN(n10689) );
  NOR2_X1 U13625 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17963), .ZN(n17951) );
  OR2_X1 U13626 ( .A1(n20105), .A2(n10681), .ZN(n18212) );
  NOR2_X1 U13627 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18096), .ZN(n18086) );
  NOR2_X1 U13628 ( .A1(n19968), .A2(n10677), .ZN(n18169) );
  NOR2_X1 U13629 ( .A1(n21460), .A2(n18144), .ZN(n18140) );
  INV_X1 U13630 ( .A(n18219), .ZN(n18193) );
  INV_X1 U13631 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21576) );
  INV_X1 U13632 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18123) );
  NOR3_X1 U13633 ( .A1(n18697), .A2(n18731), .A3(n18861), .ZN(n18723) );
  OR2_X1 U13634 ( .A1(n18655), .A2(n18697), .ZN(n18739) );
  INV_X1 U13635 ( .A(n19059), .ZN(n19103) );
  OAI211_X1 U13636 ( .C1(n20083), .C2(n19496), .A(n18856), .B(n18855), .ZN(
        n18882) );
  OR2_X1 U13637 ( .A1(n11831), .A2(n11830), .ZN(n13245) );
  AND2_X1 U13638 ( .A1(n19252), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13502) );
  NOR2_X2 U13639 ( .A1(n19151), .A2(n19481), .ZN(n19124) );
  NAND2_X1 U13640 ( .A1(n19783), .A2(n19837), .ZN(n19507) );
  INV_X1 U13641 ( .A(n19210), .ZN(n19220) );
  NOR2_X1 U13642 ( .A1(n19477), .A2(n17578), .ZN(n13240) );
  INV_X1 U13643 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19235) );
  INV_X1 U13644 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19257) );
  INV_X1 U13645 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19303) );
  NOR2_X1 U13646 ( .A1(n19373), .A2(n19459), .ZN(n19404) );
  AND2_X1 U13647 ( .A1(n19470), .A2(n13243), .ZN(n19443) );
  NOR2_X1 U13648 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n20103) );
  CLKBUF_X1 U13649 ( .A(n19556), .Z(n19580) );
  INV_X1 U13650 ( .A(n19609), .ZN(n19600) );
  INV_X1 U13651 ( .A(n19627), .ZN(n19628) );
  INV_X1 U13652 ( .A(n19650), .ZN(n19651) );
  INV_X1 U13653 ( .A(n19704), .ZN(n19685) );
  INV_X1 U13654 ( .A(n19723), .ZN(n19718) );
  INV_X1 U13655 ( .A(n19772), .ZN(n19773) );
  INV_X1 U13656 ( .A(n19888), .ZN(n19812) );
  NOR2_X1 U13657 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19942), .ZN(
        n19779) );
  NOR2_X1 U13658 ( .A1(n19493), .A2(n19520), .ZN(n19872) );
  AND2_X1 U13659 ( .A1(n19783), .A2(BUF2_REG_3__SCAN_IN), .ZN(n19889) );
  NOR2_X1 U13660 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20070), .ZN(n19978) );
  INV_X1 U13661 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19988) );
  INV_X1 U13662 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21428) );
  INV_X1 U13663 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21681) );
  NAND2_X1 U13664 ( .A1(n15544), .A2(n14057), .ZN(n15556) );
  NAND2_X1 U13665 ( .A1(n15544), .A2(n15558), .ZN(n15545) );
  AND2_X1 U13666 ( .A1(n13903), .A2(n13902), .ZN(n14292) );
  NAND2_X1 U13667 ( .A1(n21206), .A2(n14697), .ZN(n21191) );
  OR2_X1 U13668 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17704), .ZN(n21218) );
  NOR2_X1 U13669 ( .A1(n15196), .A2(n14284), .ZN(n14327) );
  INV_X1 U13670 ( .A(n11722), .ZN(n11723) );
  NAND2_X1 U13671 ( .A1(n21094), .A2(n11717), .ZN(n17671) );
  INV_X1 U13672 ( .A(n21250), .ZN(n16051) );
  INV_X1 U13673 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U13674 ( .A1(n16126), .A2(n16124), .B1(n16203), .B2(n16122), .ZN(
        n16157) );
  NAND2_X1 U13675 ( .A1(n14541), .A2(n16346), .ZN(n16167) );
  AOI22_X1 U13676 ( .A1(n16163), .A2(n16160), .B1(n16203), .B2(n16249), .ZN(
        n16196) );
  NAND2_X1 U13677 ( .A1(n14541), .A2(n16118), .ZN(n16237) );
  NOR2_X1 U13678 ( .A1(n16205), .A2(n16204), .ZN(n16245) );
  INV_X1 U13679 ( .A(n14351), .ZN(n14369) );
  AOI22_X1 U13680 ( .A1(n16255), .A2(n16250), .B1(n16249), .B2(n16342), .ZN(
        n16286) );
  AOI22_X1 U13681 ( .A1(n14154), .A2(n21274), .B1(n16251), .B2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14187) );
  NAND3_X1 U13682 ( .A1(n14024), .A2(n16287), .A3(n11176), .ZN(n21270) );
  AOI22_X1 U13683 ( .A1(n14437), .A2(n14445), .B1(n16203), .B2(n16343), .ZN(
        n14473) );
  INV_X1 U13684 ( .A(n16336), .ZN(n21757) );
  AOI22_X1 U13685 ( .A1(n16293), .A2(n16300), .B1(n16342), .B2(n16292), .ZN(
        n16340) );
  NAND2_X1 U13686 ( .A1(n21280), .A2(n16287), .ZN(n21333) );
  AOI22_X1 U13687 ( .A1(n16344), .A2(n21274), .B1(n16343), .B2(n16342), .ZN(
        n16380) );
  INV_X1 U13688 ( .A(n21306), .ZN(n16412) );
  NOR2_X1 U13689 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17708) );
  NOR2_X1 U13690 ( .A1(n21438), .A2(n21348), .ZN(n21339) );
  INV_X1 U13691 ( .A(n21339), .ZN(n21416) );
  INV_X1 U13692 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21363) );
  NAND2_X1 U13693 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21438), .ZN(n21402) );
  INV_X1 U13694 ( .A(n21438), .ZN(n21425) );
  INV_X1 U13695 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20937) );
  NAND2_X1 U13696 ( .A1(n13178), .A2(n13177), .ZN(n13522) );
  OR3_X1 U13697 ( .A1(n21069), .A2(n12388), .A3(n15166), .ZN(n20251) );
  OR2_X1 U13698 ( .A1(n20184), .A2(n20183), .ZN(n20195) );
  INV_X1 U13699 ( .A(n20235), .ZN(n20267) );
  OR2_X1 U13700 ( .A1(n14625), .A2(n14529), .ZN(n20191) );
  AND2_X1 U13701 ( .A1(n13636), .A2(n20929), .ZN(n20291) );
  INV_X1 U13702 ( .A(n20307), .ZN(n16868) );
  INV_X1 U13703 ( .A(n16819), .ZN(n20402) );
  AND2_X1 U13704 ( .A1(n13581), .A2(n13580), .ZN(n20305) );
  NAND2_X1 U13705 ( .A1(n20321), .A2(n9888), .ZN(n13720) );
  INV_X1 U13706 ( .A(n20321), .ZN(n20348) );
  OR2_X1 U13707 ( .A1(n13532), .A2(n21078), .ZN(n15096) );
  NAND2_X1 U13708 ( .A1(n13522), .A2(n13180), .ZN(n17723) );
  NAND2_X1 U13709 ( .A1(n13186), .A2(n14904), .ZN(n17116) );
  INV_X1 U13710 ( .A(n13270), .ZN(n13271) );
  NAND2_X1 U13711 ( .A1(n12998), .A2(n21056), .ZN(n20358) );
  INV_X1 U13712 ( .A(n17574), .ZN(n21022) );
  OR2_X1 U13713 ( .A1(n20674), .A2(n20569), .ZN(n20442) );
  INV_X1 U13714 ( .A(n20443), .ZN(n20472) );
  AND2_X1 U13715 ( .A1(n20479), .A2(n20478), .ZN(n20492) );
  INV_X1 U13716 ( .A(n20535), .ZN(n20513) );
  INV_X1 U13717 ( .A(n20564), .ZN(n20562) );
  INV_X1 U13718 ( .A(n20588), .ZN(n20597) );
  OR2_X1 U13719 ( .A1(n20869), .A2(n20598), .ZN(n20670) );
  OR2_X1 U13720 ( .A1(n20813), .A2(n20674), .ZN(n20705) );
  INV_X1 U13721 ( .A(n20711), .ZN(n20734) );
  INV_X1 U13722 ( .A(n20894), .ZN(n20757) );
  AOI21_X1 U13723 ( .B1(n14599), .B2(n14598), .A(n14597), .ZN(n20790) );
  INV_X1 U13724 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21637) );
  OR2_X1 U13725 ( .A1(n20671), .A2(n20869), .ZN(n20925) );
  AND2_X1 U13726 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13516), .ZN(n17411) );
  INV_X1 U13727 ( .A(n21016), .ZN(n20935) );
  INV_X1 U13728 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20957) );
  INV_X1 U13729 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U13730 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20937), .ZN(n21085) );
  INV_X1 U13731 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17849) );
  NOR4_X1 U13732 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13376) );
  INV_X1 U13733 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17924) );
  INV_X1 U13734 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18987) );
  NAND2_X1 U13735 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18212), .ZN(n18219) );
  INV_X1 U13736 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18155) );
  NOR2_X1 U13737 ( .A1(n18832), .A2(n18758), .ZN(n18755) );
  NOR2_X1 U13738 ( .A1(n18836), .A2(n18761), .ZN(n18764) );
  INV_X1 U13739 ( .A(n18786), .ZN(n18794) );
  INV_X1 U13740 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18797) );
  OR2_X1 U13741 ( .A1(n20084), .A2(n18841), .ZN(n18821) );
  NAND2_X1 U13742 ( .A1(n18841), .A2(n18798), .ZN(n18823) );
  OR2_X1 U13743 ( .A1(n19481), .A2(n19103), .ZN(n18843) );
  INV_X1 U13744 ( .A(n18841), .ZN(n18853) );
  INV_X1 U13745 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19489) );
  INV_X1 U13746 ( .A(n18905), .ZN(n18900) );
  INV_X1 U13747 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18908) );
  OR2_X2 U13748 ( .A1(n19217), .A2(n13245), .ZN(n19177) );
  INV_X1 U13749 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n19142) );
  INV_X1 U13750 ( .A(n19477), .ZN(n19216) );
  INV_X1 U13751 ( .A(n19190), .ZN(n19223) );
  NAND2_X1 U13752 ( .A1(n13241), .A2(n13240), .ZN(n13250) );
  INV_X1 U13753 ( .A(n19477), .ZN(n19428) );
  INV_X1 U13754 ( .A(n19377), .ZN(n19416) );
  OR2_X1 U13755 ( .A1(n19470), .A2(n19477), .ZN(n19466) );
  INV_X1 U13756 ( .A(n19476), .ZN(n19430) );
  INV_X1 U13757 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19961) );
  NAND2_X1 U13758 ( .A1(n19657), .A2(n19705), .ZN(n19704) );
  INV_X1 U13759 ( .A(n19750), .ZN(n19749) );
  INV_X1 U13760 ( .A(n19872), .ZN(n19786) );
  INV_X1 U13761 ( .A(n19885), .ZN(n19815) );
  INV_X1 U13762 ( .A(n19891), .ZN(n19849) );
  NAND2_X1 U13763 ( .A1(n19871), .A2(BUF2_REG_23__SCAN_IN), .ZN(n19864) );
  NAND2_X1 U13764 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19871), .ZN(n19888) );
  INV_X1 U13765 ( .A(n20087), .ZN(n19976) );
  AOI22_X1 U13766 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19994), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n20001), .ZN(n20067) );
  INV_X1 U13767 ( .A(HOLD), .ZN(n21355) );
  INV_X1 U13768 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20020) );
  INV_X1 U13769 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20048) );
  INV_X2 U13770 ( .A(n20099), .ZN(n20101) );
  INV_X1 U13771 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n21470) );
  INV_X1 U13772 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19518) );
  INV_X1 U13773 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19499) );
  INV_X1 U13774 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20960) );
  INV_X1 U13775 ( .A(n17843), .ZN(n17844) );
  OAI21_X1 U13776 ( .B1(n14729), .B2(n20360), .A(n10448), .ZN(P2_U3025) );
  NAND2_X1 U13777 ( .A1(n13250), .A2(n13249), .ZN(P3_U2834) );
  AND3_X1 U13778 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18075) );
  NAND3_X1 U13779 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18075), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18059) );
  INV_X1 U13780 ( .A(n18059), .ZN(n19106) );
  INV_X1 U13781 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n19120) );
  NAND2_X1 U13782 ( .A1(n19102), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19063) );
  NAND4_X1 U13783 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10483) );
  INV_X1 U13784 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18951) );
  INV_X1 U13785 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13369) );
  XNOR2_X1 U13786 ( .A(n10490), .B(n13369), .ZN(n13365) );
  INV_X1 U13787 ( .A(n10482), .ZN(n19017) );
  NAND2_X1 U13788 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19017), .ZN(
        n10488) );
  INV_X1 U13789 ( .A(n10498), .ZN(n10486) );
  NAND2_X1 U13790 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18937), .ZN(
        n10501) );
  INV_X1 U13791 ( .A(n10501), .ZN(n10502) );
  NAND2_X1 U13792 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n10502), .ZN(
        n10484) );
  NAND2_X1 U13793 ( .A1(n18936), .A2(n10502), .ZN(n13508) );
  INV_X1 U13794 ( .A(n13508), .ZN(n10504) );
  AOI21_X1 U13795 ( .B1(n21563), .B2(n10484), .A(n10504), .ZN(n18940) );
  NAND2_X1 U13796 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10498), .ZN(
        n10485) );
  AOI21_X1 U13797 ( .B1(n18987), .B2(n10485), .A(n18937), .ZN(n18985) );
  AOI22_X1 U13798 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10498), .B1(
        n10486), .B2(n18993), .ZN(n18996) );
  INV_X1 U13799 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19018) );
  NOR2_X1 U13800 ( .A1(n19018), .A2(n10488), .ZN(n10495) );
  AOI21_X1 U13801 ( .B1(n19018), .B2(n10488), .A(n10495), .ZN(n19046) );
  INV_X1 U13802 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19065) );
  INV_X1 U13803 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19078) );
  NAND2_X1 U13804 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n10487), .ZN(
        n19058) );
  NOR2_X1 U13805 ( .A1(n19078), .A2(n19058), .ZN(n10492) );
  INV_X1 U13806 ( .A(n10492), .ZN(n18020) );
  INV_X1 U13807 ( .A(n10488), .ZN(n10489) );
  AOI21_X1 U13808 ( .B1(n19065), .B2(n18020), .A(n10489), .ZN(n19060) );
  INV_X1 U13809 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18221) );
  NAND2_X1 U13810 ( .A1(n10490), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10491) );
  XNOR2_X2 U13811 ( .A(n10491), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10512) );
  NOR2_X1 U13812 ( .A1(n19046), .A2(n18004), .ZN(n18003) );
  NOR2_X1 U13813 ( .A1(n18003), .A2(n9750), .ZN(n17993) );
  INV_X1 U13814 ( .A(n17993), .ZN(n10494) );
  INV_X1 U13815 ( .A(n10495), .ZN(n19020) );
  INV_X1 U13816 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21731) );
  AOI22_X1 U13817 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n10495), .B1(
        n19020), .B2(n21731), .ZN(n19036) );
  INV_X1 U13818 ( .A(n19036), .ZN(n10493) );
  INV_X1 U13819 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19021) );
  NAND2_X1 U13820 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n10495), .ZN(
        n10497) );
  NAND3_X1 U13821 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n10495), .ZN(n18983) );
  INV_X1 U13822 ( .A(n18983), .ZN(n10496) );
  AOI21_X1 U13823 ( .B1(n19021), .B2(n10497), .A(n10496), .ZN(n19024) );
  INV_X1 U13824 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n19002) );
  AOI21_X1 U13825 ( .B1(n19002), .B2(n18983), .A(n10498), .ZN(n19005) );
  NOR2_X1 U13826 ( .A1(n17969), .A2(n19005), .ZN(n17968) );
  NOR2_X1 U13827 ( .A1(n17968), .A2(n9750), .ZN(n17961) );
  NOR2_X1 U13828 ( .A1(n18996), .A2(n17961), .ZN(n17960) );
  NOR2_X1 U13829 ( .A1(n17960), .A2(n9750), .ZN(n17953) );
  NOR2_X1 U13830 ( .A1(n18985), .A2(n17953), .ZN(n17952) );
  NOR2_X1 U13831 ( .A1(n17952), .A2(n9750), .ZN(n17936) );
  INV_X1 U13832 ( .A(n17936), .ZN(n10500) );
  OAI21_X1 U13833 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18937), .A(
        n10501), .ZN(n10499) );
  INV_X1 U13834 ( .A(n10499), .ZN(n18968) );
  NAND2_X1 U13835 ( .A1(n10500), .A2(n10499), .ZN(n17934) );
  AND2_X2 U13836 ( .A1(n17934), .A2(n18132), .ZN(n17928) );
  AOI22_X1 U13837 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n10502), .B1(
        n10501), .B2(n18951), .ZN(n18960) );
  NOR2_X1 U13838 ( .A1(n17928), .A2(n18960), .ZN(n17927) );
  NOR2_X1 U13839 ( .A1(n17927), .A2(n9750), .ZN(n17915) );
  NOR2_X1 U13840 ( .A1(n18940), .A2(n17915), .ZN(n17914) );
  NOR2_X1 U13841 ( .A1(n17914), .A2(n9750), .ZN(n17906) );
  OAI21_X1 U13842 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n10504), .A(
        n10503), .ZN(n10505) );
  INV_X1 U13843 ( .A(n10505), .ZN(n18928) );
  NOR2_X1 U13844 ( .A1(n17906), .A2(n18928), .ZN(n17904) );
  OR2_X1 U13845 ( .A1(n17904), .A2(n9750), .ZN(n17890) );
  NOR2_X1 U13846 ( .A1(n18916), .A2(n10503), .ZN(n10508) );
  AOI21_X1 U13847 ( .B1(n18916), .B2(n10503), .A(n10508), .ZN(n18913) );
  AND2_X2 U13848 ( .A1(n17891), .A2(n18132), .ZN(n17883) );
  NOR2_X1 U13849 ( .A1(n10508), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10509) );
  NOR2_X1 U13850 ( .A1(n17883), .A2(n10510), .ZN(n17882) );
  NOR2_X1 U13851 ( .A1(n17882), .A2(n9750), .ZN(n17870) );
  INV_X1 U13852 ( .A(n10507), .ZN(n10511) );
  AOI21_X1 U13853 ( .B1(n17872), .B2(n10511), .A(n10490), .ZN(n17871) );
  NOR2_X1 U13854 ( .A1(n17870), .A2(n17871), .ZN(n17869) );
  NOR2_X1 U13855 ( .A1(n17869), .A2(n9750), .ZN(n13364) );
  INV_X1 U13856 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20092) );
  NAND3_X1 U13857 ( .A1(n20092), .A2(n20102), .A3(n17849), .ZN(n19984) );
  NAND2_X1 U13858 ( .A1(n18132), .A2(n18189), .ZN(n18220) );
  NOR3_X1 U13859 ( .A1(n13365), .A2(n13364), .A3(n18220), .ZN(n10691) );
  INV_X1 U13860 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10515) );
  INV_X2 U13861 ( .A(n10611), .ZN(n11802) );
  NAND2_X1 U13862 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10514) );
  NAND2_X1 U13863 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10513) );
  OAI211_X1 U13864 ( .C1(n10515), .C2(n9745), .A(n10514), .B(n10513), .ZN(
        n10516) );
  INV_X1 U13865 ( .A(n10516), .ZN(n10520) );
  AOI22_X1 U13866 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10519) );
  AND2_X2 U13867 ( .A1(n10523), .A2(n10522), .ZN(n17550) );
  AOI22_X1 U13868 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U13869 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10517) );
  NAND4_X1 U13870 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10530) );
  AOI22_X1 U13871 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10528) );
  AND2_X2 U13872 ( .A1(n10522), .A2(n13935), .ZN(n10603) );
  AOI22_X1 U13873 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10527) );
  AND2_X2 U13874 ( .A1(n10523), .A2(n14113), .ZN(n18606) );
  AND2_X2 U13875 ( .A1(n10522), .A2(n14667), .ZN(n11842) );
  AOI22_X1 U13876 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13877 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10525) );
  NAND4_X1 U13878 ( .A1(n10528), .A2(n10527), .A3(n10526), .A4(n10525), .ZN(
        n10529) );
  OR2_X2 U13879 ( .A1(n10530), .A2(n10529), .ZN(n18798) );
  INV_X1 U13880 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13881 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10531) );
  OAI211_X1 U13882 ( .C1(n10533), .C2(n9745), .A(n10532), .B(n10531), .ZN(
        n10534) );
  INV_X1 U13883 ( .A(n10534), .ZN(n10538) );
  AOI22_X1 U13884 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13885 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10536) );
  NAND2_X1 U13886 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10535) );
  AOI22_X1 U13887 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13888 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13889 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13890 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10541) );
  INV_X1 U13891 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13892 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10548) );
  NAND2_X1 U13893 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10547) );
  OAI211_X1 U13894 ( .C1(n10549), .C2(n9744), .A(n10548), .B(n10547), .ZN(
        n10550) );
  INV_X1 U13895 ( .A(n10550), .ZN(n10554) );
  AOI22_X1 U13896 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13897 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U13898 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10551) );
  NAND4_X1 U13899 ( .A1(n10554), .A2(n10553), .A3(n10552), .A4(n10551), .ZN(
        n10560) );
  AOI22_X1 U13900 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13901 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13902 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13903 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10555) );
  NAND4_X1 U13904 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10559) );
  INV_X1 U13905 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U13906 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10562) );
  NAND2_X1 U13907 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10561) );
  OAI211_X1 U13908 ( .C1(n10563), .C2(n9726), .A(n10562), .B(n10561), .ZN(
        n10564) );
  INV_X1 U13909 ( .A(n10564), .ZN(n10568) );
  AOI22_X1 U13910 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13911 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10566) );
  NAND2_X1 U13912 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10565) );
  NAND4_X1 U13913 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n10574) );
  AOI22_X1 U13914 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13915 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13916 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13917 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10569) );
  NAND4_X1 U13918 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10573) );
  INV_X1 U13919 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U13920 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13921 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10575) );
  OAI211_X1 U13922 ( .C1(n10577), .C2(n9745), .A(n10576), .B(n10575), .ZN(
        n10578) );
  INV_X1 U13923 ( .A(n10578), .ZN(n10582) );
  AOI22_X1 U13924 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13925 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13926 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10579) );
  NAND4_X1 U13927 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10588) );
  AOI22_X1 U13928 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13929 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13930 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13931 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10583) );
  NAND4_X1 U13932 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10587) );
  INV_X1 U13933 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U13934 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10590) );
  NAND2_X1 U13935 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10589) );
  OAI211_X1 U13936 ( .C1(n10591), .C2(n9745), .A(n10590), .B(n10589), .ZN(
        n10592) );
  INV_X1 U13937 ( .A(n10592), .ZN(n10596) );
  AOI22_X1 U13938 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13939 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10594) );
  NAND2_X1 U13940 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10593) );
  NAND4_X1 U13941 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n10602) );
  AOI22_X1 U13942 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13943 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13944 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13945 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10597) );
  NAND4_X1 U13946 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .ZN(
        n10601) );
  NAND2_X1 U13947 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10606) );
  NAND2_X1 U13948 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10605) );
  NAND2_X1 U13949 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10604) );
  AOI22_X1 U13950 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13951 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13952 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10607) );
  NAND4_X1 U13953 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10607), .ZN(
        n10617) );
  AOI22_X1 U13954 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13955 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18613), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13956 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11802), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13957 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13958 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10616) );
  NAND2_X1 U13959 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10621) );
  NAND2_X1 U13960 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10620) );
  NAND2_X1 U13961 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13962 ( .A1(n11843), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U13963 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13964 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13965 ( .A1(n18611), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13966 ( .A1(n17549), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13967 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10629) );
  INV_X2 U13968 ( .A(n10611), .ZN(n18570) );
  NAND2_X1 U13969 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10628) );
  NAND2_X1 U13970 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10627) );
  NAND2_X1 U13971 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10634) );
  NAND2_X1 U13972 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10633) );
  NAND2_X1 U13973 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13974 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10631) );
  NOR2_X1 U13975 ( .A1(n18798), .A2(n19521), .ZN(n10644) );
  NOR2_X1 U13976 ( .A1(n20089), .A2(n18798), .ZN(n13996) );
  NAND2_X1 U13977 ( .A1(n19500), .A2(n19503), .ZN(n13920) );
  NAND2_X1 U13978 ( .A1(n19511), .A2(n11922), .ZN(n11920) );
  INV_X1 U13979 ( .A(n13993), .ZN(n10640) );
  NAND3_X1 U13980 ( .A1(n13996), .A2(n18697), .A3(n10640), .ZN(n10641) );
  NAND2_X1 U13981 ( .A1(n19500), .A2(n18659), .ZN(n13229) );
  AOI211_X1 U13982 ( .C1(n18697), .C2(n14115), .A(n19493), .B(n20089), .ZN(
        n13219) );
  AOI21_X1 U13983 ( .B1(n10649), .B2(n13229), .A(n13219), .ZN(n10653) );
  INV_X1 U13984 ( .A(n11919), .ZN(n10642) );
  AOI211_X1 U13985 ( .C1(n19508), .C2(n18659), .A(n10642), .B(n11898), .ZN(
        n10643) );
  NOR2_X1 U13986 ( .A1(n19521), .A2(n10648), .ZN(n10647) );
  INV_X1 U13987 ( .A(n10644), .ZN(n10645) );
  NAND2_X1 U13988 ( .A1(n19500), .A2(n10648), .ZN(n13221) );
  AOI21_X1 U13989 ( .B1(n10649), .B2(n13221), .A(n18798), .ZN(n10650) );
  INV_X1 U13990 ( .A(n11902), .ZN(n10655) );
  MUX2_X1 U13991 ( .A(n19755), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11907) );
  NAND2_X1 U13992 ( .A1(n11907), .A2(n11908), .ZN(n10669) );
  NAND2_X1 U13993 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19755), .ZN(
        n10657) );
  NAND2_X1 U13994 ( .A1(n10669), .A2(n10657), .ZN(n10667) );
  MUX2_X1 U13995 ( .A(n19938), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10665) );
  INV_X1 U13996 ( .A(n10673), .ZN(n10659) );
  NAND2_X1 U13997 ( .A1(n10659), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10664) );
  INV_X1 U13998 ( .A(n10660), .ZN(n10661) );
  NAND2_X1 U13999 ( .A1(n10661), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10670) );
  NAND2_X1 U14000 ( .A1(n10670), .A2(n10662), .ZN(n10663) );
  NAND2_X1 U14001 ( .A1(n10664), .A2(n10663), .ZN(n11916) );
  INV_X1 U14002 ( .A(n10665), .ZN(n10666) );
  XNOR2_X1 U14003 ( .A(n10667), .B(n10666), .ZN(n11914) );
  INV_X1 U14004 ( .A(n11914), .ZN(n10668) );
  OAI21_X1 U14005 ( .B1(n11908), .B2(n11907), .A(n10669), .ZN(n10674) );
  NAND2_X1 U14006 ( .A1(n10670), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10672) );
  NAND2_X1 U14007 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20089), .ZN(n10675) );
  AOI211_X4 U14008 ( .C1(n17849), .C2(n20083), .A(n10677), .B(n10675), .ZN(
        n18171) );
  INV_X1 U14009 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18181) );
  NAND2_X1 U14010 ( .A1(n18194), .A2(n18181), .ZN(n18170) );
  NOR2_X1 U14011 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18170), .ZN(n18149) );
  NAND2_X1 U14012 ( .A1(n18149), .A2(n18155), .ZN(n18148) );
  NAND2_X1 U14013 ( .A1(n18133), .A2(n18123), .ZN(n18122) );
  INV_X1 U14014 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18097) );
  NAND2_X1 U14015 ( .A1(n18108), .A2(n18097), .ZN(n18096) );
  NAND2_X1 U14016 ( .A1(n18086), .A2(n21456), .ZN(n18074) );
  NAND2_X1 U14017 ( .A1(n18061), .A2(n18050), .ZN(n18049) );
  NAND2_X1 U14018 ( .A1(n18031), .A2(n18514), .ZN(n18022) );
  INV_X1 U14019 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21723) );
  NAND2_X1 U14020 ( .A1(n18014), .A2(n21723), .ZN(n18001) );
  INV_X1 U14021 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17981) );
  NAND2_X1 U14022 ( .A1(n17989), .A2(n17981), .ZN(n17979) );
  INV_X1 U14023 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18419) );
  NAND2_X1 U14024 ( .A1(n17970), .A2(n18419), .ZN(n17963) );
  INV_X1 U14025 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17943) );
  NAND2_X1 U14026 ( .A1(n17951), .A2(n17943), .ZN(n17942) );
  NAND2_X1 U14027 ( .A1(n17913), .A2(n17924), .ZN(n17903) );
  INV_X1 U14028 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17898) );
  NAND2_X1 U14029 ( .A1(n17902), .A2(n17898), .ZN(n17897) );
  INV_X1 U14030 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17868) );
  NAND2_X1 U14031 ( .A1(n17881), .A2(n17868), .ZN(n13368) );
  NOR2_X1 U14032 ( .A1(n18226), .A2(n13368), .ZN(n13370) );
  INV_X1 U14033 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18228) );
  AND2_X1 U14034 ( .A1(n13370), .A2(n18228), .ZN(n10690) );
  INV_X1 U14035 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20001) );
  NAND2_X2 U14036 ( .A1(n20101), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n20062) );
  OAI211_X1 U14037 ( .C1(n20088), .C2(n20089), .A(n20083), .B(n17849), .ZN(
        n19968) );
  INV_X1 U14038 ( .A(n19968), .ZN(n10676) );
  AOI211_X4 U14039 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20089), .A(n10676), .B(
        n10677), .ZN(n18217) );
  INV_X1 U14040 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20061) );
  INV_X1 U14041 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20050) );
  INV_X1 U14042 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20044) );
  INV_X1 U14043 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20027) );
  INV_X1 U14044 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20024) );
  INV_X1 U14045 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20006) );
  NAND2_X1 U14046 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_3__SCAN_IN), 
        .ZN(n18157) );
  NOR2_X1 U14047 ( .A1(n20006), .A2(n18157), .ZN(n18168) );
  NAND3_X1 U14048 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .A3(n18168), .ZN(n18088) );
  NAND3_X1 U14049 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n18069) );
  NAND2_X1 U14050 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n18070) );
  NOR4_X1 U14051 ( .A1(n20020), .A2(n18088), .A3(n18069), .A4(n18070), .ZN(
        n18065) );
  NAND2_X1 U14052 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18065), .ZN(n18030) );
  NOR3_X1 U14053 ( .A1(n20027), .A2(n20024), .A3(n18030), .ZN(n17949) );
  INV_X1 U14054 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20040) );
  NAND3_X1 U14055 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n17985) );
  NAND2_X1 U14056 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17986) );
  NOR2_X1 U14057 ( .A1(n17985), .A2(n17986), .ZN(n17974) );
  NAND2_X1 U14058 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17974), .ZN(n17950) );
  NOR2_X1 U14059 ( .A1(n20040), .A2(n17950), .ZN(n17948) );
  NAND3_X1 U14060 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17949), .A3(n17948), 
        .ZN(n17939) );
  NOR2_X1 U14061 ( .A1(n20044), .A2(n17939), .ZN(n17937) );
  NAND2_X1 U14062 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17937), .ZN(n17916) );
  NOR2_X1 U14063 ( .A1(n20048), .A2(n17916), .ZN(n10683) );
  NAND2_X1 U14064 ( .A1(n18169), .A2(n10683), .ZN(n17912) );
  NAND4_X1 U14065 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17880), .ZN(n10685) );
  NOR3_X1 U14066 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20061), .A3(n10685), 
        .ZN(n10678) );
  AOI21_X1 U14067 ( .B1(n18217), .B2(P3_EBX_REG_31__SCAN_IN), .A(n10678), .ZN(
        n10682) );
  INV_X1 U14068 ( .A(n19978), .ZN(n19865) );
  NOR2_X1 U14069 ( .A1(n19980), .A2(n19865), .ZN(n19973) );
  NOR2_X1 U14070 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n10679) );
  AND2_X2 U14071 ( .A1(n20103), .A2(n10679), .ZN(n19477) );
  OR2_X1 U14072 ( .A1(n18189), .A2(n19477), .ZN(n10680) );
  OR2_X1 U14073 ( .A1(n19973), .A2(n10680), .ZN(n10681) );
  INV_X1 U14074 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17437) );
  NAND3_X1 U14075 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n10684) );
  OAI221_X1 U14076 ( .B1(n18205), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n18205), 
        .C2(n10683), .A(n18212), .ZN(n17909) );
  AOI21_X1 U14077 ( .B1(n18156), .B2(n10684), .A(n17909), .ZN(n17873) );
  NOR2_X1 U14078 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n10685), .ZN(n13374) );
  INV_X1 U14079 ( .A(n13374), .ZN(n10686) );
  INV_X1 U14080 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20059) );
  AOI21_X1 U14081 ( .B1(n17873), .B2(n10686), .A(n20059), .ZN(n10687) );
  INV_X1 U14084 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10693) );
  INV_X1 U14085 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10694) );
  INV_X4 U14086 ( .A(n10846), .ZN(n11697) );
  AOI22_X1 U14087 ( .A1(n10837), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10700) );
  AND2_X2 U14088 ( .A1(n10695), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15001) );
  AND2_X2 U14089 ( .A1(n15001), .A2(n10703), .ZN(n10973) );
  NAND2_X2 U14090 ( .A1(n10703), .A2(n10701), .ZN(n10833) );
  AOI22_X1 U14091 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10923), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10699) );
  AND2_X2 U14092 ( .A1(n14997), .A2(n10696), .ZN(n11528) );
  AOI22_X1 U14093 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10698) );
  NOR2_X4 U14094 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U14095 ( .A1(n10818), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U14096 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11004), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10707) );
  AND2_X2 U14097 ( .A1(n15001), .A2(n15011), .ZN(n11012) );
  AOI22_X1 U14098 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11623), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U14099 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10705) );
  AND2_X2 U14100 ( .A1(n10703), .A2(n10702), .ZN(n10931) );
  AOI22_X1 U14101 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U14102 ( .A1(n10923), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10713) );
  NAND2_X1 U14103 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U14104 ( .A1(n10837), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U14105 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10718) );
  NAND2_X1 U14106 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U14107 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10716) );
  NAND2_X1 U14108 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10715) );
  NAND2_X1 U14109 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U14110 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U14111 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10720) );
  NAND2_X1 U14112 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10719) );
  INV_X2 U14113 ( .A(n10723), .ZN(n11690) );
  NAND2_X1 U14114 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10727) );
  NAND2_X1 U14115 ( .A1(n10931), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10726) );
  NAND2_X1 U14116 ( .A1(n10818), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10725) );
  NAND2_X1 U14117 ( .A1(n10960), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10724) );
  NAND2_X1 U14119 ( .A1(n10881), .A2(n14697), .ZN(n10740) );
  AOI22_X1 U14120 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10818), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U14121 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U14122 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U14123 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U14124 ( .A1(n10923), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U14125 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U14126 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U14127 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10736) );
  NAND2_X4 U14128 ( .A1(n9752), .A2(n10480), .ZN(n14691) );
  NAND2_X1 U14129 ( .A1(n10740), .A2(n14287), .ZN(n10779) );
  NAND2_X1 U14130 ( .A1(n13032), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U14131 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10744) );
  NAND2_X1 U14132 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10743) );
  NAND2_X1 U14133 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10742) );
  NAND2_X1 U14134 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10741) );
  NAND2_X1 U14135 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U14136 ( .A1(n10837), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10747) );
  NAND2_X1 U14137 ( .A1(n10923), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10746) );
  NAND2_X1 U14138 ( .A1(n11623), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10745) );
  NAND2_X1 U14139 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10752) );
  NAND2_X1 U14140 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U14141 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10750) );
  NAND2_X1 U14142 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10749) );
  NAND2_X1 U14143 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10756) );
  NAND2_X1 U14144 ( .A1(n10931), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U14145 ( .A1(n10818), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10754) );
  NAND2_X1 U14146 ( .A1(n10960), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10753) );
  NAND2_X1 U14147 ( .A1(n16294), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10762) );
  NAND2_X1 U14148 ( .A1(n14983), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U14149 ( .A1(n10762), .A2(n10761), .ZN(n10771) );
  NAND2_X1 U14150 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21271), .ZN(
        n10774) );
  NAND2_X1 U14151 ( .A1(n15029), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U14152 ( .A1(n14992), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10763) );
  NAND2_X1 U14153 ( .A1(n10791), .A2(n10763), .ZN(n10765) );
  NAND2_X1 U14154 ( .A1(n10764), .A2(n10765), .ZN(n10768) );
  INV_X1 U14155 ( .A(n10765), .ZN(n10766) );
  NAND2_X1 U14156 ( .A1(n10767), .A2(n10766), .ZN(n10792) );
  NAND2_X1 U14157 ( .A1(n10768), .A2(n10792), .ZN(n13002) );
  MUX2_X1 U14158 ( .A(n11133), .B(n11132), .S(n13002), .Z(n10786) );
  NAND2_X1 U14159 ( .A1(n11133), .A2(n14691), .ZN(n10770) );
  NAND2_X1 U14160 ( .A1(n10881), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10769) );
  NAND2_X1 U14161 ( .A1(n10770), .A2(n10769), .ZN(n10781) );
  NAND2_X1 U14162 ( .A1(n10038), .A2(n14691), .ZN(n10798) );
  NAND2_X1 U14163 ( .A1(n10771), .A2(n10774), .ZN(n10772) );
  NAND2_X1 U14164 ( .A1(n10773), .A2(n10772), .ZN(n13003) );
  INV_X1 U14165 ( .A(n13003), .ZN(n10784) );
  NAND2_X1 U14166 ( .A1(n10781), .A2(n10784), .ZN(n10783) );
  OAI21_X1 U14167 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21271), .A(
        n10774), .ZN(n10775) );
  INV_X1 U14168 ( .A(n10775), .ZN(n10778) );
  NAND2_X1 U14169 ( .A1(n11133), .A2(n10778), .ZN(n10776) );
  OAI211_X1 U14170 ( .C1(n10864), .C2(n13032), .A(n10779), .B(n10778), .ZN(
        n10780) );
  OAI211_X1 U14171 ( .C1(n10798), .C2(n10784), .A(n10783), .B(n10782), .ZN(
        n10785) );
  OAI21_X1 U14172 ( .B1(n10788), .B2(n10786), .A(n10785), .ZN(n10790) );
  INV_X1 U14173 ( .A(n13002), .ZN(n10787) );
  NAND3_X1 U14174 ( .A1(n10788), .A2(n10787), .A3(n11133), .ZN(n10789) );
  NAND2_X1 U14175 ( .A1(n10790), .A2(n10789), .ZN(n10802) );
  NAND2_X1 U14176 ( .A1(n10792), .A2(n10791), .ZN(n10795) );
  XNOR2_X1 U14177 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10794) );
  AND2_X1 U14178 ( .A1(n15015), .A2(n10800), .ZN(n10793) );
  NOR2_X1 U14179 ( .A1(n10795), .A2(n10794), .ZN(n10796) );
  INV_X1 U14180 ( .A(n11146), .ZN(n13783) );
  OAI22_X1 U14181 ( .A1(n10798), .A2(n13005), .B1(n10801), .B2(n13783), .ZN(
        n10799) );
  OAI21_X1 U14182 ( .B1(n10802), .B2(n10799), .A(n11132), .ZN(n10804) );
  AOI222_X1 U14183 ( .A1(n10800), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n10800), .B2(n15015), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n15015), .ZN(n13006) );
  NAND3_X1 U14184 ( .A1(n10802), .A2(n10801), .A3(n13005), .ZN(n10803) );
  INV_X1 U14185 ( .A(n10805), .ZN(n10806) );
  NAND2_X1 U14186 ( .A1(n13006), .A2(n10806), .ZN(n10807) );
  AOI22_X1 U14187 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U14188 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10818), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U14189 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U14190 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U14191 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U14192 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10815) );
  INV_X2 U14193 ( .A(n10830), .ZN(n10903) );
  NAND2_X2 U14194 ( .A1(n10903), .A2(n15557), .ZN(n10829) );
  INV_X1 U14195 ( .A(n10829), .ZN(n10828) );
  AOI22_X1 U14196 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11004), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U14197 ( .A1(n10931), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U14198 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10818), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U14199 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U14200 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U14201 ( .A1(n10837), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10923), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U14202 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U14203 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U14204 ( .A1(n10828), .A2(n10827), .ZN(n10870) );
  INV_X1 U14205 ( .A(n10829), .ZN(n10873) );
  NAND2_X1 U14206 ( .A1(n10873), .A2(n13409), .ZN(n10832) );
  NAND2_X1 U14207 ( .A1(n10881), .A2(n10879), .ZN(n10831) );
  INV_X1 U14208 ( .A(n10895), .ZN(n10860) );
  INV_X1 U14209 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10997) );
  INV_X1 U14210 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10835) );
  OAI22_X1 U14211 ( .A1(n10833), .A2(n10997), .B1(n11650), .B2(n10835), .ZN(
        n10836) );
  INV_X1 U14212 ( .A(n10836), .ZN(n10841) );
  AOI22_X1 U14213 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U14214 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U14215 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U14216 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10818), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U14217 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U14218 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U14219 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10842) );
  INV_X1 U14220 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10848) );
  INV_X1 U14221 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10847) );
  OAI22_X1 U14222 ( .A1(n10846), .A2(n10848), .B1(n11650), .B2(n10847), .ZN(
        n10849) );
  INV_X1 U14223 ( .A(n10849), .ZN(n10853) );
  AOI22_X1 U14224 ( .A1(n10923), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11012), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U14225 ( .A1(n11004), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U14226 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10818), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10850) );
  NAND4_X1 U14227 ( .A1(n10853), .A2(n10852), .A3(n10851), .A4(n10850), .ZN(
        n10859) );
  AOI22_X1 U14228 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U14229 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U14230 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U14231 ( .A1(n10837), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10854) );
  NAND4_X1 U14232 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10858) );
  OAI211_X1 U14233 ( .C1(n13146), .C2(n14697), .A(n10860), .B(n10015), .ZN(
        n13018) );
  OR2_X1 U14234 ( .A1(n13018), .A2(n10864), .ZN(n13026) );
  INV_X1 U14235 ( .A(n10878), .ZN(n10862) );
  NAND2_X1 U14236 ( .A1(n14090), .A2(n10883), .ZN(n14974) );
  NAND2_X1 U14237 ( .A1(n10862), .A2(n14974), .ZN(n10863) );
  NOR2_X1 U14238 ( .A1(n10895), .A2(n10863), .ZN(n10876) );
  NAND2_X1 U14239 ( .A1(n15557), .A2(n10879), .ZN(n10865) );
  OAI21_X1 U14240 ( .B1(n10868), .B2(n10879), .A(n14057), .ZN(n10869) );
  NAND2_X1 U14241 ( .A1(n10872), .A2(n10871), .ZN(n10894) );
  NAND2_X1 U14242 ( .A1(n10894), .A2(n13032), .ZN(n10875) );
  NAND2_X1 U14243 ( .A1(n13032), .A2(n14691), .ZN(n15466) );
  NAND2_X1 U14244 ( .A1(n10873), .A2(n14283), .ZN(n13016) );
  NAND2_X1 U14245 ( .A1(n13016), .A2(n14051), .ZN(n10874) );
  NAND4_X1 U14246 ( .A1(n10876), .A2(n10875), .A3(n10901), .A4(n10874), .ZN(
        n10877) );
  NAND2_X1 U14247 ( .A1(n10877), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10888) );
  NOR2_X2 U14248 ( .A1(n10883), .A2(n14691), .ZN(n10898) );
  NAND2_X1 U14249 ( .A1(n13134), .A2(n10898), .ZN(n10880) );
  OAI21_X1 U14250 ( .B1(n10894), .B2(n10880), .A(n13027), .ZN(n10887) );
  NAND4_X1 U14251 ( .A1(n10903), .A2(n13409), .A3(n10881), .A4(n14057), .ZN(
        n10882) );
  XNOR2_X1 U14252 ( .A(n21357), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U14253 ( .B1(n10887), .B2(n10886), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10891) );
  NAND2_X1 U14254 ( .A1(n10888), .A2(n10891), .ZN(n10910) );
  NAND2_X1 U14255 ( .A1(n10910), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10890) );
  NAND2_X1 U14256 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10913) );
  OAI21_X1 U14257 ( .B1(n11720), .B2(n16164), .A(n10906), .ZN(n10889) );
  NAND2_X1 U14258 ( .A1(n10910), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10893) );
  MUX2_X1 U14259 ( .A(n11720), .B(n17620), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10892) );
  NAND2_X1 U14260 ( .A1(n10894), .A2(n10898), .ZN(n10897) );
  NAND2_X1 U14261 ( .A1(n10895), .A2(n14691), .ZN(n10896) );
  INV_X1 U14262 ( .A(n10898), .ZN(n15477) );
  AND2_X1 U14263 ( .A1(n15477), .A2(n13196), .ZN(n15197) );
  NAND2_X1 U14264 ( .A1(n10829), .A2(n14045), .ZN(n10899) );
  NAND3_X1 U14265 ( .A1(n13016), .A2(n14697), .A3(n14051), .ZN(n10900) );
  INV_X1 U14266 ( .A(n13013), .ZN(n10902) );
  INV_X2 U14267 ( .A(n14283), .ZN(n11047) );
  NAND2_X1 U14268 ( .A1(n15092), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21092) );
  AOI21_X1 U14269 ( .B1(n10902), .B2(n11047), .A(n21092), .ZN(n10905) );
  INV_X1 U14270 ( .A(n14974), .ZN(n10904) );
  AOI21_X1 U14271 ( .B1(n10878), .B2(n10903), .A(n10904), .ZN(n13139) );
  INV_X1 U14272 ( .A(n10906), .ZN(n10908) );
  OAI21_X1 U14273 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n10908), .A(
        n10907), .ZN(n10909) );
  NAND2_X1 U14274 ( .A1(n10911), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10918) );
  INV_X1 U14275 ( .A(n11720), .ZN(n10916) );
  INV_X1 U14276 ( .A(n10913), .ZN(n10912) );
  NAND2_X1 U14277 ( .A1(n10912), .A2(n15029), .ZN(n14535) );
  NAND2_X1 U14278 ( .A1(n10913), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10914) );
  NAND2_X1 U14279 ( .A1(n14535), .A2(n10914), .ZN(n14443) );
  INV_X1 U14280 ( .A(n17620), .ZN(n10915) );
  AOI22_X1 U14281 ( .A1(n10916), .A2(n14443), .B1(n10915), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U14282 ( .A1(n10918), .A2(n10917), .ZN(n10996) );
  NAND2_X1 U14283 ( .A1(n10911), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10922) );
  NAND2_X1 U14284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16251), .ZN(
        n14155) );
  NAND2_X1 U14285 ( .A1(n17600), .A2(n14155), .ZN(n10919) );
  NAND3_X1 U14286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16386) );
  INV_X1 U14287 ( .A(n16386), .ZN(n16383) );
  NAND2_X1 U14288 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16383), .ZN(
        n16381) );
  NAND2_X1 U14289 ( .A1(n10919), .A2(n16381), .ZN(n16121) );
  OAI22_X1 U14290 ( .A1(n11720), .A2(n16121), .B1(n17620), .B2(n17600), .ZN(
        n10920) );
  INV_X1 U14291 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U14292 ( .A1(n14028), .A2(n21654), .ZN(n10939) );
  AOI22_X1 U14293 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U14294 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10929) );
  INV_X1 U14295 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10925) );
  INV_X1 U14296 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10924) );
  OAI22_X1 U14297 ( .A1(n11652), .A2(n10925), .B1(n11650), .B2(n10924), .ZN(
        n10926) );
  INV_X1 U14298 ( .A(n10926), .ZN(n10928) );
  AOI22_X1 U14299 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U14300 ( .A1(n10930), .A2(n10929), .A3(n10928), .A4(n10927), .ZN(
        n10937) );
  AOI22_X1 U14301 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10935) );
  INV_X1 U14302 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n21619) );
  AOI22_X1 U14303 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10934) );
  INV_X2 U14304 ( .A(n10723), .ZN(n11413) );
  AOI22_X1 U14305 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10933) );
  BUF_X1 U14306 ( .A(n11528), .Z(n11692) );
  AOI22_X1 U14307 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10932) );
  NAND4_X1 U14308 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10932), .ZN(
        n10936) );
  AOI22_X1 U14309 ( .A1(n11133), .A2(n11055), .B1(n11132), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U14310 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14311 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14312 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14313 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U14314 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10954) );
  AOI22_X1 U14315 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10952) );
  INV_X1 U14316 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10947) );
  INV_X1 U14317 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10946) );
  OAI22_X1 U14318 ( .A1(n9722), .A2(n10947), .B1(n10833), .B2(n10946), .ZN(
        n10948) );
  INV_X1 U14319 ( .A(n10948), .ZN(n10951) );
  AOI22_X1 U14320 ( .A1(n11700), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14321 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10949) );
  NAND4_X1 U14322 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n10953) );
  NAND2_X1 U14323 ( .A1(n10984), .A2(n11084), .ZN(n10955) );
  AOI22_X1 U14324 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14325 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14326 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14327 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14328 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10967) );
  AOI22_X1 U14329 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U14330 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U14331 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U14332 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U14333 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10966) );
  INV_X1 U14334 ( .A(n11150), .ZN(n10980) );
  AOI22_X1 U14335 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11606), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14336 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11413), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U14337 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11701), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14338 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11533), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U14339 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10979) );
  AOI22_X1 U14340 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11699), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14341 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U14342 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11700), .B1(
        n10960), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14343 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n11629), .ZN(n10974) );
  NAND4_X1 U14344 ( .A1(n10977), .A2(n10976), .A3(n10975), .A4(n10974), .ZN(
        n10978) );
  XNOR2_X1 U14345 ( .A(n10980), .B(n11085), .ZN(n10981) );
  NAND2_X1 U14346 ( .A1(n10981), .A2(n10984), .ZN(n11071) );
  AOI21_X1 U14347 ( .B1(n13032), .B2(n11085), .A(n21654), .ZN(n11075) );
  AOI21_X1 U14348 ( .B1(n11071), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11075), 
        .ZN(n10982) );
  NAND2_X1 U14349 ( .A1(n10983), .A2(n10982), .ZN(n10986) );
  NAND2_X1 U14350 ( .A1(n10984), .A2(n11150), .ZN(n10985) );
  NAND2_X1 U14351 ( .A1(n10986), .A2(n10985), .ZN(n10993) );
  NAND2_X1 U14352 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10990) );
  INV_X1 U14353 ( .A(n10987), .ZN(n10988) );
  NAND2_X1 U14354 ( .A1(n10988), .A2(n11084), .ZN(n10989) );
  OAI211_X1 U14355 ( .C1(n10991), .C2(n11150), .A(n10990), .B(n10989), .ZN(
        n10992) );
  NAND2_X1 U14356 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  AOI22_X1 U14357 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14358 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11002) );
  INV_X1 U14359 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10998) );
  OAI22_X1 U14360 ( .A1(n11652), .A2(n10998), .B1(n11650), .B2(n10997), .ZN(
        n10999) );
  INV_X1 U14361 ( .A(n10999), .ZN(n11001) );
  AOI22_X1 U14362 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11000) );
  NAND4_X1 U14363 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11010) );
  AOI22_X1 U14364 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14365 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U14366 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14367 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11005) );
  NAND4_X1 U14368 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n11009) );
  AOI22_X1 U14369 ( .A1(n11133), .A2(n11045), .B1(n11132), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U14370 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14371 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11018) );
  INV_X1 U14372 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11014) );
  INV_X1 U14373 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11013) );
  OAI22_X1 U14374 ( .A1(n11652), .A2(n11014), .B1(n11650), .B2(n11013), .ZN(
        n11015) );
  INV_X1 U14375 ( .A(n11015), .ZN(n11017) );
  AOI22_X1 U14376 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U14377 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11025) );
  AOI22_X1 U14378 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14379 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11022) );
  AOI22_X1 U14380 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14381 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11020) );
  NAND4_X1 U14382 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11024) );
  AOI22_X1 U14383 ( .A1(n11133), .A2(n11062), .B1(n11132), .B2(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14384 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14385 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11032) );
  INV_X1 U14386 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11028) );
  INV_X1 U14387 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11027) );
  OAI22_X1 U14388 ( .A1(n11652), .A2(n11028), .B1(n11650), .B2(n11027), .ZN(
        n11029) );
  INV_X1 U14389 ( .A(n11029), .ZN(n11031) );
  INV_X1 U14390 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14391 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11030) );
  NAND4_X1 U14392 ( .A1(n11033), .A2(n11032), .A3(n11031), .A4(n11030), .ZN(
        n11039) );
  AOI22_X1 U14393 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14394 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14395 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14396 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11034) );
  NAND4_X1 U14397 ( .A1(n11037), .A2(n11036), .A3(n11035), .A4(n11034), .ZN(
        n11038) );
  NAND2_X1 U14398 ( .A1(n11133), .A2(n11048), .ZN(n11041) );
  NAND2_X1 U14399 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14400 ( .A1(n11041), .A2(n11040), .ZN(n11043) );
  NAND2_X1 U14401 ( .A1(n11061), .A2(n10232), .ZN(n11044) );
  NAND2_X1 U14402 ( .A1(n11085), .A2(n11084), .ZN(n11100) );
  INV_X1 U14403 ( .A(n11045), .ZN(n11101) );
  NAND2_X1 U14404 ( .A1(n11100), .A2(n11101), .ZN(n11099) );
  NAND2_X1 U14405 ( .A1(n11099), .A2(n11055), .ZN(n11063) );
  INV_X1 U14406 ( .A(n11062), .ZN(n11046) );
  NOR2_X1 U14407 ( .A1(n11063), .A2(n11046), .ZN(n11049) );
  NAND2_X1 U14408 ( .A1(n11049), .A2(n11048), .ZN(n11138) );
  OAI211_X1 U14409 ( .C1(n11049), .C2(n11048), .A(n11138), .B(n11047), .ZN(
        n11050) );
  INV_X1 U14410 ( .A(n11113), .ZN(n17662) );
  NAND2_X1 U14411 ( .A1(n17662), .A2(n17695), .ZN(n11109) );
  NAND2_X1 U14412 ( .A1(n14024), .A2(n11146), .ZN(n11057) );
  OAI211_X1 U14413 ( .C1(n11055), .C2(n11099), .A(n11063), .B(n11047), .ZN(
        n11056) );
  NAND2_X1 U14414 ( .A1(n11057), .A2(n11056), .ZN(n14374) );
  NAND2_X1 U14415 ( .A1(n11059), .A2(n11058), .ZN(n11060) );
  NAND2_X1 U14416 ( .A1(n11214), .A2(n11146), .ZN(n11066) );
  XNOR2_X1 U14417 ( .A(n11063), .B(n11062), .ZN(n11064) );
  NAND2_X1 U14418 ( .A1(n11064), .A2(n11047), .ZN(n11065) );
  AND2_X2 U14419 ( .A1(n11066), .A2(n11065), .ZN(n17660) );
  INV_X1 U14420 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17658) );
  NAND2_X1 U14421 ( .A1(n17660), .A2(n17658), .ZN(n11067) );
  INV_X1 U14422 ( .A(n11069), .ZN(n11070) );
  NAND2_X1 U14423 ( .A1(n11072), .A2(n11071), .ZN(n11077) );
  NAND2_X1 U14424 ( .A1(n11132), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U14425 ( .A1(n13409), .A2(n11150), .ZN(n11073) );
  NAND3_X1 U14426 ( .A1(n11075), .A2(n11074), .A3(n11073), .ZN(n11076) );
  OR2_X1 U14427 ( .A1(n14283), .A2(n11085), .ZN(n13784) );
  INV_X1 U14428 ( .A(n13784), .ZN(n11079) );
  NAND2_X1 U14429 ( .A1(n13032), .A2(n14045), .ZN(n13785) );
  NOR2_X1 U14430 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  AND2_X1 U14431 ( .A1(n13783), .A2(n13785), .ZN(n11081) );
  INV_X1 U14432 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15090) );
  AOI21_X1 U14433 ( .B1(n11081), .B2(n13784), .A(n15090), .ZN(n11082) );
  XNOR2_X1 U14434 ( .A(n11085), .B(n11084), .ZN(n11087) );
  OAI211_X1 U14435 ( .C1(n11087), .C2(n14283), .A(n11086), .B(n15557), .ZN(
        n11088) );
  INV_X1 U14436 ( .A(n11088), .ZN(n11089) );
  INV_X1 U14437 ( .A(n13788), .ZN(n11092) );
  NAND2_X1 U14438 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  INV_X1 U14439 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13041) );
  INV_X1 U14440 ( .A(n11094), .ZN(n11096) );
  NAND2_X1 U14441 ( .A1(n11096), .A2(n11095), .ZN(n11098) );
  NAND2_X1 U14442 ( .A1(n11098), .A2(n11097), .ZN(n11176) );
  OAI21_X1 U14443 ( .B1(n11101), .B2(n11100), .A(n11099), .ZN(n11102) );
  AOI21_X1 U14444 ( .B1(n11102), .B2(n11047), .A(n11078), .ZN(n11103) );
  OAI21_X1 U14445 ( .B1(n11176), .B2(n13783), .A(n11103), .ZN(n13868) );
  AND2_X1 U14446 ( .A1(n11104), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11105) );
  NAND2_X1 U14447 ( .A1(n14374), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11106) );
  AND2_X1 U14448 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11111) );
  INV_X1 U14449 ( .A(n17660), .ZN(n11110) );
  AOI22_X1 U14450 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14451 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14452 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14453 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11115) );
  NAND4_X1 U14454 ( .A1(n11118), .A2(n11117), .A3(n11116), .A4(n11115), .ZN(
        n11124) );
  AOI22_X1 U14455 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14456 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14457 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11120) );
  AOI22_X1 U14458 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11119) );
  NAND4_X1 U14459 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(
        n11123) );
  AOI22_X1 U14460 ( .A1(n11133), .A2(n11139), .B1(n11132), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11125) );
  NAND3_X1 U14461 ( .A1(n11148), .A2(n11226), .A3(n11146), .ZN(n11129) );
  XNOR2_X1 U14462 ( .A(n11138), .B(n11139), .ZN(n11127) );
  NAND2_X1 U14463 ( .A1(n11127), .A2(n11047), .ZN(n11128) );
  NAND2_X1 U14464 ( .A1(n11129), .A2(n11128), .ZN(n11130) );
  INV_X1 U14465 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21461) );
  XNOR2_X1 U14466 ( .A(n11130), .B(n21461), .ZN(n14423) );
  OR2_X1 U14467 ( .A1(n11130), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11131) );
  INV_X1 U14468 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11136) );
  INV_X1 U14469 ( .A(n11132), .ZN(n11135) );
  NAND2_X1 U14470 ( .A1(n11133), .A2(n11150), .ZN(n11134) );
  OAI21_X1 U14471 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n11137) );
  NAND2_X1 U14472 ( .A1(n11233), .A2(n11146), .ZN(n11143) );
  INV_X1 U14473 ( .A(n11138), .ZN(n11140) );
  NAND2_X1 U14474 ( .A1(n11140), .A2(n11139), .ZN(n11149) );
  XNOR2_X1 U14475 ( .A(n11149), .B(n11150), .ZN(n11141) );
  NAND2_X1 U14476 ( .A1(n11141), .A2(n11047), .ZN(n11142) );
  INV_X1 U14477 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17690) );
  OR2_X1 U14478 ( .A1(n11144), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11145) );
  INV_X1 U14479 ( .A(n11149), .ZN(n11151) );
  NAND3_X1 U14480 ( .A1(n11151), .A2(n11047), .A3(n11150), .ZN(n11152) );
  NAND2_X1 U14481 ( .A1(n15831), .A2(n11152), .ZN(n11153) );
  NAND2_X1 U14482 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U14483 ( .A1(n15831), .A2(n11154), .ZN(n11160) );
  INV_X1 U14484 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16010) );
  NAND2_X1 U14485 ( .A1(n15831), .A2(n16010), .ZN(n11155) );
  NAND2_X1 U14486 ( .A1(n15801), .A2(n11155), .ZN(n15816) );
  INV_X1 U14487 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U14488 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U14489 ( .A1(n15831), .A2(n11156), .ZN(n15811) );
  NAND2_X1 U14490 ( .A1(n15822), .A2(n15811), .ZN(n11157) );
  INV_X1 U14491 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U14492 ( .A1(n15729), .A2(n15970), .ZN(n11158) );
  NAND2_X1 U14493 ( .A1(n15664), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11159) );
  NAND2_X1 U14494 ( .A1(n11159), .A2(n15801), .ZN(n11161) );
  XNOR2_X1 U14495 ( .A(n15729), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15784) );
  INV_X1 U14496 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16007) );
  NAND2_X1 U14497 ( .A1(n15831), .A2(n16007), .ZN(n15794) );
  INV_X1 U14498 ( .A(n11161), .ZN(n11163) );
  NOR2_X1 U14499 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11162) );
  OR2_X1 U14500 ( .A1(n15729), .A2(n11162), .ZN(n15812) );
  INV_X1 U14501 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15771) );
  INV_X1 U14502 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15983) );
  NAND3_X1 U14503 ( .A1(n16007), .A2(n15771), .A3(n15983), .ZN(n11164) );
  NAND2_X1 U14504 ( .A1(n15840), .A2(n11164), .ZN(n11165) );
  INV_X1 U14505 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16069) );
  NAND2_X1 U14506 ( .A1(n11165), .A2(n15766), .ZN(n11166) );
  NOR2_X1 U14507 ( .A1(n15780), .A2(n11166), .ZN(n11167) );
  XNOR2_X1 U14508 ( .A(n15729), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15757) );
  AND2_X1 U14509 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15943) );
  INV_X1 U14510 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15947) );
  INV_X1 U14511 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15938) );
  INV_X1 U14512 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15946) );
  NAND3_X1 U14513 ( .A1(n15947), .A2(n15938), .A3(n15946), .ZN(n11168) );
  NAND3_X1 U14514 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15891) );
  INV_X1 U14515 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15690) );
  NOR2_X1 U14516 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15661) );
  INV_X1 U14517 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15677) );
  INV_X1 U14518 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U14519 ( .A1(n15677), .A2(n13123), .ZN(n15872) );
  INV_X1 U14520 ( .A(n15872), .ZN(n11170) );
  NAND2_X1 U14521 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15871) );
  NAND2_X1 U14522 ( .A1(n13191), .A2(n13192), .ZN(n11171) );
  XNOR2_X1 U14523 ( .A(n11171), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13174) );
  NAND2_X1 U14524 ( .A1(n13417), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11207) );
  INV_X1 U14525 ( .A(n11207), .ZN(n11202) );
  INV_X1 U14526 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11173) );
  XNOR2_X1 U14527 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15481) );
  AOI21_X1 U14528 ( .B1(n11190), .B2(n15481), .A(n13405), .ZN(n11172) );
  OAI21_X1 U14529 ( .B1(n11711), .B2(n11173), .A(n11172), .ZN(n11174) );
  AOI21_X1 U14530 ( .B1(n11202), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11174), .ZN(n11175) );
  NAND2_X1 U14531 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11194) );
  NAND2_X1 U14532 ( .A1(n11177), .A2(n11194), .ZN(n13973) );
  INV_X1 U14533 ( .A(n13973), .ZN(n11193) );
  NAND2_X1 U14534 ( .A1(n11179), .A2(n11178), .ZN(n11180) );
  NAND2_X1 U14535 ( .A1(n16079), .A2(n11383), .ZN(n11184) );
  INV_X1 U14536 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15485) );
  OAI22_X1 U14537 ( .A1(n11711), .A2(n21217), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15485), .ZN(n11182) );
  AOI21_X1 U14538 ( .B1(n11202), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11182), .ZN(n11183) );
  NAND2_X1 U14539 ( .A1(n9720), .A2(n10903), .ZN(n11185) );
  NAND2_X1 U14540 ( .A1(n11185), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13780) );
  NAND2_X1 U14541 ( .A1(n13406), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11187) );
  NAND2_X1 U14542 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11186) );
  OAI211_X1 U14543 ( .C1(n11207), .C2(n15095), .A(n11187), .B(n11186), .ZN(
        n11188) );
  OR2_X1 U14544 ( .A1(n10104), .A2(n11715), .ZN(n13795) );
  NAND2_X1 U14545 ( .A1(n13796), .A2(n13795), .ZN(n11191) );
  NAND2_X1 U14546 ( .A1(n13794), .A2(n11191), .ZN(n13972) );
  INV_X1 U14547 ( .A(n13972), .ZN(n11192) );
  NAND2_X1 U14548 ( .A1(n11193), .A2(n11192), .ZN(n13970) );
  NAND2_X1 U14549 ( .A1(n14024), .A2(n11383), .ZN(n11204) );
  INV_X1 U14550 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U14551 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11196) );
  INV_X1 U14552 ( .A(n11196), .ZN(n11195) );
  INV_X1 U14553 ( .A(n11208), .ZN(n11210) );
  INV_X1 U14554 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U14555 ( .A1(n11197), .A2(n11196), .ZN(n11198) );
  NAND2_X1 U14556 ( .A1(n11210), .A2(n11198), .ZN(n21183) );
  AOI22_X1 U14557 ( .A1(n21183), .A2(n14683), .B1(n13405), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11199) );
  OAI21_X1 U14558 ( .B1(n11711), .B2(n11200), .A(n11199), .ZN(n11201) );
  AOI21_X1 U14559 ( .B1(n11202), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11201), .ZN(n11203) );
  NAND2_X1 U14560 ( .A1(n11204), .A2(n11203), .ZN(n13962) );
  NAND2_X1 U14561 ( .A1(n13963), .A2(n13962), .ZN(n13961) );
  INV_X1 U14562 ( .A(n13961), .ZN(n11216) );
  NAND2_X1 U14563 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U14564 ( .A1(n13406), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11205) );
  OAI211_X1 U14565 ( .C1(n11207), .C2(n15015), .A(n11206), .B(n11205), .ZN(
        n11212) );
  INV_X1 U14566 ( .A(n11217), .ZN(n11218) );
  INV_X1 U14567 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14568 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  NAND2_X1 U14569 ( .A1(n11218), .A2(n11211), .ZN(n21171) );
  MUX2_X1 U14570 ( .A(n11212), .B(n21171), .S(n14683), .Z(n11213) );
  AOI21_X1 U14571 ( .B1(n11214), .B2(n11383), .A(n11213), .ZN(n14370) );
  NAND2_X1 U14572 ( .A1(n11216), .A2(n11215), .ZN(n14329) );
  INV_X1 U14573 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11222) );
  INV_X1 U14574 ( .A(n11227), .ZN(n11220) );
  INV_X1 U14575 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21695) );
  NAND2_X1 U14576 ( .A1(n11218), .A2(n21695), .ZN(n11219) );
  NAND2_X1 U14577 ( .A1(n11220), .A2(n11219), .ZN(n21156) );
  AOI22_X1 U14578 ( .A1(n21156), .A2(n14683), .B1(n13405), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11221) );
  OAI21_X1 U14579 ( .B1(n11711), .B2(n11222), .A(n11221), .ZN(n11223) );
  INV_X1 U14580 ( .A(n11223), .ZN(n11224) );
  NAND2_X1 U14581 ( .A1(n11226), .A2(n11383), .ZN(n11232) );
  INV_X1 U14582 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14583 ( .A1(n11227), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11234) );
  OAI21_X1 U14584 ( .B1(n11227), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11234), .ZN(n21136) );
  AOI22_X1 U14585 ( .A1(n21136), .A2(n14683), .B1(n13405), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11228) );
  OAI21_X1 U14586 ( .B1(n11711), .B2(n11229), .A(n11228), .ZN(n11230) );
  INV_X1 U14587 ( .A(n11230), .ZN(n11231) );
  NAND2_X1 U14588 ( .A1(n11232), .A2(n11231), .ZN(n14514) );
  NAND2_X1 U14589 ( .A1(n11233), .A2(n11383), .ZN(n11240) );
  INV_X1 U14590 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11237) );
  OAI21_X1 U14591 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11235), .A(
        n11269), .ZN(n21123) );
  AOI22_X1 U14592 ( .A1(n14683), .A2(n21123), .B1(n13405), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11236) );
  OAI21_X1 U14593 ( .B1(n11711), .B2(n11237), .A(n11236), .ZN(n11238) );
  INV_X1 U14594 ( .A(n11238), .ZN(n11239) );
  NAND2_X1 U14595 ( .A1(n11240), .A2(n11239), .ZN(n15546) );
  INV_X1 U14596 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15641) );
  INV_X1 U14597 ( .A(n11269), .ZN(n11241) );
  XNOR2_X1 U14598 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11241), .ZN(
        n15859) );
  AOI22_X1 U14599 ( .A1(n14683), .A2(n15859), .B1(n13405), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11242) );
  OAI21_X1 U14600 ( .B1(n11711), .B2(n15641), .A(n11242), .ZN(n11243) );
  INV_X1 U14601 ( .A(n11243), .ZN(n11257) );
  AOI22_X1 U14602 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11575), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14603 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14604 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11699), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14605 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11244) );
  NAND4_X1 U14606 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11255) );
  AOI22_X1 U14607 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11701), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11253) );
  INV_X1 U14608 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16213) );
  INV_X1 U14609 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11248) );
  OAI22_X1 U14610 ( .A1(n16213), .A2(n11652), .B1(n11650), .B2(n11248), .ZN(
        n11249) );
  INV_X1 U14611 ( .A(n11249), .ZN(n11252) );
  AOI22_X1 U14612 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14613 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11250) );
  NAND4_X1 U14614 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11254) );
  OAI21_X1 U14615 ( .B1(n11255), .B2(n11254), .A(n11383), .ZN(n11256) );
  AOI22_X1 U14616 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14617 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14618 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14619 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11259) );
  NAND4_X1 U14620 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11268) );
  AOI22_X1 U14621 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11606), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14622 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14623 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14624 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14625 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11267) );
  OAI21_X1 U14626 ( .B1(n11268), .B2(n11267), .A(n11383), .ZN(n11273) );
  XNOR2_X1 U14627 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11274), .ZN(
        n21118) );
  INV_X1 U14628 ( .A(n21118), .ZN(n11270) );
  AOI22_X1 U14629 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n13405), .B1(
        n14683), .B2(n11270), .ZN(n11272) );
  NAND2_X1 U14630 ( .A1(n13406), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11271) );
  XNOR2_X1 U14631 ( .A(n11293), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17644) );
  NAND2_X1 U14632 ( .A1(n17644), .A2(n14683), .ZN(n11292) );
  AOI22_X1 U14633 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14634 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11279) );
  INV_X1 U14635 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16221) );
  INV_X1 U14636 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11275) );
  OAI22_X1 U14637 ( .A1(n11652), .A2(n16221), .B1(n11650), .B2(n11275), .ZN(
        n11276) );
  INV_X1 U14638 ( .A(n11276), .ZN(n11278) );
  AOI22_X1 U14639 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11277) );
  NAND4_X1 U14640 ( .A1(n11280), .A2(n11279), .A3(n11278), .A4(n11277), .ZN(
        n11286) );
  AOI22_X1 U14641 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14642 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14643 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14644 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11281) );
  NAND4_X1 U14645 ( .A1(n11284), .A2(n11283), .A3(n11282), .A4(n11281), .ZN(
        n11285) );
  NOR2_X1 U14646 ( .A1(n11286), .A2(n11285), .ZN(n11289) );
  NAND2_X1 U14647 ( .A1(n13406), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U14648 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11287) );
  OAI211_X1 U14649 ( .C1(n11364), .C2(n11289), .A(n11288), .B(n11287), .ZN(
        n11290) );
  INV_X1 U14650 ( .A(n11290), .ZN(n11291) );
  NAND2_X1 U14651 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11294) );
  NOR2_X2 U14652 ( .A1(n11368), .A2(n11294), .ZN(n11311) );
  NAND2_X1 U14653 ( .A1(n11311), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11387) );
  XNOR2_X1 U14654 ( .A(n11387), .B(n15397), .ZN(n15791) );
  AOI22_X1 U14655 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14656 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11299) );
  INV_X1 U14657 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16244) );
  INV_X1 U14658 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11295) );
  OAI22_X1 U14659 ( .A1(n11652), .A2(n16244), .B1(n11650), .B2(n11295), .ZN(
        n11296) );
  INV_X1 U14660 ( .A(n11296), .ZN(n11298) );
  AOI22_X1 U14661 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11297) );
  NAND4_X1 U14662 ( .A1(n11300), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(
        n11306) );
  AOI22_X1 U14663 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14664 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14665 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14666 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11301) );
  NAND4_X1 U14667 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11305) );
  NOR2_X1 U14668 ( .A1(n11306), .A2(n11305), .ZN(n11309) );
  NAND2_X1 U14669 ( .A1(n13406), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U14670 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11307) );
  OAI211_X1 U14671 ( .C1(n11364), .C2(n11309), .A(n11308), .B(n11307), .ZN(
        n11310) );
  AOI21_X1 U14672 ( .B1(n15791), .B2(n14683), .A(n11310), .ZN(n15392) );
  XNOR2_X1 U14673 ( .A(n11311), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15807) );
  NAND2_X1 U14674 ( .A1(n15807), .A2(n14683), .ZN(n11329) );
  AOI22_X1 U14675 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14676 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11316) );
  INV_X1 U14677 ( .A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16236) );
  INV_X1 U14678 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11312) );
  OAI22_X1 U14679 ( .A1(n11652), .A2(n16236), .B1(n11650), .B2(n11312), .ZN(
        n11313) );
  INV_X1 U14680 ( .A(n11313), .ZN(n11315) );
  AOI22_X1 U14681 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11314) );
  NAND4_X1 U14682 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11323) );
  AOI22_X1 U14683 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14684 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14685 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14686 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11318) );
  NAND4_X1 U14687 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11322) );
  NOR2_X1 U14688 ( .A1(n11323), .A2(n11322), .ZN(n11326) );
  NAND2_X1 U14689 ( .A1(n13406), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U14690 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11324) );
  OAI211_X1 U14691 ( .C1(n11364), .C2(n11326), .A(n11325), .B(n11324), .ZN(
        n11327) );
  INV_X1 U14692 ( .A(n11327), .ZN(n11328) );
  NAND2_X1 U14693 ( .A1(n11329), .A2(n11328), .ZN(n15405) );
  INV_X1 U14694 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15442) );
  NOR2_X1 U14695 ( .A1(n11368), .A2(n15442), .ZN(n11330) );
  XNOR2_X1 U14696 ( .A(n11330), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15818) );
  NAND2_X1 U14697 ( .A1(n15818), .A2(n14683), .ZN(n11348) );
  AOI22_X1 U14698 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14699 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14700 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14701 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14702 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11342) );
  AOI22_X1 U14703 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11340) );
  INV_X1 U14704 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16232) );
  INV_X1 U14705 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11335) );
  OAI22_X1 U14706 ( .A1(n11652), .A2(n16232), .B1(n11650), .B2(n11335), .ZN(
        n11336) );
  INV_X1 U14707 ( .A(n11336), .ZN(n11339) );
  AOI22_X1 U14708 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14709 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U14710 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11341) );
  NOR2_X1 U14711 ( .A1(n11342), .A2(n11341), .ZN(n11345) );
  NAND2_X1 U14712 ( .A1(n13406), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11344) );
  NAND2_X1 U14713 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11343) );
  OAI211_X1 U14714 ( .C1(n11364), .C2(n11345), .A(n11344), .B(n11343), .ZN(
        n11346) );
  INV_X1 U14715 ( .A(n11346), .ZN(n11347) );
  NAND2_X1 U14716 ( .A1(n11348), .A2(n11347), .ZN(n15421) );
  XNOR2_X1 U14717 ( .A(n11368), .B(n15442), .ZN(n15826) );
  NAND2_X1 U14718 ( .A1(n15826), .A2(n14683), .ZN(n11367) );
  AOI22_X1 U14719 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14720 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11353) );
  INV_X1 U14721 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11466) );
  INV_X1 U14722 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11349) );
  OAI22_X1 U14723 ( .A1(n10833), .A2(n11466), .B1(n11650), .B2(n11349), .ZN(
        n11350) );
  INV_X1 U14724 ( .A(n11350), .ZN(n11352) );
  AOI22_X1 U14725 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14726 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11360) );
  AOI22_X1 U14727 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14728 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14729 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14730 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14731 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  NOR2_X1 U14732 ( .A1(n11360), .A2(n11359), .ZN(n11363) );
  NAND2_X1 U14733 ( .A1(n13406), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11362) );
  NAND2_X1 U14734 ( .A1(n13405), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11361) );
  OAI211_X1 U14735 ( .C1(n11364), .C2(n11363), .A(n11362), .B(n11361), .ZN(
        n11365) );
  INV_X1 U14736 ( .A(n11365), .ZN(n11366) );
  NAND2_X1 U14737 ( .A1(n11367), .A2(n11366), .ZN(n15438) );
  OAI21_X1 U14738 ( .B1(n11369), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n11368), .ZN(n17638) );
  INV_X1 U14739 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15631) );
  INV_X1 U14740 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11370) );
  INV_X1 U14741 ( .A(n13405), .ZN(n11420) );
  OAI22_X1 U14742 ( .A1(n11711), .A2(n15631), .B1(n11370), .B2(n11420), .ZN(
        n11371) );
  AOI21_X1 U14743 ( .B1(n17638), .B2(n14683), .A(n11371), .ZN(n15389) );
  AOI22_X1 U14744 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14745 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14746 ( .A1(n11575), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14747 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U14748 ( .A1(n11375), .A2(n11374), .A3(n11373), .A4(n11372), .ZN(
        n11381) );
  AOI22_X1 U14749 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14750 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14751 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14752 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14753 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11380) );
  OR2_X1 U14754 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  NAND2_X1 U14755 ( .A1(n11383), .A2(n11382), .ZN(n15525) );
  NAND2_X1 U14756 ( .A1(n15389), .A2(n15525), .ZN(n11384) );
  NAND4_X1 U14757 ( .A1(n15405), .A2(n15421), .A3(n15438), .A4(n11384), .ZN(
        n11385) );
  NOR2_X1 U14758 ( .A1(n15392), .A2(n11385), .ZN(n11386) );
  NAND2_X1 U14759 ( .A1(n15387), .A2(n11386), .ZN(n15373) );
  OR2_X2 U14760 ( .A1(n11387), .A2(n15397), .ZN(n11404) );
  XNOR2_X1 U14761 ( .A(n11404), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15785) );
  NAND2_X1 U14762 ( .A1(n15785), .A2(n14683), .ZN(n11402) );
  AOI22_X1 U14763 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n9719), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14764 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11655), .B1(
        n11606), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14765 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14766 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14767 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11397) );
  AOI22_X1 U14768 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11701), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14769 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11699), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14770 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14771 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14772 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  NOR2_X1 U14773 ( .A1(n11397), .A2(n11396), .ZN(n11400) );
  INV_X1 U14774 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15787) );
  AOI21_X1 U14775 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15787), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11398) );
  AOI21_X1 U14776 ( .B1(n13406), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11398), .ZN(
        n11399) );
  OAI21_X1 U14777 ( .B1(n11685), .B2(n11400), .A(n11399), .ZN(n11401) );
  NAND2_X1 U14778 ( .A1(n11402), .A2(n11401), .ZN(n15375) );
  XNOR2_X1 U14779 ( .A(n11426), .B(n15364), .ZN(n15776) );
  AOI22_X1 U14780 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14781 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14782 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14783 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11406) );
  NAND4_X1 U14784 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11419) );
  INV_X1 U14785 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11411) );
  INV_X1 U14786 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11410) );
  OAI22_X1 U14787 ( .A1(n11652), .A2(n11411), .B1(n10833), .B2(n11410), .ZN(
        n11412) );
  INV_X1 U14788 ( .A(n11412), .ZN(n11417) );
  AOI22_X1 U14789 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14790 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14791 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11414) );
  NAND4_X1 U14792 ( .A1(n11417), .A2(n11416), .A3(n11415), .A4(n11414), .ZN(
        n11418) );
  NOR2_X1 U14793 ( .A1(n11419), .A2(n11418), .ZN(n11423) );
  INV_X1 U14794 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15610) );
  OAI22_X1 U14795 ( .A1(n11711), .A2(n15610), .B1(n15364), .B2(n11420), .ZN(
        n11421) );
  INV_X1 U14796 ( .A(n11421), .ZN(n11422) );
  OAI21_X1 U14797 ( .B1(n11685), .B2(n11423), .A(n11422), .ZN(n11424) );
  AOI21_X1 U14798 ( .B1(n15776), .B2(n14683), .A(n11424), .ZN(n15361) );
  INV_X1 U14799 ( .A(n15361), .ZN(n11425) );
  OR2_X2 U14800 ( .A1(n11426), .A2(n15364), .ZN(n11445) );
  XNOR2_X1 U14801 ( .A(n11445), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15759) );
  NAND2_X1 U14802 ( .A1(n15759), .A2(n14683), .ZN(n11444) );
  AOI22_X1 U14803 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14804 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11432) );
  INV_X1 U14805 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11428) );
  INV_X1 U14806 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11427) );
  OAI22_X1 U14807 ( .A1(n11652), .A2(n11428), .B1(n11650), .B2(n11427), .ZN(
        n11429) );
  INV_X1 U14808 ( .A(n11429), .ZN(n11431) );
  AOI22_X1 U14809 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11430) );
  NAND4_X1 U14810 ( .A1(n11433), .A2(n11432), .A3(n11431), .A4(n11430), .ZN(
        n11439) );
  AOI22_X1 U14811 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14812 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14813 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11435) );
  INV_X1 U14814 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n21443) );
  AOI22_X1 U14815 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11434) );
  NAND4_X1 U14816 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11438) );
  NOR2_X1 U14817 ( .A1(n11439), .A2(n11438), .ZN(n11442) );
  NAND2_X1 U14818 ( .A1(n13406), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n11441) );
  OAI21_X1 U14819 ( .B1(n21428), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14687), .ZN(n11440) );
  OAI211_X1 U14820 ( .C1(n11685), .C2(n11442), .A(n11441), .B(n11440), .ZN(
        n11443) );
  NAND2_X1 U14821 ( .A1(n11444), .A2(n11443), .ZN(n15349) );
  OR2_X2 U14822 ( .A1(n11445), .A2(n15761), .ZN(n11446) );
  NAND2_X1 U14823 ( .A1(n11446), .A2(n15340), .ZN(n11447) );
  NAND2_X1 U14824 ( .A1(n11484), .A2(n11447), .ZN(n15748) );
  AOI22_X1 U14825 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14826 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14827 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14828 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14829 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11460) );
  AOI22_X1 U14830 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11458) );
  INV_X1 U14831 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11453) );
  INV_X1 U14832 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11452) );
  OAI22_X1 U14833 ( .A1(n11652), .A2(n11453), .B1(n11650), .B2(n11452), .ZN(
        n11454) );
  INV_X1 U14834 ( .A(n11454), .ZN(n11457) );
  AOI22_X1 U14835 ( .A1(n11700), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14836 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14837 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11459) );
  NOR2_X1 U14838 ( .A1(n11460), .A2(n11459), .ZN(n11464) );
  INV_X1 U14839 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n11461) );
  OAI22_X1 U14840 ( .A1(n11711), .A2(n11461), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15340), .ZN(n11462) );
  INV_X1 U14841 ( .A(n11462), .ZN(n11463) );
  OAI21_X1 U14842 ( .B1(n11685), .B2(n11464), .A(n11463), .ZN(n11465) );
  MUX2_X1 U14843 ( .A(n15748), .B(n11465), .S(n11715), .Z(n15334) );
  XNOR2_X1 U14844 ( .A(n11484), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15741) );
  NAND2_X1 U14845 ( .A1(n15741), .A2(n11190), .ZN(n11483) );
  AOI22_X1 U14846 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14847 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11471) );
  INV_X1 U14848 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11467) );
  OAI22_X1 U14849 ( .A1(n11652), .A2(n11467), .B1(n11650), .B2(n11466), .ZN(
        n11468) );
  INV_X1 U14850 ( .A(n11468), .ZN(n11470) );
  AOI22_X1 U14851 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11469) );
  NAND4_X1 U14852 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n11478) );
  AOI22_X1 U14853 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14854 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14855 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14856 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11473) );
  NAND4_X1 U14857 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11477) );
  NOR2_X1 U14858 ( .A1(n11478), .A2(n11477), .ZN(n11481) );
  NAND2_X1 U14859 ( .A1(n13406), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n11480) );
  OAI21_X1 U14860 ( .B1(n21428), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14687), .ZN(n11479) );
  OAI211_X1 U14861 ( .C1(n11685), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  NAND2_X1 U14862 ( .A1(n11483), .A2(n11482), .ZN(n15323) );
  INV_X1 U14863 ( .A(n11485), .ZN(n11486) );
  INV_X1 U14864 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15733) );
  NAND2_X1 U14865 ( .A1(n11486), .A2(n15733), .ZN(n11487) );
  AND2_X1 U14866 ( .A1(n11574), .A2(n11487), .ZN(n15735) );
  INV_X1 U14867 ( .A(n11685), .ZN(n11713) );
  AOI22_X1 U14868 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14869 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14870 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14871 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11489) );
  NAND4_X1 U14872 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11498) );
  AOI22_X1 U14873 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14874 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14875 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14876 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11493) );
  NAND4_X1 U14877 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(
        n11497) );
  OR2_X1 U14878 ( .A1(n11498), .A2(n11497), .ZN(n11501) );
  INV_X1 U14879 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n11499) );
  OAI22_X1 U14880 ( .A1(n11711), .A2(n11499), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15733), .ZN(n11500) );
  AOI21_X1 U14881 ( .B1(n11713), .B2(n11501), .A(n11500), .ZN(n11502) );
  MUX2_X1 U14882 ( .A(n15735), .B(n11502), .S(n11715), .Z(n15315) );
  NAND2_X1 U14883 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11503) );
  INV_X1 U14884 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11505) );
  OR2_X2 U14885 ( .A1(n11557), .A2(n11505), .ZN(n11617) );
  NAND2_X1 U14886 ( .A1(n11557), .A2(n11505), .ZN(n11506) );
  NAND2_X1 U14887 ( .A1(n11617), .A2(n11506), .ZN(n15700) );
  AOI22_X1 U14888 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14889 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14890 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14891 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11507) );
  NAND4_X1 U14892 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11516) );
  AOI22_X1 U14893 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14894 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14895 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14896 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U14897 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11515) );
  NOR2_X1 U14898 ( .A1(n11516), .A2(n11515), .ZN(n11598) );
  AOI22_X1 U14899 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14900 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14901 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14902 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11517) );
  NAND4_X1 U14903 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11527) );
  AOI22_X1 U14904 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14905 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14906 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14907 ( .A1(n11700), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14908 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11526) );
  NOR2_X1 U14909 ( .A1(n11527), .A2(n11526), .ZN(n11568) );
  AOI22_X1 U14910 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10931), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14911 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14912 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14913 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U14914 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11539) );
  AOI22_X1 U14915 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11697), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14916 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11701), .B1(
        n10837), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14917 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14918 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14919 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  NOR2_X1 U14920 ( .A1(n11539), .A2(n11538), .ZN(n11569) );
  NOR2_X1 U14921 ( .A1(n11568), .A2(n11569), .ZN(n11560) );
  AOI22_X1 U14922 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14923 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11544) );
  INV_X1 U14924 ( .A(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11540) );
  OAI22_X1 U14925 ( .A1(n11652), .A2(n11540), .B1(n11650), .B2(n11410), .ZN(
        n11541) );
  INV_X1 U14926 ( .A(n11541), .ZN(n11543) );
  AOI22_X1 U14927 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11542) );
  NAND4_X1 U14928 ( .A1(n11545), .A2(n11544), .A3(n11543), .A4(n11542), .ZN(
        n11551) );
  AOI22_X1 U14929 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14930 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14931 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14932 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11546) );
  NAND4_X1 U14933 ( .A1(n11549), .A2(n11548), .A3(n11547), .A4(n11546), .ZN(
        n11550) );
  OR2_X1 U14934 ( .A1(n11551), .A2(n11550), .ZN(n11558) );
  NAND2_X1 U14935 ( .A1(n11560), .A2(n11558), .ZN(n11597) );
  XNOR2_X1 U14936 ( .A(n11598), .B(n11597), .ZN(n11554) );
  OAI21_X1 U14937 ( .B1(n21428), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14687), .ZN(n11553) );
  NAND2_X1 U14938 ( .A1(n13406), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14939 ( .C1(n11554), .C2(n11685), .A(n11553), .B(n11552), .ZN(
        n11555) );
  OAI21_X1 U14940 ( .B1(n15700), .B2(n11715), .A(n11555), .ZN(n15265) );
  INV_X1 U14941 ( .A(n15265), .ZN(n11595) );
  INV_X1 U14942 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21549) );
  NAND2_X1 U14943 ( .A1(n11566), .A2(n21549), .ZN(n11556) );
  AND2_X1 U14944 ( .A1(n11557), .A2(n11556), .ZN(n15707) );
  INV_X1 U14945 ( .A(n11558), .ZN(n11559) );
  XNOR2_X1 U14946 ( .A(n11560), .B(n11559), .ZN(n11563) );
  INV_X1 U14947 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11561) );
  OAI22_X1 U14948 ( .A1(n11711), .A2(n11561), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21549), .ZN(n11562) );
  AOI21_X1 U14949 ( .B1(n11563), .B2(n11713), .A(n11562), .ZN(n11564) );
  MUX2_X1 U14950 ( .A(n15707), .B(n11564), .S(n11715), .Z(n15278) );
  INV_X1 U14951 ( .A(n15278), .ZN(n11594) );
  INV_X1 U14952 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15719) );
  INV_X1 U14953 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11565) );
  OAI21_X1 U14954 ( .B1(n11574), .B2(n15719), .A(n11565), .ZN(n11567) );
  NAND2_X1 U14955 ( .A1(n11567), .A2(n11566), .ZN(n15713) );
  XNOR2_X1 U14956 ( .A(n11569), .B(n11568), .ZN(n11572) );
  NAND2_X1 U14957 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14958 ( .A1(n13406), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n11570) );
  OAI211_X1 U14959 ( .C1(n11685), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        n11573) );
  MUX2_X1 U14960 ( .A(n15713), .B(n11573), .S(n11715), .Z(n15288) );
  XNOR2_X1 U14961 ( .A(n11574), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15721) );
  AOI22_X1 U14962 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14963 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11581) );
  INV_X1 U14964 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11577) );
  INV_X1 U14965 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11576) );
  OAI22_X1 U14966 ( .A1(n11652), .A2(n11577), .B1(n11650), .B2(n11576), .ZN(
        n11578) );
  INV_X1 U14967 ( .A(n11578), .ZN(n11580) );
  AOI22_X1 U14968 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14969 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11588) );
  AOI22_X1 U14970 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14971 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11585) );
  INV_X1 U14972 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n21467) );
  AOI22_X1 U14973 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14974 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U14975 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11587) );
  OR2_X1 U14976 ( .A1(n11588), .A2(n11587), .ZN(n11592) );
  INV_X1 U14977 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n11590) );
  OAI21_X1 U14978 ( .B1(n21428), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14687), .ZN(n11589) );
  OAI21_X1 U14979 ( .B1(n11711), .B2(n11590), .A(n11589), .ZN(n11591) );
  AOI21_X1 U14980 ( .B1(n11713), .B2(n11592), .A(n11591), .ZN(n11593) );
  AOI21_X1 U14981 ( .B1(n15721), .B2(n11190), .A(n11593), .ZN(n15304) );
  AND2_X1 U14982 ( .A1(n15288), .A2(n15304), .ZN(n15275) );
  INV_X1 U14983 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15254) );
  XNOR2_X1 U14984 ( .A(n11617), .B(n15254), .ZN(n15685) );
  NOR2_X1 U14985 ( .A1(n11598), .A2(n11597), .ZN(n11622) );
  AOI22_X1 U14986 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11533), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14987 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11604) );
  INV_X1 U14988 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11600) );
  INV_X1 U14989 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11599) );
  OAI22_X1 U14990 ( .A1(n11652), .A2(n11600), .B1(n11650), .B2(n11599), .ZN(
        n11601) );
  INV_X1 U14991 ( .A(n11601), .ZN(n11603) );
  AOI22_X1 U14992 ( .A1(n11628), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14993 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11612) );
  AOI22_X1 U14994 ( .A1(n11606), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14995 ( .A1(n10931), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14996 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14997 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U14998 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  OR2_X1 U14999 ( .A1(n11612), .A2(n11611), .ZN(n11621) );
  XNOR2_X1 U15000 ( .A(n11622), .B(n11621), .ZN(n11615) );
  NAND2_X1 U15001 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U15002 ( .A1(n13406), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n11613) );
  OAI211_X1 U15003 ( .C1(n11615), .C2(n11685), .A(n11614), .B(n11613), .ZN(
        n11616) );
  MUX2_X1 U15004 ( .A(n15685), .B(n11616), .S(n11715), .Z(n15251) );
  NAND2_X1 U15005 ( .A1(n15250), .A2(n15251), .ZN(n15236) );
  INV_X1 U15006 ( .A(n15236), .ZN(n11641) );
  OR2_X2 U15007 ( .A1(n11619), .A2(n15243), .ZN(n11644) );
  NAND2_X1 U15008 ( .A1(n11619), .A2(n15243), .ZN(n11620) );
  NAND2_X1 U15009 ( .A1(n11644), .A2(n11620), .ZN(n15680) );
  NAND2_X1 U15010 ( .A1(n11622), .A2(n11621), .ZN(n11646) );
  AOI22_X1 U15011 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U15012 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U15013 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U15014 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11624) );
  NAND4_X1 U15015 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11635) );
  AOI22_X1 U15016 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11628), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U15017 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U15018 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U15019 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11630) );
  NAND4_X1 U15020 ( .A1(n11633), .A2(n11632), .A3(n11631), .A4(n11630), .ZN(
        n11634) );
  NOR2_X1 U15021 ( .A1(n11635), .A2(n11634), .ZN(n11647) );
  XNOR2_X1 U15022 ( .A(n11646), .B(n11647), .ZN(n11638) );
  NAND2_X1 U15023 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11637) );
  NAND2_X1 U15024 ( .A1(n13406), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11636) );
  OAI211_X1 U15025 ( .C1(n11638), .C2(n11685), .A(n11637), .B(n11636), .ZN(
        n11639) );
  MUX2_X1 U15026 ( .A(n15680), .B(n11639), .S(n11715), .Z(n11640) );
  NAND2_X1 U15027 ( .A1(n11641), .A2(n11640), .ZN(n15223) );
  INV_X1 U15028 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11643) );
  NAND2_X1 U15029 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  NAND2_X1 U15030 ( .A1(n11668), .A2(n11645), .ZN(n15669) );
  NOR2_X1 U15031 ( .A1(n11647), .A2(n11646), .ZN(n11682) );
  INV_X1 U15032 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11648) );
  NOR2_X1 U15033 ( .A1(n10833), .A2(n11648), .ZN(n11654) );
  INV_X1 U15034 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11651) );
  OAI22_X1 U15035 ( .A1(n11652), .A2(n11651), .B1(n11650), .B2(n11649), .ZN(
        n11653) );
  AOI211_X1 U15036 ( .C1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .C2(n11575), .A(
        n11654), .B(n11653), .ZN(n11663) );
  AOI22_X1 U15037 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11655), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U15038 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U15039 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U15040 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11656) );
  AND4_X1 U15041 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11662) );
  AOI22_X1 U15042 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U15043 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U15044 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11681) );
  XNOR2_X1 U15045 ( .A(n11682), .B(n11681), .ZN(n11666) );
  NAND2_X1 U15046 ( .A1(n13406), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11665) );
  OAI21_X1 U15047 ( .B1(n21428), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14687), .ZN(n11664) );
  OAI211_X1 U15048 ( .C1(n11666), .C2(n11685), .A(n11665), .B(n11664), .ZN(
        n11667) );
  OAI21_X1 U15049 ( .B1(n15669), .B2(n11715), .A(n11667), .ZN(n15225) );
  INV_X1 U15050 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U15051 ( .A1(n11668), .A2(n15218), .ZN(n11669) );
  NAND2_X1 U15052 ( .A1(n13464), .A2(n11669), .ZN(n15648) );
  AOI22_X1 U15053 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U15054 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U15055 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11670), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U15056 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U15057 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11680) );
  AOI22_X1 U15058 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U15059 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U15060 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U15061 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U15062 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  NOR2_X1 U15063 ( .A1(n11680), .A2(n11679), .ZN(n11689) );
  NAND2_X1 U15064 ( .A1(n11682), .A2(n11681), .ZN(n11688) );
  XNOR2_X1 U15065 ( .A(n11689), .B(n11688), .ZN(n11686) );
  NAND2_X1 U15066 ( .A1(n14687), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11684) );
  NAND2_X1 U15067 ( .A1(n13406), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11683) );
  OAI211_X1 U15068 ( .C1(n11686), .C2(n11685), .A(n11684), .B(n11683), .ZN(
        n11687) );
  MUX2_X1 U15069 ( .A(n15648), .B(n11687), .S(n11715), .Z(n15213) );
  XNOR2_X1 U15070 ( .A(n13464), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15209) );
  NOR2_X1 U15071 ( .A1(n11689), .A2(n11688), .ZN(n11709) );
  AOI22_X1 U15072 ( .A1(n11655), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U15073 ( .A1(n11012), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11575), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U15074 ( .A1(n11670), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11692), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U15075 ( .A1(n11533), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U15076 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n11707) );
  AOI22_X1 U15077 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U15078 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U15079 ( .A1(n10808), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U15080 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11629), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U15081 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NOR2_X1 U15082 ( .A1(n11707), .A2(n11706), .ZN(n11708) );
  XNOR2_X1 U15083 ( .A(n11709), .B(n11708), .ZN(n11714) );
  INV_X1 U15084 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n11710) );
  INV_X1 U15085 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13463) );
  OAI22_X1 U15086 ( .A1(n11711), .A2(n11710), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13463), .ZN(n11712) );
  AOI21_X1 U15087 ( .B1(n11714), .B2(n11713), .A(n11712), .ZN(n11716) );
  MUX2_X1 U15088 ( .A(n15209), .B(n11716), .S(n11715), .Z(n13403) );
  AND2_X1 U15089 ( .A1(n21654), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21430) );
  NAND2_X1 U15090 ( .A1(n15200), .A2(n17654), .ZN(n11724) );
  NAND2_X1 U15091 ( .A1(n11720), .A2(n16385), .ZN(n21433) );
  NAND2_X1 U15092 ( .A1(n21433), .A2(n21654), .ZN(n11717) );
  NAND2_X1 U15093 ( .A1(n21428), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11719) );
  NOR2_X1 U15094 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14687), .ZN(n21429) );
  INV_X1 U15095 ( .A(n21429), .ZN(n11718) );
  NAND2_X1 U15096 ( .A1(n11719), .A2(n11718), .ZN(n13789) );
  NAND2_X1 U15097 ( .A1(n15209), .A2(n17655), .ZN(n11721) );
  OR2_X2 U15098 ( .A1(n11720), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17669) );
  NAND2_X1 U15099 ( .A1(n15856), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13171) );
  OAI211_X1 U15100 ( .C1(n13463), .C2(n17671), .A(n11721), .B(n13171), .ZN(
        n11722) );
  OAI211_X1 U15101 ( .C1(n21094), .C2(n13174), .A(n11724), .B(n11723), .ZN(
        P1_U2969) );
  AOI22_X1 U15102 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U15103 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U15104 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U15105 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11726) );
  NAND4_X1 U15106 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11739) );
  NAND2_X1 U15107 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U15108 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U15109 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11730) );
  AOI22_X1 U15110 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11769), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11736) );
  INV_X1 U15111 ( .A(n11733), .ZN(n18498) );
  AOI22_X1 U15112 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U15113 ( .A1(n11740), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11734) );
  NAND4_X1 U15114 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11738) );
  OR2_X2 U15115 ( .A1(n11739), .A2(n11738), .ZN(n11930) );
  AOI22_X1 U15116 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U15117 ( .A1(n11740), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11742) );
  AOI22_X1 U15118 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U15119 ( .A1(n11769), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U15120 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U15121 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U15122 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11744) );
  INV_X1 U15123 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U15124 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U15125 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11748) );
  OAI211_X1 U15126 ( .C1(n11750), .C2(n9744), .A(n11749), .B(n11748), .ZN(
        n11751) );
  INV_X1 U15127 ( .A(n11751), .ZN(n11752) );
  NAND3_X2 U15128 ( .A1(n10453), .A2(n11753), .A3(n11752), .ZN(n13998) );
  INV_X1 U15129 ( .A(n11857), .ZN(n11768) );
  INV_X1 U15130 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U15131 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U15132 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11754) );
  OAI211_X1 U15133 ( .C1(n11756), .C2(n9726), .A(n11755), .B(n11754), .ZN(
        n11757) );
  INV_X1 U15134 ( .A(n11757), .ZN(n11761) );
  AOI22_X1 U15135 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15136 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11759) );
  NAND2_X1 U15137 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11758) );
  NAND4_X1 U15138 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11767) );
  AOI22_X1 U15139 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U15140 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11764) );
  INV_X2 U15141 ( .A(n18592), .ZN(n18564) );
  AOI22_X1 U15142 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U15143 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11762) );
  NAND4_X1 U15144 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n11766) );
  OR2_X2 U15145 ( .A1(n11767), .A2(n11766), .ZN(n18785) );
  NAND2_X1 U15146 ( .A1(n11768), .A2(n18785), .ZN(n11860) );
  INV_X1 U15147 ( .A(n11860), .ZN(n11787) );
  AOI22_X1 U15148 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n17550), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U15149 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U15150 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U15151 ( .A1(n18439), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11770) );
  NAND2_X1 U15152 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U15153 ( .A1(n17549), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U15154 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11775) );
  NAND2_X1 U15155 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11774) );
  NAND4_X1 U15156 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11784) );
  INV_X1 U15157 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11778) );
  OR2_X1 U15158 ( .A1(n9726), .A2(n11778), .ZN(n11782) );
  NAND2_X1 U15159 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15160 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U15161 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11779) );
  NAND4_X1 U15162 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  NOR2_X1 U15163 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U15164 ( .A1(n11786), .A2(n11785), .ZN(n11943) );
  NAND2_X1 U15165 ( .A1(n11787), .A2(n11943), .ZN(n11865) );
  INV_X1 U15166 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U15167 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U15168 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11788) );
  OAI211_X1 U15169 ( .C1(n11790), .C2(n9726), .A(n11789), .B(n11788), .ZN(
        n11791) );
  INV_X1 U15170 ( .A(n11791), .ZN(n11795) );
  AOI22_X1 U15171 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U15172 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U15173 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11792) );
  NAND4_X1 U15174 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11801) );
  AOI22_X1 U15175 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U15176 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U15177 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15178 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U15179 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  INV_X1 U15180 ( .A(n11870), .ZN(n11817) );
  INV_X1 U15181 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U15182 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U15183 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11803) );
  OAI211_X1 U15184 ( .C1(n11805), .C2(n9745), .A(n11804), .B(n11803), .ZN(
        n11806) );
  INV_X1 U15185 ( .A(n11806), .ZN(n11810) );
  AOI22_X1 U15186 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U15187 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11808) );
  NAND2_X1 U15188 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11807) );
  NAND4_X1 U15189 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11816) );
  AOI22_X1 U15190 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15191 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U15192 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15193 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U15194 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11815) );
  NAND2_X1 U15195 ( .A1(n11817), .A2(n11950), .ZN(n11874) );
  INV_X1 U15196 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18506) );
  NAND2_X1 U15197 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U15198 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11818) );
  OAI211_X1 U15199 ( .C1(n18506), .C2(n9745), .A(n11819), .B(n11818), .ZN(
        n11820) );
  INV_X1 U15200 ( .A(n11820), .ZN(n11824) );
  AOI22_X1 U15201 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U15202 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U15203 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11821) );
  NAND4_X1 U15204 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11831) );
  AOI22_X1 U15205 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U15206 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U15207 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U15208 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U15209 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11830) );
  OR2_X2 U15210 ( .A1(n11874), .A2(n18769), .ZN(n19174) );
  XNOR2_X1 U15211 ( .A(n13998), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13862) );
  INV_X1 U15212 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U15213 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11833) );
  NAND2_X1 U15214 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11832) );
  OAI211_X1 U15215 ( .C1(n11834), .C2(n9726), .A(n11833), .B(n11832), .ZN(
        n11835) );
  INV_X1 U15216 ( .A(n11835), .ZN(n11840) );
  AOI22_X1 U15217 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15218 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11838) );
  NAND2_X1 U15219 ( .A1(n11740), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11837) );
  NAND4_X1 U15220 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11849) );
  AOI22_X1 U15221 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15222 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15223 ( .A1(n11725), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11844) );
  NAND4_X1 U15224 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11848) );
  NAND2_X1 U15225 ( .A1(n14007), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13861) );
  INV_X1 U15226 ( .A(n13861), .ZN(n13956) );
  NAND2_X1 U15227 ( .A1(n13862), .A2(n13956), .ZN(n11851) );
  INV_X1 U15228 ( .A(n13998), .ZN(n11935) );
  NAND2_X1 U15229 ( .A1(n11935), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U15230 ( .A1(n11851), .A2(n11850), .ZN(n19214) );
  OAI21_X1 U15231 ( .B1(n11930), .B2(n13998), .A(n11857), .ZN(n11852) );
  XNOR2_X1 U15232 ( .A(n11852), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19215) );
  NAND2_X1 U15233 ( .A1(n19214), .A2(n19215), .ZN(n11855) );
  INV_X1 U15234 ( .A(n11852), .ZN(n11853) );
  NAND2_X1 U15235 ( .A1(n11853), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11854) );
  INV_X1 U15236 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11856) );
  XNOR2_X1 U15237 ( .A(n11857), .B(n18785), .ZN(n13884) );
  NAND2_X1 U15238 ( .A1(n11858), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11859) );
  INV_X1 U15239 ( .A(n11943), .ZN(n18781) );
  XNOR2_X1 U15240 ( .A(n11860), .B(n18781), .ZN(n11861) );
  XNOR2_X1 U15241 ( .A(n11861), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17462) );
  INV_X1 U15242 ( .A(n11861), .ZN(n11862) );
  NAND2_X1 U15243 ( .A1(n11862), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11863) );
  NAND2_X2 U15244 ( .A1(n11864), .A2(n11863), .ZN(n11868) );
  XNOR2_X1 U15245 ( .A(n11865), .B(n11927), .ZN(n11866) );
  XNOR2_X2 U15246 ( .A(n11868), .B(n11866), .ZN(n13810) );
  INV_X1 U15247 ( .A(n11866), .ZN(n11867) );
  NAND2_X1 U15248 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  XNOR2_X1 U15249 ( .A(n11870), .B(n18772), .ZN(n11871) );
  XNOR2_X1 U15250 ( .A(n11871), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13822) );
  INV_X1 U15251 ( .A(n11871), .ZN(n11872) );
  NAND2_X1 U15252 ( .A1(n11872), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U15253 ( .A1(n11874), .A2(n18769), .ZN(n11875) );
  NAND2_X1 U15254 ( .A1(n19174), .A2(n11875), .ZN(n11876) );
  INV_X1 U15255 ( .A(n11876), .ZN(n11877) );
  NAND2_X1 U15256 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  INV_X1 U15257 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19389) );
  INV_X1 U15258 ( .A(n19092), .ZN(n11881) );
  INV_X1 U15259 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11880) );
  INV_X1 U15260 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19093) );
  AND2_X2 U15261 ( .A1(n11882), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19382) );
  INV_X1 U15262 ( .A(n19382), .ZN(n19081) );
  NAND2_X1 U15263 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19386) );
  NOR2_X1 U15264 ( .A1(n19386), .A2(n19142), .ZN(n19358) );
  NAND3_X1 U15265 ( .A1(n19358), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19068) );
  INV_X1 U15266 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19310) );
  NAND2_X1 U15267 ( .A1(n19056), .A2(n19037), .ZN(n11886) );
  NOR2_X1 U15268 ( .A1(n19012), .A2(n19257), .ZN(n19273) );
  AND2_X1 U15269 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11888) );
  AND2_X1 U15270 ( .A1(n11888), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11887) );
  AND2_X1 U15271 ( .A1(n19273), .A2(n11887), .ZN(n13233) );
  AND2_X1 U15272 ( .A1(n19037), .A2(n11888), .ZN(n11889) );
  AND2_X1 U15273 ( .A1(n19273), .A2(n11889), .ZN(n19252) );
  AND2_X1 U15274 ( .A1(n19174), .A2(n19303), .ZN(n19025) );
  NAND2_X1 U15275 ( .A1(n19025), .A2(n19012), .ZN(n11890) );
  NOR2_X1 U15276 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11890), .ZN(
        n18997) );
  INV_X1 U15277 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19268) );
  INV_X1 U15278 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19250) );
  INV_X1 U15279 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19261) );
  NAND3_X1 U15280 ( .A1(n18977), .A2(n19250), .A3(n19261), .ZN(n11891) );
  NAND2_X1 U15281 ( .A1(n11892), .A2(n11891), .ZN(n11893) );
  OR2_X2 U15282 ( .A1(n17521), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17522) );
  NAND3_X1 U15283 ( .A1(n17522), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n18965), .ZN(n11894) );
  INV_X1 U15284 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17516) );
  NAND2_X1 U15285 ( .A1(n11894), .A2(n19113), .ZN(n18945) );
  NAND2_X1 U15286 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17481) );
  NAND2_X1 U15287 ( .A1(n19113), .A2(n17481), .ZN(n11895) );
  AND2_X2 U15288 ( .A1(n18945), .A2(n11895), .ZN(n11896) );
  AND2_X1 U15289 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17584) );
  AND2_X1 U15290 ( .A1(n17584), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17483) );
  NAND2_X1 U15291 ( .A1(n17425), .A2(n19113), .ZN(n17423) );
  INV_X1 U15292 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n19225) );
  INV_X1 U15293 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17578) );
  NOR2_X1 U15294 ( .A1(n13996), .A2(n17536), .ZN(n20106) );
  NOR2_X1 U15295 ( .A1(n11898), .A2(n11903), .ZN(n11901) );
  NAND2_X1 U15296 ( .A1(n11899), .A2(n14115), .ZN(n11900) );
  NOR2_X1 U15297 ( .A1(n19508), .A2(n11922), .ZN(n13918) );
  OAI21_X2 U15298 ( .B1(n13920), .B2(n11905), .A(n13919), .ZN(n19390) );
  NOR2_X2 U15299 ( .A1(n11906), .A2(n11905), .ZN(n19253) );
  INV_X1 U15300 ( .A(n11907), .ZN(n11912) );
  INV_X1 U15301 ( .A(n11908), .ZN(n11911) );
  NAND2_X1 U15302 ( .A1(n11909), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11910) );
  NAND2_X1 U15303 ( .A1(n11911), .A2(n11910), .ZN(n11923) );
  NOR2_X1 U15304 ( .A1(n11912), .A2(n11923), .ZN(n11913) );
  NOR2_X1 U15305 ( .A1(n11914), .A2(n11913), .ZN(n11915) );
  OR2_X1 U15306 ( .A1(n11916), .A2(n11915), .ZN(n11918) );
  AND3_X1 U15307 ( .A1(n11921), .A2(n11920), .A3(n11919), .ZN(n13217) );
  AND2_X1 U15308 ( .A1(n19500), .A2(n20089), .ZN(n13227) );
  NOR2_X1 U15309 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  OR2_X1 U15310 ( .A1(n17850), .A2(n11925), .ZN(n19947) );
  OR2_X2 U15311 ( .A1(n17853), .A2(n19496), .ZN(n19217) );
  NAND2_X1 U15312 ( .A1(n17491), .A2(n19128), .ZN(n11973) );
  INV_X1 U15313 ( .A(n17483), .ZN(n17476) );
  NAND2_X1 U15314 ( .A1(n19177), .A2(n19210), .ZN(n13501) );
  INV_X1 U15315 ( .A(n11930), .ZN(n18793) );
  NAND2_X1 U15316 ( .A1(n11933), .A2(n18793), .ZN(n11929) );
  NAND2_X1 U15317 ( .A1(n11929), .A2(n18785), .ZN(n11944) );
  NOR2_X1 U15318 ( .A1(n18781), .A2(n11944), .ZN(n11928) );
  NAND2_X1 U15319 ( .A1(n11928), .A2(n18775), .ZN(n11951) );
  NOR2_X1 U15320 ( .A1(n18772), .A2(n11951), .ZN(n11954) );
  NAND2_X1 U15321 ( .A1(n11954), .A2(n13245), .ZN(n11955) );
  XNOR2_X1 U15322 ( .A(n11928), .B(n11927), .ZN(n11948) );
  AND2_X1 U15323 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11948), .ZN(
        n11949) );
  XNOR2_X1 U15324 ( .A(n11929), .B(n18785), .ZN(n11940) );
  NOR2_X1 U15325 ( .A1(n11856), .A2(n11940), .ZN(n11942) );
  INV_X1 U15326 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19465) );
  NOR2_X1 U15327 ( .A1(n11931), .A2(n19465), .ZN(n11939) );
  NOR2_X1 U15328 ( .A1(n14007), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13957) );
  INV_X1 U15329 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11932) );
  OR2_X1 U15330 ( .A1(n13957), .A2(n11932), .ZN(n11936) );
  OAI21_X1 U15331 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n11933), .ZN(n11934) );
  AOI21_X1 U15332 ( .B1(n11936), .B2(n11935), .A(n11934), .ZN(n19211) );
  INV_X1 U15333 ( .A(n19211), .ZN(n11937) );
  NOR2_X1 U15334 ( .A1(n19212), .A2(n11937), .ZN(n11938) );
  NOR2_X1 U15335 ( .A1(n11939), .A2(n11938), .ZN(n13891) );
  XNOR2_X1 U15336 ( .A(n11856), .B(n11940), .ZN(n13890) );
  NOR2_X1 U15337 ( .A1(n13891), .A2(n13890), .ZN(n11941) );
  XOR2_X1 U15338 ( .A(n11944), .B(n11943), .Z(n11946) );
  NOR2_X1 U15339 ( .A1(n11945), .A2(n11946), .ZN(n11947) );
  INV_X1 U15340 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19449) );
  XNOR2_X1 U15341 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11948), .ZN(
        n13816) );
  NOR2_X1 U15342 ( .A1(n11949), .A2(n13815), .ZN(n11952) );
  XOR2_X1 U15343 ( .A(n11951), .B(n11950), .Z(n11953) );
  INV_X1 U15344 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19420) );
  XNOR2_X1 U15345 ( .A(n11954), .B(n13245), .ZN(n11957) );
  NAND2_X1 U15346 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n19185), .ZN(
        n11959) );
  NOR2_X1 U15347 ( .A1(n11955), .A2(n11959), .ZN(n11961) );
  INV_X1 U15348 ( .A(n11955), .ZN(n11960) );
  OR2_X1 U15349 ( .A1(n11957), .A2(n11956), .ZN(n19186) );
  OAI21_X1 U15350 ( .B1(n11960), .B2(n11959), .A(n19186), .ZN(n11958) );
  AOI21_X1 U15351 ( .B1(n11960), .B2(n11959), .A(n11958), .ZN(n19173) );
  NOR2_X2 U15352 ( .A1(n19173), .A2(n9983), .ZN(n19172) );
  INV_X1 U15353 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U15354 ( .A1(n18941), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17515) );
  INV_X1 U15355 ( .A(n17515), .ZN(n13216) );
  NAND3_X1 U15356 ( .A1(n13502), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18942) );
  NOR2_X1 U15357 ( .A1(n17481), .A2(n18942), .ZN(n13236) );
  AOI21_X1 U15358 ( .B1(n17476), .B2(n13501), .A(n18925), .ZN(n11970) );
  INV_X1 U15359 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17497) );
  OR2_X1 U15360 ( .A1(n19095), .A2(n19210), .ZN(n11963) );
  NAND2_X1 U15361 ( .A1(n18981), .A2(n19382), .ZN(n11962) );
  NAND2_X2 U15362 ( .A1(n11963), .A2(n11962), .ZN(n19164) );
  AND2_X2 U15363 ( .A1(n19164), .A2(n19296), .ZN(n19048) );
  INV_X1 U15364 ( .A(n13236), .ZN(n19224) );
  NOR2_X1 U15365 ( .A1(n19067), .A2(n19224), .ZN(n18919) );
  NOR2_X1 U15366 ( .A1(n17476), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17501) );
  INV_X1 U15367 ( .A(n20103), .ZN(n14134) );
  NAND2_X1 U15368 ( .A1(n20102), .A2(n20070), .ZN(n17846) );
  NAND2_X1 U15369 ( .A1(n14134), .A2(n17846), .ZN(n17560) );
  NOR2_X1 U15370 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17452), .ZN(
        n17743) );
  NAND3_X1 U15371 ( .A1(n11964), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17746) );
  NOR2_X1 U15372 ( .A1(n17872), .A2(n17746), .ZN(n11965) );
  OR2_X1 U15373 ( .A1(n19507), .A2(n11965), .ZN(n17747) );
  OAI211_X1 U15374 ( .C1(n10507), .C2(n19103), .A(n19202), .B(n17747), .ZN(
        n17742) );
  NOR2_X1 U15375 ( .A1(n17743), .A2(n17742), .ZN(n17438) );
  NOR2_X1 U15376 ( .A1(n17438), .A2(n13369), .ZN(n11968) );
  INV_X1 U15377 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18177) );
  NAND2_X1 U15378 ( .A1(n11965), .A2(n19062), .ZN(n17442) );
  NAND2_X1 U15379 ( .A1(n19477), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17495) );
  NAND2_X1 U15380 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n19105) );
  NAND2_X2 U15381 ( .A1(n19202), .A2(n19105), .ZN(n19151) );
  NAND2_X1 U15382 ( .A1(n19124), .A2(n13365), .ZN(n11966) );
  OAI211_X1 U15383 ( .C1(n17442), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17495), .B(n11966), .ZN(n11967) );
  AOI211_X1 U15384 ( .C1(n18919), .C2(n17501), .A(n11968), .B(n11967), .ZN(
        n11969) );
  OAI21_X1 U15385 ( .B1(n11970), .B2(n17497), .A(n11969), .ZN(n11971) );
  INV_X1 U15386 ( .A(n11971), .ZN(n11972) );
  NAND2_X1 U15387 ( .A1(n11973), .A2(n11972), .ZN(P3_U2800) );
  INV_X2 U15388 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14248) );
  AOI22_X1 U15389 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11977) );
  INV_X1 U15390 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11974) );
  AND2_X2 U15391 ( .A1(n11974), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12186) );
  AND2_X4 U15392 ( .A1(n12186), .A2(n14209), .ZN(n14783) );
  AOI22_X1 U15393 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11976) );
  AND2_X2 U15394 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12455) );
  AND2_X4 U15395 ( .A1(n12455), .A2(n14248), .ZN(n14789) );
  AOI22_X1 U15396 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15397 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  NAND2_X1 U15398 ( .A1(n11979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11987) );
  AOI22_X1 U15399 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15400 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15401 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11981) );
  NAND4_X1 U15402 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11985) );
  NAND2_X1 U15403 ( .A1(n11985), .A2(n11984), .ZN(n11986) );
  AOI22_X1 U15404 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15405 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15406 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15407 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11988) );
  NAND4_X1 U15408 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11992) );
  NAND2_X1 U15409 ( .A1(n11992), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11999) );
  AOI22_X1 U15410 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15411 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U15412 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11997) );
  NAND2_X1 U15413 ( .A1(n11997), .A2(n11984), .ZN(n11998) );
  INV_X2 U15414 ( .A(n12080), .ZN(n12083) );
  AOI22_X1 U15415 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15416 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15417 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15418 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U15419 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12013) );
  AOI22_X1 U15420 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15421 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15422 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12008) );
  NAND4_X1 U15423 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12012) );
  NAND2_X2 U15424 ( .A1(n12013), .A2(n12012), .ZN(n12091) );
  AOI22_X1 U15425 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12043), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15426 ( .A1(n12181), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15427 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14783), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15428 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U15429 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12018) );
  NAND2_X1 U15430 ( .A1(n12018), .A2(n11984), .ZN(n12025) );
  AOI22_X1 U15431 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15432 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14783), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15433 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15434 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15435 ( .A1(n12021), .A2(n12022), .A3(n12020), .A4(n12019), .ZN(
        n12023) );
  NAND2_X1 U15436 ( .A1(n12023), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12024) );
  NAND4_X2 U15437 ( .A1(n12602), .A2(n12083), .A3(n12091), .A4(n12103), .ZN(
        n12051) );
  AOI22_X1 U15438 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15439 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15440 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15441 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12030) );
  NAND2_X1 U15442 ( .A1(n12030), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12037) );
  AOI22_X1 U15443 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15444 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15445 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U15446 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12035) );
  NAND2_X1 U15447 ( .A1(n12035), .A2(n11984), .ZN(n12036) );
  AOI22_X1 U15448 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15449 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15450 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15451 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9747), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U15452 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12042) );
  NAND2_X1 U15453 ( .A1(n12042), .A2(n11984), .ZN(n12050) );
  AOI22_X1 U15454 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15455 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15456 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U15457 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12048) );
  NAND2_X1 U15458 ( .A1(n12048), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12049) );
  INV_X1 U15459 ( .A(n12437), .ZN(n12067) );
  NOR2_X2 U15460 ( .A1(n12051), .A2(n12095), .ZN(n12447) );
  AOI22_X1 U15461 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15462 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9748), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15463 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12052) );
  NAND3_X1 U15464 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12058) );
  OR2_X2 U15465 ( .A1(n12056), .A2(n12055), .ZN(n12057) );
  OAI21_X2 U15466 ( .B1(n12058), .B2(n12057), .A(n11984), .ZN(n12065) );
  AOI22_X1 U15467 ( .A1(n12180), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12043), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15468 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15469 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15470 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9747), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U15471 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12063) );
  NAND2_X2 U15472 ( .A1(n12065), .A2(n12064), .ZN(n12605) );
  AOI22_X1 U15473 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15474 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15475 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15476 ( .A1(n14789), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9748), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15477 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12072) );
  NAND2_X1 U15478 ( .A1(n12072), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12079) );
  AOI22_X1 U15479 ( .A1(n12043), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15480 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12181), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15481 ( .A1(n14788), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12180), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15482 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9747), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U15483 ( .A1(n12076), .A2(n12075), .A3(n12074), .A4(n12073), .ZN(
        n12077) );
  NAND2_X1 U15484 ( .A1(n12077), .A2(n11984), .ZN(n12078) );
  INV_X1 U15485 ( .A(n12103), .ZN(n12081) );
  NAND4_X1 U15486 ( .A1(n12081), .A2(n12602), .A3(n12080), .A4(n12091), .ZN(
        n12082) );
  INV_X1 U15487 ( .A(n14263), .ZN(n12088) );
  AND2_X1 U15488 ( .A1(n12095), .A2(n12083), .ZN(n12086) );
  OAI21_X1 U15489 ( .B1(n9874), .B2(n13769), .A(n12084), .ZN(n12085) );
  NAND3_X1 U15490 ( .A1(n12105), .A2(n12086), .A3(n12085), .ZN(n12087) );
  NAND3_X1 U15491 ( .A1(n12088), .A2(n12087), .A3(n9725), .ZN(n12573) );
  NAND2_X1 U15492 ( .A1(n12127), .A2(n9725), .ZN(n12092) );
  NAND2_X1 U15493 ( .A1(n12573), .A2(n12092), .ZN(n12093) );
  NAND2_X1 U15494 ( .A1(n12093), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12094) );
  INV_X1 U15495 ( .A(n12121), .ZN(n12102) );
  NAND2_X1 U15496 ( .A1(n12609), .A2(n9874), .ZN(n12426) );
  AND2_X1 U15497 ( .A1(n12426), .A2(n12602), .ZN(n12098) );
  NAND2_X1 U15498 ( .A1(n12096), .A2(n12095), .ZN(n12432) );
  NAND2_X1 U15499 ( .A1(n12098), .A2(n12424), .ZN(n12565) );
  NAND2_X1 U15500 ( .A1(n12565), .A2(n14604), .ZN(n12100) );
  NAND2_X1 U15501 ( .A1(n12100), .A2(n12099), .ZN(n12128) );
  NAND2_X1 U15502 ( .A1(n12128), .A2(n12116), .ZN(n12101) );
  NAND2_X2 U15503 ( .A1(n12102), .A2(n12101), .ZN(n12156) );
  NAND2_X1 U15504 ( .A1(n12156), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U15505 ( .A1(n9735), .A2(n12388), .ZN(n13738) );
  NAND3_X1 U15506 ( .A1(n13738), .A2(n9874), .A3(n12602), .ZN(n12108) );
  NAND3_X1 U15507 ( .A1(n12419), .A2(n12123), .A3(n13769), .ZN(n12104) );
  NAND2_X1 U15508 ( .A1(n12104), .A2(n12081), .ZN(n12106) );
  NAND2_X1 U15509 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  NOR2_X2 U15510 ( .A1(n12108), .A2(n12107), .ZN(n12563) );
  NAND2_X1 U15511 ( .A1(n12563), .A2(n12576), .ZN(n14206) );
  INV_X1 U15512 ( .A(n14206), .ZN(n12113) );
  INV_X1 U15513 ( .A(n12576), .ZN(n12423) );
  NOR2_X1 U15514 ( .A1(n12109), .A2(n12423), .ZN(n12110) );
  AND2_X2 U15515 ( .A1(n12110), .A2(n12116), .ZN(n12139) );
  NAND2_X1 U15516 ( .A1(n17409), .A2(n21075), .ZN(n21066) );
  INV_X1 U15517 ( .A(n21066), .ZN(n12133) );
  NAND2_X1 U15518 ( .A1(n12133), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U15519 ( .A1(n12150), .A2(n12111), .ZN(n12112) );
  AOI21_X1 U15520 ( .B1(n12113), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12112), 
        .ZN(n12114) );
  INV_X1 U15521 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n20123) );
  NAND2_X1 U15522 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12117) );
  AND2_X1 U15523 ( .A1(n21066), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U15524 ( .A1(n12139), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12118) );
  OAI211_X1 U15525 ( .C1(n12499), .C2(n20123), .A(n12119), .B(n12118), .ZN(
        n12120) );
  NOR2_X1 U15526 ( .A1(n12121), .A2(n12120), .ZN(n12131) );
  AND2_X2 U15527 ( .A1(n12123), .A2(n12602), .ZN(n13744) );
  NAND2_X1 U15528 ( .A1(n13744), .A2(n20400), .ZN(n12124) );
  NAND2_X1 U15529 ( .A1(n12132), .A2(n14904), .ZN(n12126) );
  NAND2_X1 U15530 ( .A1(n12562), .A2(n10473), .ZN(n12130) );
  NAND2_X1 U15531 ( .A1(n10463), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12129) );
  NAND3_X1 U15532 ( .A1(n12131), .A2(n12130), .A3(n12129), .ZN(n12162) );
  NAND2_X1 U15533 ( .A1(n12156), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12135) );
  AOI22_X1 U15534 ( .A1(n12132), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12133), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U15535 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U15536 ( .A1(n12139), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n12136) );
  OAI211_X1 U15537 ( .C1(n12499), .C2(n20957), .A(n12137), .B(n12136), .ZN(
        n12138) );
  NAND2_X1 U15538 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12141) );
  NAND2_X1 U15539 ( .A1(n12139), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12140) );
  OAI211_X1 U15540 ( .C1(n12499), .C2(n20959), .A(n12141), .B(n12140), .ZN(
        n12142) );
  INV_X1 U15541 ( .A(n12142), .ZN(n12143) );
  OAI21_X1 U15542 ( .B1(n21692), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n17409), 
        .ZN(n12145) );
  AOI21_X2 U15543 ( .B1(n12156), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12145), .ZN(n12147) );
  XNOR2_X2 U15544 ( .A(n12146), .B(n12147), .ZN(n12158) );
  INV_X1 U15545 ( .A(n12146), .ZN(n12148) );
  NAND2_X1 U15546 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  INV_X1 U15547 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12152) );
  NAND2_X1 U15548 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12151) );
  NAND2_X2 U15549 ( .A1(n12155), .A2(n12154), .ZN(n12481) );
  NOR2_X1 U15550 ( .A1(n21066), .A2(n21494), .ZN(n12157) );
  XNOR2_X2 U15551 ( .A(n12481), .B(n12482), .ZN(n12479) );
  INV_X1 U15552 ( .A(n12163), .ZN(n12164) );
  NAND2_X1 U15553 ( .A1(n9739), .A2(n12164), .ZN(n12165) );
  INV_X1 U15554 ( .A(n12167), .ZN(n12168) );
  AND2_X2 U15555 ( .A1(n12176), .A2(n12177), .ZN(n12290) );
  AND2_X2 U15556 ( .A1(n12176), .A2(n12171), .ZN(n12299) );
  AOI22_X1 U15557 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n12290), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12169) );
  INV_X1 U15558 ( .A(n13952), .ZN(n12170) );
  AOI22_X1 U15559 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12298), .B1(
        n12291), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U15560 ( .A1(n12178), .A2(n12177), .ZN(n12210) );
  AND2_X2 U15561 ( .A1(n14783), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12352) );
  AOI22_X1 U15562 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14803), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12185) );
  AND2_X2 U15563 ( .A1(n14788), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12349) );
  AOI22_X1 U15564 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n12349), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12183) );
  AND2_X2 U15565 ( .A1(n9749), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12252) );
  AOI22_X1 U15566 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12273), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15567 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12194) );
  AND2_X2 U15568 ( .A1(n14789), .A2(n11984), .ZN(n14804) );
  AOI22_X1 U15569 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12278), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12192) );
  AND2_X2 U15570 ( .A1(n12001), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12257) );
  AND2_X2 U15571 ( .A1(n12001), .A2(n11984), .ZN(n12245) );
  AOI22_X1 U15572 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12257), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15573 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12231), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12190) );
  NOR2_X1 U15574 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15575 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12233), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12189) );
  NAND4_X1 U15576 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12193) );
  NAND2_X1 U15577 ( .A1(n12635), .A2(n14904), .ZN(n12195) );
  INV_X1 U15578 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12196) );
  INV_X1 U15579 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12199) );
  INV_X1 U15580 ( .A(n12291), .ZN(n12198) );
  INV_X1 U15581 ( .A(n12299), .ZN(n20675) );
  INV_X1 U15582 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12197) );
  OAI22_X1 U15583 ( .A1(n12199), .A2(n12198), .B1(n20675), .B2(n12197), .ZN(
        n12200) );
  NOR2_X1 U15584 ( .A1(n12201), .A2(n12200), .ZN(n12227) );
  INV_X1 U15585 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12203) );
  INV_X1 U15586 ( .A(n12296), .ZN(n12202) );
  INV_X1 U15587 ( .A(n12290), .ZN(n20743) );
  INV_X1 U15588 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21575) );
  OAI22_X1 U15589 ( .A1(n12203), .A2(n12202), .B1(n20743), .B2(n21575), .ZN(
        n12206) );
  INV_X1 U15590 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12204) );
  NOR2_X1 U15591 ( .A1(n12206), .A2(n12205), .ZN(n12226) );
  INV_X1 U15592 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12212) );
  INV_X1 U15593 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12209) );
  OAI211_X1 U15594 ( .C1(n12213), .C2(n12212), .A(n12211), .B(n21078), .ZN(
        n12214) );
  INV_X1 U15595 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12217) );
  INV_X1 U15596 ( .A(n14396), .ZN(n12300) );
  INV_X1 U15597 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12216) );
  OAI22_X1 U15598 ( .A1(n12217), .A2(n12300), .B1(n14594), .B2(n12216), .ZN(
        n12223) );
  INV_X1 U15599 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12221) );
  INV_X1 U15600 ( .A(n12297), .ZN(n12220) );
  INV_X1 U15601 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12219) );
  OAI22_X1 U15602 ( .A1(n12221), .A2(n12220), .B1(n12218), .B2(n12219), .ZN(
        n12222) );
  NOR2_X1 U15603 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  AOI22_X1 U15604 ( .A1(n12240), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15605 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15606 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15607 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15608 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15609 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15610 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12349), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15611 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14803), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15612 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n12352), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15613 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15614 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12273), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12241) );
  NAND4_X1 U15615 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .ZN(
        n12251) );
  AOI22_X1 U15616 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12278), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15617 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12245), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15618 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12231), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15619 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12233), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15620 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12250) );
  NAND3_X1 U15621 ( .A1(n14904), .A2(n13563), .A3(n12611), .ZN(n12267) );
  AOI22_X1 U15622 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15623 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15624 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15625 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12253) );
  NAND4_X1 U15626 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12263) );
  AOI22_X1 U15627 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15628 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15629 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15630 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15631 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  NAND2_X1 U15632 ( .A1(n12267), .A2(n12621), .ZN(n12264) );
  NOR2_X1 U15633 ( .A1(n13563), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12265) );
  XNOR2_X1 U15634 ( .A(n12265), .B(n12611), .ZN(n13665) );
  NAND2_X1 U15635 ( .A1(n13665), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13667) );
  INV_X1 U15636 ( .A(n13563), .ZN(n12604) );
  NAND3_X1 U15637 ( .A1(n12604), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n12611), .ZN(n12266) );
  NAND2_X1 U15638 ( .A1(n13667), .A2(n12266), .ZN(n12268) );
  INV_X1 U15639 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14653) );
  XNOR2_X1 U15640 ( .A(n12268), .B(n14653), .ZN(n13648) );
  XNOR2_X1 U15641 ( .A(n12267), .B(n12621), .ZN(n13647) );
  NAND2_X1 U15642 ( .A1(n13648), .A2(n13647), .ZN(n13650) );
  NAND2_X1 U15643 ( .A1(n12268), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15644 ( .A1(n13650), .A2(n12269), .ZN(n12271) );
  XNOR2_X1 U15645 ( .A(n12271), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17132) );
  INV_X1 U15646 ( .A(n17132), .ZN(n12270) );
  NAND2_X1 U15647 ( .A1(n12271), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12272) );
  AOI22_X1 U15648 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15649 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15650 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15651 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15652 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12284) );
  AOI22_X1 U15653 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15654 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15655 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15656 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12279) );
  NAND4_X1 U15657 ( .A1(n12282), .A2(n12281), .A3(n12280), .A4(n12279), .ZN(
        n12283) );
  INV_X1 U15658 ( .A(n12395), .ZN(n12285) );
  NAND2_X1 U15659 ( .A1(n12286), .A2(n12285), .ZN(n12287) );
  INV_X1 U15660 ( .A(n17113), .ZN(n12288) );
  INV_X1 U15661 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20363) );
  AOI22_X1 U15662 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20374), .B1(
        n20599), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15663 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n12290), .B1(
        n20635), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15664 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12291), .B1(
        n20446), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15665 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12296), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15666 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12297), .B1(
        n20862), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15667 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12298), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12304) );
  INV_X1 U15668 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12301) );
  INV_X1 U15669 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21707) );
  OAI22_X1 U15670 ( .A1(n12301), .A2(n9905), .B1(n12300), .B2(n21707), .ZN(
        n12302) );
  INV_X1 U15671 ( .A(n12302), .ZN(n12303) );
  AOI22_X1 U15672 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15673 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15674 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15675 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15676 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12316) );
  AOI22_X1 U15677 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15678 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15679 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15680 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15681 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12315) );
  NOR2_X1 U15682 ( .A1(n12316), .A2(n12315), .ZN(n12817) );
  NAND2_X1 U15683 ( .A1(n12817), .A2(n14904), .ZN(n12317) );
  INV_X1 U15684 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U15685 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12296), .B1(
        n14601), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15686 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20374), .B1(
        n12297), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15687 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20599), .B1(
        n20862), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15688 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12320), .B1(
        n14396), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15689 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12290), .B1(
        n12299), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15690 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20446), .B1(
        n20709), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15691 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12298), .B1(
        n12291), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15692 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12349), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15693 ( .A1(n12240), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15694 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15695 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12329) );
  NAND4_X1 U15696 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12338) );
  AOI22_X1 U15697 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15698 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15699 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15700 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12333) );
  NAND4_X1 U15701 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12337) );
  NAND2_X1 U15702 ( .A1(n12844), .A2(n14904), .ZN(n12339) );
  NAND2_X1 U15703 ( .A1(n12341), .A2(n12843), .ZN(n12346) );
  INV_X1 U15704 ( .A(n12348), .ZN(n12344) );
  INV_X1 U15705 ( .A(n12349), .ZN(n12456) );
  INV_X1 U15706 ( .A(n14802), .ZN(n12351) );
  INV_X1 U15707 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12350) );
  OAI22_X1 U15708 ( .A1(n12456), .A2(n21637), .B1(n12351), .B2(n12350), .ZN(
        n12358) );
  INV_X1 U15709 ( .A(n12352), .ZN(n12356) );
  INV_X1 U15710 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14945) );
  INV_X1 U15711 ( .A(n12353), .ZN(n12355) );
  INV_X1 U15712 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12354) );
  OAI22_X1 U15713 ( .A1(n12356), .A2(n14945), .B1(n12355), .B2(n12354), .ZN(
        n12357) );
  NOR2_X1 U15714 ( .A1(n12358), .A2(n12357), .ZN(n12370) );
  AOI22_X1 U15715 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15716 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12361) );
  NAND2_X1 U15717 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12360) );
  NAND2_X1 U15718 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12359) );
  NAND2_X1 U15719 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U15720 ( .A1(n12240), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12365) );
  NAND2_X1 U15721 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12364) );
  NAND2_X1 U15722 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12363) );
  AOI22_X1 U15723 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12367) );
  NAND4_X2 U15724 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12822) );
  INV_X1 U15725 ( .A(n12371), .ZN(n12372) );
  NAND2_X1 U15726 ( .A1(n12372), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12373) );
  INV_X1 U15727 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17341) );
  NAND2_X1 U15728 ( .A1(n14716), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13334) );
  NAND2_X1 U15729 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12378) );
  NOR2_X1 U15730 ( .A1(n13334), .A2(n12378), .ZN(n13454) );
  AND2_X1 U15731 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13301) );
  AND2_X1 U15732 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17262) );
  AND2_X1 U15733 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12379) );
  NAND3_X1 U15734 ( .A1(n13301), .A2(n17262), .A3(n12379), .ZN(n13299) );
  INV_X1 U15735 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13307) );
  NOR2_X1 U15736 ( .A1(n13299), .A2(n13307), .ZN(n12380) );
  NAND2_X1 U15737 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17194) );
  NAND2_X1 U15738 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17151) );
  AND2_X1 U15739 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13175) );
  AND2_X1 U15740 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n13175), .ZN(
        n12381) );
  NAND2_X1 U15741 ( .A1(n16870), .A2(n12381), .ZN(n12383) );
  INV_X1 U15742 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12382) );
  INV_X1 U15743 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20936) );
  NOR2_X1 U15744 ( .A1(n20936), .A2(n20955), .ZN(n20947) );
  NAND2_X1 U15745 ( .A1(n14609), .A2(n14204), .ZN(n12418) );
  XNOR2_X1 U15746 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15747 ( .A1(n12402), .A2(n12399), .ZN(n12385) );
  NAND2_X1 U15748 ( .A1(n21050), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12384) );
  NAND2_X1 U15749 ( .A1(n12385), .A2(n12384), .ZN(n12397) );
  XNOR2_X1 U15750 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15751 ( .A1(n12397), .A2(n12396), .ZN(n12387) );
  NAND2_X1 U15752 ( .A1(n21692), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12386) );
  NAND2_X1 U15753 ( .A1(n12387), .A2(n12386), .ZN(n12391) );
  XNOR2_X1 U15754 ( .A(n12391), .B(n12389), .ZN(n12408) );
  INV_X1 U15755 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U15756 ( .A1(n12391), .A2(n12390), .ZN(n12393) );
  NAND2_X1 U15757 ( .A1(n21494), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12392) );
  NAND2_X1 U15758 ( .A1(n12393), .A2(n12392), .ZN(n12411) );
  OR2_X1 U15759 ( .A1(n12411), .A2(n12412), .ZN(n12409) );
  MUX2_X1 U15760 ( .A(n12395), .B(n12409), .S(n12388), .Z(n12816) );
  NAND2_X1 U15761 ( .A1(n21074), .A2(n21078), .ZN(n12398) );
  XNOR2_X1 U15762 ( .A(n12397), .B(n12396), .ZN(n12441) );
  INV_X1 U15763 ( .A(n12441), .ZN(n12451) );
  MUX2_X1 U15764 ( .A(n12398), .B(n12388), .S(n12451), .Z(n12407) );
  NAND2_X1 U15765 ( .A1(n12122), .A2(n12451), .ZN(n12405) );
  INV_X1 U15766 ( .A(n12402), .ZN(n12444) );
  INV_X1 U15767 ( .A(n12399), .ZN(n12401) );
  NAND2_X1 U15768 ( .A1(n14248), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12400) );
  NAND2_X1 U15769 ( .A1(n12401), .A2(n12400), .ZN(n12440) );
  OAI21_X1 U15770 ( .B1(n12444), .B2(n12440), .A(n12997), .ZN(n12404) );
  INV_X1 U15771 ( .A(n12440), .ZN(n12450) );
  XNOR2_X1 U15772 ( .A(n12402), .B(n12401), .ZN(n12428) );
  OAI211_X1 U15773 ( .C1(n12450), .C2(n21078), .A(n9725), .B(n12428), .ZN(
        n12403) );
  NAND3_X1 U15774 ( .A1(n12405), .A2(n12404), .A3(n12403), .ZN(n12406) );
  NAND2_X1 U15775 ( .A1(n12407), .A2(n12406), .ZN(n12410) );
  NAND2_X1 U15776 ( .A1(n12409), .A2(n12408), .ZN(n12430) );
  INV_X1 U15777 ( .A(n12430), .ZN(n12453) );
  NAND2_X1 U15778 ( .A1(n12416), .A2(n9725), .ZN(n12414) );
  NAND2_X1 U15779 ( .A1(n12414), .A2(n9874), .ZN(n12417) );
  INV_X1 U15780 ( .A(n12449), .ZN(n21057) );
  OAI21_X1 U15781 ( .B1(n12091), .B2(n21078), .A(n9725), .ZN(n12420) );
  NAND2_X1 U15782 ( .A1(n12420), .A2(n12602), .ZN(n12421) );
  NAND2_X1 U15783 ( .A1(n12421), .A2(n12083), .ZN(n12422) );
  AND3_X1 U15784 ( .A1(n12424), .A2(n12423), .A3(n12422), .ZN(n12436) );
  NAND2_X1 U15785 ( .A1(n12426), .A2(n12083), .ZN(n12427) );
  NAND2_X1 U15786 ( .A1(n12425), .A2(n12427), .ZN(n12435) );
  NAND2_X1 U15787 ( .A1(n12451), .A2(n12428), .ZN(n12429) );
  NAND3_X1 U15788 ( .A1(n12437), .A2(n13523), .A3(n14204), .ZN(n12434) );
  NAND2_X1 U15789 ( .A1(n12432), .A2(n12602), .ZN(n12433) );
  AND2_X1 U15790 ( .A1(n14904), .A2(n21077), .ZN(n12448) );
  NAND2_X1 U15791 ( .A1(n12433), .A2(n12448), .ZN(n12566) );
  MUX2_X1 U15792 ( .A(n12437), .B(n14609), .S(n14904), .Z(n12438) );
  AND2_X1 U15793 ( .A1(n13523), .A2(n21073), .ZN(n13739) );
  NAND2_X1 U15794 ( .A1(n12438), .A2(n13739), .ZN(n12439) );
  NAND2_X1 U15795 ( .A1(n14225), .A2(n12439), .ZN(n12463) );
  MUX2_X1 U15796 ( .A(n12604), .B(n12440), .S(n12388), .Z(n12832) );
  OAI21_X1 U15797 ( .B1(n12443), .B2(n12388), .A(n12442), .ZN(n12805) );
  OAI21_X1 U15798 ( .B1(n12832), .B2(n12444), .A(n12805), .ZN(n12446) );
  NAND2_X1 U15799 ( .A1(n12446), .A2(n12445), .ZN(n21055) );
  NAND3_X1 U15800 ( .A1(n21055), .A2(n21056), .A3(n12449), .ZN(n12462) );
  AND2_X1 U15801 ( .A1(n12451), .A2(n12450), .ZN(n12452) );
  AOI21_X1 U15802 ( .B1(n12453), .B2(n12452), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n12454) );
  NAND2_X1 U15803 ( .A1(n13523), .A2(n12454), .ZN(n12460) );
  AOI21_X1 U15804 ( .B1(n14229), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14264) );
  NAND2_X1 U15805 ( .A1(n12456), .A2(n14264), .ZN(n12458) );
  INV_X1 U15806 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12457) );
  NAND2_X1 U15807 ( .A1(n12458), .A2(n12457), .ZN(n12459) );
  NAND2_X1 U15808 ( .A1(n12459), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17403) );
  NAND2_X1 U15809 ( .A1(n12460), .A2(n17403), .ZN(n21061) );
  NAND3_X1 U15810 ( .A1(n21061), .A2(n12447), .A3(n21078), .ZN(n12461) );
  INV_X1 U15811 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20975) );
  CLKBUF_X3 U15812 ( .A(n12466), .Z(n12559) );
  OR2_X1 U15813 ( .A1(n12552), .A2(n17250), .ZN(n12468) );
  INV_X2 U15814 ( .A(n12150), .ZN(n12555) );
  AOI22_X1 U15815 ( .A1(n12555), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12467) );
  OAI211_X1 U15816 ( .C1(n12557), .C2(n20975), .A(n12468), .B(n12467), .ZN(
        n14624) );
  INV_X1 U15817 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17268) );
  OR2_X1 U15818 ( .A1(n12552), .A2(n17268), .ZN(n12470) );
  AOI22_X1 U15819 ( .A1(n12555), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12469) );
  OAI211_X1 U15820 ( .C1(n12557), .C2(n20973), .A(n12470), .B(n12469), .ZN(
        n14528) );
  INV_X1 U15821 ( .A(n14528), .ZN(n12478) );
  INV_X1 U15822 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n21471) );
  NAND2_X1 U15823 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12472) );
  NAND2_X1 U15824 ( .A1(n12555), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12471) );
  OAI211_X1 U15825 ( .C1(n12557), .C2(n21471), .A(n12472), .B(n12471), .ZN(
        n12473) );
  AOI21_X1 U15826 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12473), .ZN(n14587) );
  INV_X1 U15827 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U15828 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U15829 ( .A1(n12555), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12474) );
  OAI211_X1 U15830 ( .C1(n12557), .C2(n12476), .A(n12475), .B(n12474), .ZN(
        n12477) );
  AOI21_X1 U15831 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12477), .ZN(n16753) );
  OR2_X1 U15832 ( .A1(n14587), .A2(n16753), .ZN(n14527) );
  NOR2_X1 U15833 ( .A1(n12478), .A2(n14527), .ZN(n14525) );
  AND2_X1 U15834 ( .A1(n14624), .A2(n14525), .ZN(n12515) );
  NAND2_X1 U15835 ( .A1(n12480), .A2(n12479), .ZN(n12485) );
  INV_X1 U15836 ( .A(n12481), .ZN(n12483) );
  NAND2_X1 U15837 ( .A1(n12483), .A2(n12482), .ZN(n12484) );
  NAND2_X1 U15838 ( .A1(n12485), .A2(n12484), .ZN(n17107) );
  INV_X1 U15839 ( .A(n17107), .ZN(n12491) );
  INV_X1 U15840 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12488) );
  NAND2_X1 U15841 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12487) );
  NAND2_X1 U15842 ( .A1(n12555), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12486) );
  OAI211_X1 U15843 ( .C1(n12499), .C2(n12488), .A(n12487), .B(n12486), .ZN(
        n12489) );
  AOI21_X1 U15844 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12489), .ZN(n17106) );
  INV_X1 U15845 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15846 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15847 ( .A1(n12555), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12492) );
  OAI211_X1 U15848 ( .C1(n12499), .C2(n12494), .A(n12493), .B(n12492), .ZN(
        n12495) );
  AOI21_X1 U15849 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12495), .ZN(n14015) );
  INV_X1 U15850 ( .A(n14015), .ZN(n12496) );
  INV_X1 U15851 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20961) );
  NAND2_X1 U15852 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12498) );
  NAND2_X1 U15853 ( .A1(n12555), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12497) );
  OAI211_X1 U15854 ( .C1(n12499), .C2(n20961), .A(n12498), .B(n12497), .ZN(
        n12500) );
  AOI21_X1 U15855 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12500), .ZN(n13487) );
  INV_X1 U15856 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20963) );
  INV_X1 U15857 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17357) );
  OR2_X1 U15858 ( .A1(n12552), .A2(n17357), .ZN(n12502) );
  AOI22_X1 U15859 ( .A1(n12555), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12501) );
  OAI211_X1 U15860 ( .C1(n12557), .C2(n20963), .A(n12502), .B(n12501), .ZN(
        n14128) );
  INV_X1 U15861 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17077) );
  NAND2_X1 U15862 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U15863 ( .A1(n12555), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12503) );
  OAI211_X1 U15864 ( .C1(n12557), .C2(n17077), .A(n12504), .B(n12503), .ZN(
        n12505) );
  AOI21_X1 U15865 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12505), .ZN(n14415) );
  INV_X1 U15866 ( .A(n14415), .ZN(n12506) );
  INV_X1 U15867 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20966) );
  NAND2_X1 U15868 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12509) );
  NAND2_X1 U15869 ( .A1(n12555), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12508) );
  OAI211_X1 U15870 ( .C1(n12557), .C2(n20966), .A(n12509), .B(n12508), .ZN(
        n12510) );
  AOI21_X1 U15871 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12510), .ZN(n14409) );
  INV_X1 U15872 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20968) );
  OR2_X1 U15873 ( .A1(n12552), .A2(n17319), .ZN(n12512) );
  AOI22_X1 U15874 ( .A1(n12555), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12511) );
  OAI211_X1 U15875 ( .C1(n12557), .C2(n20968), .A(n12512), .B(n12511), .ZN(
        n17050) );
  INV_X1 U15876 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12707) );
  INV_X1 U15877 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17302) );
  OR2_X1 U15878 ( .A1(n12552), .A2(n17302), .ZN(n12514) );
  AOI22_X1 U15879 ( .A1(n12555), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12513) );
  OAI211_X1 U15880 ( .C1(n12557), .C2(n12707), .A(n12514), .B(n12513), .ZN(
        n14619) );
  NAND2_X1 U15881 ( .A1(n12515), .A2(n14526), .ZN(n14645) );
  INV_X1 U15882 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20977) );
  NAND2_X1 U15883 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U15884 ( .A1(n12555), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12516) );
  OAI211_X1 U15885 ( .C1(n12557), .C2(n20977), .A(n12517), .B(n12516), .ZN(
        n12518) );
  AOI21_X1 U15886 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12518), .ZN(n14644) );
  INV_X1 U15887 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20979) );
  NAND2_X1 U15888 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12520) );
  NAND2_X1 U15889 ( .A1(n12555), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12519) );
  OAI211_X1 U15890 ( .C1(n12557), .C2(n20979), .A(n12520), .B(n12519), .ZN(
        n12521) );
  AOI21_X1 U15891 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12521), .ZN(n14629) );
  INV_X1 U15892 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20981) );
  NAND2_X1 U15893 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U15894 ( .A1(n12555), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12522) );
  OAI211_X1 U15895 ( .C1(n12557), .C2(n20981), .A(n12523), .B(n12522), .ZN(
        n12524) );
  AOI21_X1 U15896 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n12524), .ZN(n13318) );
  INV_X1 U15897 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20983) );
  OR2_X1 U15898 ( .A1(n12552), .A2(n16952), .ZN(n12526) );
  AOI22_X1 U15899 ( .A1(n12555), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n12525) );
  OAI211_X1 U15900 ( .C1(n12557), .C2(n20983), .A(n12526), .B(n12525), .ZN(
        n16743) );
  INV_X1 U15901 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20985) );
  NAND2_X1 U15902 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12528) );
  NAND2_X1 U15903 ( .A1(n12555), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12527) );
  OAI211_X1 U15904 ( .C1(n12557), .C2(n20985), .A(n12528), .B(n12527), .ZN(
        n12529) );
  AOI21_X1 U15905 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12529), .ZN(n13294) );
  INV_X1 U15906 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20987) );
  NAND2_X1 U15907 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U15908 ( .A1(n12555), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12530) );
  OAI211_X1 U15909 ( .C1(n12557), .C2(n20987), .A(n12531), .B(n12530), .ZN(
        n12532) );
  AOI21_X1 U15910 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12532), .ZN(n13448) );
  INV_X1 U15911 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20989) );
  OR2_X1 U15912 ( .A1(n12552), .A2(n17214), .ZN(n12534) );
  AOI22_X1 U15913 ( .A1(n12555), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12533) );
  OAI211_X1 U15914 ( .C1(n12557), .C2(n20989), .A(n12534), .B(n12533), .ZN(
        n16530) );
  INV_X1 U15915 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20991) );
  INV_X1 U15916 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12952) );
  OR2_X1 U15917 ( .A1(n12552), .A2(n12952), .ZN(n12536) );
  AOI22_X1 U15918 ( .A1(n12555), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12535) );
  OAI211_X1 U15919 ( .C1(n12557), .C2(n20991), .A(n12536), .B(n12535), .ZN(
        n16522) );
  NAND2_X1 U15920 ( .A1(n16521), .A2(n16522), .ZN(n16498) );
  INV_X1 U15921 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20993) );
  NAND2_X1 U15922 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15923 ( .A1(n12555), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12537) );
  OAI211_X1 U15924 ( .C1(n12557), .C2(n20993), .A(n12538), .B(n12537), .ZN(
        n12539) );
  AOI21_X1 U15925 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12539), .ZN(n16499) );
  OR2_X2 U15926 ( .A1(n16498), .A2(n16499), .ZN(n16501) );
  INV_X1 U15927 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20995) );
  NAND2_X1 U15928 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15929 ( .A1(n12555), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12540) );
  OAI211_X1 U15930 ( .C1(n12557), .C2(n20995), .A(n12541), .B(n12540), .ZN(
        n12542) );
  AOI21_X1 U15931 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n12542), .ZN(n16485) );
  NOR2_X4 U15932 ( .A1(n16501), .A2(n16485), .ZN(n16484) );
  INV_X1 U15933 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20997) );
  INV_X1 U15934 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13253) );
  OR2_X1 U15935 ( .A1(n12552), .A2(n13253), .ZN(n12544) );
  AOI22_X1 U15936 ( .A1(n12555), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12543) );
  OAI211_X1 U15937 ( .C1(n12557), .C2(n20997), .A(n12544), .B(n12543), .ZN(
        n13257) );
  INV_X1 U15938 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n21001) );
  OR2_X1 U15939 ( .A1(n12552), .A2(n17152), .ZN(n12546) );
  AOI22_X1 U15940 ( .A1(n12555), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12545) );
  OAI211_X1 U15941 ( .C1(n12557), .C2(n21001), .A(n12546), .B(n12545), .ZN(
        n16463) );
  INV_X1 U15942 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U15943 ( .A1(n12555), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12549) );
  NAND2_X1 U15944 ( .A1(n12547), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12548) );
  OAI211_X1 U15945 ( .C1(n12552), .C2(n17140), .A(n12549), .B(n12548), .ZN(
        n16449) );
  INV_X1 U15946 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n21004) );
  AOI22_X1 U15947 ( .A1(n12555), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12550) );
  OAI21_X1 U15948 ( .B1(n12557), .B2(n21004), .A(n12550), .ZN(n12551) );
  AOI21_X1 U15949 ( .B1(n12466), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12551), .ZN(n13179) );
  INV_X1 U15950 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15174) );
  INV_X1 U15951 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12582) );
  OR2_X1 U15952 ( .A1(n12552), .A2(n12582), .ZN(n12554) );
  AOI22_X1 U15953 ( .A1(n12555), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12553) );
  OAI211_X1 U15954 ( .C1(n12557), .C2(n15174), .A(n12554), .B(n12553), .ZN(
        n13360) );
  NAND2_X1 U15955 ( .A1(n13361), .A2(n13360), .ZN(n12561) );
  INV_X1 U15956 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15957 ( .A1(n12555), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12556) );
  OAI21_X1 U15958 ( .B1(n12557), .B2(n12800), .A(n12556), .ZN(n12558) );
  AOI21_X1 U15959 ( .B1(n12559), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12558), .ZN(n12560) );
  NAND2_X1 U15960 ( .A1(n12998), .A2(n9740), .ZN(n17352) );
  AND3_X1 U15961 ( .A1(n14904), .A2(n12083), .A3(n12991), .ZN(n12564) );
  AND2_X1 U15962 ( .A1(n12563), .A2(n12564), .ZN(n14213) );
  NAND2_X1 U15963 ( .A1(n12998), .A2(n14213), .ZN(n14707) );
  NAND2_X1 U15964 ( .A1(n12565), .A2(n21078), .ZN(n14239) );
  NAND2_X1 U15965 ( .A1(n14239), .A2(n12566), .ZN(n12567) );
  NAND2_X1 U15966 ( .A1(n12567), .A2(n14604), .ZN(n12575) );
  INV_X1 U15967 ( .A(n12568), .ZN(n12570) );
  INV_X1 U15968 ( .A(n13634), .ZN(n12569) );
  NAND2_X1 U15969 ( .A1(n12570), .A2(n12569), .ZN(n13741) );
  INV_X1 U15970 ( .A(n13738), .ZN(n13528) );
  OAI21_X1 U15971 ( .B1(n12576), .B2(n9874), .A(n13528), .ZN(n12572) );
  NAND2_X1 U15972 ( .A1(n14609), .A2(n21077), .ZN(n12571) );
  AND4_X1 U15973 ( .A1(n12573), .A2(n13741), .A3(n12572), .A4(n12571), .ZN(
        n12574) );
  NAND2_X1 U15974 ( .A1(n12575), .A2(n12574), .ZN(n13635) );
  AOI21_X1 U15975 ( .B1(n10463), .B2(n12576), .A(n13635), .ZN(n14238) );
  NAND2_X1 U15976 ( .A1(n14238), .A2(n13634), .ZN(n12577) );
  NAND2_X1 U15977 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17379) );
  INV_X1 U15978 ( .A(n17379), .ZN(n14651) );
  AND2_X1 U15979 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14651), .ZN(
        n12588) );
  INV_X1 U15980 ( .A(n12588), .ZN(n12578) );
  NAND2_X1 U15981 ( .A1(n14707), .A2(n12578), .ZN(n12579) );
  NAND2_X1 U15982 ( .A1(n14653), .A2(n17379), .ZN(n12587) );
  NAND2_X1 U15983 ( .A1(n12579), .A2(n12587), .ZN(n12580) );
  NAND3_X1 U15984 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U15985 ( .A1(n13451), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12581) );
  INV_X1 U15986 ( .A(n17194), .ZN(n12594) );
  NAND2_X1 U15987 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n12585), .ZN(
        n13259) );
  INV_X1 U15988 ( .A(n13175), .ZN(n13384) );
  NOR3_X1 U15989 ( .A1(n13384), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12582), .ZN(n12583) );
  NAND2_X1 U15990 ( .A1(n17409), .A2(n20821), .ZN(n21025) );
  NAND2_X1 U15991 ( .A1(n20864), .A2(n21075), .ZN(n15155) );
  NOR2_X1 U15992 ( .A1(n12586), .A2(n12800), .ZN(n13394) );
  AOI21_X1 U15993 ( .B1(n17137), .B2(n12583), .A(n13394), .ZN(n12584) );
  INV_X1 U15994 ( .A(n12584), .ZN(n12599) );
  INV_X1 U15995 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17181) );
  NAND2_X1 U15996 ( .A1(n12585), .A2(n17181), .ZN(n17180) );
  OR2_X1 U15997 ( .A1(n12998), .A2(n20263), .ZN(n17396) );
  AND2_X1 U15998 ( .A1(n17396), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12590) );
  OR2_X1 U15999 ( .A1(n14707), .A2(n12587), .ZN(n14662) );
  OR2_X1 U16000 ( .A1(n14709), .A2(n12588), .ZN(n12589) );
  INV_X1 U16001 ( .A(n12591), .ZN(n12592) );
  AND2_X1 U16002 ( .A1(n17367), .A2(n12592), .ZN(n12593) );
  NAND2_X1 U16003 ( .A1(n17730), .A2(n12593), .ZN(n17258) );
  NAND3_X1 U16004 ( .A1(n13451), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12594), .ZN(n12595) );
  OAI21_X1 U16005 ( .B1(n17258), .B2(n12595), .A(n17259), .ZN(n17182) );
  NAND2_X1 U16006 ( .A1(n17180), .A2(n17182), .ZN(n17164) );
  AND2_X1 U16007 ( .A1(n17380), .A2(n17151), .ZN(n12596) );
  OR2_X1 U16008 ( .A1(n17164), .A2(n12596), .ZN(n17157) );
  AOI21_X1 U16009 ( .B1(n17380), .B2(n17152), .A(n17157), .ZN(n17141) );
  OAI211_X1 U16010 ( .C1(n17397), .C2(n13175), .A(n17141), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13349) );
  OAI211_X1 U16011 ( .C1(n17380), .C2(n17164), .A(n13349), .B(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12597) );
  INV_X1 U16012 ( .A(n12597), .ZN(n12598) );
  OAI21_X1 U16013 ( .B1(n15183), .B2(n17352), .A(n12600), .ZN(n12601) );
  INV_X1 U16014 ( .A(n12601), .ZN(n13000) );
  NAND2_X1 U16015 ( .A1(n13749), .A2(n12632), .ZN(n12622) );
  MUX2_X1 U16016 ( .A(n12602), .B(n14390), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12603) );
  AOI21_X1 U16017 ( .B1(n12605), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U16018 ( .A1(n13751), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12606) );
  NAND2_X1 U16019 ( .A1(n13746), .A2(n13745), .ZN(n12616) );
  NOR2_X1 U16020 ( .A1(n12602), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U16021 ( .A1(n12625), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12608) );
  OAI21_X1 U16022 ( .B1(n12624), .B2(n20957), .A(n12608), .ZN(n12617) );
  XNOR2_X1 U16023 ( .A(n12616), .B(n12617), .ZN(n14193) );
  NAND2_X1 U16024 ( .A1(n12609), .A2(n12602), .ZN(n12610) );
  MUX2_X1 U16025 ( .A(n12610), .B(n21050), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12615) );
  NAND2_X1 U16026 ( .A1(n12611), .A2(n12991), .ZN(n12809) );
  INV_X1 U16027 ( .A(n12809), .ZN(n12613) );
  NAND2_X1 U16028 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  AND2_X1 U16029 ( .A1(n12615), .A2(n12614), .ZN(n14192) );
  INV_X1 U16030 ( .A(n12617), .ZN(n12618) );
  NAND2_X1 U16031 ( .A1(n12616), .A2(n12618), .ZN(n12619) );
  NAND2_X1 U16032 ( .A1(n14195), .A2(n12619), .ZN(n12630) );
  OR2_X1 U16033 ( .A1(n12620), .A2(n12621), .ZN(n12623) );
  OAI211_X1 U16034 ( .C1(n20821), .C2(n21692), .A(n12623), .B(n12622), .ZN(
        n12628) );
  XNOR2_X1 U16035 ( .A(n12630), .B(n12628), .ZN(n14189) );
  NAND2_X1 U16036 ( .A1(n12793), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U16037 ( .A1(n12794), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12626) );
  AND2_X1 U16038 ( .A1(n12627), .A2(n12626), .ZN(n14188) );
  INV_X1 U16039 ( .A(n12628), .ZN(n12629) );
  NAND2_X1 U16040 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  NAND2_X1 U16041 ( .A1(n12793), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U16042 ( .A1(n12632), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12634) );
  NAND2_X1 U16043 ( .A1(n12794), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12633) );
  AND2_X1 U16044 ( .A1(n12634), .A2(n12633), .ZN(n12638) );
  INV_X1 U16045 ( .A(n12620), .ZN(n12636) );
  NAND2_X1 U16046 ( .A1(n12636), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U16047 ( .A1(n12793), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U16048 ( .A1(n12794), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12642) );
  OR2_X1 U16049 ( .A1(n12620), .A2(n12285), .ZN(n12641) );
  NAND2_X1 U16050 ( .A1(n12793), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U16051 ( .A1(n12794), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12647) );
  OR2_X1 U16052 ( .A1(n12620), .A2(n12817), .ZN(n12646) );
  AOI22_X1 U16053 ( .A1(n12794), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12649) );
  OAI21_X1 U16054 ( .B1(n12624), .B2(n20961), .A(n12649), .ZN(n13760) );
  AOI22_X1 U16055 ( .A1(n12794), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12650) );
  OAI21_X1 U16056 ( .B1(n12624), .B2(n20963), .A(n12650), .ZN(n13763) );
  AND2_X1 U16057 ( .A1(n13760), .A2(n13763), .ZN(n12652) );
  INV_X1 U16058 ( .A(n13763), .ZN(n12651) );
  OR2_X1 U16059 ( .A1(n12620), .A2(n12994), .ZN(n13761) );
  AOI21_X1 U16060 ( .B1(n13489), .B2(n12652), .A(n10450), .ZN(n13756) );
  INV_X1 U16061 ( .A(n13756), .ZN(n12667) );
  NAND2_X1 U16062 ( .A1(n12793), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U16063 ( .A1(n12794), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U16064 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12349), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U16065 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U16066 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U16067 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12653) );
  NAND4_X1 U16068 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n12662) );
  AOI22_X1 U16069 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U16070 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U16071 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U16072 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12657) );
  NAND4_X1 U16073 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12661) );
  INV_X1 U16074 ( .A(n14474), .ZN(n14407) );
  OR2_X1 U16075 ( .A1(n12620), .A2(n14407), .ZN(n12663) );
  NAND2_X1 U16076 ( .A1(n12667), .A2(n12666), .ZN(n13754) );
  NAND2_X1 U16077 ( .A1(n12793), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U16078 ( .A1(n12794), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12632), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U16079 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14803), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U16080 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U16081 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12349), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U16082 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12273), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12668) );
  NAND4_X1 U16083 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        n12677) );
  AOI22_X1 U16084 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14804), .B1(
        n12278), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U16085 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12245), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U16086 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12232), .B1(
        n12231), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U16087 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12233), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12672) );
  NAND4_X1 U16088 ( .A1(n12675), .A2(n12674), .A3(n12673), .A4(n12672), .ZN(
        n12676) );
  INV_X1 U16089 ( .A(n14616), .ZN(n12678) );
  OR2_X1 U16090 ( .A1(n12620), .A2(n12678), .ZN(n12679) );
  NAND2_X1 U16091 ( .A1(n12793), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U16092 ( .A1(n12794), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U16093 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U16094 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U16095 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U16096 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12682) );
  NAND4_X1 U16097 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12691) );
  AOI22_X1 U16098 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U16099 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U16100 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U16101 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U16102 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12690) );
  INV_X1 U16103 ( .A(n14477), .ZN(n20285) );
  OR2_X1 U16104 ( .A1(n12620), .A2(n20285), .ZN(n12692) );
  AOI22_X1 U16105 ( .A1(n12794), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U16106 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14803), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U16107 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U16108 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U16109 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12273), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12695) );
  NAND4_X1 U16110 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        n12704) );
  AOI22_X1 U16111 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14804), .B1(
        n12278), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U16112 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U16113 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12232), .B1(
        n12231), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U16114 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12233), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12699) );
  NAND4_X1 U16115 ( .A1(n12702), .A2(n12701), .A3(n12700), .A4(n12699), .ZN(
        n12703) );
  INV_X1 U16116 ( .A(n14618), .ZN(n16758) );
  OR2_X1 U16117 ( .A1(n12620), .A2(n16758), .ZN(n12705) );
  OAI211_X1 U16118 ( .C1(n12624), .C2(n12707), .A(n12706), .B(n12705), .ZN(
        n13859) );
  NAND2_X1 U16119 ( .A1(n12793), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U16120 ( .A1(n12794), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U16121 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12349), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U16122 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U16123 ( .A1(n12240), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U16124 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12708) );
  NAND4_X1 U16125 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n12708), .ZN(
        n12717) );
  AOI22_X1 U16126 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U16127 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U16128 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U16129 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12712) );
  NAND4_X1 U16130 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n12716) );
  NOR2_X1 U16131 ( .A1(n12717), .A2(n12716), .ZN(n16757) );
  OR2_X1 U16132 ( .A1(n12620), .A2(n16757), .ZN(n12718) );
  NAND2_X1 U16133 ( .A1(n12793), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U16134 ( .A1(n12794), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U16135 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U16136 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U16137 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U16138 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12723) );
  NAND4_X1 U16139 ( .A1(n12726), .A2(n12725), .A3(n12724), .A4(n12723), .ZN(
        n12732) );
  AOI22_X1 U16140 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U16141 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U16142 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U16143 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U16144 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12731) );
  OR2_X1 U16145 ( .A1(n12732), .A2(n12731), .ZN(n14492) );
  INV_X1 U16146 ( .A(n14492), .ZN(n14583) );
  OR2_X1 U16147 ( .A1(n12620), .A2(n14583), .ZN(n12733) );
  AOI22_X1 U16148 ( .A1(n12794), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U16149 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12349), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U16150 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U16151 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12737) );
  AOI22_X1 U16152 ( .A1(n14804), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12736) );
  NAND4_X1 U16153 ( .A1(n12739), .A2(n12738), .A3(n12737), .A4(n12736), .ZN(
        n12745) );
  AOI22_X1 U16154 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U16155 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U16156 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U16157 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12740) );
  NAND4_X1 U16158 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n12740), .ZN(
        n12744) );
  INV_X1 U16159 ( .A(n14530), .ZN(n12746) );
  OR2_X1 U16160 ( .A1(n12620), .A2(n12746), .ZN(n12747) );
  OAI211_X1 U16161 ( .C1(n12624), .C2(n20973), .A(n12748), .B(n12747), .ZN(
        n14002) );
  AOI22_X1 U16162 ( .A1(n12794), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16163 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U16164 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16165 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U16166 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12749) );
  NAND4_X1 U16167 ( .A1(n12752), .A2(n12751), .A3(n12750), .A4(n12749), .ZN(
        n12758) );
  AOI22_X1 U16168 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16169 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16170 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U16171 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U16172 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12757) );
  OR2_X1 U16173 ( .A1(n12758), .A2(n12757), .ZN(n14493) );
  INV_X1 U16174 ( .A(n14493), .ZN(n14622) );
  OR2_X1 U16175 ( .A1(n12620), .A2(n14622), .ZN(n12759) );
  OAI211_X1 U16176 ( .C1(n12624), .C2(n20975), .A(n12760), .B(n12759), .ZN(
        n14280) );
  NAND2_X1 U16177 ( .A1(n12793), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U16178 ( .A1(n12794), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U16179 ( .A1(n12793), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U16180 ( .A1(n12794), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16181 ( .A1(n12794), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12767) );
  OAI21_X1 U16182 ( .B1(n12624), .B2(n20981), .A(n12767), .ZN(n13333) );
  NAND2_X1 U16183 ( .A1(n12793), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16184 ( .A1(n12794), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U16185 ( .A1(n12793), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16186 ( .A1(n12794), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12772) );
  NAND2_X1 U16187 ( .A1(n12793), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U16188 ( .A1(n12794), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U16189 ( .A1(n12794), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12778) );
  OAI21_X1 U16190 ( .B1(n12624), .B2(n20989), .A(n12778), .ZN(n16529) );
  NAND2_X1 U16191 ( .A1(n12793), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U16192 ( .A1(n12794), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12779) );
  AND2_X1 U16193 ( .A1(n12780), .A2(n12779), .ZN(n16513) );
  NAND2_X1 U16194 ( .A1(n12793), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16195 ( .A1(n12794), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U16196 ( .A1(n12794), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12785) );
  OAI21_X1 U16197 ( .B1(n12624), .B2(n20995), .A(n12785), .ZN(n16483) );
  AOI22_X1 U16198 ( .A1(n12794), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12786) );
  OAI21_X1 U16199 ( .B1(n12624), .B2(n20997), .A(n12786), .ZN(n13265) );
  NAND2_X1 U16200 ( .A1(n12793), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16201 ( .A1(n12794), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12787) );
  NAND2_X1 U16202 ( .A1(n12793), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U16203 ( .A1(n12794), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12789) );
  AND2_X1 U16204 ( .A1(n12790), .A2(n12789), .ZN(n16445) );
  INV_X1 U16205 ( .A(n16445), .ZN(n12791) );
  AOI22_X1 U16206 ( .A1(n12794), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12792) );
  OAI21_X1 U16207 ( .B1(n12624), .B2(n21004), .A(n12792), .ZN(n13381) );
  INV_X1 U16208 ( .A(n13383), .ZN(n12798) );
  NAND2_X1 U16209 ( .A1(n12793), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16210 ( .A1(n12794), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12795) );
  AND2_X1 U16211 ( .A1(n12796), .A2(n12795), .ZN(n13345) );
  INV_X1 U16212 ( .A(n13345), .ZN(n12797) );
  NAND2_X1 U16213 ( .A1(n12798), .A2(n12797), .ZN(n13347) );
  AOI22_X1 U16214 ( .A1(n12794), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12632), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12799) );
  OAI21_X1 U16215 ( .B1(n12624), .B2(n12800), .A(n12799), .ZN(n12801) );
  NAND2_X1 U16216 ( .A1(n12802), .A2(n21078), .ZN(n12803) );
  NAND2_X1 U16217 ( .A1(n12803), .A2(n14258), .ZN(n12804) );
  INV_X1 U16218 ( .A(n12805), .ZN(n12807) );
  INV_X1 U16219 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12806) );
  NOR2_X1 U16220 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n12808) );
  NAND2_X1 U16221 ( .A1(n12123), .A2(n12808), .ZN(n12810) );
  NAND2_X1 U16222 ( .A1(n12810), .A2(n12809), .ZN(n12828) );
  NAND2_X1 U16223 ( .A1(n12827), .A2(n12828), .ZN(n12831) );
  INV_X1 U16224 ( .A(n12811), .ZN(n12813) );
  NOR2_X2 U16225 ( .A1(n12831), .A2(n12824), .ZN(n12823) );
  INV_X1 U16226 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n20265) );
  MUX2_X1 U16227 ( .A(n12816), .B(n20265), .S(n12123), .Z(n12840) );
  INV_X1 U16228 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14017) );
  INV_X1 U16229 ( .A(n12817), .ZN(n12818) );
  MUX2_X1 U16230 ( .A(n14017), .B(n12818), .S(n12991), .Z(n12819) );
  NAND2_X1 U16231 ( .A1(n12820), .A2(n9918), .ZN(n12821) );
  NAND2_X1 U16232 ( .A1(n12849), .A2(n12821), .ZN(n16631) );
  INV_X1 U16233 ( .A(n12823), .ZN(n12841) );
  NAND2_X1 U16234 ( .A1(n12831), .A2(n12824), .ZN(n12825) );
  NAND2_X1 U16235 ( .A1(n12841), .A2(n12825), .ZN(n16641) );
  INV_X1 U16236 ( .A(n12827), .ZN(n12829) );
  INV_X1 U16237 ( .A(n12828), .ZN(n12835) );
  NAND2_X1 U16238 ( .A1(n12829), .A2(n12835), .ZN(n12830) );
  NAND2_X1 U16239 ( .A1(n12831), .A2(n12830), .ZN(n16659) );
  XNOR2_X1 U16240 ( .A(n16659), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13655) );
  INV_X1 U16241 ( .A(n12832), .ZN(n12833) );
  MUX2_X1 U16242 ( .A(P2_EBX_REG_0__SCAN_IN), .B(n12833), .S(n12812), .Z(
        n16679) );
  NAND2_X1 U16243 ( .A1(n16679), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13664) );
  INV_X1 U16244 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13774) );
  NAND3_X1 U16245 ( .A1(n12985), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12834) );
  AND2_X1 U16246 ( .A1(n12835), .A2(n12834), .ZN(n13662) );
  NAND2_X1 U16247 ( .A1(n13662), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12837) );
  INV_X1 U16248 ( .A(n13662), .ZN(n16671) );
  INV_X1 U16249 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21596) );
  AND2_X1 U16250 ( .A1(n16671), .A2(n21596), .ZN(n12836) );
  AOI21_X1 U16251 ( .B1(n13664), .B2(n12837), .A(n12836), .ZN(n13656) );
  NAND2_X1 U16252 ( .A1(n13655), .A2(n13656), .ZN(n14658) );
  INV_X1 U16253 ( .A(n16659), .ZN(n12838) );
  NAND2_X1 U16254 ( .A1(n12838), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12839) );
  AND2_X1 U16255 ( .A1(n14658), .A2(n12839), .ZN(n17122) );
  XNOR2_X1 U16256 ( .A(n12841), .B(n12840), .ZN(n12842) );
  XNOR2_X1 U16257 ( .A(n12842), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17104) );
  INV_X1 U16258 ( .A(n12842), .ZN(n20261) );
  NAND2_X1 U16259 ( .A1(n12843), .A2(n12994), .ZN(n12845) );
  MUX2_X1 U16260 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12844), .S(n12812), .Z(
        n12848) );
  XNOR2_X1 U16261 ( .A(n12849), .B(n12848), .ZN(n16620) );
  INV_X1 U16262 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16263 ( .A1(n12847), .A2(n13492), .ZN(n12846) );
  INV_X1 U16264 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12850) );
  MUX2_X1 U16265 ( .A(n12850), .B(n12822), .S(n12812), .Z(n12855) );
  NAND2_X1 U16266 ( .A1(n12854), .A2(n12855), .ZN(n12851) );
  INV_X1 U16267 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n20231) );
  NOR2_X1 U16268 ( .A1(n12812), .A2(n20231), .ZN(n12852) );
  NAND2_X1 U16269 ( .A1(n12851), .A2(n12852), .ZN(n12853) );
  NAND2_X1 U16270 ( .A1(n12860), .A2(n12853), .ZN(n20230) );
  NOR2_X1 U16271 ( .A1(n20230), .A2(n12994), .ZN(n12895) );
  NAND2_X1 U16272 ( .A1(n12895), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17074) );
  INV_X1 U16273 ( .A(n17074), .ZN(n12858) );
  INV_X1 U16274 ( .A(n12854), .ZN(n12856) );
  XNOR2_X1 U16275 ( .A(n12856), .B(n12855), .ZN(n20247) );
  NAND2_X1 U16276 ( .A1(n20247), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17086) );
  INV_X1 U16277 ( .A(n17086), .ZN(n12857) );
  NOR2_X1 U16278 ( .A1(n12858), .A2(n12857), .ZN(n12859) );
  INV_X1 U16279 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16280 ( .A1(n12905), .A2(n12906), .ZN(n12901) );
  NAND2_X1 U16281 ( .A1(n12985), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12899) );
  INV_X1 U16282 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12861) );
  NOR2_X1 U16283 ( .A1(n12812), .A2(n12861), .ZN(n12889) );
  NOR2_X1 U16284 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n12863) );
  NOR2_X1 U16285 ( .A1(n12812), .A2(n12863), .ZN(n12864) );
  NOR2_X2 U16286 ( .A1(n12888), .A2(n12864), .ZN(n12880) );
  OAI21_X1 U16287 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n12985), .ZN(n12865) );
  NAND2_X1 U16288 ( .A1(n12880), .A2(n12865), .ZN(n12877) );
  INV_X1 U16289 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12866) );
  NOR2_X1 U16290 ( .A1(n12812), .A2(n12866), .ZN(n12878) );
  INV_X1 U16291 ( .A(n12878), .ZN(n12867) );
  INV_X1 U16292 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12869) );
  NOR2_X1 U16293 ( .A1(n12812), .A2(n12869), .ZN(n12874) );
  INV_X1 U16294 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16544) );
  NAND2_X2 U16295 ( .A1(n12949), .A2(n12972), .ZN(n12947) );
  NAND3_X1 U16296 ( .A1(n9761), .A2(n12985), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n12870) );
  AND2_X1 U16297 ( .A1(n12871), .A2(n12870), .ZN(n16551) );
  NAND2_X1 U16298 ( .A1(n16551), .A2(n12822), .ZN(n12925) );
  NAND2_X1 U16299 ( .A1(n12925), .A2(n13453), .ZN(n13444) );
  NAND2_X1 U16300 ( .A1(n12985), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12872) );
  XNOR2_X1 U16301 ( .A(n12876), .B(n12872), .ZN(n16563) );
  NAND2_X1 U16302 ( .A1(n16563), .A2(n12822), .ZN(n12943) );
  NAND2_X1 U16303 ( .A1(n12943), .A2(n13307), .ZN(n13284) );
  NAND2_X1 U16304 ( .A1(n12873), .A2(n12874), .ZN(n12875) );
  AND2_X1 U16305 ( .A1(n12876), .A2(n12875), .ZN(n20139) );
  NAND2_X1 U16306 ( .A1(n20139), .A2(n12822), .ZN(n12927) );
  NAND2_X1 U16307 ( .A1(n12927), .A2(n16952), .ZN(n16955) );
  NAND2_X1 U16308 ( .A1(n12877), .A2(n12878), .ZN(n12879) );
  NAND2_X1 U16309 ( .A1(n12873), .A2(n12879), .ZN(n20154) );
  OR2_X1 U16310 ( .A1(n20154), .A2(n12994), .ZN(n12929) );
  INV_X1 U16311 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21651) );
  NAND2_X1 U16312 ( .A1(n12929), .A2(n21651), .ZN(n16954) );
  NAND2_X1 U16313 ( .A1(n16955), .A2(n16954), .ZN(n13282) );
  INV_X1 U16314 ( .A(n12880), .ZN(n12915) );
  INV_X1 U16315 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n20172) );
  NOR2_X1 U16316 ( .A1(n12991), .A2(n20172), .ZN(n12881) );
  INV_X1 U16317 ( .A(n12972), .ZN(n12959) );
  AOI21_X1 U16318 ( .B1(n12915), .B2(n12881), .A(n12959), .ZN(n12882) );
  NAND2_X1 U16319 ( .A1(n20174), .A2(n12822), .ZN(n12939) );
  INV_X1 U16320 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17243) );
  XNOR2_X1 U16321 ( .A(n12939), .B(n17243), .ZN(n16974) );
  INV_X1 U16322 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12883) );
  NOR2_X1 U16323 ( .A1(n12812), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U16324 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  NAND2_X1 U16325 ( .A1(n12886), .A2(n12877), .ZN(n16569) );
  OR2_X1 U16326 ( .A1(n16569), .A2(n12994), .ZN(n12887) );
  INV_X1 U16327 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U16328 ( .A1(n12887), .A2(n14718), .ZN(n13280) );
  NAND2_X1 U16329 ( .A1(n12903), .A2(n12889), .ZN(n12890) );
  AND2_X1 U16330 ( .A1(n12888), .A2(n12890), .ZN(n16590) );
  NAND2_X1 U16331 ( .A1(n16590), .A2(n12822), .ZN(n12937) );
  INV_X1 U16332 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17274) );
  NAND2_X1 U16333 ( .A1(n12937), .A2(n17274), .ZN(n17008) );
  NAND2_X1 U16334 ( .A1(n12933), .A2(n17319), .ZN(n17045) );
  NAND2_X1 U16335 ( .A1(n12985), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12891) );
  MUX2_X1 U16336 ( .A(n12985), .B(n12891), .S(n12860), .Z(n12893) );
  AND2_X1 U16337 ( .A1(n12893), .A2(n12892), .ZN(n16608) );
  NAND2_X1 U16338 ( .A1(n16608), .A2(n12822), .ZN(n12894) );
  INV_X1 U16339 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17329) );
  NAND2_X1 U16340 ( .A1(n12894), .A2(n17329), .ZN(n17029) );
  INV_X1 U16341 ( .A(n12895), .ZN(n12896) );
  NAND2_X1 U16342 ( .A1(n12896), .A2(n17341), .ZN(n17073) );
  INV_X1 U16343 ( .A(n20247), .ZN(n12897) );
  NAND2_X1 U16344 ( .A1(n12897), .A2(n17357), .ZN(n17085) );
  AND2_X1 U16345 ( .A1(n17073), .A2(n17085), .ZN(n17028) );
  AND2_X1 U16346 ( .A1(n17029), .A2(n17028), .ZN(n12898) );
  AND2_X1 U16347 ( .A1(n17045), .A2(n12898), .ZN(n13273) );
  INV_X1 U16348 ( .A(n12899), .ZN(n12900) );
  NAND2_X1 U16349 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U16350 ( .A1(n12903), .A2(n12902), .ZN(n20200) );
  OR2_X1 U16351 ( .A1(n20200), .A2(n12994), .ZN(n12904) );
  INV_X1 U16352 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17277) );
  NAND2_X1 U16353 ( .A1(n12904), .A2(n17277), .ZN(n17019) );
  INV_X1 U16354 ( .A(n12905), .ZN(n12908) );
  NOR2_X1 U16355 ( .A1(n12812), .A2(n12906), .ZN(n12907) );
  AND2_X1 U16356 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  OR2_X1 U16357 ( .A1(n12910), .A2(n12909), .ZN(n16600) );
  OAI21_X1 U16358 ( .B1(n16600), .B2(n12994), .A(n17302), .ZN(n17031) );
  AND4_X1 U16359 ( .A1(n17008), .A2(n13273), .A3(n17019), .A4(n17031), .ZN(
        n12922) );
  INV_X1 U16360 ( .A(n12888), .ZN(n12912) );
  INV_X1 U16361 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12911) );
  NAND2_X1 U16362 ( .A1(n12912), .A2(n12911), .ZN(n12919) );
  INV_X1 U16363 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12913) );
  NOR2_X1 U16364 ( .A1(n12812), .A2(n12913), .ZN(n12914) );
  NAND2_X1 U16365 ( .A1(n12919), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U16366 ( .A1(n12916), .A2(n12915), .ZN(n16577) );
  OR2_X1 U16367 ( .A1(n16577), .A2(n12994), .ZN(n12917) );
  NAND2_X1 U16368 ( .A1(n12917), .A2(n17250), .ZN(n16984) );
  NAND2_X1 U16369 ( .A1(n12985), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12918) );
  MUX2_X1 U16370 ( .A(n12985), .B(n12918), .S(n12888), .Z(n12920) );
  NAND2_X1 U16371 ( .A1(n20189), .A2(n12822), .ZN(n12921) );
  NAND2_X1 U16372 ( .A1(n12921), .A2(n17268), .ZN(n13276) );
  NAND4_X1 U16373 ( .A1(n13280), .A2(n12922), .A3(n16984), .A4(n13276), .ZN(
        n12923) );
  NOR3_X1 U16374 ( .A1(n13282), .A2(n16974), .A3(n12923), .ZN(n12924) );
  INV_X1 U16375 ( .A(n12925), .ZN(n12926) );
  NAND2_X1 U16376 ( .A1(n12926), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13445) );
  INV_X1 U16377 ( .A(n12927), .ZN(n12928) );
  INV_X1 U16378 ( .A(n12929), .ZN(n12930) );
  NAND2_X1 U16379 ( .A1(n12930), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13328) );
  AND2_X1 U16380 ( .A1(n12822), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12931) );
  NAND2_X1 U16381 ( .A1(n20189), .A2(n12931), .ZN(n16985) );
  OR3_X1 U16382 ( .A1(n16577), .A2(n12994), .A3(n17250), .ZN(n16983) );
  AND2_X1 U16383 ( .A1(n16985), .A2(n16983), .ZN(n13277) );
  NAND2_X1 U16384 ( .A1(n12822), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12932) );
  OR2_X1 U16385 ( .A1(n16569), .A2(n12932), .ZN(n13279) );
  INV_X1 U16386 ( .A(n12933), .ZN(n12934) );
  NAND2_X1 U16387 ( .A1(n12934), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17046) );
  AND2_X1 U16388 ( .A1(n12822), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12935) );
  NAND2_X1 U16389 ( .A1(n16608), .A2(n12935), .ZN(n17043) );
  NAND2_X1 U16390 ( .A1(n17046), .A2(n17043), .ZN(n17030) );
  NAND2_X1 U16391 ( .A1(n12822), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12936) );
  NOR2_X1 U16392 ( .A1(n16600), .A2(n12936), .ZN(n17032) );
  OR3_X1 U16393 ( .A1(n20200), .A2(n12994), .A3(n17277), .ZN(n17018) );
  INV_X1 U16394 ( .A(n12937), .ZN(n12938) );
  NAND2_X1 U16395 ( .A1(n12938), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17009) );
  AND4_X1 U16396 ( .A1(n13279), .A2(n17017), .A3(n17018), .A4(n17009), .ZN(
        n12941) );
  INV_X1 U16397 ( .A(n12939), .ZN(n12940) );
  NAND2_X1 U16398 ( .A1(n12940), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13278) );
  NAND4_X1 U16399 ( .A1(n13328), .A2(n13277), .A3(n12941), .A4(n13278), .ZN(
        n12942) );
  NOR2_X1 U16400 ( .A1(n13281), .A2(n12942), .ZN(n12945) );
  INV_X1 U16401 ( .A(n12943), .ZN(n12944) );
  NAND2_X1 U16402 ( .A1(n12944), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13442) );
  AND3_X1 U16403 ( .A1(n13445), .A2(n12945), .A3(n13442), .ZN(n12946) );
  NAND2_X1 U16404 ( .A1(n12985), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12948) );
  NAND2_X1 U16405 ( .A1(n12949), .A2(n10379), .ZN(n12950) );
  NAND2_X1 U16406 ( .A1(n12957), .A2(n12950), .ZN(n16533) );
  OR2_X1 U16407 ( .A1(n16533), .A2(n12994), .ZN(n12951) );
  NAND2_X1 U16408 ( .A1(n12951), .A2(n17214), .ZN(n16933) );
  NAND2_X1 U16409 ( .A1(n12985), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12955) );
  XNOR2_X1 U16410 ( .A(n12957), .B(n12955), .ZN(n16526) );
  NAND2_X1 U16411 ( .A1(n16526), .A2(n12822), .ZN(n12953) );
  XNOR2_X1 U16412 ( .A(n12953), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16930) );
  OR2_X1 U16413 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  INV_X1 U16414 ( .A(n12955), .ZN(n12956) );
  INV_X1 U16415 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12958) );
  NOR2_X1 U16416 ( .A1(n12991), .A2(n12958), .ZN(n12960) );
  AOI21_X1 U16417 ( .B1(n9811), .B2(n12960), .A(n12959), .ZN(n12961) );
  NAND2_X1 U16418 ( .A1(n12961), .A2(n16489), .ZN(n16508) );
  NOR2_X1 U16419 ( .A1(n16508), .A2(n12994), .ZN(n12962) );
  AND2_X1 U16420 ( .A1(n12962), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16919) );
  INV_X1 U16421 ( .A(n12962), .ZN(n12963) );
  NAND2_X1 U16422 ( .A1(n12963), .A2(n17181), .ZN(n16920) );
  NOR2_X1 U16423 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n12964) );
  NAND2_X1 U16424 ( .A1(n12965), .A2(n12964), .ZN(n12968) );
  NAND2_X1 U16425 ( .A1(n12985), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12966) );
  INV_X1 U16426 ( .A(n12966), .ZN(n12967) );
  NAND2_X1 U16427 ( .A1(n12968), .A2(n12967), .ZN(n12969) );
  NAND2_X1 U16428 ( .A1(n12979), .A2(n12969), .ZN(n16872) );
  NOR2_X1 U16429 ( .A1(n16872), .A2(n12994), .ZN(n16885) );
  NOR2_X1 U16430 ( .A1(n17140), .A2(n17152), .ZN(n12973) );
  INV_X1 U16431 ( .A(n12992), .ZN(n12971) );
  OAI211_X1 U16432 ( .C1(n16489), .C2(P2_EBX_REG_25__SCAN_IN), .A(n12985), .B(
        P2_EBX_REG_26__SCAN_IN), .ZN(n12970) );
  NAND2_X1 U16433 ( .A1(n12971), .A2(n12970), .ZN(n16479) );
  NAND2_X1 U16434 ( .A1(n12972), .A2(n12822), .ZN(n12975) );
  INV_X1 U16435 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17168) );
  NAND2_X1 U16436 ( .A1(n12975), .A2(n17168), .ZN(n16904) );
  OAI211_X1 U16437 ( .C1(n16885), .C2(n12973), .A(n13255), .B(n16904), .ZN(
        n12978) );
  NAND2_X1 U16438 ( .A1(n12974), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13254) );
  INV_X1 U16439 ( .A(n12975), .ZN(n12976) );
  NAND2_X1 U16440 ( .A1(n12976), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16905) );
  OAI21_X1 U16441 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16874), .ZN(n12977) );
  INV_X1 U16442 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12980) );
  NOR2_X1 U16443 ( .A1(n12812), .A2(n12980), .ZN(n12982) );
  XNOR2_X1 U16444 ( .A(n12981), .B(n12982), .ZN(n16440) );
  INV_X1 U16445 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13387) );
  OAI21_X1 U16446 ( .B1(n16440), .B2(n12994), .A(n13387), .ZN(n13185) );
  INV_X1 U16447 ( .A(n12982), .ZN(n12983) );
  NAND2_X1 U16448 ( .A1(n12984), .A2(n12983), .ZN(n12989) );
  NAND2_X1 U16449 ( .A1(n12985), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12986) );
  XNOR2_X1 U16450 ( .A(n12989), .B(n12986), .ZN(n15162) );
  AOI21_X1 U16451 ( .B1(n15162), .B2(n12822), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13355) );
  AND2_X1 U16452 ( .A1(n12822), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12987) );
  NAND2_X1 U16453 ( .A1(n15162), .A2(n12987), .ZN(n13356) );
  INV_X1 U16454 ( .A(n16440), .ZN(n12988) );
  NAND3_X1 U16455 ( .A1(n12988), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12822), .ZN(n13353) );
  INV_X1 U16456 ( .A(n12989), .ZN(n12990) );
  INV_X1 U16457 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14971) );
  NAND2_X1 U16458 ( .A1(n12990), .A2(n14971), .ZN(n12993) );
  MUX2_X1 U16459 ( .A(n12993), .B(n12992), .S(n12991), .Z(n15189) );
  XNOR2_X1 U16460 ( .A(n12995), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12996) );
  AND2_X1 U16461 ( .A1(n12447), .A2(n12997), .ZN(n21053) );
  OAI211_X1 U16462 ( .C1(n13402), .C2(n20358), .A(n13000), .B(n12999), .ZN(
        P2_U3015) );
  NAND2_X1 U16463 ( .A1(n13001), .A2(n21345), .ZN(n17626) );
  NOR3_X1 U16464 ( .A1(n13004), .A2(n13003), .A3(n13002), .ZN(n13007) );
  OAI21_X1 U16465 ( .B1(n13007), .B2(n13006), .A(n13005), .ZN(n14682) );
  NAND2_X1 U16466 ( .A1(n21434), .A2(n14682), .ZN(n13413) );
  AOI21_X1 U16467 ( .B1(n14691), .B2(n17626), .A(n13413), .ZN(n13012) );
  NAND2_X1 U16468 ( .A1(n14976), .A2(n21434), .ZN(n13008) );
  NAND2_X1 U16469 ( .A1(n13008), .A2(n14697), .ZN(n13010) );
  INV_X1 U16470 ( .A(n17626), .ZN(n14690) );
  OR2_X1 U16471 ( .A1(n14283), .A2(n14690), .ZN(n13009) );
  AOI21_X1 U16472 ( .B1(n13010), .B2(n13009), .A(n13417), .ZN(n13011) );
  NAND3_X1 U16473 ( .A1(n17587), .A2(n13146), .A3(n14691), .ZN(n13021) );
  NAND2_X1 U16474 ( .A1(n13013), .A2(n13409), .ZN(n13014) );
  NAND2_X1 U16475 ( .A1(n13014), .A2(n14697), .ZN(n13015) );
  NAND2_X1 U16476 ( .A1(n13015), .A2(n10829), .ZN(n13017) );
  AND2_X1 U16477 ( .A1(n13017), .A2(n13016), .ZN(n13136) );
  NOR2_X1 U16478 ( .A1(n13136), .A2(n13018), .ZN(n13020) );
  OR2_X1 U16479 ( .A1(n10864), .A2(n14697), .ZN(n13019) );
  OR2_X1 U16480 ( .A1(n13020), .A2(n14680), .ZN(n13722) );
  NAND2_X1 U16481 ( .A1(n13021), .A2(n13722), .ZN(n13022) );
  NOR2_X1 U16482 ( .A1(n15477), .A2(n13144), .ZN(n13025) );
  NAND2_X1 U16483 ( .A1(n13146), .A2(n13025), .ZN(n14984) );
  AND2_X1 U16484 ( .A1(n13026), .A2(n14984), .ZN(n13556) );
  INV_X1 U16485 ( .A(n13027), .ZN(n13029) );
  AOI22_X1 U16486 ( .A1(n13029), .A2(n14051), .B1(n13559), .B2(n14691), .ZN(
        n13030) );
  NAND2_X1 U16487 ( .A1(n14680), .A2(n14287), .ZN(n15013) );
  NAND3_X1 U16488 ( .A1(n13556), .A2(n13030), .A3(n15013), .ZN(n13031) );
  NAND2_X1 U16489 ( .A1(n13196), .A2(n13124), .ZN(n13044) );
  AOI22_X1 U16490 ( .A1(n13044), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13040), .ZN(n13195) );
  INV_X1 U16491 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13033) );
  NAND2_X1 U16492 ( .A1(n13047), .A2(n13033), .ZN(n13036) );
  NAND2_X1 U16493 ( .A1(n13124), .A2(n16099), .ZN(n13034) );
  NAND2_X1 U16494 ( .A1(n13036), .A2(n13035), .ZN(n13038) );
  NAND2_X1 U16495 ( .A1(n13124), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13037) );
  OAI21_X1 U16496 ( .B1(n13119), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13037), .ZN(
        n13802) );
  XNOR2_X1 U16497 ( .A(n13038), .B(n13802), .ZN(n13799) );
  INV_X1 U16498 ( .A(n13038), .ZN(n13039) );
  NAND2_X1 U16499 ( .A1(n13124), .A2(n13041), .ZN(n13042) );
  OAI211_X1 U16500 ( .C1(n13040), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13042), .B(
        n13196), .ZN(n13043) );
  OAI21_X1 U16501 ( .B1(n13127), .B2(P1_EBX_REG_2__SCAN_IN), .A(n13043), .ZN(
        n13876) );
  MUX2_X1 U16502 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13046) );
  NOR2_X1 U16503 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13045) );
  NOR2_X1 U16504 ( .A1(n13046), .A2(n13045), .ZN(n13965) );
  NAND2_X1 U16505 ( .A1(n13874), .A2(n13965), .ZN(n13964) );
  INV_X2 U16506 ( .A(n13964), .ZN(n13053) );
  INV_X1 U16507 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U16508 ( .A1(n13047), .A2(n13048), .ZN(n13051) );
  OAI21_X1 U16509 ( .B1(n13119), .B2(n17658), .A(n13124), .ZN(n13049) );
  OAI21_X1 U16510 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n13040), .A(n13049), .ZN(
        n13050) );
  AND2_X1 U16511 ( .A1(n13051), .A2(n13050), .ZN(n14376) );
  INV_X1 U16512 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16513 ( .A1(n13120), .A2(n13054), .ZN(n13057) );
  NAND2_X1 U16514 ( .A1(n13196), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13055) );
  OAI211_X1 U16515 ( .C1(n13040), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13055), .B(
        n13124), .ZN(n13056) );
  NAND2_X1 U16516 ( .A1(n13057), .A2(n13056), .ZN(n14334) );
  INV_X1 U16517 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21646) );
  NAND2_X1 U16518 ( .A1(n13120), .A2(n21646), .ZN(n13060) );
  NAND2_X1 U16519 ( .A1(n13196), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13058) );
  OAI211_X1 U16520 ( .C1(n13040), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13058), .B(
        n13124), .ZN(n13059) );
  AND2_X1 U16521 ( .A1(n13060), .A2(n13059), .ZN(n15548) );
  OAI21_X1 U16522 ( .B1(n13119), .B2(n21461), .A(n13124), .ZN(n13061) );
  OAI21_X1 U16523 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n13040), .A(n13061), .ZN(
        n13062) );
  OAI21_X1 U16524 ( .B1(n13127), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13062), .ZN(
        n15549) );
  INV_X1 U16525 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17682) );
  OAI21_X1 U16526 ( .B1(n13119), .B2(n17682), .A(n13124), .ZN(n13063) );
  OAI21_X1 U16527 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n13040), .A(n13063), .ZN(
        n13064) );
  OAI21_X1 U16528 ( .B1(n13127), .B2(P1_EBX_REG_8__SCAN_IN), .A(n13064), .ZN(
        n15458) );
  INV_X1 U16529 ( .A(n15456), .ZN(n13070) );
  INV_X1 U16530 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U16531 ( .A1(n13120), .A2(n13065), .ZN(n13068) );
  NAND2_X1 U16532 ( .A1(n13196), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13066) );
  OAI211_X1 U16533 ( .C1(n13040), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13066), .B(
        n13124), .ZN(n13067) );
  NAND2_X1 U16534 ( .A1(n13068), .A2(n13067), .ZN(n15540) );
  NAND2_X1 U16535 ( .A1(n13070), .A2(n13069), .ZN(n15532) );
  INV_X1 U16536 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n17642) );
  NAND2_X1 U16537 ( .A1(n13047), .A2(n17642), .ZN(n13073) );
  INV_X1 U16538 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U16539 ( .A1(n13124), .A2(n16059), .ZN(n13071) );
  OAI211_X1 U16540 ( .C1(n13040), .C2(P1_EBX_REG_10__SCAN_IN), .A(n13071), .B(
        n13196), .ZN(n13072) );
  AND2_X1 U16541 ( .A1(n13073), .A2(n13072), .ZN(n15533) );
  MUX2_X1 U16542 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13075) );
  NOR2_X1 U16543 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13074) );
  NOR2_X1 U16544 ( .A1(n13075), .A2(n13074), .ZN(n15527) );
  MUX2_X1 U16545 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13077) );
  NOR2_X1 U16546 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13076) );
  NOR2_X1 U16547 ( .A1(n13077), .A2(n13076), .ZN(n15425) );
  NAND2_X1 U16548 ( .A1(n13124), .A2(n16040), .ZN(n13078) );
  OAI211_X1 U16549 ( .C1(n13040), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13078), .B(
        n13196), .ZN(n13079) );
  OAI21_X1 U16550 ( .B1(n13127), .B2(P1_EBX_REG_12__SCAN_IN), .A(n13079), .ZN(
        n15440) );
  AND2_X1 U16551 ( .A1(n15425), .A2(n15440), .ZN(n13080) );
  INV_X1 U16552 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15518) );
  NAND2_X1 U16553 ( .A1(n13047), .A2(n15518), .ZN(n13083) );
  NAND2_X1 U16554 ( .A1(n13124), .A2(n15970), .ZN(n13081) );
  OAI211_X1 U16555 ( .C1(n13040), .C2(P1_EBX_REG_14__SCAN_IN), .A(n13081), .B(
        n13196), .ZN(n13082) );
  AND2_X1 U16556 ( .A1(n13083), .A2(n13082), .ZN(n15409) );
  MUX2_X1 U16557 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13084) );
  INV_X1 U16558 ( .A(n13084), .ZN(n13086) );
  INV_X1 U16559 ( .A(n13044), .ZN(n13804) );
  NAND2_X1 U16560 ( .A1(n13804), .A2(n16007), .ZN(n13085) );
  NAND2_X1 U16561 ( .A1(n13086), .A2(n13085), .ZN(n15395) );
  NAND2_X1 U16562 ( .A1(n13124), .A2(n15771), .ZN(n13088) );
  OAI211_X1 U16563 ( .C1(n13040), .C2(P1_EBX_REG_16__SCAN_IN), .A(n13088), .B(
        n13196), .ZN(n13089) );
  OAI21_X1 U16564 ( .B1(n13127), .B2(P1_EBX_REG_16__SCAN_IN), .A(n13089), .ZN(
        n15379) );
  MUX2_X1 U16565 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13091) );
  NOR2_X1 U16566 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13090) );
  NOR2_X1 U16567 ( .A1(n13091), .A2(n13090), .ZN(n15363) );
  NAND2_X1 U16568 ( .A1(n15362), .A2(n15363), .ZN(n15350) );
  INV_X1 U16569 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n13092) );
  NAND2_X1 U16570 ( .A1(n13047), .A2(n13092), .ZN(n13095) );
  INV_X1 U16571 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U16572 ( .A1(n13124), .A2(n15977), .ZN(n13093) );
  OAI211_X1 U16573 ( .C1(n13040), .C2(P1_EBX_REG_18__SCAN_IN), .A(n13093), .B(
        n13196), .ZN(n13094) );
  MUX2_X1 U16574 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13096) );
  INV_X1 U16575 ( .A(n13096), .ZN(n13098) );
  NAND2_X1 U16576 ( .A1(n13804), .A2(n15947), .ZN(n13097) );
  NAND2_X1 U16577 ( .A1(n13098), .A2(n13097), .ZN(n15338) );
  INV_X1 U16578 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U16579 ( .A1(n13047), .A2(n15510), .ZN(n13102) );
  OAI21_X1 U16580 ( .B1(n13119), .B2(n15946), .A(n13124), .ZN(n13100) );
  OAI21_X1 U16581 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n13040), .A(n13100), .ZN(
        n13101) );
  MUX2_X1 U16582 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13104) );
  NOR2_X1 U16583 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13103) );
  NOR2_X1 U16584 ( .A1(n13104), .A2(n13103), .ZN(n15313) );
  INV_X1 U16585 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U16586 ( .A1(n13047), .A2(n13105), .ZN(n13109) );
  INV_X1 U16587 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U16588 ( .A1(n13124), .A2(n13106), .ZN(n13107) );
  OAI211_X1 U16589 ( .C1(n13040), .C2(P1_EBX_REG_22__SCAN_IN), .A(n13107), .B(
        n13196), .ZN(n13108) );
  MUX2_X1 U16590 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13110) );
  INV_X1 U16591 ( .A(n13110), .ZN(n13111) );
  OAI21_X1 U16592 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13044), .A(
        n13111), .ZN(n15290) );
  INV_X1 U16593 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21683) );
  NAND2_X1 U16594 ( .A1(n13124), .A2(n21683), .ZN(n13112) );
  OAI211_X1 U16595 ( .C1(n13040), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13112), .B(
        n13196), .ZN(n13113) );
  OAI21_X1 U16596 ( .B1(n13127), .B2(P1_EBX_REG_24__SCAN_IN), .A(n13113), .ZN(
        n15282) );
  NAND2_X1 U16597 ( .A1(n15291), .A2(n15282), .ZN(n15266) );
  MUX2_X1 U16598 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13114) );
  INV_X1 U16599 ( .A(n13114), .ZN(n13115) );
  OAI21_X1 U16600 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13044), .A(
        n13115), .ZN(n15267) );
  NAND2_X1 U16601 ( .A1(n13047), .A2(n21681), .ZN(n13118) );
  NAND2_X1 U16602 ( .A1(n13124), .A2(n15690), .ZN(n13116) );
  OAI211_X1 U16603 ( .C1(n13040), .C2(P1_EBX_REG_26__SCAN_IN), .A(n13116), .B(
        n13196), .ZN(n13117) );
  MUX2_X1 U16604 ( .A(n13120), .B(n13119), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13122) );
  NOR2_X1 U16605 ( .A1(n13044), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13121) );
  NOR2_X1 U16606 ( .A1(n13122), .A2(n13121), .ZN(n15241) );
  NAND2_X1 U16607 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  OAI211_X1 U16608 ( .C1(n13040), .C2(P1_EBX_REG_28__SCAN_IN), .A(n13125), .B(
        n13196), .ZN(n13126) );
  OAI21_X1 U16609 ( .B1(n13127), .B2(P1_EBX_REG_28__SCAN_IN), .A(n13126), .ZN(
        n15227) );
  INV_X1 U16610 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U16611 ( .A1(n13800), .A2(n15500), .ZN(n13128) );
  OAI21_X1 U16612 ( .B1(n13044), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13128), .ZN(n13129) );
  MUX2_X1 U16613 ( .A(n13129), .B(n13128), .S(n13119), .Z(n15214) );
  NOR2_X4 U16614 ( .A1(n9773), .A2(n15214), .ZN(n15216) );
  OAI22_X1 U16615 ( .A1(n15216), .A2(n13196), .B1(n13129), .B2(n9773), .ZN(
        n13130) );
  NAND2_X1 U16616 ( .A1(n14976), .A2(n11047), .ZN(n13672) );
  OAI21_X1 U16617 ( .B1(n13027), .B2(n14051), .A(n13672), .ZN(n13131) );
  NAND2_X1 U16618 ( .A1(n13044), .A2(n13144), .ZN(n13133) );
  NAND2_X1 U16619 ( .A1(n10878), .A2(n14691), .ZN(n13132) );
  OAI211_X1 U16620 ( .C1(n13134), .C2(n15466), .A(n13133), .B(n13132), .ZN(
        n13135) );
  NOR2_X1 U16621 ( .A1(n13136), .A2(n13135), .ZN(n13138) );
  AND2_X1 U16622 ( .A1(n13138), .A2(n13137), .ZN(n14981) );
  OAI211_X1 U16623 ( .C1(n14697), .C2(n14975), .A(n14981), .B(n13139), .ZN(
        n13140) );
  NAND2_X1 U16624 ( .A1(n13151), .A2(n13140), .ZN(n13166) );
  NAND2_X1 U16625 ( .A1(n13151), .A2(n16090), .ZN(n13906) );
  NAND2_X1 U16626 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17674) );
  NOR2_X1 U16627 ( .A1(n17674), .A2(n21461), .ZN(n16054) );
  AND2_X1 U16628 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13141) );
  AND2_X1 U16629 ( .A1(n16054), .A2(n13141), .ZN(n16033) );
  NAND2_X1 U16630 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14427) );
  NOR2_X1 U16631 ( .A1(n17695), .A2(n14427), .ZN(n14429) );
  NAND2_X1 U16632 ( .A1(n16033), .A2(n14429), .ZN(n16024) );
  AND2_X1 U16633 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13147) );
  NOR2_X1 U16634 ( .A1(n13041), .A2(n16099), .ZN(n13983) );
  NAND2_X1 U16635 ( .A1(n13147), .A2(n13983), .ZN(n13142) );
  OR2_X1 U16636 ( .A1(n16024), .A2(n13142), .ZN(n15966) );
  INV_X1 U16637 ( .A(n15966), .ZN(n13143) );
  NAND2_X1 U16638 ( .A1(n16031), .A2(n13143), .ZN(n13148) );
  NOR2_X1 U16639 ( .A1(n13040), .A2(n13144), .ZN(n13145) );
  NAND2_X1 U16640 ( .A1(n13146), .A2(n13145), .ZN(n14985) );
  INV_X1 U16641 ( .A(n14985), .ZN(n13727) );
  NAND2_X1 U16642 ( .A1(n16033), .A2(n13147), .ZN(n16009) );
  OAI21_X1 U16643 ( .B1(n15090), .B2(n16099), .A(n13041), .ZN(n16025) );
  NAND2_X1 U16644 ( .A1(n14429), .A2(n16025), .ZN(n16052) );
  NOR2_X1 U16645 ( .A1(n16009), .A2(n16052), .ZN(n13153) );
  NAND2_X1 U16646 ( .A1(n16027), .A2(n13153), .ZN(n15944) );
  NAND2_X1 U16647 ( .A1(n13148), .A2(n15944), .ZN(n16020) );
  NAND2_X1 U16648 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15971) );
  NOR2_X1 U16649 ( .A1(n15971), .A2(n15977), .ZN(n13149) );
  AND3_X1 U16650 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15973) );
  AND2_X1 U16651 ( .A1(n13149), .A2(n15973), .ZN(n13157) );
  NAND2_X1 U16652 ( .A1(n16020), .A2(n13157), .ZN(n15958) );
  INV_X1 U16653 ( .A(n15943), .ZN(n13158) );
  NAND2_X1 U16654 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13161) );
  INV_X1 U16655 ( .A(n15891), .ZN(n15687) );
  NAND2_X1 U16656 ( .A1(n15687), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13150) );
  NOR2_X1 U16657 ( .A1(n15908), .A2(n13150), .ZN(n15873) );
  NAND3_X1 U16658 ( .A1(n15873), .A2(n10100), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13204) );
  INV_X1 U16659 ( .A(n13204), .ZN(n13169) );
  AND2_X2 U16660 ( .A1(n13155), .A2(n15969), .ZN(n16030) );
  INV_X1 U16661 ( .A(n13151), .ZN(n13152) );
  NAND2_X1 U16662 ( .A1(n13152), .A2(n17669), .ZN(n13904) );
  OAI21_X1 U16663 ( .B1(n13166), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13904), .ZN(n13159) );
  NOR2_X1 U16664 ( .A1(n15969), .A2(n13153), .ZN(n13154) );
  NOR2_X1 U16665 ( .A1(n13159), .A2(n13154), .ZN(n15968) );
  NAND2_X1 U16666 ( .A1(n15965), .A2(n15966), .ZN(n13156) );
  OAI211_X1 U16667 ( .C1(n16030), .C2(n13157), .A(n15968), .B(n13156), .ZN(
        n15961) );
  OR2_X1 U16668 ( .A1(n15961), .A2(n13158), .ZN(n13160) );
  INV_X1 U16669 ( .A(n13159), .ZN(n13871) );
  NAND2_X1 U16670 ( .A1(n16030), .A2(n13871), .ZN(n16056) );
  NAND2_X1 U16671 ( .A1(n17673), .A2(n13161), .ZN(n13162) );
  NAND2_X1 U16672 ( .A1(n16027), .A2(n10347), .ZN(n13163) );
  NAND2_X1 U16673 ( .A1(n15969), .A2(n13166), .ZN(n21253) );
  NAND2_X1 U16674 ( .A1(n21253), .A2(n21683), .ZN(n13165) );
  INV_X1 U16675 ( .A(n13906), .ZN(n21255) );
  NAND2_X1 U16676 ( .A1(n21255), .A2(n15891), .ZN(n13164) );
  OAI211_X1 U16677 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n13166), .A(
        n13165), .B(n13164), .ZN(n13167) );
  NOR2_X1 U16678 ( .A1(n15901), .A2(n17673), .ZN(n13203) );
  INV_X1 U16679 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15889) );
  NOR3_X1 U16680 ( .A1(n15901), .A2(n15889), .A3(n15690), .ZN(n13168) );
  OAI21_X1 U16681 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13169), .A(
        n13207), .ZN(n13170) );
  OAI211_X1 U16682 ( .C1(n15212), .C2(n16051), .A(n13171), .B(n13170), .ZN(
        n13172) );
  INV_X1 U16683 ( .A(n13172), .ZN(n13173) );
  OAI21_X1 U16684 ( .B1(n13174), .B2(n16064), .A(n13173), .ZN(P1_U3001) );
  AOI21_X1 U16685 ( .B1(n16870), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13176) );
  NOR2_X2 U16686 ( .A1(n13176), .A2(n13344), .ZN(n13378) );
  AND2_X1 U16687 ( .A1(n21077), .A2(n20929), .ZN(n13177) );
  INV_X1 U16688 ( .A(n13522), .ZN(n13186) );
  NAND2_X1 U16689 ( .A1(n13378), .A2(n17718), .ZN(n13189) );
  NAND2_X1 U16690 ( .A1(n21025), .A2(n21065), .ZN(n21040) );
  NAND2_X1 U16691 ( .A1(n21040), .A2(n21075), .ZN(n13180) );
  NOR2_X1 U16692 ( .A1(n17409), .A2(n20814), .ZN(n21041) );
  NAND2_X1 U16693 ( .A1(n15113), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15118) );
  NAND2_X1 U16694 ( .A1(n15119), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15121) );
  NAND2_X1 U16695 ( .A1(n15146), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15145) );
  OR2_X1 U16696 ( .A1(n15152), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13182) );
  NAND2_X1 U16697 ( .A1(n9814), .A2(n13182), .ZN(n16434) );
  NAND2_X1 U16698 ( .A1(n20814), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15154) );
  NAND2_X1 U16699 ( .A1(n13833), .A2(n15154), .ZN(n13564) );
  NAND2_X1 U16700 ( .A1(n20263), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n13386) );
  NAND2_X1 U16701 ( .A1(n17109), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13183) );
  OAI211_X1 U16702 ( .C1(n16434), .C2(n17112), .A(n13386), .B(n13183), .ZN(
        n13184) );
  AOI21_X1 U16703 ( .B1(n16690), .B2(n17716), .A(n13184), .ZN(n13187) );
  INV_X1 U16704 ( .A(n17719), .ZN(n17136) );
  NAND2_X1 U16705 ( .A1(n13189), .A2(n13188), .ZN(P2_U2985) );
  NAND2_X1 U16706 ( .A1(n13191), .A2(n13190), .ZN(n13194) );
  NAND2_X1 U16707 ( .A1(n13192), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13193) );
  NAND2_X1 U16708 ( .A1(n13469), .A2(n21251), .ZN(n13211) );
  NAND2_X1 U16709 ( .A1(n15216), .A2(n13195), .ZN(n13198) );
  AOI22_X1 U16710 ( .A1(n13044), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13040), .ZN(n13199) );
  INV_X1 U16711 ( .A(n13199), .ZN(n13200) );
  INV_X1 U16712 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13202) );
  NOR2_X1 U16713 ( .A1(n13203), .A2(n13202), .ZN(n13206) );
  NOR3_X1 U16714 ( .A1(n13204), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13190), .ZN(n13205) );
  INV_X1 U16715 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21409) );
  NOR2_X1 U16716 ( .A1(n17669), .A2(n21409), .ZN(n13466) );
  NOR2_X1 U16717 ( .A1(n10445), .A2(n13209), .ZN(n13210) );
  NAND2_X1 U16718 ( .A1(n13211), .A2(n13210), .ZN(P1_U3000) );
  XNOR2_X1 U16719 ( .A(n19174), .B(n17578), .ZN(n13500) );
  NAND2_X1 U16720 ( .A1(n17512), .A2(n17584), .ZN(n17738) );
  NAND2_X1 U16721 ( .A1(n13215), .A2(n13243), .ZN(n13239) );
  NAND2_X1 U16722 ( .A1(n13216), .A2(n17584), .ZN(n17740) );
  NAND2_X1 U16723 ( .A1(n13218), .A2(n13217), .ZN(n13220) );
  AOI21_X1 U16724 ( .B1(n13220), .B2(n17852), .A(n13219), .ZN(n13930) );
  AOI21_X1 U16725 ( .B1(n19508), .B2(n13221), .A(n13994), .ZN(n13225) );
  INV_X1 U16726 ( .A(n13222), .ZN(n13223) );
  NOR2_X1 U16727 ( .A1(n19947), .A2(n13223), .ZN(n13224) );
  NOR2_X1 U16728 ( .A1(n13225), .A2(n13224), .ZN(n13230) );
  OAI21_X1 U16729 ( .B1(n19500), .B2(n20089), .A(n19992), .ZN(n13226) );
  OAI21_X1 U16730 ( .B1(n13227), .B2(n13226), .A(n20083), .ZN(n13228) );
  INV_X1 U16731 ( .A(n13228), .ZN(n17851) );
  NAND3_X1 U16732 ( .A1(n13930), .A2(n13230), .A3(n10456), .ZN(n13231) );
  INV_X1 U16733 ( .A(n19253), .ZN(n19469) );
  NOR2_X1 U16734 ( .A1(n19949), .A2(n19469), .ZN(n19398) );
  NAND3_X1 U16735 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U16736 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13888) );
  NOR2_X1 U16737 ( .A1(n13819), .A2(n13888), .ZN(n13812) );
  NAND4_X1 U16738 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n13812), .ZN(n19318) );
  NOR2_X1 U16739 ( .A1(n19055), .A2(n19318), .ZN(n19254) );
  NOR3_X1 U16740 ( .A1(n19250), .A2(n18957), .A3(n19235), .ZN(n18921) );
  NAND2_X1 U16741 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18921), .ZN(
        n17508) );
  INV_X1 U16742 ( .A(n13502), .ZN(n19245) );
  INV_X1 U16743 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19472) );
  NOR2_X1 U16744 ( .A1(n19472), .A2(n19318), .ZN(n19407) );
  NAND2_X1 U16745 ( .A1(n19296), .A2(n19407), .ZN(n19321) );
  NOR2_X1 U16746 ( .A1(n19245), .A2(n19321), .ZN(n17510) );
  NOR2_X1 U16747 ( .A1(n17508), .A2(n19225), .ZN(n13503) );
  AOI21_X1 U16748 ( .B1(n17510), .B2(n13503), .A(n19406), .ZN(n13234) );
  INV_X1 U16749 ( .A(n19949), .ZN(n14106) );
  INV_X1 U16750 ( .A(n19037), .ZN(n19302) );
  AOI21_X1 U16751 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13886) );
  INV_X1 U16752 ( .A(n13819), .ZN(n13232) );
  NAND4_X1 U16753 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n13232), .ZN(n19294) );
  NOR2_X1 U16754 ( .A1(n13886), .A2(n19294), .ZN(n19317) );
  NAND2_X1 U16755 ( .A1(n19296), .A2(n19317), .ZN(n13242) );
  OAI21_X1 U16756 ( .B1(n19302), .B2(n13242), .A(n19949), .ZN(n19255) );
  OAI21_X1 U16757 ( .B1(n13233), .B2(n14106), .A(n19255), .ZN(n17530) );
  AOI211_X1 U16758 ( .C1(n19949), .C2(n17508), .A(n13234), .B(n17530), .ZN(
        n13235) );
  OAI221_X1 U16759 ( .B1(n19253), .B2(n13236), .C1(n19253), .C2(n19254), .A(
        n13235), .ZN(n17475) );
  INV_X1 U16760 ( .A(n17475), .ZN(n13237) );
  OAI21_X1 U16761 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n19398), .A(
        n13237), .ZN(n17579) );
  AOI211_X1 U16762 ( .C1(n17740), .C2(n19948), .A(n19468), .B(n17579), .ZN(
        n13238) );
  INV_X1 U16763 ( .A(n19948), .ZN(n19384) );
  NAND2_X1 U16764 ( .A1(n13243), .A2(n18769), .ZN(n19381) );
  OAI22_X1 U16765 ( .A1(n19095), .A2(n19384), .B1(n19081), .B2(n19381), .ZN(
        n19295) );
  INV_X1 U16766 ( .A(n19254), .ZN(n19297) );
  AOI21_X1 U16767 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19390), .A(
        n19469), .ZN(n19451) );
  OAI22_X1 U16768 ( .A1(n14106), .A2(n13242), .B1(n19297), .B2(n19451), .ZN(
        n17480) );
  AOI21_X1 U16769 ( .B1(n19295), .B2(n19296), .A(n17480), .ZN(n19262) );
  NOR2_X1 U16770 ( .A1(n19262), .A2(n19459), .ZN(n19267) );
  NAND2_X1 U16771 ( .A1(n19267), .A2(n13502), .ZN(n17506) );
  INV_X1 U16772 ( .A(n17506), .ZN(n13244) );
  AOI22_X1 U16773 ( .A1(n13244), .A2(n13503), .B1(n17575), .B2(n19443), .ZN(
        n13247) );
  NAND3_X1 U16774 ( .A1(n18909), .A2(n19377), .A3(n13500), .ZN(n13246) );
  NAND2_X1 U16775 ( .A1(n19477), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n13506) );
  OAI211_X1 U16776 ( .C1(n13247), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n13246), .B(n13506), .ZN(n13248) );
  INV_X1 U16777 ( .A(n13248), .ZN(n13249) );
  NAND2_X1 U16778 ( .A1(n13252), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17175) );
  NAND2_X1 U16779 ( .A1(n16901), .A2(n17726), .ZN(n13272) );
  INV_X1 U16780 ( .A(n16904), .ZN(n16871) );
  NOR2_X1 U16781 ( .A1(n16484), .A2(n13257), .ZN(n13258) );
  OR2_X1 U16782 ( .A1(n13256), .A2(n13258), .ZN(n16899) );
  NAND2_X1 U16783 ( .A1(n20263), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16894) );
  INV_X1 U16784 ( .A(n13259), .ZN(n17166) );
  OAI211_X1 U16785 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17151), .B(n17166), .ZN(
        n13260) );
  NAND2_X1 U16786 ( .A1(n16894), .A2(n13260), .ZN(n13261) );
  AOI21_X1 U16787 ( .B1(n17164), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13261), .ZN(n13262) );
  OAI21_X1 U16788 ( .B1(n16899), .B2(n17352), .A(n13262), .ZN(n13268) );
  OR2_X1 U16789 ( .A1(n13264), .A2(n13265), .ZN(n13266) );
  NAND2_X1 U16790 ( .A1(n13263), .A2(n13266), .ZN(n16793) );
  NOR2_X1 U16791 ( .A1(n16793), .A2(n17372), .ZN(n13267) );
  NAND2_X1 U16792 ( .A1(n13272), .A2(n13271), .ZN(P2_U3020) );
  AND2_X1 U16793 ( .A1(n13273), .A2(n17031), .ZN(n13274) );
  INV_X1 U16794 ( .A(n17019), .ZN(n17006) );
  INV_X1 U16795 ( .A(n13276), .ZN(n16997) );
  NAND2_X1 U16796 ( .A1(n13280), .A2(n13279), .ZN(n14713) );
  INV_X1 U16797 ( .A(n13443), .ZN(n13286) );
  NAND2_X1 U16798 ( .A1(n16943), .A2(n17383), .ZN(n13315) );
  INV_X1 U16799 ( .A(n17262), .ZN(n13302) );
  INV_X1 U16800 ( .A(n14716), .ZN(n13288) );
  NAND2_X1 U16801 ( .A1(n13290), .A2(n13289), .ZN(n16951) );
  INV_X1 U16802 ( .A(n13292), .ZN(n13293) );
  AOI21_X1 U16803 ( .B1(n13294), .B2(n13291), .A(n13293), .ZN(n16948) );
  NAND2_X1 U16804 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  NAND2_X1 U16805 ( .A1(n13295), .A2(n13298), .ZN(n16839) );
  NOR2_X1 U16806 ( .A1(n16839), .A2(n17372), .ZN(n13310) );
  OAI21_X1 U16807 ( .B1(n17258), .B2(n13299), .A(n17259), .ZN(n17246) );
  AOI21_X1 U16808 ( .B1(n17380), .B2(n13334), .A(n21651), .ZN(n13300) );
  NAND2_X1 U16809 ( .A1(n17246), .A2(n13300), .ZN(n17222) );
  NOR2_X1 U16810 ( .A1(n17333), .A2(n17329), .ZN(n17320) );
  NAND2_X1 U16811 ( .A1(n17320), .A2(n13301), .ZN(n17278) );
  INV_X1 U16812 ( .A(n13334), .ZN(n13303) );
  NAND3_X1 U16813 ( .A1(n13303), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16952), .ZN(n13304) );
  NOR2_X1 U16814 ( .A1(n17238), .A2(n13304), .ZN(n17226) );
  AOI21_X1 U16815 ( .B1(n17259), .B2(n17222), .A(n17226), .ZN(n13308) );
  NOR2_X1 U16816 ( .A1(n12586), .A2(n20985), .ZN(n16944) );
  INV_X1 U16817 ( .A(n16944), .ZN(n13306) );
  NAND3_X1 U16818 ( .A1(n17251), .A2(n13454), .A3(n13307), .ZN(n13305) );
  OAI211_X1 U16819 ( .C1(n13308), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13309) );
  AOI211_X1 U16820 ( .C1(n16948), .C2(n20356), .A(n13310), .B(n13309), .ZN(
        n13311) );
  INV_X1 U16821 ( .A(n13311), .ZN(n13312) );
  NOR2_X1 U16822 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  NAND2_X1 U16823 ( .A1(n13315), .A2(n13314), .ZN(P2_U3026) );
  INV_X1 U16824 ( .A(n16953), .ZN(n13317) );
  AOI21_X1 U16825 ( .B1(n16963), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13316) );
  AND2_X1 U16826 ( .A1(n14630), .A2(n13318), .ZN(n13319) );
  OR2_X1 U16827 ( .A1(n13319), .A2(n16744), .ZN(n20156) );
  NAND2_X1 U16828 ( .A1(n13320), .A2(n13323), .ZN(n13321) );
  AND2_X1 U16829 ( .A1(n15131), .A2(n13321), .ZN(n20148) );
  NOR2_X1 U16830 ( .A1(n12586), .A2(n20981), .ZN(n13336) );
  INV_X1 U16831 ( .A(n13336), .ZN(n13322) );
  OAI21_X1 U16832 ( .B1(n17723), .B2(n13323), .A(n13322), .ZN(n13324) );
  AOI21_X1 U16833 ( .B1(n20148), .B2(n17714), .A(n13324), .ZN(n13325) );
  OAI21_X1 U16834 ( .B1(n20156), .B2(n17098), .A(n13325), .ZN(n13326) );
  AOI21_X1 U16835 ( .B1(n13340), .B2(n17718), .A(n13326), .ZN(n13331) );
  NAND2_X1 U16836 ( .A1(n13328), .A2(n16954), .ZN(n13329) );
  XNOR2_X1 U16837 ( .A(n13327), .B(n13329), .ZN(n13341) );
  NAND2_X1 U16838 ( .A1(n13331), .A2(n13330), .ZN(P2_U2996) );
  OAI21_X1 U16839 ( .B1(n9758), .B2(n13333), .A(n16841), .ZN(n20157) );
  OAI21_X1 U16840 ( .B1(n17238), .B2(n13334), .A(n21651), .ZN(n13337) );
  NOR2_X1 U16841 ( .A1(n20156), .A2(n17352), .ZN(n13335) );
  AOI211_X1 U16842 ( .C1(n17222), .C2(n13337), .A(n13336), .B(n13335), .ZN(
        n13338) );
  OAI21_X1 U16843 ( .B1(n17372), .B2(n20157), .A(n13338), .ZN(n13339) );
  AOI21_X1 U16844 ( .B1(n13340), .B2(n17726), .A(n13339), .ZN(n13343) );
  NAND2_X1 U16845 ( .A1(n13343), .A2(n13342), .ZN(P2_U3028) );
  NAND2_X1 U16846 ( .A1(n13383), .A2(n13345), .ZN(n13346) );
  NAND2_X1 U16847 ( .A1(n20263), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14672) );
  INV_X1 U16848 ( .A(n14672), .ZN(n13350) );
  INV_X1 U16849 ( .A(n17137), .ZN(n13348) );
  OAI21_X1 U16850 ( .B1(n14964), .B2(n17372), .A(n13351), .ZN(n13352) );
  INV_X1 U16851 ( .A(n13352), .ZN(n13363) );
  NAND2_X1 U16852 ( .A1(n13354), .A2(n13353), .ZN(n13359) );
  INV_X1 U16853 ( .A(n13355), .ZN(n13357) );
  NAND2_X1 U16854 ( .A1(n13357), .A2(n13356), .ZN(n13358) );
  OR2_X1 U16855 ( .A1(n15182), .A2(n17352), .ZN(n13362) );
  XNOR2_X1 U16856 ( .A(n13365), .B(n13364), .ZN(n13367) );
  OR2_X1 U16857 ( .A1(n13367), .A2(n13366), .ZN(n13377) );
  NAND2_X1 U16858 ( .A1(n18171), .A2(n13368), .ZN(n17878) );
  NOR2_X1 U16859 ( .A1(n17878), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n13375) );
  OAI22_X1 U16860 ( .A1(n17873), .A2(n20061), .B1(n13369), .B2(n18219), .ZN(
        n13373) );
  OAI21_X1 U16861 ( .B1(n18217), .B2(n13370), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n13371) );
  INV_X1 U16862 ( .A(n13371), .ZN(n13372) );
  NAND2_X1 U16863 ( .A1(n13377), .A2(n13376), .ZN(P3_U2641) );
  NAND2_X1 U16864 ( .A1(n13378), .A2(n17726), .ZN(n13391) );
  INV_X1 U16865 ( .A(n13379), .ZN(n13380) );
  NAND2_X1 U16866 ( .A1(n13380), .A2(n17383), .ZN(n13390) );
  OAI211_X1 U16867 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n17137), .B(n13384), .ZN(
        n13385) );
  OAI211_X1 U16868 ( .C1(n17141), .C2(n13387), .A(n13386), .B(n13385), .ZN(
        n13388) );
  INV_X1 U16869 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13392) );
  NAND2_X1 U16870 ( .A1(n15097), .A2(n17714), .ZN(n13396) );
  AOI21_X1 U16871 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13394), .ZN(n13395) );
  OAI21_X1 U16872 ( .B1(n15183), .B2(n17098), .A(n13397), .ZN(n13398) );
  INV_X1 U16873 ( .A(n13398), .ZN(n13401) );
  NAND2_X1 U16874 ( .A1(n13399), .A2(n17719), .ZN(n13400) );
  OAI211_X1 U16875 ( .C1(n13402), .C2(n17116), .A(n13401), .B(n13400), .ZN(
        P2_U2983) );
  AOI22_X1 U16876 ( .A1(n13406), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13405), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13407) );
  INV_X1 U16877 ( .A(n13559), .ZN(n13408) );
  NAND2_X1 U16878 ( .A1(n14691), .A2(n21434), .ZN(n13411) );
  INV_X1 U16879 ( .A(n14979), .ZN(n13410) );
  NAND4_X1 U16880 ( .A1(n15558), .A2(n13409), .A3(n14679), .A4(n10879), .ZN(
        n13437) );
  OAI22_X1 U16881 ( .A1(n15196), .A2(n13411), .B1(n13410), .B2(n13437), .ZN(
        n13412) );
  INV_X1 U16882 ( .A(n13412), .ZN(n13415) );
  OAI22_X1 U16883 ( .A1(n17587), .A2(n14984), .B1(n13413), .B2(n15013), .ZN(
        n13724) );
  NAND2_X1 U16884 ( .A1(n13724), .A2(n14679), .ZN(n13414) );
  NAND2_X1 U16885 ( .A1(n14678), .A2(n13416), .ZN(n13435) );
  INV_X1 U16886 ( .A(n13417), .ZN(n13429) );
  NOR4_X1 U16887 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13421) );
  NOR4_X1 U16888 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n13420) );
  NOR4_X1 U16889 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13419) );
  NOR4_X1 U16890 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13418) );
  AND4_X1 U16891 ( .A1(n13421), .A2(n13420), .A3(n13419), .A4(n13418), .ZN(
        n13426) );
  NOR4_X1 U16892 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13424) );
  NOR4_X1 U16893 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n13423) );
  NOR4_X1 U16894 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_28__SCAN_IN), .A3(P1_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_ADDRESS_REG_26__SCAN_IN), .ZN(n13422) );
  AND4_X1 U16895 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n21359), .ZN(
        n13425) );
  NAND2_X1 U16896 ( .A1(n13426), .A2(n13425), .ZN(n13427) );
  NOR2_X1 U16897 ( .A1(n13429), .A2(n14022), .ZN(n13428) );
  NAND2_X1 U16898 ( .A1(n15644), .A2(n13428), .ZN(n15611) );
  INV_X1 U16899 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17756) );
  NOR2_X1 U16900 ( .A1(n15611), .A2(n17756), .ZN(n13433) );
  NOR3_X1 U16901 ( .A1(n15637), .A2(n15585), .A3(n13429), .ZN(n13430) );
  AOI22_X1 U16902 ( .A1(n15618), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15637), .ZN(n13431) );
  INV_X1 U16903 ( .A(n13431), .ZN(n13432) );
  NOR2_X1 U16904 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  NAND2_X1 U16905 ( .A1(n13435), .A2(n13434), .ZN(P1_U2873) );
  NOR2_X1 U16906 ( .A1(n14985), .A2(n21089), .ZN(n13436) );
  NAND2_X1 U16907 ( .A1(n17587), .A2(n13436), .ZN(n13440) );
  INV_X1 U16908 ( .A(n13437), .ZN(n13438) );
  INV_X1 U16909 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U16910 ( .A1(n13443), .A2(n13442), .ZN(n13446) );
  NAND2_X1 U16911 ( .A1(n13289), .A2(n13453), .ZN(n14726) );
  NAND3_X1 U16912 ( .A1(n13447), .A2(n17726), .A3(n14726), .ZN(n13462) );
  AND2_X1 U16913 ( .A1(n13292), .A2(n13448), .ZN(n13450) );
  NAND2_X1 U16914 ( .A1(n17258), .A2(n17259), .ZN(n17328) );
  OR2_X1 U16915 ( .A1(n17397), .A2(n13451), .ZN(n13452) );
  NAND2_X1 U16916 ( .A1(n17328), .A2(n13452), .ZN(n17191) );
  NOR2_X1 U16917 ( .A1(n12586), .A2(n20987), .ZN(n14722) );
  AOI21_X1 U16918 ( .B1(n17191), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14722), .ZN(n13456) );
  AND3_X1 U16919 ( .A1(n13454), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n13453), .ZN(n13455) );
  NAND2_X1 U16920 ( .A1(n17251), .A2(n13455), .ZN(n17193) );
  OAI211_X1 U16921 ( .C1(n16738), .C2(n17352), .A(n13456), .B(n17193), .ZN(
        n13457) );
  INV_X1 U16922 ( .A(n13457), .ZN(n13461) );
  NOR2_X1 U16923 ( .A1(n13458), .A2(n10470), .ZN(n16826) );
  NAND2_X1 U16924 ( .A1(n16826), .A2(n20355), .ZN(n13460) );
  AOI21_X1 U16925 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13466), .ZN(n13467) );
  OAI21_X1 U16926 ( .B1(n15203), .B2(n17665), .A(n13467), .ZN(n13468) );
  AOI21_X1 U16927 ( .B1(n14678), .B2(n17654), .A(n13468), .ZN(n13470) );
  NOR2_X1 U16928 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13472) );
  NOR4_X1 U16929 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13471) );
  NAND4_X1 U16930 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13472), .A4(n13471), .ZN(n13485) );
  NOR2_X4 U16931 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13485), .ZN(n17833)
         );
  NOR3_X1 U16932 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21426), .ZN(n13474) );
  NOR4_X1 U16933 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_D_C_N_REG_SCAN_IN), .ZN(n13473) );
  NAND4_X1 U16934 ( .A1(n15585), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13474), .A4(
        n13473), .ZN(U214) );
  NOR4_X1 U16935 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n13478) );
  NOR4_X1 U16936 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n13477) );
  NOR4_X1 U16937 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n13476) );
  NOR4_X1 U16938 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n13475) );
  AND4_X1 U16939 ( .A1(n13478), .A2(n13477), .A3(n13476), .A4(n13475), .ZN(
        n13483) );
  NOR4_X1 U16940 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_3__SCAN_IN), .A4(
        P2_ADDRESS_REG_2__SCAN_IN), .ZN(n13481) );
  NOR4_X1 U16941 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n13480) );
  NOR4_X1 U16942 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U16943 ( .A1(n17755), .A2(U214), .ZN(U212) );
  NOR2_X1 U16944 ( .A1(n20961), .A2(n12586), .ZN(n13498) );
  AOI21_X1 U16945 ( .B1(n13487), .B2(n13486), .A(n14129), .ZN(n16622) );
  INV_X1 U16946 ( .A(n16622), .ZN(n17099) );
  NAND3_X1 U16947 ( .A1(n17730), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17367), .ZN(n13488) );
  NAND2_X1 U16948 ( .A1(n13488), .A2(n17259), .ZN(n17356) );
  OAI22_X1 U16949 ( .A1(n17099), .A2(n17352), .B1(n13492), .B2(n17356), .ZN(
        n13497) );
  XNOR2_X1 U16950 ( .A(n13489), .B(n13760), .ZN(n16625) );
  OAI22_X1 U16951 ( .A1(n17340), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16625), .B2(n17372), .ZN(n13496) );
  OR2_X1 U16952 ( .A1(n13491), .A2(n13490), .ZN(n17071) );
  XNOR2_X1 U16953 ( .A(n17069), .B(n13492), .ZN(n17070) );
  XOR2_X1 U16954 ( .A(n17071), .B(n17070), .Z(n17101) );
  INV_X1 U16955 ( .A(n17101), .ZN(n13494) );
  XNOR2_X1 U16956 ( .A(n13493), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17103) );
  OAI22_X1 U16957 ( .A1(n13494), .A2(n20360), .B1(n17103), .B2(n20358), .ZN(
        n13495) );
  OR4_X1 U16958 ( .A1(n13498), .A2(n13497), .A3(n13496), .A4(n13495), .ZN(
        P2_U3040) );
  INV_X1 U16959 ( .A(n13501), .ZN(n19010) );
  NAND2_X1 U16960 ( .A1(n19048), .A2(n13502), .ZN(n18976) );
  INV_X1 U16961 ( .A(n13503), .ZN(n13504) );
  NOR3_X1 U16962 ( .A1(n18976), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n13504), .ZN(n13515) );
  NAND4_X1 U16963 ( .A1(n19062), .A2(n13505), .A3(n18936), .A4(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18917) );
  XNOR2_X1 U16964 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13513) );
  INV_X1 U16965 ( .A(n13506), .ZN(n13507) );
  AOI21_X1 U16966 ( .B1(n19124), .B2(n10510), .A(n13507), .ZN(n13512) );
  NAND2_X1 U16967 ( .A1(n19059), .A2(n13508), .ZN(n13509) );
  OAI211_X1 U16968 ( .C1(n11964), .C2(n19105), .A(n19202), .B(n13509), .ZN(
        n18926) );
  NOR2_X1 U16969 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17452), .ZN(
        n18929) );
  NOR2_X1 U16970 ( .A1(n18926), .A2(n18929), .ZN(n18915) );
  OR2_X1 U16971 ( .A1(n18915), .A2(n13510), .ZN(n13511) );
  OAI211_X1 U16972 ( .C1(n18917), .C2(n13513), .A(n13512), .B(n13511), .ZN(
        n13514) );
  OAI21_X1 U16973 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13518)
         );
  INV_X1 U16974 ( .A(n14393), .ZN(n13516) );
  NOR2_X1 U16975 ( .A1(n21075), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U16976 ( .A1(n21071), .A2(n13517), .ZN(n14317) );
  INV_X1 U16977 ( .A(n14317), .ZN(n20930) );
  AOI211_X1 U16978 ( .C1(n20864), .C2(n13518), .A(n17411), .B(n20930), .ZN(
        P2_U3178) );
  NOR2_X1 U16979 ( .A1(n9741), .A2(n13521), .ZN(n13687) );
  NAND2_X1 U16980 ( .A1(n13687), .A2(n13523), .ZN(n16664) );
  INV_X1 U16981 ( .A(n16664), .ZN(n20270) );
  INV_X1 U16982 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n21087) );
  NOR2_X1 U16983 ( .A1(n21065), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13526) );
  INV_X1 U16984 ( .A(n13526), .ZN(n13524) );
  OAI211_X1 U16985 ( .C1(n20270), .C2(n21087), .A(n13532), .B(n13524), .ZN(
        P2_U2814) );
  INV_X1 U16986 ( .A(n14204), .ZN(n14220) );
  OAI211_X1 U16987 ( .C1(n13528), .C2(n21071), .A(n12802), .B(n14220), .ZN(
        n13520) );
  NOR2_X1 U16988 ( .A1(n13520), .A2(n14260), .ZN(n14265) );
  NOR2_X1 U16989 ( .A1(n14265), .A2(n13521), .ZN(n21063) );
  OAI21_X1 U16990 ( .B1(n21063), .B2(n12457), .A(n13522), .ZN(P2_U2819) );
  NAND3_X1 U16991 ( .A1(n12802), .A2(n20929), .A3(n13523), .ZN(n21069) );
  INV_X1 U16992 ( .A(n21069), .ZN(n13525) );
  INV_X1 U16993 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n21530) );
  OAI22_X1 U16994 ( .A1(n13525), .A2(n21530), .B1(n21075), .B2(n13524), .ZN(
        P2_U2816) );
  OAI21_X1 U16995 ( .B1(n13526), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n21069), 
        .ZN(n13527) );
  OAI21_X1 U16996 ( .B1(n13528), .B2(n21069), .A(n13527), .ZN(P2_U3612) );
  INV_X1 U16997 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13717) );
  NOR3_X4 U16998 ( .A1(n13532), .A2(n14904), .A3(n21071), .ZN(n13626) );
  INV_X1 U16999 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13529) );
  OR2_X1 U17000 ( .A1(n14505), .A2(n13529), .ZN(n13531) );
  NAND2_X1 U17001 ( .A1(n14505), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13530) );
  NAND2_X1 U17002 ( .A1(n13531), .A2(n13530), .ZN(n16777) );
  NAND2_X1 U17003 ( .A1(n13626), .A2(n16777), .ZN(n20352) );
  INV_X1 U17004 ( .A(n13532), .ZN(n15168) );
  OAI21_X2 U17005 ( .B1(n14904), .B2(n21073), .A(n15168), .ZN(n13623) );
  NAND2_X1 U17006 ( .A1(n13623), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13533) );
  OAI211_X1 U17007 ( .C1(n13717), .C2(n15096), .A(n20352), .B(n13533), .ZN(
        P2_U2964) );
  INV_X1 U17008 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13709) );
  INV_X1 U17009 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13534) );
  OR2_X1 U17010 ( .A1(n14505), .A2(n13534), .ZN(n13536) );
  NAND2_X1 U17011 ( .A1(n14505), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13535) );
  NAND2_X1 U17012 ( .A1(n13536), .A2(n13535), .ZN(n14508) );
  NAND2_X1 U17013 ( .A1(n13626), .A2(n14508), .ZN(n13589) );
  NAND2_X1 U17014 ( .A1(n13623), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13537) );
  OAI211_X1 U17015 ( .C1(n13709), .C2(n15096), .A(n13589), .B(n13537), .ZN(
        P2_U2952) );
  INV_X1 U17016 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13701) );
  INV_X1 U17017 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17789) );
  OR2_X1 U17018 ( .A1(n14505), .A2(n17789), .ZN(n13539) );
  NAND2_X1 U17019 ( .A1(n14505), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U17020 ( .A1(n13539), .A2(n13538), .ZN(n16791) );
  NAND2_X1 U17021 ( .A1(n13626), .A2(n16791), .ZN(n13542) );
  NAND2_X1 U17022 ( .A1(n13623), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13540) );
  OAI211_X1 U17023 ( .C1(n13701), .C2(n15096), .A(n13542), .B(n13540), .ZN(
        P2_U2962) );
  INV_X1 U17024 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20327) );
  NAND2_X1 U17025 ( .A1(n13623), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13541) );
  OAI211_X1 U17026 ( .C1(n20327), .C2(n15096), .A(n13542), .B(n13541), .ZN(
        P2_U2977) );
  INV_X1 U17027 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13695) );
  INV_X1 U17028 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13543) );
  OR2_X1 U17029 ( .A1(n14505), .A2(n13543), .ZN(n13545) );
  NAND2_X1 U17030 ( .A1(n14505), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13544) );
  NAND2_X1 U17031 ( .A1(n13545), .A2(n13544), .ZN(n14965) );
  NAND2_X1 U17032 ( .A1(n13626), .A2(n14965), .ZN(n13548) );
  NAND2_X1 U17033 ( .A1(n13623), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13546) );
  OAI211_X1 U17034 ( .C1(n13695), .C2(n15096), .A(n13548), .B(n13546), .ZN(
        P2_U2966) );
  INV_X1 U17035 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20318) );
  NAND2_X1 U17036 ( .A1(n13623), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13547) );
  OAI211_X1 U17037 ( .C1(n20318), .C2(n15096), .A(n13548), .B(n13547), .ZN(
        P2_U2981) );
  INV_X1 U17038 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13553) );
  INV_X1 U17039 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13552) );
  INV_X1 U17040 ( .A(n13623), .ZN(n13570) );
  INV_X1 U17041 ( .A(n13626), .ZN(n13551) );
  INV_X1 U17042 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13549) );
  NOR2_X1 U17043 ( .A1(n14399), .A2(n13549), .ZN(n13550) );
  AOI21_X1 U17044 ( .B1(BUF1_REG_15__SCAN_IN), .B2(n14399), .A(n13550), .ZN(
        n14281) );
  OAI222_X1 U17045 ( .A1(n15096), .A2(n13553), .B1(n13552), .B2(n13570), .C1(
        n13551), .C2(n14281), .ZN(P2_U2982) );
  AOI21_X1 U17046 ( .B1(n14682), .B2(n14680), .A(n13559), .ZN(n13554) );
  AOI21_X1 U17047 ( .B1(n17587), .B2(n15477), .A(n13554), .ZN(n21088) );
  NAND3_X1 U17048 ( .A1(n15477), .A2(n17626), .A3(n13040), .ZN(n13555) );
  NAND2_X1 U17049 ( .A1(n13555), .A2(n21434), .ZN(n21427) );
  NAND2_X1 U17050 ( .A1(n21088), .A2(n21427), .ZN(n17603) );
  AND2_X1 U17051 ( .A1(n17603), .A2(n14679), .ZN(n21096) );
  INV_X1 U17052 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17604) );
  MUX2_X1 U17053 ( .A(n14985), .B(n13556), .S(n17587), .Z(n13561) );
  INV_X1 U17054 ( .A(n14680), .ZN(n13557) );
  NOR2_X1 U17055 ( .A1(n14682), .A2(n13557), .ZN(n13558) );
  AOI21_X1 U17056 ( .B1(n17587), .B2(n13559), .A(n13558), .ZN(n13560) );
  NAND2_X1 U17057 ( .A1(n13561), .A2(n13560), .ZN(n17605) );
  NAND2_X1 U17058 ( .A1(n21096), .A2(n17605), .ZN(n13562) );
  OAI21_X1 U17059 ( .B1(n21096), .B2(n17604), .A(n13562), .ZN(P1_U3484) );
  XNOR2_X1 U17060 ( .A(n13563), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17395) );
  INV_X1 U17061 ( .A(n17395), .ZN(n13569) );
  OR2_X1 U17062 ( .A1(n17109), .A2(n13564), .ZN(n13565) );
  AOI22_X1 U17063 ( .A1(n17393), .A2(n17716), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13565), .ZN(n13568) );
  OAI21_X1 U17064 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16679), .A(
        n13664), .ZN(n17390) );
  INV_X1 U17065 ( .A(n17390), .ZN(n13566) );
  NOR2_X1 U17066 ( .A1(n20169), .A2(n20123), .ZN(n17392) );
  AOI21_X1 U17067 ( .B1(n17719), .B2(n13566), .A(n17392), .ZN(n13567) );
  OAI211_X1 U17068 ( .C1(n17116), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        P2_U3014) );
  AOI22_X1 U17069 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13574) );
  INV_X1 U17070 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13571) );
  OR2_X1 U17071 ( .A1(n14505), .A2(n13571), .ZN(n13573) );
  NAND2_X1 U17072 ( .A1(n14505), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13572) );
  NAND2_X1 U17073 ( .A1(n13573), .A2(n13572), .ZN(n16769) );
  NAND2_X1 U17074 ( .A1(n13626), .A2(n16769), .ZN(n13598) );
  NAND2_X1 U17075 ( .A1(n13574), .A2(n13598), .ZN(P2_U2965) );
  AOI22_X1 U17076 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13578) );
  INV_X1 U17077 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13575) );
  OR2_X1 U17078 ( .A1(n14505), .A2(n13575), .ZN(n13577) );
  NAND2_X1 U17079 ( .A1(n14505), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13576) );
  AND2_X1 U17080 ( .A1(n13577), .A2(n13576), .ZN(n20388) );
  INV_X1 U17081 ( .A(n20388), .ZN(n16833) );
  NAND2_X1 U17082 ( .A1(n13626), .A2(n16833), .ZN(n13628) );
  NAND2_X1 U17083 ( .A1(n13578), .A2(n13628), .ZN(P2_U2971) );
  AOI22_X1 U17084 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13582) );
  INV_X1 U17085 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13579) );
  OR2_X1 U17086 ( .A1(n14505), .A2(n13579), .ZN(n13581) );
  NAND2_X1 U17087 ( .A1(n14505), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13580) );
  INV_X1 U17088 ( .A(n20305), .ZN(n16842) );
  NAND2_X1 U17089 ( .A1(n13626), .A2(n16842), .ZN(n13591) );
  NAND2_X1 U17090 ( .A1(n13582), .A2(n13591), .ZN(P2_U2970) );
  AOI22_X1 U17091 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13584) );
  INV_X1 U17092 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17801) );
  NOR2_X1 U17093 ( .A1(n14505), .A2(n17801), .ZN(n13583) );
  AOI21_X1 U17094 ( .B1(BUF2_REG_2__SCAN_IN), .B2(n14505), .A(n13583), .ZN(
        n14608) );
  INV_X1 U17095 ( .A(n14608), .ZN(n16849) );
  NAND2_X1 U17096 ( .A1(n13626), .A2(n16849), .ZN(n13593) );
  NAND2_X1 U17097 ( .A1(n13584), .A2(n13593), .ZN(P2_U2969) );
  AOI22_X1 U17098 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13588) );
  INV_X1 U17099 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13585) );
  OR2_X1 U17100 ( .A1(n14505), .A2(n13585), .ZN(n13587) );
  NAND2_X1 U17101 ( .A1(n14505), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13586) );
  AND2_X1 U17102 ( .A1(n13587), .A2(n13586), .ZN(n20380) );
  INV_X1 U17103 ( .A(n20380), .ZN(n16857) );
  NAND2_X1 U17104 ( .A1(n13626), .A2(n16857), .ZN(n13595) );
  NAND2_X1 U17105 ( .A1(n13588), .A2(n13595), .ZN(P2_U2968) );
  AOI22_X1 U17106 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U17107 ( .A1(n13590), .A2(n13589), .ZN(P2_U2967) );
  AOI22_X1 U17108 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13592) );
  NAND2_X1 U17109 ( .A1(n13592), .A2(n13591), .ZN(P2_U2955) );
  AOI22_X1 U17110 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13594) );
  NAND2_X1 U17111 ( .A1(n13594), .A2(n13593), .ZN(P2_U2954) );
  AOI22_X1 U17112 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U17113 ( .A1(n13596), .A2(n13595), .ZN(P2_U2953) );
  AOI22_X1 U17114 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13597) );
  MUX2_X1 U17115 ( .A(BUF1_REG_6__SCAN_IN), .B(BUF2_REG_6__SCAN_IN), .S(n14505), .Z(n16819) );
  NAND2_X1 U17116 ( .A1(n13626), .A2(n16819), .ZN(n13624) );
  NAND2_X1 U17117 ( .A1(n13597), .A2(n13624), .ZN(P2_U2973) );
  AOI22_X1 U17118 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13599) );
  NAND2_X1 U17119 ( .A1(n13599), .A2(n13598), .ZN(P2_U2980) );
  AOI22_X1 U17120 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13603) );
  INV_X1 U17121 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13600) );
  OR2_X1 U17122 ( .A1(n14505), .A2(n13600), .ZN(n13602) );
  NAND2_X1 U17123 ( .A1(n14505), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13601) );
  NAND2_X1 U17124 ( .A1(n13602), .A2(n13601), .ZN(n16812) );
  NAND2_X1 U17125 ( .A1(n13626), .A2(n16812), .ZN(n13621) );
  NAND2_X1 U17126 ( .A1(n13603), .A2(n13621), .ZN(P2_U2974) );
  AOI22_X1 U17127 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13606) );
  INV_X1 U17128 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17791) );
  OR2_X1 U17129 ( .A1(n14505), .A2(n17791), .ZN(n13605) );
  NAND2_X1 U17130 ( .A1(n14505), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13604) );
  NAND2_X1 U17131 ( .A1(n13605), .A2(n13604), .ZN(n16805) );
  NAND2_X1 U17132 ( .A1(n13626), .A2(n16805), .ZN(n13617) );
  NAND2_X1 U17133 ( .A1(n13606), .A2(n13617), .ZN(P2_U2975) );
  AOI22_X1 U17134 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13610) );
  INV_X1 U17135 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13607) );
  OR2_X1 U17136 ( .A1(n14505), .A2(n13607), .ZN(n13609) );
  NAND2_X1 U17137 ( .A1(n14505), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U17138 ( .A1(n13609), .A2(n13608), .ZN(n16785) );
  NAND2_X1 U17139 ( .A1(n13626), .A2(n16785), .ZN(n13619) );
  NAND2_X1 U17140 ( .A1(n13610), .A2(n13619), .ZN(P2_U2963) );
  AOI22_X1 U17141 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13614) );
  INV_X1 U17142 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13611) );
  OR2_X1 U17143 ( .A1(n14505), .A2(n13611), .ZN(n13613) );
  NAND2_X1 U17144 ( .A1(n14505), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U17145 ( .A1(n13613), .A2(n13612), .ZN(n16798) );
  NAND2_X1 U17146 ( .A1(n13626), .A2(n16798), .ZN(n13615) );
  NAND2_X1 U17147 ( .A1(n13614), .A2(n13615), .ZN(P2_U2976) );
  AOI22_X1 U17148 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U17149 ( .A1(n13616), .A2(n13615), .ZN(P2_U2961) );
  AOI22_X1 U17150 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13618) );
  NAND2_X1 U17151 ( .A1(n13618), .A2(n13617), .ZN(P2_U2960) );
  AOI22_X1 U17152 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U17153 ( .A1(n13620), .A2(n13619), .ZN(P2_U2978) );
  AOI22_X1 U17154 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13622) );
  NAND2_X1 U17155 ( .A1(n13622), .A2(n13621), .ZN(P2_U2959) );
  AOI22_X1 U17156 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13623), .B1(n20350), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U17157 ( .A1(n13625), .A2(n13624), .ZN(P2_U2958) );
  AOI22_X1 U17158 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13627) );
  MUX2_X1 U17159 ( .A(BUF1_REG_5__SCAN_IN), .B(BUF2_REG_5__SCAN_IN), .S(n14505), .Z(n20396) );
  NAND2_X1 U17160 ( .A1(n13626), .A2(n20396), .ZN(n13630) );
  NAND2_X1 U17161 ( .A1(n13627), .A2(n13630), .ZN(P2_U2957) );
  AOI22_X1 U17162 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13629) );
  NAND2_X1 U17163 ( .A1(n13629), .A2(n13628), .ZN(P2_U2956) );
  AOI22_X1 U17164 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13631) );
  NAND2_X1 U17165 ( .A1(n13631), .A2(n13630), .ZN(P2_U2972) );
  INV_X1 U17166 ( .A(n14314), .ZN(n13633) );
  INV_X1 U17167 ( .A(n14258), .ZN(n13632) );
  NAND2_X1 U17168 ( .A1(n13633), .A2(n13632), .ZN(n14223) );
  OR2_X1 U17169 ( .A1(n13635), .A2(n13634), .ZN(n14207) );
  NAND2_X1 U17170 ( .A1(n14223), .A2(n14207), .ZN(n13636) );
  NAND2_X1 U17171 ( .A1(n20400), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13637) );
  NOR2_X1 U17172 ( .A1(n21065), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13638) );
  NAND2_X1 U17173 ( .A1(n21078), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13640) );
  AND4_X1 U17174 ( .A1(n13769), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13640), 
        .A4(n20821), .ZN(n13641) );
  INV_X1 U17175 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13642) );
  MUX2_X1 U17176 ( .A(n13642), .B(n16684), .S(n20291), .Z(n13643) );
  OAI21_X1 U17177 ( .B1(n20283), .B2(n20368), .A(n13643), .ZN(P2_U2887) );
  INV_X1 U17178 ( .A(n15099), .ZN(n13646) );
  INV_X1 U17179 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13644) );
  NAND2_X1 U17180 ( .A1(n15098), .A2(n13644), .ZN(n13645) );
  NAND2_X1 U17181 ( .A1(n13646), .A2(n13645), .ZN(n16652) );
  INV_X1 U17182 ( .A(n16652), .ZN(n13654) );
  OR2_X1 U17183 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  AND2_X1 U17184 ( .A1(n13650), .A2(n13649), .ZN(n14656) );
  NAND2_X1 U17185 ( .A1(n17718), .A2(n14656), .ZN(n13652) );
  NOR2_X1 U17186 ( .A1(n20169), .A2(n20959), .ZN(n14657) );
  INV_X1 U17187 ( .A(n14657), .ZN(n13651) );
  OAI211_X1 U17188 ( .C1(n13644), .C2(n17723), .A(n13652), .B(n13651), .ZN(
        n13653) );
  AOI21_X1 U17189 ( .B1(n17714), .B2(n13654), .A(n13653), .ZN(n13660) );
  INV_X1 U17190 ( .A(n13655), .ZN(n13658) );
  INV_X1 U17191 ( .A(n13656), .ZN(n13657) );
  NAND2_X1 U17192 ( .A1(n13658), .A2(n13657), .ZN(n14659) );
  NAND3_X1 U17193 ( .A1(n14659), .A2(n17719), .A3(n14658), .ZN(n13659) );
  OAI211_X1 U17194 ( .C1(n13661), .C2(n17098), .A(n13660), .B(n13659), .ZN(
        P2_U3012) );
  XNOR2_X1 U17195 ( .A(n13662), .B(n21596), .ZN(n13663) );
  XNOR2_X1 U17196 ( .A(n13664), .B(n13663), .ZN(n17382) );
  AOI22_X1 U17197 ( .A1(n17714), .A2(n15098), .B1(n17719), .B2(n17382), .ZN(
        n13669) );
  OR2_X1 U17198 ( .A1(n13665), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13666) );
  AND2_X1 U17199 ( .A1(n13667), .A2(n13666), .ZN(n17381) );
  NOR2_X1 U17200 ( .A1(n20169), .A2(n20957), .ZN(n17385) );
  AOI21_X1 U17201 ( .B1(n17718), .B2(n17381), .A(n17385), .ZN(n13668) );
  OAI211_X1 U17202 ( .C1(n15098), .C2(n17723), .A(n13669), .B(n13668), .ZN(
        n13670) );
  AOI21_X1 U17203 ( .B1(n13767), .B2(n17716), .A(n13670), .ZN(n13671) );
  INV_X1 U17204 ( .A(n13671), .ZN(P2_U3013) );
  INV_X1 U17205 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13675) );
  NOR2_X1 U17206 ( .A1(n13672), .A2(n17626), .ZN(n17613) );
  INV_X1 U17207 ( .A(n16074), .ZN(n17704) );
  NOR2_X4 U17208 ( .A1(n21206), .A2(n21435), .ZN(n13845) );
  AOI22_X1 U17209 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13674) );
  OAI21_X1 U17210 ( .B1(n13675), .B2(n21191), .A(n13674), .ZN(P1_U2907) );
  INV_X1 U17211 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U17212 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13676) );
  OAI21_X1 U17213 ( .B1(n13677), .B2(n21191), .A(n13676), .ZN(P1_U2908) );
  AOI22_X1 U17214 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13678) );
  OAI21_X1 U17215 ( .B1(n11590), .B2(n21191), .A(n13678), .ZN(P1_U2914) );
  INV_X1 U17216 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U17217 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13679) );
  OAI21_X1 U17218 ( .B1(n13680), .B2(n21191), .A(n13679), .ZN(P1_U2911) );
  AOI22_X1 U17219 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13681) );
  OAI21_X1 U17220 ( .B1(n11561), .B2(n21191), .A(n13681), .ZN(P1_U2912) );
  AOI22_X1 U17221 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13682) );
  OAI21_X1 U17222 ( .B1(n11710), .B2(n21191), .A(n13682), .ZN(P1_U2906) );
  INV_X1 U17223 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U17224 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13683) );
  OAI21_X1 U17225 ( .B1(n13684), .B2(n21191), .A(n13683), .ZN(P1_U2913) );
  INV_X1 U17226 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U17227 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13685) );
  OAI21_X1 U17228 ( .B1(n13686), .B2(n21191), .A(n13685), .ZN(P1_U2909) );
  INV_X1 U17229 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13691) );
  INV_X1 U17230 ( .A(n13687), .ZN(n13688) );
  OAI21_X1 U17231 ( .B1(n14219), .B2(n13688), .A(n15096), .ZN(n13689) );
  NOR2_X4 U17232 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14393), .ZN(n13718) );
  AOI22_X1 U17233 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20344), .B1(n13718), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13690) );
  OAI21_X1 U17234 ( .B1(n13691), .B2(n13720), .A(n13690), .ZN(P2_U2926) );
  INV_X1 U17235 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13693) );
  AOI22_X1 U17236 ( .A1(n13718), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U17237 ( .B1(n13693), .B2(n13720), .A(n13692), .ZN(P2_U2927) );
  AOI22_X1 U17238 ( .A1(n13718), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13694) );
  OAI21_X1 U17239 ( .B1(n13695), .B2(n13720), .A(n13694), .ZN(P2_U2921) );
  INV_X1 U17240 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U17241 ( .A1(n13718), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13696) );
  OAI21_X1 U17242 ( .B1(n13697), .B2(n13720), .A(n13696), .ZN(P2_U2922) );
  INV_X1 U17243 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U17244 ( .A1(n13718), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13698) );
  OAI21_X1 U17245 ( .B1(n13699), .B2(n13720), .A(n13698), .ZN(P2_U2924) );
  AOI22_X1 U17246 ( .A1(n13718), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U17247 ( .B1(n13701), .B2(n13720), .A(n13700), .ZN(P2_U2925) );
  INV_X1 U17248 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U17249 ( .A1(n13718), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13702) );
  OAI21_X1 U17250 ( .B1(n13703), .B2(n13720), .A(n13702), .ZN(P2_U2928) );
  INV_X1 U17251 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U17252 ( .A1(n13718), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13704) );
  OAI21_X1 U17253 ( .B1(n13705), .B2(n13720), .A(n13704), .ZN(P2_U2933) );
  INV_X1 U17254 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13707) );
  AOI22_X1 U17255 ( .A1(n13718), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13706) );
  OAI21_X1 U17256 ( .B1(n13707), .B2(n13720), .A(n13706), .ZN(P2_U2929) );
  AOI22_X1 U17257 ( .A1(n13718), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13708) );
  OAI21_X1 U17258 ( .B1(n13709), .B2(n13720), .A(n13708), .ZN(P2_U2935) );
  INV_X1 U17259 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U17260 ( .A1(n13718), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13710) );
  OAI21_X1 U17261 ( .B1(n13711), .B2(n13720), .A(n13710), .ZN(P2_U2930) );
  INV_X1 U17262 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17263 ( .A1(n13718), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U17264 ( .B1(n13713), .B2(n13720), .A(n13712), .ZN(P2_U2931) );
  INV_X1 U17265 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17266 ( .A1(n13718), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13714) );
  OAI21_X1 U17267 ( .B1(n13715), .B2(n13720), .A(n13714), .ZN(P2_U2932) );
  AOI22_X1 U17268 ( .A1(n13718), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U17269 ( .B1(n13717), .B2(n13720), .A(n13716), .ZN(P2_U2923) );
  INV_X1 U17270 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U17271 ( .A1(n13718), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13719) );
  OAI21_X1 U17272 ( .B1(n13721), .B2(n13720), .A(n13719), .ZN(P2_U2934) );
  OAI21_X1 U17273 ( .B1(n15466), .B2(n14090), .A(n13722), .ZN(n13723) );
  OR2_X1 U17274 ( .A1(n13724), .A2(n13723), .ZN(n13730) );
  OAI21_X1 U17275 ( .B1(n16090), .B2(n14976), .A(n14690), .ZN(n13726) );
  NAND2_X1 U17276 ( .A1(n14976), .A2(n13800), .ZN(n13725) );
  INV_X1 U17277 ( .A(n21434), .ZN(n21340) );
  AOI21_X1 U17278 ( .B1(n13726), .B2(n13725), .A(n21340), .ZN(n13728) );
  MUX2_X1 U17279 ( .A(n13728), .B(n13727), .S(n17587), .Z(n13729) );
  NAND2_X1 U17280 ( .A1(n15012), .A2(n14679), .ZN(n13734) );
  INV_X1 U17281 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21095) );
  NAND2_X1 U17282 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16074), .ZN(n17709) );
  OR2_X1 U17283 ( .A1(n21095), .A2(n17709), .ZN(n13732) );
  NAND2_X1 U17284 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21654), .ZN(n13731) );
  AND2_X1 U17285 ( .A1(n13732), .A2(n13731), .ZN(n13733) );
  INV_X1 U17286 ( .A(n14152), .ZN(n16290) );
  XNOR2_X1 U17287 ( .A(n13735), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15014) );
  INV_X1 U17288 ( .A(n15014), .ZN(n21158) );
  INV_X1 U17289 ( .A(n15013), .ZN(n13736) );
  NAND4_X1 U17290 ( .A1(n21158), .A2(n13736), .A3(n15092), .A4(n16116), .ZN(
        n13737) );
  OAI21_X1 U17291 ( .B1(n15015), .B2(n16116), .A(n13737), .ZN(P1_U3468) );
  INV_X1 U17292 ( .A(n14508), .ZN(n14402) );
  AND3_X1 U17293 ( .A1(n12802), .A2(n13739), .A3(n9734), .ZN(n13740) );
  AOI21_X1 U17294 ( .B1(n14314), .B2(n14213), .A(n13740), .ZN(n14224) );
  NAND2_X1 U17295 ( .A1(n14224), .A2(n13741), .ZN(n13742) );
  NAND2_X1 U17296 ( .A1(n12602), .A2(n20400), .ZN(n13743) );
  OR2_X1 U17297 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  NAND2_X1 U17298 ( .A1(n12616), .A2(n13747), .ZN(n13748) );
  INV_X1 U17299 ( .A(n13748), .ZN(n17394) );
  NOR2_X1 U17300 ( .A1(n20368), .A2(n13748), .ZN(n20310) );
  INV_X1 U17301 ( .A(n20310), .ZN(n13750) );
  NAND2_X1 U17302 ( .A1(n14282), .A2(n13749), .ZN(n20311) );
  OAI211_X1 U17303 ( .C1(n20421), .C2(n17394), .A(n13750), .B(n20295), .ZN(
        n13753) );
  AOI22_X1 U17304 ( .A1(n20307), .A2(n17394), .B1(n20306), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13752) );
  OAI211_X1 U17305 ( .C1(n14402), .C2(n20315), .A(n13753), .B(n13752), .ZN(
        P2_U2919) );
  NAND2_X1 U17306 ( .A1(n13756), .A2(n13757), .ZN(n13758) );
  NAND2_X1 U17307 ( .A1(n13755), .A2(n13758), .ZN(n20234) );
  INV_X1 U17308 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20331) );
  INV_X1 U17309 ( .A(n16805), .ZN(n13759) );
  OAI222_X1 U17310 ( .A1(n20234), .A2(n14582), .B1(n14282), .B2(n20331), .C1(
        n20315), .C2(n13759), .ZN(P2_U2911) );
  NAND2_X1 U17311 ( .A1(n13489), .A2(n13760), .ZN(n13762) );
  NAND2_X1 U17312 ( .A1(n13762), .A2(n13761), .ZN(n13764) );
  OR2_X1 U17313 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  NAND2_X1 U17314 ( .A1(n13756), .A2(n13765), .ZN(n20250) );
  INV_X1 U17315 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20333) );
  INV_X1 U17316 ( .A(n16812), .ZN(n20410) );
  OAI222_X1 U17317 ( .A1(n20250), .A2(n14582), .B1(n20333), .B2(n14282), .C1(
        n20315), .C2(n20410), .ZN(P2_U2912) );
  INV_X1 U17318 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20335) );
  OAI222_X1 U17319 ( .A1(n16625), .A2(n14582), .B1(n20335), .B2(n14282), .C1(
        n20315), .C2(n20402), .ZN(P2_U2913) );
  INV_X1 U17320 ( .A(n13833), .ZN(n13766) );
  NAND2_X1 U17321 ( .A1(n20820), .A2(n20672), .ZN(n20818) );
  AOI21_X1 U17322 ( .B1(n13941), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20706), .ZN(n13768) );
  MUX2_X1 U17323 ( .A(n13774), .B(n16674), .S(n20291), .Z(n13775) );
  OAI21_X1 U17324 ( .B1(n20369), .B2(n20283), .A(n13775), .ZN(P2_U2886) );
  INV_X1 U17325 ( .A(n13806), .ZN(n13776) );
  AOI21_X1 U17326 ( .B1(n13777), .B2(n13755), .A(n13776), .ZN(n17331) );
  INV_X1 U17327 ( .A(n17331), .ZN(n13779) );
  INV_X1 U17328 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20329) );
  INV_X1 U17329 ( .A(n16798), .ZN(n13778) );
  OAI222_X1 U17330 ( .A1(n13779), .A2(n14582), .B1(n14282), .B2(n20329), .C1(
        n20315), .C2(n13778), .ZN(P2_U2910) );
  INV_X1 U17331 ( .A(n13780), .ZN(n13781) );
  OAI21_X1 U17332 ( .B1(n13781), .B2(n10104), .A(n13796), .ZN(n15495) );
  OR2_X1 U17333 ( .A1(n9720), .A2(n13783), .ZN(n13786) );
  NAND4_X1 U17334 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n15090), .ZN(
        n13787) );
  AND2_X1 U17335 ( .A1(n13788), .A2(n13787), .ZN(n21252) );
  INV_X1 U17336 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13791) );
  OAI21_X1 U17337 ( .B1(n15857), .B2(n13789), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13790) );
  OAI21_X1 U17338 ( .B1(n13791), .B2(n17669), .A(n13790), .ZN(n13792) );
  AOI21_X1 U17339 ( .B1(n17668), .B2(n21252), .A(n13792), .ZN(n13793) );
  OAI21_X1 U17340 ( .B1(n15495), .B2(n17666), .A(n13793), .ZN(P1_U2999) );
  INV_X1 U17341 ( .A(n13794), .ZN(n13797) );
  NAND3_X1 U17342 ( .A1(n13797), .A2(n13796), .A3(n13795), .ZN(n13798) );
  NAND2_X1 U17343 ( .A1(n13798), .A2(n13972), .ZN(n15488) );
  XNOR2_X1 U17344 ( .A(n13799), .B(n13800), .ZN(n13910) );
  AOI22_X1 U17345 ( .A1(n15554), .A2(n13910), .B1(n15553), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13801) );
  OAI21_X1 U17346 ( .B1(n15488), .B2(n15556), .A(n13801), .ZN(P1_U2871) );
  INV_X1 U17347 ( .A(n13802), .ZN(n13803) );
  AOI21_X1 U17348 ( .B1(n13804), .B2(n15090), .A(n13803), .ZN(n21249) );
  INV_X1 U17349 ( .A(n21249), .ZN(n13805) );
  INV_X1 U17350 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n15490) );
  OAI222_X1 U17351 ( .A1(n13805), .A2(n15545), .B1(n15544), .B2(n15490), .C1(
        n15495), .C2(n15530), .ZN(P1_U2872) );
  AOI21_X1 U17352 ( .B1(n13807), .B2(n13806), .A(n9815), .ZN(n20221) );
  INV_X1 U17353 ( .A(n20221), .ZN(n13809) );
  AOI22_X1 U17354 ( .A1(n14579), .A2(n16791), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n20306), .ZN(n13808) );
  OAI21_X1 U17355 ( .B1(n13809), .B2(n14582), .A(n13808), .ZN(P2_U2909) );
  XNOR2_X1 U17356 ( .A(n13810), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19194) );
  INV_X1 U17357 ( .A(n19443), .ZN(n19471) );
  OAI22_X1 U17358 ( .A1(n14106), .A2(n13886), .B1(n13888), .B2(n19451), .ZN(
        n13893) );
  INV_X1 U17359 ( .A(n13893), .ZN(n19438) );
  NOR4_X1 U17360 ( .A1(n19438), .A2(n19449), .A3(n11856), .A4(n19459), .ZN(
        n13814) );
  NOR2_X1 U17361 ( .A1(n19390), .A2(n19469), .ZN(n19454) );
  OAI21_X1 U17362 ( .B1(n13886), .B2(n13819), .A(n19949), .ZN(n13811) );
  NOR2_X1 U17363 ( .A1(n19406), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19298) );
  INV_X1 U17364 ( .A(n19298), .ZN(n19452) );
  OAI211_X1 U17365 ( .C1(n13812), .C2(n19454), .A(n13811), .B(n19452), .ZN(
        n13813) );
  INV_X1 U17366 ( .A(n13813), .ZN(n19419) );
  OAI21_X1 U17367 ( .B1(n19419), .B2(n19459), .A(n19466), .ZN(n13824) );
  INV_X1 U17368 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n21460) );
  NOR2_X1 U17369 ( .A1(n19428), .A2(n21460), .ZN(n19197) );
  AOI221_X1 U17370 ( .B1(n13814), .B2(n10333), .C1(n13824), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n19197), .ZN(n13818) );
  AOI21_X1 U17371 ( .B1(n9850), .B2(n13816), .A(n13815), .ZN(n19198) );
  NAND2_X1 U17372 ( .A1(n19476), .A2(n19198), .ZN(n13817) );
  OAI211_X1 U17373 ( .C1(n19194), .C2(n19471), .A(n13818), .B(n13817), .ZN(
        P3_U2857) );
  NOR3_X1 U17374 ( .A1(n19438), .A2(n13819), .A3(n19459), .ZN(n19427) );
  INV_X1 U17375 ( .A(n19427), .ZN(n13828) );
  AOI21_X1 U17376 ( .B1(n13821), .B2(n19420), .A(n13820), .ZN(n17455) );
  XNOR2_X1 U17377 ( .A(n13823), .B(n13822), .ZN(n17451) );
  NAND2_X1 U17378 ( .A1(n13824), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13825) );
  NAND2_X1 U17379 ( .A1(n19477), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n17450) );
  OAI211_X1 U17380 ( .C1(n17451), .C2(n19471), .A(n13825), .B(n17450), .ZN(
        n13826) );
  AOI21_X1 U17381 ( .B1(n19476), .B2(n17455), .A(n13826), .ZN(n13827) );
  OAI21_X1 U17382 ( .B1(n13828), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13827), .ZN(P3_U2856) );
  INV_X1 U17383 ( .A(n13829), .ZN(n13830) );
  XNOR2_X1 U17384 ( .A(n20475), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14592) );
  AOI22_X1 U17385 ( .A1(n13941), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21028), .B2(n14592), .ZN(n13835) );
  NAND2_X1 U17386 ( .A1(n13836), .A2(n13835), .ZN(n13839) );
  OAI21_X1 U17387 ( .B1(n13839), .B2(n13838), .A(n13947), .ZN(n13840) );
  MUX2_X1 U17388 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n16661), .S(n20291), .Z(
        n13843) );
  INV_X1 U17389 ( .A(n13843), .ZN(n13844) );
  OAI21_X1 U17390 ( .B1(n21036), .B2(n20283), .A(n13844), .ZN(P2_U2885) );
  INV_X1 U17391 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17392 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13846) );
  OAI21_X1 U17393 ( .B1(n13847), .B2(n21191), .A(n13846), .ZN(P1_U2920) );
  AOI22_X1 U17394 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13848) );
  OAI21_X1 U17395 ( .B1(n15610), .B2(n21191), .A(n13848), .ZN(P1_U2919) );
  INV_X1 U17396 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21648) );
  AOI22_X1 U17397 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13849) );
  OAI21_X1 U17398 ( .B1(n21648), .B2(n21191), .A(n13849), .ZN(P1_U2910) );
  AOI22_X1 U17399 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13850) );
  OAI21_X1 U17400 ( .B1(n11499), .B2(n21191), .A(n13850), .ZN(P1_U2915) );
  AOI22_X1 U17401 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13851) );
  OAI21_X1 U17402 ( .B1(n11461), .B2(n21191), .A(n13851), .ZN(P1_U2917) );
  XNOR2_X1 U17403 ( .A(n13852), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13912) );
  INV_X1 U17404 ( .A(n15488), .ZN(n13855) );
  AOI22_X1 U17405 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15856), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13853) );
  OAI21_X1 U17406 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17665), .A(
        n13853), .ZN(n13854) );
  AOI21_X1 U17407 ( .B1(n13855), .B2(n17654), .A(n13854), .ZN(n13856) );
  OAI21_X1 U17408 ( .B1(n13912), .B2(n21094), .A(n13856), .ZN(P1_U2998) );
  OAI21_X1 U17409 ( .B1(n9815), .B2(n13859), .A(n13858), .ZN(n17308) );
  INV_X1 U17410 ( .A(n16785), .ZN(n13860) );
  INV_X1 U17411 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20325) );
  OAI222_X1 U17412 ( .A1(n17308), .A2(n14582), .B1(n13860), .B2(n20315), .C1(
        n20325), .C2(n14282), .ZN(P2_U2908) );
  XNOR2_X1 U17413 ( .A(n13862), .B(n13957), .ZN(n17474) );
  XNOR2_X1 U17414 ( .A(n13862), .B(n13861), .ZN(n17470) );
  INV_X1 U17415 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n13863) );
  NOR2_X1 U17416 ( .A1(n19216), .A2(n13863), .ZN(n17469) );
  INV_X1 U17417 ( .A(n19440), .ZN(n19323) );
  NOR2_X1 U17418 ( .A1(n19323), .A2(n19459), .ZN(n19421) );
  INV_X1 U17419 ( .A(n19421), .ZN(n17477) );
  AOI211_X1 U17420 ( .C1(n19253), .C2(n19472), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17477), .ZN(n13864) );
  AOI211_X1 U17421 ( .C1(n19443), .C2(n17470), .A(n17469), .B(n13864), .ZN(
        n13867) );
  OR3_X1 U17422 ( .A1(n19459), .A2(n19346), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19478) );
  AOI21_X1 U17423 ( .B1(n19478), .B2(n19466), .A(n11932), .ZN(n13865) );
  INV_X1 U17424 ( .A(n13865), .ZN(n13866) );
  OAI211_X1 U17425 ( .C1(n17474), .C2(n19430), .A(n13867), .B(n13866), .ZN(
        P3_U2861) );
  XNOR2_X1 U17426 ( .A(n13869), .B(n13868), .ZN(n13981) );
  NAND2_X1 U17427 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13873) );
  INV_X1 U17428 ( .A(n13983), .ZN(n13870) );
  NAND2_X1 U17429 ( .A1(n15965), .A2(n13870), .ZN(n13872) );
  OAI21_X1 U17430 ( .B1(n15969), .B2(n13873), .A(n16055), .ZN(n13882) );
  NOR2_X1 U17431 ( .A1(n13875), .A2(n13876), .ZN(n13877) );
  OR2_X1 U17432 ( .A1(n13874), .A2(n13877), .ZN(n15467) );
  NAND3_X1 U17433 ( .A1(n16031), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13041), .ZN(n13880) );
  NOR2_X1 U17434 ( .A1(n15969), .A2(n16025), .ZN(n13878) );
  AOI21_X1 U17435 ( .B1(n15856), .B2(P1_REIP_REG_2__SCAN_IN), .A(n13878), .ZN(
        n13879) );
  OAI211_X1 U17436 ( .C1(n16051), .C2(n15467), .A(n13880), .B(n13879), .ZN(
        n13881) );
  AOI21_X1 U17437 ( .B1(n13882), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13881), .ZN(n13883) );
  OAI21_X1 U17438 ( .B1(n16064), .B2(n13981), .A(n13883), .ZN(P1_U3029) );
  XNOR2_X1 U17439 ( .A(n13885), .B(n13884), .ZN(n19203) );
  INV_X1 U17440 ( .A(n19454), .ZN(n13887) );
  AND2_X1 U17441 ( .A1(n19949), .A2(n13886), .ZN(n19455) );
  AOI211_X1 U17442 ( .C1(n13888), .C2(n13887), .A(n19455), .B(n19298), .ZN(
        n13889) );
  AOI21_X1 U17443 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13889), .A(
        n19459), .ZN(n19441) );
  XNOR2_X1 U17444 ( .A(n13891), .B(n13890), .ZN(n19209) );
  OAI22_X1 U17445 ( .A1(n11856), .A2(n19466), .B1(n19430), .B2(n19209), .ZN(
        n13892) );
  AOI221_X1 U17446 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19441), .C1(
        n13893), .C2(n19441), .A(n13892), .ZN(n13894) );
  NAND2_X1 U17447 ( .A1(n19477), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19207) );
  OAI211_X1 U17448 ( .C1(n19203), .C2(n19471), .A(n13894), .B(n19207), .ZN(
        P3_U2859) );
  NAND2_X1 U17449 ( .A1(n13858), .A2(n13896), .ZN(n13897) );
  NAND2_X1 U17450 ( .A1(n13895), .A2(n13897), .ZN(n20205) );
  AOI22_X1 U17451 ( .A1(n14579), .A2(n16777), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n20306), .ZN(n13898) );
  OAI21_X1 U17452 ( .B1(n20205), .B2(n14582), .A(n13898), .ZN(P2_U2907) );
  NAND2_X1 U17453 ( .A1(n10829), .A2(n14057), .ZN(n13899) );
  INV_X1 U17454 ( .A(DATAI_1_), .ZN(n13901) );
  NAND2_X1 U17455 ( .A1(n15585), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13900) );
  OAI21_X1 U17456 ( .B1(n15585), .B2(n13901), .A(n13900), .ZN(n15613) );
  INV_X1 U17457 ( .A(n15613), .ZN(n14040) );
  INV_X1 U17458 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21217) );
  OAI222_X1 U17459 ( .A1(n15488), .A2(n15643), .B1(n15646), .B2(n14040), .C1(
        n15644), .C2(n21217), .ZN(P1_U2903) );
  NAND2_X1 U17460 ( .A1(n14022), .A2(DATAI_0_), .ZN(n13903) );
  NAND2_X1 U17461 ( .A1(n15585), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13902) );
  INV_X1 U17462 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21219) );
  OAI222_X1 U17463 ( .A1(n15495), .A2(n15643), .B1(n15646), .B2(n14292), .C1(
        n15644), .C2(n21219), .ZN(P1_U2904) );
  INV_X1 U17464 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21358) );
  INV_X1 U17465 ( .A(n21253), .ZN(n13905) );
  OAI21_X1 U17466 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13905), .A(
        n13904), .ZN(n21254) );
  AOI21_X1 U17467 ( .B1(n15090), .B2(n13906), .A(n16030), .ZN(n13907) );
  AOI22_X1 U17468 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21254), .B1(
        n13907), .B2(n16099), .ZN(n13908) );
  OAI21_X1 U17469 ( .B1(n17669), .B2(n21358), .A(n13908), .ZN(n13909) );
  AOI21_X1 U17470 ( .B1(n21250), .B2(n13910), .A(n13909), .ZN(n13911) );
  OAI21_X1 U17471 ( .B1(n13912), .B2(n16064), .A(n13911), .ZN(P1_U3030) );
  NOR2_X1 U17472 ( .A1(n18217), .A2(n18171), .ZN(n13916) );
  INV_X1 U17473 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18650) );
  AND2_X1 U17474 ( .A1(n20105), .A2(n19493), .ZN(n20107) );
  INV_X1 U17475 ( .A(n20107), .ZN(n18214) );
  NAND3_X1 U17476 ( .A1(n18212), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14134), .ZN(n13913) );
  OAI21_X1 U17477 ( .B1(n18214), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13913), .ZN(n13914) );
  AOI21_X1 U17478 ( .B1(n18156), .B2(P3_REIP_REG_0__SCAN_IN), .A(n13914), .ZN(
        n13915) );
  OAI21_X1 U17479 ( .B1(n13916), .B2(n18650), .A(n13915), .ZN(P3_U2671) );
  INV_X1 U17480 ( .A(n13917), .ZN(n18182) );
  AND2_X1 U17481 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13923) );
  INV_X1 U17482 ( .A(n13918), .ZN(n13921) );
  OAI21_X1 U17483 ( .B1(n13921), .B2(n13920), .A(n13919), .ZN(n14100) );
  INV_X1 U17484 ( .A(n14100), .ZN(n13922) );
  OAI21_X1 U17485 ( .B1(n19253), .B2(n13923), .A(n13922), .ZN(n13926) );
  INV_X1 U17486 ( .A(n14113), .ZN(n14099) );
  NAND2_X1 U17487 ( .A1(n14099), .A2(n13924), .ZN(n14098) );
  INV_X1 U17488 ( .A(n14098), .ZN(n13925) );
  AOI21_X1 U17489 ( .B1(n13926), .B2(n18182), .A(n13925), .ZN(n19927) );
  NOR2_X1 U17490 ( .A1(n19927), .A2(n14134), .ZN(n13933) );
  NOR2_X1 U17491 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n20070), .ZN(n19492) );
  INV_X1 U17492 ( .A(n18856), .ZN(n18858) );
  NOR2_X1 U17493 ( .A1(n20089), .A2(n18858), .ZN(n19967) );
  NAND2_X1 U17494 ( .A1(n19953), .A2(n20083), .ZN(n13931) );
  NOR2_X1 U17495 ( .A1(n13994), .A2(n13995), .ZN(n13928) );
  NOR2_X1 U17496 ( .A1(n13928), .A2(n13997), .ZN(n13929) );
  OAI211_X1 U17497 ( .C1(n18796), .C2(n13931), .A(n13930), .B(n13929), .ZN(
        n19960) );
  INV_X1 U17498 ( .A(n19960), .ZN(n19936) );
  INV_X1 U17499 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19482) );
  NAND3_X1 U17500 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n20068)
         );
  OAI22_X1 U17501 ( .A1(n19936), .A2(n19976), .B1(n19482), .B2(n20068), .ZN(
        n13932) );
  AOI211_X1 U17502 ( .C1(n19965), .C2(n18182), .A(n13933), .B(n14139), .ZN(
        n13939) );
  NAND2_X1 U17503 ( .A1(n19390), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13934) );
  NAND2_X1 U17504 ( .A1(n13934), .A2(n19253), .ZN(n14112) );
  NAND3_X1 U17505 ( .A1(n14112), .A2(n13935), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13937) );
  NAND3_X1 U17506 ( .A1(n19949), .A2(n19926), .A3(n14098), .ZN(n13936) );
  NAND2_X1 U17507 ( .A1(n13937), .A2(n13936), .ZN(n19928) );
  AOI22_X1 U17508 ( .A1(n19928), .A2(n20103), .B1(n9723), .B2(n19965), .ZN(
        n13938) );
  OAI22_X1 U17509 ( .A1(n13939), .A2(n19926), .B1(n14139), .B2(n13938), .ZN(
        P3_U3285) );
  NAND2_X1 U17510 ( .A1(n13952), .A2(n13766), .ZN(n13943) );
  OAI21_X1 U17511 ( .B1(n20475), .B2(n21692), .A(n21494), .ZN(n13940) );
  INV_X1 U17512 ( .A(n20475), .ZN(n20737) );
  NAND2_X1 U17513 ( .A1(n20737), .A2(n20863), .ZN(n20871) );
  AOI21_X1 U17514 ( .B1(n13941), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14600), .ZN(n13942) );
  NAND2_X1 U17515 ( .A1(n13943), .A2(n13942), .ZN(n14013) );
  NAND2_X1 U17516 ( .A1(n14013), .A2(n13945), .ZN(n14574) );
  NAND2_X1 U17517 ( .A1(n13948), .A2(n13947), .ZN(n13950) );
  MUX2_X1 U17518 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n13953), .S(n20291), .Z(
        n13954) );
  AOI21_X1 U17519 ( .B1(n21030), .B2(n20288), .A(n13954), .ZN(n13955) );
  INV_X1 U17520 ( .A(n13955), .ZN(P2_U2884) );
  NOR2_X1 U17521 ( .A1(n13957), .A2(n13956), .ZN(n19467) );
  INV_X1 U17522 ( .A(n19217), .ZN(n17471) );
  AOI22_X1 U17523 ( .A1(n17471), .A2(n19467), .B1(n19477), .B2(
        P3_REIP_REG_0__SCAN_IN), .ZN(n13960) );
  NAND3_X1 U17524 ( .A1(n19481), .A2(n19103), .A3(n19202), .ZN(n13958) );
  NAND2_X1 U17525 ( .A1(n13958), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13959) );
  OAI211_X1 U17526 ( .C1(n19467), .C2(n19210), .A(n13960), .B(n13959), .ZN(
        P3_U2830) );
  OAI21_X1 U17527 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n14140) );
  OR2_X1 U17528 ( .A1(n13874), .A2(n13965), .ZN(n13966) );
  AND2_X1 U17529 ( .A1(n13964), .A2(n13966), .ZN(n21175) );
  AOI22_X1 U17530 ( .A1(n15554), .A2(n21175), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15553), .ZN(n13967) );
  OAI21_X1 U17531 ( .B1(n14140), .B2(n15530), .A(n13967), .ZN(P1_U2869) );
  INV_X1 U17532 ( .A(DATAI_3_), .ZN(n13969) );
  NAND2_X1 U17533 ( .A1(n15585), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13968) );
  OAI21_X1 U17534 ( .B1(n15585), .B2(n13969), .A(n13968), .ZN(n15603) );
  INV_X1 U17535 ( .A(n15603), .ZN(n14044) );
  OAI222_X1 U17536 ( .A1(n14140), .A2(n15643), .B1(n15646), .B2(n14044), .C1(
        n15644), .C2(n11200), .ZN(P1_U2901) );
  INV_X1 U17537 ( .A(n13970), .ZN(n13971) );
  AOI21_X1 U17538 ( .B1(n13973), .B2(n13972), .A(n13971), .ZN(n15478) );
  INV_X1 U17539 ( .A(n15478), .ZN(n13991) );
  INV_X1 U17540 ( .A(n15467), .ZN(n13974) );
  AOI22_X1 U17541 ( .A1(n15554), .A2(n13974), .B1(n15553), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13975) );
  OAI21_X1 U17542 ( .B1(n13991), .B2(n15530), .A(n13975), .ZN(P1_U2870) );
  INV_X1 U17543 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20320) );
  INV_X1 U17544 ( .A(n16769), .ZN(n13977) );
  XNOR2_X1 U17545 ( .A(n13895), .B(n9846), .ZN(n17284) );
  INV_X1 U17546 ( .A(n17284), .ZN(n13976) );
  OAI222_X1 U17547 ( .A1(n14282), .A2(n20320), .B1(n13977), .B2(n20315), .C1(
        n13976), .C2(n14582), .ZN(P2_U2906) );
  AOI22_X1 U17548 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n15856), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13978) );
  OAI21_X1 U17549 ( .B1(n15481), .B2(n17665), .A(n13978), .ZN(n13979) );
  AOI21_X1 U17550 ( .B1(n15478), .B2(n17654), .A(n13979), .ZN(n13980) );
  OAI21_X1 U17551 ( .B1(n21094), .B2(n13981), .A(n13980), .ZN(P1_U2997) );
  XNOR2_X1 U17552 ( .A(n14372), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14375) );
  XNOR2_X1 U17553 ( .A(n14375), .B(n14374), .ZN(n14145) );
  INV_X1 U17554 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13982) );
  OR2_X1 U17555 ( .A1(n17669), .A2(n13982), .ZN(n14141) );
  OAI21_X1 U17556 ( .B1(n15969), .B2(n16025), .A(n16055), .ZN(n14378) );
  NAND2_X1 U17557 ( .A1(n13983), .A2(n16031), .ZN(n14428) );
  NAND2_X1 U17558 ( .A1(n15969), .A2(n14428), .ZN(n13984) );
  INV_X1 U17559 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U17560 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14378), .B1(
        n17692), .B2(n13985), .ZN(n13986) );
  NAND2_X1 U17561 ( .A1(n14141), .A2(n13986), .ZN(n13987) );
  AOI21_X1 U17562 ( .B1(n21250), .B2(n21175), .A(n13987), .ZN(n13988) );
  OAI21_X1 U17563 ( .B1(n14145), .B2(n16064), .A(n13988), .ZN(P1_U3028) );
  INV_X1 U17564 ( .A(DATAI_2_), .ZN(n13990) );
  NAND2_X1 U17565 ( .A1(n15585), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13989) );
  OAI21_X1 U17566 ( .B1(n15585), .B2(n13990), .A(n13989), .ZN(n15606) );
  INV_X1 U17567 ( .A(n15606), .ZN(n14092) );
  OAI222_X1 U17568 ( .A1(n13991), .A2(n15643), .B1(n15646), .B2(n14092), .C1(
        n15644), .C2(n11173), .ZN(P1_U2902) );
  NAND2_X1 U17569 ( .A1(n19521), .A2(n19508), .ZN(n13992) );
  OAI22_X2 U17570 ( .A1(n13995), .A2(n13994), .B1(n13993), .B2(n13992), .ZN(
        n17535) );
  INV_X1 U17571 ( .A(n18739), .ZN(n14006) );
  OAI221_X1 U17572 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(P3_EAX_REG_0__SCAN_IN), 
        .C1(P3_EAX_REG_1__SCAN_IN), .C2(n14006), .A(n18784), .ZN(n14000) );
  NAND2_X1 U17573 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18652) );
  NOR2_X1 U17574 ( .A1(n18655), .A2(n18652), .ZN(n18790) );
  NAND2_X1 U17575 ( .A1(n14115), .A2(n18777), .ZN(n18795) );
  AOI22_X1 U17576 ( .A1(n13998), .A2(n18786), .B1(BUF2_REG_1__SCAN_IN), .B2(
        n18787), .ZN(n13999) );
  OAI21_X1 U17577 ( .B1(n14000), .B2(n18790), .A(n13999), .ZN(P3_U2734) );
  NOR2_X1 U17578 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  OR2_X1 U17579 ( .A1(n14001), .A2(n14004), .ZN(n20190) );
  AOI22_X1 U17580 ( .A1(n14579), .A2(n14965), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n20306), .ZN(n14005) );
  OAI21_X1 U17581 ( .B1(n20190), .B2(n14582), .A(n14005), .ZN(P2_U2905) );
  INV_X1 U17582 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18854) );
  INV_X1 U17583 ( .A(n18655), .ZN(n14010) );
  NAND2_X1 U17584 ( .A1(n14006), .A2(n18854), .ZN(n14009) );
  AOI22_X1 U17585 ( .A1(n14007), .A2(n18786), .B1(BUF2_REG_0__SCAN_IN), .B2(
        n18787), .ZN(n14008) );
  OAI211_X1 U17586 ( .C1(n18854), .C2(n14010), .A(n14009), .B(n14008), .ZN(
        P3_U2735) );
  NAND2_X1 U17587 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20400), .ZN(
        n14011) );
  XOR2_X1 U17588 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14578), .Z(n14020)
         );
  NAND2_X1 U17589 ( .A1(n14014), .A2(n14015), .ZN(n14016) );
  AND2_X1 U17590 ( .A1(n13486), .A2(n14016), .ZN(n17715) );
  INV_X1 U17591 ( .A(n17715), .ZN(n14018) );
  MUX2_X1 U17592 ( .A(n14018), .B(n14017), .S(n16764), .Z(n14019) );
  OAI21_X1 U17593 ( .B1(n14020), .B2(n20283), .A(n14019), .ZN(P2_U2882) );
  AND2_X1 U17594 ( .A1(n11176), .A2(n16079), .ZN(n14025) );
  AOI22_X1 U17595 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9716), .B1(DATAI_30_), 
        .B2(n9715), .ZN(n21323) );
  INV_X1 U17596 ( .A(n21323), .ZN(n16329) );
  INV_X1 U17597 ( .A(DATAI_6_), .ZN(n14027) );
  NAND2_X1 U17598 ( .A1(n15585), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14026) );
  OAI21_X1 U17599 ( .B1(n15585), .B2(n14027), .A(n14026), .ZN(n15592) );
  INV_X1 U17600 ( .A(n15592), .ZN(n14534) );
  INV_X1 U17601 ( .A(n15053), .ZN(n14030) );
  NOR2_X1 U17602 ( .A1(n15489), .A2(n14029), .ZN(n16382) );
  INV_X1 U17603 ( .A(n16382), .ZN(n14153) );
  OR2_X1 U17604 ( .A1(n14535), .A2(n17600), .ZN(n21747) );
  OAI21_X1 U17605 ( .B1(n14030), .B2(n14153), .A(n21747), .ZN(n14031) );
  NAND3_X1 U17606 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n15029), .ZN(n14438) );
  INV_X1 U17607 ( .A(n14438), .ZN(n14036) );
  AOI22_X1 U17608 ( .A1(n14031), .A2(n21274), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14036), .ZN(n21749) );
  NAND2_X1 U17609 ( .A1(n14091), .A2(n10879), .ZN(n16327) );
  OAI22_X1 U17610 ( .A1(n16422), .A2(n21749), .B1(n16327), .B2(n21747), .ZN(
        n14033) );
  AOI21_X1 U17611 ( .B1(n21753), .B2(n16329), .A(n14033), .ZN(n14039) );
  INV_X1 U17612 ( .A(n14034), .ZN(n14035) );
  INV_X1 U17613 ( .A(n14159), .ZN(n16081) );
  NOR2_X1 U17614 ( .A1(n14035), .A2(n16081), .ZN(n14037) );
  AOI21_X1 U17615 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21271), .A(n16202), 
        .ZN(n21281) );
  NAND2_X1 U17616 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14038) );
  OAI211_X1 U17617 ( .C1(n16418), .C2(n21757), .A(n14039), .B(n14038), .ZN(
        P1_U3127) );
  AOI22_X1 U17618 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9716), .B1(DATAI_25_), 
        .B2(n9715), .ZN(n21293) );
  INV_X1 U17619 ( .A(n21293), .ZN(n16306) );
  NAND2_X1 U17620 ( .A1(n14091), .A2(n14691), .ZN(n16304) );
  OAI22_X1 U17621 ( .A1(n16399), .A2(n21749), .B1(n16304), .B2(n21747), .ZN(
        n14041) );
  AOI21_X1 U17622 ( .B1(n21753), .B2(n16306), .A(n14041), .ZN(n14043) );
  NAND2_X1 U17623 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14042) );
  OAI211_X1 U17624 ( .C1(n16395), .C2(n21757), .A(n14043), .B(n14042), .ZN(
        P1_U3122) );
  AOI22_X1 U17625 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9716), .B1(DATAI_27_), 
        .B2(n9715), .ZN(n21305) );
  INV_X1 U17626 ( .A(n21305), .ZN(n16314) );
  NAND2_X1 U17627 ( .A1(n14091), .A2(n14045), .ZN(n16312) );
  OAI22_X1 U17628 ( .A1(n16407), .A2(n21749), .B1(n16312), .B2(n21747), .ZN(
        n14046) );
  AOI21_X1 U17629 ( .B1(n21753), .B2(n16314), .A(n14046), .ZN(n14048) );
  NAND2_X1 U17630 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14047) );
  OAI211_X1 U17631 ( .C1(n16403), .C2(n21757), .A(n14048), .B(n14047), .ZN(
        P1_U3124) );
  AOI22_X1 U17632 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9716), .B1(DATAI_28_), 
        .B2(n9715), .ZN(n21311) );
  INV_X1 U17633 ( .A(n21311), .ZN(n16319) );
  INV_X1 U17634 ( .A(DATAI_4_), .ZN(n14050) );
  NAND2_X1 U17635 ( .A1(n15585), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14049) );
  OAI21_X1 U17636 ( .B1(n15585), .B2(n14050), .A(n14049), .ZN(n15599) );
  INV_X1 U17637 ( .A(n15599), .ZN(n14371) );
  NAND2_X1 U17638 ( .A1(n14091), .A2(n14051), .ZN(n16317) );
  OAI22_X1 U17639 ( .A1(n16412), .A2(n21749), .B1(n16317), .B2(n21747), .ZN(
        n14052) );
  AOI21_X1 U17640 ( .B1(n21753), .B2(n16319), .A(n14052), .ZN(n14054) );
  NAND2_X1 U17641 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14053) );
  OAI211_X1 U17642 ( .C1(n16408), .C2(n21757), .A(n14054), .B(n14053), .ZN(
        P1_U3125) );
  AOI22_X1 U17643 ( .A1(DATAI_31_), .A2(n9715), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9716), .ZN(n21334) );
  INV_X1 U17644 ( .A(n21334), .ZN(n16335) );
  INV_X1 U17645 ( .A(DATAI_7_), .ZN(n14056) );
  NAND2_X1 U17646 ( .A1(n15585), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14055) );
  OAI21_X1 U17647 ( .B1(n15585), .B2(n14056), .A(n14055), .ZN(n15589) );
  INV_X1 U17648 ( .A(n15589), .ZN(n15645) );
  NAND2_X1 U17649 ( .A1(n14091), .A2(n14057), .ZN(n16333) );
  OAI22_X1 U17650 ( .A1(n16431), .A2(n21749), .B1(n16333), .B2(n21747), .ZN(
        n14058) );
  AOI21_X1 U17651 ( .B1(n21753), .B2(n16335), .A(n14058), .ZN(n14060) );
  NAND2_X1 U17652 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n14059) );
  OAI211_X1 U17653 ( .C1(n16426), .C2(n21757), .A(n14060), .B(n14059), .ZN(
        P1_U3128) );
  AOI22_X2 U17654 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n9716), .B1(DATAI_16_), 
        .B2(n9715), .ZN(n16390) );
  AOI22_X1 U17655 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9716), .B1(DATAI_24_), 
        .B2(n9715), .ZN(n21287) );
  INV_X1 U17656 ( .A(n21287), .ZN(n16297) );
  NAND2_X1 U17657 ( .A1(n14091), .A2(n14697), .ZN(n16295) );
  OAI22_X1 U17658 ( .A1(n16394), .A2(n21749), .B1(n16295), .B2(n21747), .ZN(
        n14061) );
  AOI21_X1 U17659 ( .B1(n21753), .B2(n16297), .A(n14061), .ZN(n14063) );
  NAND2_X1 U17660 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14062) );
  OAI211_X1 U17661 ( .C1(n16390), .C2(n21757), .A(n14063), .B(n14062), .ZN(
        P1_U3121) );
  AOI22_X1 U17662 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9716), .B1(DATAI_29_), 
        .B2(n9715), .ZN(n21317) );
  INV_X1 U17663 ( .A(n21317), .ZN(n16324) );
  INV_X1 U17664 ( .A(DATAI_5_), .ZN(n14065) );
  NAND2_X1 U17665 ( .A1(n15585), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14064) );
  OAI21_X1 U17666 ( .B1(n15585), .B2(n14065), .A(n14064), .ZN(n15595) );
  INV_X1 U17667 ( .A(n15595), .ZN(n14350) );
  NAND2_X1 U17668 ( .A1(n14091), .A2(n15557), .ZN(n16322) );
  OAI22_X1 U17669 ( .A1(n16417), .A2(n21749), .B1(n16322), .B2(n21747), .ZN(
        n14066) );
  AOI21_X1 U17670 ( .B1(n21753), .B2(n16324), .A(n14066), .ZN(n14068) );
  NAND2_X1 U17671 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14067) );
  OAI211_X1 U17672 ( .C1(n16413), .C2(n21757), .A(n14068), .B(n14067), .ZN(
        P1_U3126) );
  INV_X1 U17673 ( .A(n11176), .ZN(n14069) );
  NAND3_X1 U17674 ( .A1(n17600), .A2(n15029), .A3(n16294), .ZN(n16123) );
  NOR2_X1 U17675 ( .A1(n21271), .A2(n16123), .ZN(n14094) );
  INV_X1 U17676 ( .A(n16291), .ZN(n14070) );
  NOR2_X1 U17677 ( .A1(n14337), .A2(n16385), .ZN(n15031) );
  INV_X1 U17678 ( .A(n15031), .ZN(n21276) );
  INV_X1 U17679 ( .A(n16123), .ZN(n14072) );
  AOI22_X1 U17680 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14072), .B1(n14094), 
        .B2(n21274), .ZN(n14071) );
  AOI22_X1 U17681 ( .A1(n21289), .A2(n14094), .B1(n21288), .B2(n14093), .ZN(
        n14077) );
  NAND2_X1 U17682 ( .A1(n11176), .A2(n14159), .ZN(n15033) );
  NOR2_X1 U17683 ( .A1(n14024), .A2(n15033), .ZN(n14073) );
  INV_X1 U17684 ( .A(n16287), .ZN(n14074) );
  AOI22_X1 U17685 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16155), .B2(n16306), .ZN(n14076) );
  OAI211_X1 U17686 ( .C1(n16395), .C2(n16167), .A(n14077), .B(n14076), .ZN(
        P1_U3042) );
  AOI22_X1 U17687 ( .A1(n21319), .A2(n14094), .B1(n21318), .B2(n14093), .ZN(
        n14079) );
  AOI22_X1 U17688 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16155), .B2(n16329), .ZN(n14078) );
  OAI211_X1 U17689 ( .C1(n16418), .C2(n16167), .A(n14079), .B(n14078), .ZN(
        P1_U3047) );
  AOI22_X1 U17690 ( .A1(n21313), .A2(n14094), .B1(n21312), .B2(n14093), .ZN(
        n14081) );
  AOI22_X1 U17691 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16155), .B2(n16324), .ZN(n14080) );
  OAI211_X1 U17692 ( .C1(n16413), .C2(n16167), .A(n14081), .B(n14080), .ZN(
        P1_U3046) );
  AOI22_X1 U17693 ( .A1(n21307), .A2(n14094), .B1(n21306), .B2(n14093), .ZN(
        n14083) );
  AOI22_X1 U17694 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16155), .B2(n16319), .ZN(n14082) );
  OAI211_X1 U17695 ( .C1(n16408), .C2(n16167), .A(n14083), .B(n14082), .ZN(
        P1_U3045) );
  AOI22_X1 U17696 ( .A1(n21301), .A2(n14094), .B1(n21300), .B2(n14093), .ZN(
        n14085) );
  AOI22_X1 U17697 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16155), .B2(n16314), .ZN(n14084) );
  OAI211_X1 U17698 ( .C1(n16403), .C2(n16167), .A(n14085), .B(n14084), .ZN(
        P1_U3044) );
  AOI22_X1 U17699 ( .A1(n21279), .A2(n14094), .B1(n21278), .B2(n14093), .ZN(
        n14087) );
  AOI22_X1 U17700 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16155), .B2(n16297), .ZN(n14086) );
  OAI211_X1 U17701 ( .C1(n16390), .C2(n16167), .A(n14087), .B(n14086), .ZN(
        P1_U3041) );
  AOI22_X1 U17702 ( .A1(n21327), .A2(n14094), .B1(n21325), .B2(n14093), .ZN(
        n14089) );
  AOI22_X1 U17703 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16155), .B2(n16335), .ZN(n14088) );
  OAI211_X1 U17704 ( .C1(n16426), .C2(n16167), .A(n14089), .B(n14088), .ZN(
        P1_U3048) );
  NAND2_X1 U17705 ( .A1(n14091), .A2(n14090), .ZN(n21748) );
  AOI22_X1 U17706 ( .A1(n21295), .A2(n14094), .B1(n21294), .B2(n14093), .ZN(
        n14097) );
  AOI22_X1 U17707 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9716), .B1(DATAI_26_), 
        .B2(n9715), .ZN(n21299) );
  INV_X1 U17708 ( .A(n21299), .ZN(n21752) );
  AOI22_X1 U17709 ( .A1(n14095), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16155), .B2(n21752), .ZN(n14096) );
  OAI211_X1 U17710 ( .C1(n21758), .C2(n16167), .A(n14097), .B(n14096), .ZN(
        P1_U3043) );
  AND2_X1 U17711 ( .A1(n18182), .A2(n14098), .ZN(n18195) );
  NAND2_X1 U17712 ( .A1(n14112), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14104) );
  NAND2_X1 U17713 ( .A1(n14100), .A2(n14099), .ZN(n14101) );
  OAI21_X1 U17714 ( .B1(n19253), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n14101), .ZN(n14102) );
  INV_X1 U17715 ( .A(n14102), .ZN(n14103) );
  MUX2_X1 U17716 ( .A(n14104), .B(n14103), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n14105) );
  OAI21_X1 U17717 ( .B1(n18195), .B2(n14106), .A(n14105), .ZN(n19937) );
  INV_X1 U17718 ( .A(n18195), .ZN(n14108) );
  NOR2_X1 U17719 ( .A1(n19481), .A2(n19472), .ZN(n14122) );
  INV_X1 U17720 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U17721 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n11932), .B2(n17435), .ZN(
        n14120) );
  NAND2_X1 U17722 ( .A1(n14122), .A2(n14120), .ZN(n14107) );
  OAI211_X1 U17723 ( .C1(n14124), .C2(n14108), .A(n17569), .B(n14107), .ZN(
        n14109) );
  AOI21_X1 U17724 ( .B1(n19937), .B2(n20103), .A(n14109), .ZN(n14110) );
  AOI21_X1 U17725 ( .B1(n14139), .B2(n13924), .A(n14110), .ZN(P3_U3288) );
  NAND2_X1 U17726 ( .A1(n14112), .A2(n14111), .ZN(n14118) );
  NOR2_X1 U17727 ( .A1(n14114), .A2(n14113), .ZN(n14119) );
  AND2_X1 U17728 ( .A1(n19406), .A2(n14115), .ZN(n14133) );
  INV_X1 U17729 ( .A(n14133), .ZN(n14116) );
  NAND2_X1 U17730 ( .A1(n14119), .A2(n14116), .ZN(n14117) );
  NAND2_X1 U17731 ( .A1(n14118), .A2(n14117), .ZN(n19930) );
  INV_X1 U17732 ( .A(n14119), .ZN(n18213) );
  INV_X1 U17733 ( .A(n14120), .ZN(n14121) );
  NAND2_X1 U17734 ( .A1(n14122), .A2(n14121), .ZN(n14123) );
  OAI211_X1 U17735 ( .C1(n14124), .C2(n18213), .A(n17569), .B(n14123), .ZN(
        n14125) );
  AOI21_X1 U17736 ( .B1(n19930), .B2(n20103), .A(n14125), .ZN(n14126) );
  AOI21_X1 U17737 ( .B1(n14139), .B2(n14111), .A(n14126), .ZN(P3_U3289) );
  NAND2_X1 U17738 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14476) );
  XNOR2_X1 U17739 ( .A(n14406), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14132) );
  OR2_X1 U17740 ( .A1(n14129), .A2(n14128), .ZN(n14130) );
  NAND2_X1 U17741 ( .A1(n14127), .A2(n14130), .ZN(n20252) );
  MUX2_X1 U17742 ( .A(n20252), .B(n12850), .S(n16764), .Z(n14131) );
  OAI21_X1 U17743 ( .B1(n14132), .B2(n20283), .A(n14131), .ZN(P2_U2880) );
  NAND2_X1 U17744 ( .A1(n19965), .A2(n11909), .ZN(n14138) );
  MUX2_X1 U17745 ( .A(n19253), .B(n14133), .S(n11909), .Z(n19933) );
  NOR2_X1 U17746 ( .A1(n19933), .A2(n14134), .ZN(n14136) );
  OAI21_X1 U17747 ( .B1(n19481), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17569), .ZN(n14135) );
  OAI22_X1 U17748 ( .A1(n17569), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n14136), .B2(n14135), .ZN(n14137) );
  OAI21_X1 U17749 ( .B1(n14139), .B2(n14138), .A(n14137), .ZN(P3_U3290) );
  INV_X1 U17750 ( .A(n14140), .ZN(n21186) );
  NAND2_X1 U17751 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14142) );
  OAI211_X1 U17752 ( .C1(n17665), .C2(n21183), .A(n14142), .B(n14141), .ZN(
        n14143) );
  AOI21_X1 U17753 ( .B1(n21186), .B2(n17654), .A(n14143), .ZN(n14144) );
  OAI21_X1 U17754 ( .B1(n14145), .B2(n21094), .A(n14144), .ZN(P1_U2996) );
  INV_X1 U17755 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14151) );
  INV_X1 U17756 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14146) );
  NOR2_X1 U17757 ( .A1(n14578), .A2(n14146), .ZN(n14148) );
  INV_X1 U17758 ( .A(n14406), .ZN(n14147) );
  OAI211_X1 U17759 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14148), .A(
        n14147), .B(n20288), .ZN(n14150) );
  NAND2_X1 U17760 ( .A1(n16622), .A2(n20291), .ZN(n14149) );
  OAI211_X1 U17761 ( .C1(n20291), .C2(n14151), .A(n14150), .B(n14149), .ZN(
        P2_U2881) );
  OR2_X1 U17762 ( .A1(n16291), .A2(n14152), .ZN(n16247) );
  OAI21_X1 U17763 ( .B1(n16247), .B2(n14153), .A(n14155), .ZN(n14154) );
  INV_X1 U17764 ( .A(n14155), .ZN(n14183) );
  INV_X1 U17765 ( .A(n16118), .ZN(n14157) );
  OAI22_X1 U17766 ( .A1(n14181), .A2(n16408), .B1(n21311), .B2(n16281), .ZN(
        n14158) );
  AOI21_X1 U17767 ( .B1(n21307), .B2(n14183), .A(n14158), .ZN(n14162) );
  NAND2_X1 U17768 ( .A1(n16079), .A2(n14159), .ZN(n16085) );
  NOR2_X1 U17769 ( .A1(n14160), .A2(n16085), .ZN(n15025) );
  NAND2_X1 U17770 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14161) );
  OAI211_X1 U17771 ( .C1(n16412), .C2(n14187), .A(n14162), .B(n14161), .ZN(
        P1_U3093) );
  OAI22_X1 U17772 ( .A1(n14181), .A2(n16403), .B1(n21305), .B2(n16281), .ZN(
        n14163) );
  AOI21_X1 U17773 ( .B1(n21301), .B2(n14183), .A(n14163), .ZN(n14165) );
  NAND2_X1 U17774 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14164) );
  OAI211_X1 U17775 ( .C1(n16407), .C2(n14187), .A(n14165), .B(n14164), .ZN(
        P1_U3092) );
  OAI22_X1 U17776 ( .A1(n14181), .A2(n16418), .B1(n21323), .B2(n16281), .ZN(
        n14166) );
  AOI21_X1 U17777 ( .B1(n21319), .B2(n14183), .A(n14166), .ZN(n14168) );
  NAND2_X1 U17778 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14167) );
  OAI211_X1 U17779 ( .C1(n16422), .C2(n14187), .A(n14168), .B(n14167), .ZN(
        P1_U3095) );
  OAI22_X1 U17780 ( .A1(n14181), .A2(n16395), .B1(n21293), .B2(n16281), .ZN(
        n14169) );
  AOI21_X1 U17781 ( .B1(n21289), .B2(n14183), .A(n14169), .ZN(n14171) );
  NAND2_X1 U17782 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14170) );
  OAI211_X1 U17783 ( .C1(n16399), .C2(n14187), .A(n14171), .B(n14170), .ZN(
        P1_U3090) );
  OAI22_X1 U17784 ( .A1(n14181), .A2(n16390), .B1(n21287), .B2(n16281), .ZN(
        n14172) );
  AOI21_X1 U17785 ( .B1(n21279), .B2(n14183), .A(n14172), .ZN(n14174) );
  NAND2_X1 U17786 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14173) );
  OAI211_X1 U17787 ( .C1(n16394), .C2(n14187), .A(n14174), .B(n14173), .ZN(
        P1_U3089) );
  OAI22_X1 U17788 ( .A1(n14181), .A2(n21758), .B1(n21299), .B2(n16281), .ZN(
        n14175) );
  AOI21_X1 U17789 ( .B1(n21295), .B2(n14183), .A(n14175), .ZN(n14177) );
  NAND2_X1 U17790 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14176) );
  OAI211_X1 U17791 ( .C1(n21750), .C2(n14187), .A(n14177), .B(n14176), .ZN(
        P1_U3091) );
  OAI22_X1 U17792 ( .A1(n14181), .A2(n16426), .B1(n21334), .B2(n16281), .ZN(
        n14178) );
  AOI21_X1 U17793 ( .B1(n21327), .B2(n14183), .A(n14178), .ZN(n14180) );
  NAND2_X1 U17794 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14179) );
  OAI211_X1 U17795 ( .C1(n16431), .C2(n14187), .A(n14180), .B(n14179), .ZN(
        P1_U3096) );
  OAI22_X1 U17796 ( .A1(n14181), .A2(n16413), .B1(n21317), .B2(n16281), .ZN(
        n14182) );
  AOI21_X1 U17797 ( .B1(n21313), .B2(n14183), .A(n14182), .ZN(n14186) );
  NAND2_X1 U17798 ( .A1(n14184), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14185) );
  OAI211_X1 U17799 ( .C1(n16417), .C2(n14187), .A(n14186), .B(n14185), .ZN(
        P1_U3094) );
  OR2_X1 U17800 ( .A1(n14189), .A2(n14188), .ZN(n14190) );
  NAND2_X1 U17801 ( .A1(n14191), .A2(n14190), .ZN(n16655) );
  XOR2_X1 U17802 ( .A(n16655), .B(n21036), .Z(n14200) );
  OR2_X1 U17803 ( .A1(n14193), .A2(n14192), .ZN(n14194) );
  NAND2_X1 U17804 ( .A1(n14195), .A2(n14194), .ZN(n21047) );
  OR2_X1 U17805 ( .A1(n21043), .A2(n21047), .ZN(n14197) );
  NAND2_X1 U17806 ( .A1(n21043), .A2(n21047), .ZN(n14196) );
  NAND2_X1 U17807 ( .A1(n14197), .A2(n14196), .ZN(n20309) );
  NOR2_X1 U17808 ( .A1(n20309), .A2(n20310), .ZN(n20308) );
  INV_X1 U17809 ( .A(n14197), .ZN(n14198) );
  NOR2_X1 U17810 ( .A1(n20308), .A2(n14198), .ZN(n14199) );
  NOR2_X1 U17811 ( .A1(n14200), .A2(n14199), .ZN(n14564) );
  AOI21_X1 U17812 ( .B1(n14200), .B2(n14199), .A(n14564), .ZN(n14203) );
  INV_X1 U17813 ( .A(n16655), .ZN(n21034) );
  INV_X1 U17814 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20343) );
  OAI22_X1 U17815 ( .A1(n16868), .A2(n21034), .B1(n14282), .B2(n20343), .ZN(
        n14201) );
  AOI21_X1 U17816 ( .B1(n16849), .B2(n14579), .A(n14201), .ZN(n14202) );
  OAI21_X1 U17817 ( .B1(n14203), .B2(n20311), .A(n14202), .ZN(P2_U2917) );
  AND2_X1 U17818 ( .A1(n14204), .A2(n20814), .ZN(n15164) );
  NAND2_X1 U17819 ( .A1(n15164), .A2(n14904), .ZN(n14205) );
  OR2_X1 U17820 ( .A1(n13519), .A2(n14205), .ZN(n14275) );
  INV_X1 U17821 ( .A(n14238), .ZN(n14251) );
  NAND2_X1 U17822 ( .A1(n14207), .A2(n14206), .ZN(n14208) );
  INV_X1 U17823 ( .A(n9747), .ZN(n14946) );
  NAND2_X1 U17824 ( .A1(n14208), .A2(n14946), .ZN(n14235) );
  INV_X1 U17825 ( .A(n14229), .ZN(n14211) );
  INV_X1 U17826 ( .A(n12187), .ZN(n14210) );
  NAND2_X1 U17827 ( .A1(n14210), .A2(n14209), .ZN(n14228) );
  INV_X1 U17828 ( .A(n14228), .ZN(n14234) );
  AOI21_X1 U17829 ( .B1(n12132), .B2(n14211), .A(n14234), .ZN(n14212) );
  NAND2_X1 U17830 ( .A1(n14235), .A2(n14212), .ZN(n14217) );
  INV_X1 U17831 ( .A(n14213), .ZN(n14259) );
  NAND2_X1 U17832 ( .A1(n14259), .A2(n14258), .ZN(n14232) );
  NAND2_X1 U17833 ( .A1(n14232), .A2(n14228), .ZN(n14215) );
  INV_X1 U17834 ( .A(n14946), .ZN(n14954) );
  AOI21_X1 U17835 ( .B1(n12132), .B2(n14229), .A(n14954), .ZN(n14214) );
  NAND2_X1 U17836 ( .A1(n14215), .A2(n14214), .ZN(n14216) );
  MUX2_X1 U17837 ( .A(n14217), .B(n14216), .S(n11984), .Z(n14218) );
  AOI21_X1 U17838 ( .B1(n13953), .B2(n14251), .A(n14218), .ZN(n17421) );
  INV_X1 U17839 ( .A(n14219), .ZN(n14222) );
  NOR2_X1 U17840 ( .A1(n9741), .A2(n14220), .ZN(n14221) );
  NAND2_X1 U17841 ( .A1(n14222), .A2(n14221), .ZN(n14226) );
  NAND4_X1 U17842 ( .A1(n14226), .A2(n14225), .A3(n14224), .A4(n14223), .ZN(
        n17410) );
  NOR2_X1 U17843 ( .A1(n17410), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14227) );
  AOI21_X1 U17844 ( .B1(n17421), .B2(n17410), .A(n14227), .ZN(n14270) );
  NAND2_X1 U17845 ( .A1(n14946), .A2(n14228), .ZN(n14231) );
  AOI22_X1 U17846 ( .A1(n14232), .A2(n14231), .B1(n14230), .B2(n12132), .ZN(
        n14233) );
  OAI21_X1 U17847 ( .B1(n14235), .B2(n14234), .A(n14233), .ZN(n14236) );
  AOI21_X1 U17848 ( .B1(n16661), .B2(n14251), .A(n14236), .ZN(n21018) );
  NOR2_X1 U17849 ( .A1(n17410), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14237) );
  AOI21_X1 U17850 ( .B1(n21018), .B2(n17410), .A(n14237), .ZN(n14269) );
  AND2_X1 U17851 ( .A1(n14269), .A2(n20473), .ZN(n14257) );
  OR2_X1 U17852 ( .A1(n16674), .A2(n14238), .ZN(n14247) );
  INV_X1 U17853 ( .A(n12563), .ZN(n14240) );
  NAND2_X1 U17854 ( .A1(n14240), .A2(n14239), .ZN(n14249) );
  INV_X1 U17855 ( .A(n14241), .ZN(n14244) );
  INV_X1 U17856 ( .A(n14242), .ZN(n14243) );
  NAND2_X1 U17857 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  AOI22_X1 U17858 ( .A1(n14249), .A2(n14245), .B1(n12132), .B2(n9901), .ZN(
        n14246) );
  NAND2_X1 U17859 ( .A1(n14247), .A2(n14246), .ZN(n17417) );
  MUX2_X1 U17860 ( .A(n12132), .B(n14249), .S(n14248), .Z(n14250) );
  AOI21_X1 U17861 ( .B1(n17393), .B2(n14251), .A(n14250), .ZN(n17408) );
  AOI21_X1 U17862 ( .B1(n17408), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U17863 ( .A1(n17408), .A2(n20737), .ZN(n14252) );
  OAI211_X1 U17864 ( .C1(n17417), .C2(n14253), .A(n17410), .B(n14252), .ZN(
        n14255) );
  NOR2_X1 U17865 ( .A1(n14269), .A2(n21692), .ZN(n14254) );
  AOI211_X1 U17866 ( .C1(n17421), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n14255), .B(n14254), .ZN(n14256) );
  AOI211_X1 U17867 ( .C1(n14270), .C2(n21494), .A(n14257), .B(n14256), .ZN(
        n14272) );
  MUX2_X1 U17868 ( .A(n14259), .B(n14258), .S(n14314), .Z(n14262) );
  NAND2_X1 U17869 ( .A1(n12802), .A2(n14260), .ZN(n14261) );
  NAND2_X1 U17870 ( .A1(n14262), .A2(n14261), .ZN(n21054) );
  AND2_X1 U17871 ( .A1(n14263), .A2(n12122), .ZN(n17571) );
  INV_X1 U17872 ( .A(n14264), .ZN(n17570) );
  AOI22_X1 U17873 ( .A1(n17571), .A2(n17570), .B1(n12447), .B2(n21077), .ZN(
        n14267) );
  OAI21_X1 U17874 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n14265), .ZN(n14266) );
  OAI211_X1 U17875 ( .C1(n17410), .C2(n12394), .A(n14267), .B(n14266), .ZN(
        n14268) );
  AOI211_X1 U17876 ( .C1(n14270), .C2(n14269), .A(n21054), .B(n14268), .ZN(
        n14271) );
  OAI21_X1 U17877 ( .B1(n14272), .B2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n14271), .ZN(n14315) );
  OAI21_X1 U17878 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n14315), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14273) );
  AND3_X1 U17879 ( .A1(n21066), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n14273), 
        .ZN(n14274) );
  NAND2_X1 U17880 ( .A1(n14275), .A2(n14274), .ZN(n20927) );
  INV_X1 U17881 ( .A(n20927), .ZN(n14276) );
  OAI21_X1 U17882 ( .B1(n14276), .B2(n21075), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n14277) );
  INV_X1 U17883 ( .A(n17411), .ZN(n17404) );
  NAND2_X1 U17884 ( .A1(n14277), .A2(n17404), .ZN(P2_U3593) );
  OAI21_X1 U17885 ( .B1(n14001), .B2(n14280), .A(n14279), .ZN(n17253) );
  OAI222_X1 U17886 ( .A1(n17253), .A2(n14582), .B1(n14282), .B2(n13553), .C1(
        n14281), .C2(n20315), .ZN(P2_U2904) );
  INV_X1 U17887 ( .A(DATAI_9_), .ZN(n14286) );
  NAND2_X1 U17888 ( .A1(n15585), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14285) );
  OAI21_X1 U17889 ( .B1(n15585), .B2(n14286), .A(n14285), .ZN(n15638) );
  NAND2_X1 U17890 ( .A1(n21231), .A2(n15638), .ZN(n21235) );
  AND2_X2 U17891 ( .A1(n14327), .A2(n14287), .ZN(n21246) );
  AOI22_X1 U17892 ( .A1(n21246), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U17893 ( .A1(n21235), .A2(n14288), .ZN(P1_U2946) );
  NAND2_X1 U17894 ( .A1(n21231), .A2(n15595), .ZN(n14313) );
  AOI22_X1 U17895 ( .A1(n21246), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n14289) );
  NAND2_X1 U17896 ( .A1(n14313), .A2(n14289), .ZN(P1_U2957) );
  NAND2_X1 U17897 ( .A1(n21231), .A2(n15589), .ZN(n14300) );
  AOI22_X1 U17898 ( .A1(n21246), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U17899 ( .A1(n14300), .A2(n14290), .ZN(P1_U2959) );
  NAND2_X1 U17900 ( .A1(n21231), .A2(n15599), .ZN(n14311) );
  AOI22_X1 U17901 ( .A1(n21246), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n14291) );
  NAND2_X1 U17902 ( .A1(n14311), .A2(n14291), .ZN(P1_U2956) );
  INV_X1 U17903 ( .A(n14292), .ZN(n15619) );
  NAND2_X1 U17904 ( .A1(n21231), .A2(n15619), .ZN(n14303) );
  AOI22_X1 U17905 ( .A1(n21246), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U17906 ( .A1(n14303), .A2(n14293), .ZN(P1_U2952) );
  NAND2_X1 U17907 ( .A1(n21231), .A2(n15592), .ZN(n14305) );
  AOI22_X1 U17908 ( .A1(n21246), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n14294) );
  NAND2_X1 U17909 ( .A1(n14305), .A2(n14294), .ZN(P1_U2958) );
  NAND2_X1 U17910 ( .A1(n21231), .A2(n15606), .ZN(n14298) );
  AOI22_X1 U17911 ( .A1(n21246), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U17912 ( .A1(n14298), .A2(n14295), .ZN(P1_U2954) );
  NAND2_X1 U17913 ( .A1(n21231), .A2(n15613), .ZN(n14307) );
  AOI22_X1 U17914 ( .A1(n21246), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14296) );
  NAND2_X1 U17915 ( .A1(n14307), .A2(n14296), .ZN(P1_U2938) );
  AOI22_X1 U17916 ( .A1(n21246), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U17917 ( .A1(n14298), .A2(n14297), .ZN(P1_U2939) );
  AOI22_X1 U17918 ( .A1(n21246), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U17919 ( .A1(n14300), .A2(n14299), .ZN(P1_U2944) );
  NAND2_X1 U17920 ( .A1(n21231), .A2(n15603), .ZN(n14309) );
  AOI22_X1 U17921 ( .A1(n21246), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U17922 ( .A1(n14309), .A2(n14301), .ZN(P1_U2955) );
  AOI22_X1 U17923 ( .A1(n21246), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14302) );
  NAND2_X1 U17924 ( .A1(n14303), .A2(n14302), .ZN(P1_U2937) );
  AOI22_X1 U17925 ( .A1(n21246), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U17926 ( .A1(n14305), .A2(n14304), .ZN(P1_U2943) );
  AOI22_X1 U17927 ( .A1(n21246), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n14306) );
  NAND2_X1 U17928 ( .A1(n14307), .A2(n14306), .ZN(P1_U2953) );
  AOI22_X1 U17929 ( .A1(n21246), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U17930 ( .A1(n14309), .A2(n14308), .ZN(P1_U2940) );
  AOI22_X1 U17931 ( .A1(n21246), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U17932 ( .A1(n14311), .A2(n14310), .ZN(P1_U2941) );
  AOI22_X1 U17933 ( .A1(n21246), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U17934 ( .A1(n14313), .A2(n14312), .ZN(P1_U2942) );
  NOR2_X1 U17935 ( .A1(n20927), .A2(n21073), .ZN(n20931) );
  INV_X1 U17936 ( .A(n17418), .ZN(n21021) );
  AOI21_X1 U17937 ( .B1(n21021), .B2(n21075), .A(n21072), .ZN(n14322) );
  NAND2_X1 U17938 ( .A1(n14315), .A2(n20929), .ZN(n14321) );
  NAND2_X1 U17939 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20864), .ZN(n14400) );
  NOR2_X1 U17940 ( .A1(n14316), .A2(n14400), .ZN(n15172) );
  INV_X1 U17941 ( .A(n15172), .ZN(n14318) );
  OAI211_X1 U17942 ( .C1(n20927), .C2(n21075), .A(n14318), .B(n14317), .ZN(
        n14319) );
  AOI21_X1 U17943 ( .B1(n17411), .B2(n21061), .A(n14319), .ZN(n14320) );
  OAI211_X1 U17944 ( .C1(n20931), .C2(n14322), .A(n14321), .B(n14320), .ZN(
        P2_U3176) );
  INV_X1 U17945 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14328) );
  INV_X1 U17946 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21196) );
  INV_X1 U17947 ( .A(n21231), .ZN(n14326) );
  INV_X1 U17948 ( .A(DATAI_15_), .ZN(n14324) );
  NAND2_X1 U17949 ( .A1(n15585), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U17950 ( .B1(n15585), .B2(n14324), .A(n14323), .ZN(n15624) );
  INV_X1 U17951 ( .A(n15624), .ZN(n14325) );
  OAI222_X1 U17952 ( .A1(n14349), .A2(n14328), .B1(n14327), .B2(n21196), .C1(
        n14326), .C2(n14325), .ZN(P1_U2967) );
  AND2_X1 U17953 ( .A1(n14329), .A2(n14330), .ZN(n14332) );
  OR2_X1 U17954 ( .A1(n14332), .A2(n14331), .ZN(n21152) );
  INV_X1 U17955 ( .A(n14430), .ZN(n15550) );
  AOI21_X1 U17956 ( .B1(n14334), .B2(n14333), .A(n15550), .ZN(n21146) );
  AOI22_X1 U17957 ( .A1(n21146), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14335) );
  OAI21_X1 U17958 ( .B1(n21152), .B2(n15556), .A(n14335), .ZN(P1_U2867) );
  NAND3_X1 U17959 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17600), .A3(
        n16294), .ZN(n16200) );
  NOR2_X1 U17960 ( .A1(n21271), .A2(n16200), .ZN(n14351) );
  OAI22_X1 U17961 ( .A1(n16390), .A2(n16280), .B1(n16238), .B2(n21287), .ZN(
        n14336) );
  AOI21_X1 U17962 ( .B1(n21279), .B2(n14351), .A(n14336), .ZN(n14346) );
  INV_X1 U17963 ( .A(n16247), .ZN(n14339) );
  INV_X1 U17964 ( .A(n14337), .ZN(n14338) );
  AOI21_X1 U17965 ( .B1(n14339), .B2(n14338), .A(n14351), .ZN(n14341) );
  OAI22_X1 U17966 ( .A1(n14341), .A2(n16385), .B1(n16200), .B2(n14687), .ZN(
        n14365) );
  INV_X1 U17967 ( .A(n16200), .ZN(n14344) );
  NAND2_X1 U17968 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n14340), .ZN(n14342) );
  NAND3_X1 U17969 ( .A1(n14342), .A2(n14341), .A3(n21274), .ZN(n14343) );
  OAI211_X1 U17970 ( .C1(n14344), .C2(n21274), .A(n14343), .B(n21281), .ZN(
        n14364) );
  AOI22_X1 U17971 ( .A1(n21278), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__0__SCAN_IN), .B2(n14364), .ZN(n14345) );
  NAND2_X1 U17972 ( .A1(n14346), .A2(n14345), .ZN(P1_U3073) );
  INV_X1 U17973 ( .A(DATAI_10_), .ZN(n21566) );
  NAND2_X1 U17974 ( .A1(n15585), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14347) );
  OAI21_X1 U17975 ( .B1(n15585), .B2(n21566), .A(n14347), .ZN(n15634) );
  NAND2_X1 U17976 ( .A1(n21231), .A2(n15634), .ZN(n21237) );
  NAND2_X1 U17977 ( .A1(n21245), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14348) );
  OAI211_X1 U17978 ( .C1(n21648), .C2(n14349), .A(n21237), .B(n14348), .ZN(
        P1_U2947) );
  OAI222_X1 U17979 ( .A1(n21152), .A2(n15643), .B1(n15646), .B2(n14350), .C1(
        n15644), .C2(n11222), .ZN(P1_U2899) );
  AOI22_X1 U17980 ( .A1(n21288), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n14364), .ZN(n14353) );
  INV_X1 U17981 ( .A(n16395), .ZN(n21290) );
  AOI22_X1 U17982 ( .A1(n14366), .A2(n21290), .B1(n16197), .B2(n16306), .ZN(
        n14352) );
  OAI211_X1 U17983 ( .C1(n16304), .C2(n14369), .A(n14353), .B(n14352), .ZN(
        P1_U3074) );
  AOI22_X1 U17984 ( .A1(n21318), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n14364), .ZN(n14355) );
  INV_X1 U17985 ( .A(n16418), .ZN(n21320) );
  AOI22_X1 U17986 ( .A1(n14366), .A2(n21320), .B1(n16197), .B2(n16329), .ZN(
        n14354) );
  OAI211_X1 U17987 ( .C1(n16327), .C2(n14369), .A(n14355), .B(n14354), .ZN(
        P1_U3079) );
  AOI22_X1 U17988 ( .A1(n21312), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__5__SCAN_IN), .B2(n14364), .ZN(n14357) );
  INV_X1 U17989 ( .A(n16413), .ZN(n21314) );
  AOI22_X1 U17990 ( .A1(n14366), .A2(n21314), .B1(n16197), .B2(n16324), .ZN(
        n14356) );
  OAI211_X1 U17991 ( .C1(n16322), .C2(n14369), .A(n14357), .B(n14356), .ZN(
        P1_U3078) );
  AOI22_X1 U17992 ( .A1(n21300), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n14364), .ZN(n14359) );
  INV_X1 U17993 ( .A(n16403), .ZN(n21302) );
  AOI22_X1 U17994 ( .A1(n14366), .A2(n21302), .B1(n16197), .B2(n16314), .ZN(
        n14358) );
  OAI211_X1 U17995 ( .C1(n16312), .C2(n14369), .A(n14359), .B(n14358), .ZN(
        P1_U3076) );
  AOI22_X1 U17996 ( .A1(n21325), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n14364), .ZN(n14361) );
  INV_X1 U17997 ( .A(n16426), .ZN(n21328) );
  AOI22_X1 U17998 ( .A1(n14366), .A2(n21328), .B1(n16197), .B2(n16335), .ZN(
        n14360) );
  OAI211_X1 U17999 ( .C1(n16333), .C2(n14369), .A(n14361), .B(n14360), .ZN(
        P1_U3080) );
  AOI22_X1 U18000 ( .A1(n21294), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n14364), .ZN(n14363) );
  INV_X1 U18001 ( .A(n21758), .ZN(n21296) );
  AOI22_X1 U18002 ( .A1(n14366), .A2(n21296), .B1(n16197), .B2(n21752), .ZN(
        n14362) );
  OAI211_X1 U18003 ( .C1(n21748), .C2(n14369), .A(n14363), .B(n14362), .ZN(
        P1_U3075) );
  AOI22_X1 U18004 ( .A1(n21306), .A2(n14365), .B1(
        P1_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n14364), .ZN(n14368) );
  INV_X1 U18005 ( .A(n16408), .ZN(n21308) );
  AOI22_X1 U18006 ( .A1(n14366), .A2(n21308), .B1(n16197), .B2(n16319), .ZN(
        n14367) );
  OAI211_X1 U18007 ( .C1(n16317), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        P1_U3077) );
  AOI21_X1 U18008 ( .B1(n14370), .B2(n13961), .A(n10120), .ZN(n21167) );
  INV_X1 U18009 ( .A(n21167), .ZN(n14422) );
  INV_X1 U18010 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21213) );
  OAI222_X1 U18011 ( .A1(n14422), .A2(n15643), .B1(n15646), .B2(n14371), .C1(
        n15644), .C2(n21213), .ZN(P1_U2900) );
  INV_X1 U18012 ( .A(n14372), .ZN(n14373) );
  AOI22_X1 U18013 ( .A1(n14375), .A2(n14374), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14373), .ZN(n17659) );
  XNOR2_X1 U18014 ( .A(n17659), .B(n17658), .ZN(n17661) );
  XNOR2_X1 U18015 ( .A(n17661), .B(n17660), .ZN(n14389) );
  NAND2_X1 U18016 ( .A1(n13964), .A2(n14376), .ZN(n14377) );
  NAND2_X1 U18017 ( .A1(n14333), .A2(n14377), .ZN(n21160) );
  INV_X1 U18018 ( .A(n21160), .ZN(n14383) );
  NAND2_X1 U18019 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14378), .ZN(
        n14381) );
  OAI211_X1 U18020 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n17692), .B(n14427), .ZN(n14380) );
  NOR2_X1 U18021 ( .A1(n17669), .A2(n21363), .ZN(n14385) );
  INV_X1 U18022 ( .A(n14385), .ZN(n14379) );
  NAND3_X1 U18023 ( .A1(n14381), .A2(n14380), .A3(n14379), .ZN(n14382) );
  AOI21_X1 U18024 ( .B1(n21250), .B2(n14383), .A(n14382), .ZN(n14384) );
  OAI21_X1 U18025 ( .B1(n14389), .B2(n16064), .A(n14384), .ZN(P1_U3027) );
  AOI21_X1 U18026 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14385), .ZN(n14386) );
  OAI21_X1 U18027 ( .B1(n21171), .B2(n17665), .A(n14386), .ZN(n14387) );
  AOI21_X1 U18028 ( .B1(n21167), .B2(n17654), .A(n14387), .ZN(n14388) );
  OAI21_X1 U18029 ( .B1(n14389), .B2(n21094), .A(n14388), .ZN(P1_U2995) );
  NOR2_X1 U18030 ( .A1(n20422), .A2(n20814), .ZN(n20673) );
  NOR2_X1 U18031 ( .A1(n20539), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U18032 ( .A1(n20863), .A2(n21050), .ZN(n14595) );
  INV_X1 U18033 ( .A(n14595), .ZN(n14391) );
  NAND2_X1 U18034 ( .A1(n14390), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U18035 ( .A1(n20673), .A2(n14392), .B1(n14391), .B2(n17401), .ZN(
        n14397) );
  INV_X1 U18036 ( .A(n20863), .ZN(n20819) );
  NOR2_X1 U18037 ( .A1(n20819), .A2(n20672), .ZN(n20806) );
  NOR3_X2 U18038 ( .A1(n14397), .A2(n20823), .A3(n14401), .ZN(n20812) );
  INV_X1 U18039 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14405) );
  INV_X1 U18040 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17767) );
  INV_X1 U18041 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17829) );
  OAI22_X2 U18042 ( .A1(n17767), .A2(n20391), .B1(n17829), .B2(n20393), .ZN(
        n20876) );
  AOI22_X1 U18043 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20405), .ZN(n20879) );
  INV_X1 U18044 ( .A(n20879), .ZN(n20828) );
  AOI22_X1 U18045 ( .A1(n20808), .A2(n20876), .B1(n20857), .B2(n20828), .ZN(
        n14404) );
  NOR2_X2 U18046 ( .A1(n20823), .A2(n14402), .ZN(n20867) );
  AOI22_X1 U18047 ( .A1(n20807), .A2(n20867), .B1(n20866), .B2(n20806), .ZN(
        n14403) );
  OAI211_X1 U18048 ( .C1(n20812), .C2(n14405), .A(n14404), .B(n14403), .ZN(
        P2_U3152) );
  NAND2_X1 U18049 ( .A1(n14406), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14416) );
  XNOR2_X1 U18050 ( .A(n14617), .B(n14616), .ZN(n14413) );
  AND2_X1 U18051 ( .A1(n14408), .A2(n14409), .ZN(n14411) );
  OR2_X1 U18052 ( .A1(n14411), .A2(n14410), .ZN(n17324) );
  MUX2_X1 U18053 ( .A(n17324), .B(n10375), .S(n16764), .Z(n14412) );
  OAI21_X1 U18054 ( .B1(n14413), .B2(n20283), .A(n14412), .ZN(P2_U2878) );
  INV_X1 U18055 ( .A(n14408), .ZN(n14414) );
  AOI21_X1 U18056 ( .B1(n14415), .B2(n14127), .A(n14414), .ZN(n20237) );
  INV_X1 U18057 ( .A(n20237), .ZN(n14421) );
  INV_X1 U18058 ( .A(n14416), .ZN(n14418) );
  INV_X1 U18059 ( .A(n14617), .ZN(n14417) );
  OAI211_X1 U18060 ( .C1(n14418), .C2(n14474), .A(n14417), .B(n20288), .ZN(
        n14420) );
  NAND2_X1 U18061 ( .A1(n16764), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14419) );
  OAI211_X1 U18062 ( .C1(n14421), .C2(n16764), .A(n14420), .B(n14419), .ZN(
        P2_U2879) );
  OAI222_X1 U18063 ( .A1(n21160), .A2(n15545), .B1(n15544), .B2(n13048), .C1(
        n15530), .C2(n14422), .ZN(P1_U2868) );
  XOR2_X1 U18064 ( .A(n14424), .B(n14423), .Z(n14524) );
  OR2_X1 U18065 ( .A1(n14427), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17700) );
  AND2_X1 U18066 ( .A1(n16052), .A2(n16027), .ZN(n14426) );
  INV_X1 U18067 ( .A(n16055), .ZN(n14425) );
  AOI211_X1 U18068 ( .C1(n14427), .C2(n15965), .A(n14426), .B(n14425), .ZN(
        n17696) );
  OAI21_X1 U18069 ( .B1(n14428), .B2(n17700), .A(n17696), .ZN(n17672) );
  NAND2_X1 U18070 ( .A1(n17692), .A2(n14429), .ZN(n16049) );
  XNOR2_X1 U18071 ( .A(n14430), .B(n15549), .ZN(n21135) );
  INV_X1 U18072 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21367) );
  NOR2_X1 U18073 ( .A1(n17669), .A2(n21367), .ZN(n14519) );
  AOI21_X1 U18074 ( .B1(n21250), .B2(n21135), .A(n14519), .ZN(n14431) );
  OAI21_X1 U18075 ( .B1(n16049), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14431), .ZN(n14432) );
  AOI21_X1 U18076 ( .B1(n17672), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14432), .ZN(n14433) );
  OAI21_X1 U18077 ( .B1(n16064), .B2(n14524), .A(n14433), .ZN(P1_U3025) );
  AND2_X1 U18078 ( .A1(n11176), .A2(n16346), .ZN(n14434) );
  OAI21_X1 U18079 ( .B1(n21753), .B2(n21266), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14435) );
  NAND2_X1 U18080 ( .A1(n14435), .A2(n21274), .ZN(n14446) );
  INV_X1 U18081 ( .A(n14446), .ZN(n14437) );
  AND2_X1 U18082 ( .A1(n15053), .A2(n16341), .ZN(n14445) );
  OR2_X1 U18083 ( .A1(n16164), .A2(n17600), .ZN(n14440) );
  INV_X1 U18084 ( .A(n14440), .ZN(n16343) );
  NOR2_X1 U18085 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14438), .ZN(
        n14441) );
  INV_X1 U18086 ( .A(n14441), .ZN(n14468) );
  OAI22_X1 U18087 ( .A1(n16317), .A2(n14468), .B1(n21311), .B2(n14467), .ZN(
        n14439) );
  AOI21_X1 U18088 ( .B1(n21753), .B2(n21308), .A(n14439), .ZN(n14448) );
  NAND2_X1 U18089 ( .A1(n14440), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16350) );
  OAI21_X1 U18090 ( .B1(n17711), .B2(n14441), .A(n16350), .ZN(n14442) );
  INV_X1 U18091 ( .A(n14442), .ZN(n14444) );
  NAND2_X1 U18092 ( .A1(n14443), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16248) );
  INV_X1 U18093 ( .A(n16202), .ZN(n15019) );
  NAND2_X1 U18094 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14447) );
  OAI211_X1 U18095 ( .C1(n14473), .C2(n16412), .A(n14448), .B(n14447), .ZN(
        P1_U3117) );
  OAI22_X1 U18096 ( .A1(n16322), .A2(n14468), .B1(n21317), .B2(n14467), .ZN(
        n14449) );
  AOI21_X1 U18097 ( .B1(n21753), .B2(n21314), .A(n14449), .ZN(n14451) );
  NAND2_X1 U18098 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14450) );
  OAI211_X1 U18099 ( .C1(n14473), .C2(n16417), .A(n14451), .B(n14450), .ZN(
        P1_U3118) );
  OAI22_X1 U18100 ( .A1(n16333), .A2(n14468), .B1(n21334), .B2(n14467), .ZN(
        n14452) );
  AOI21_X1 U18101 ( .B1(n21753), .B2(n21328), .A(n14452), .ZN(n14454) );
  NAND2_X1 U18102 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n14453) );
  OAI211_X1 U18103 ( .C1(n14473), .C2(n16431), .A(n14454), .B(n14453), .ZN(
        P1_U3120) );
  OAI22_X1 U18104 ( .A1(n21748), .A2(n14468), .B1(n21299), .B2(n14467), .ZN(
        n14455) );
  AOI21_X1 U18105 ( .B1(n21753), .B2(n21296), .A(n14455), .ZN(n14457) );
  NAND2_X1 U18106 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14456) );
  OAI211_X1 U18107 ( .C1(n14473), .C2(n21750), .A(n14457), .B(n14456), .ZN(
        P1_U3115) );
  OAI22_X1 U18108 ( .A1(n16327), .A2(n14468), .B1(n21323), .B2(n14467), .ZN(
        n14458) );
  AOI21_X1 U18109 ( .B1(n21753), .B2(n21320), .A(n14458), .ZN(n14460) );
  NAND2_X1 U18110 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14459) );
  OAI211_X1 U18111 ( .C1(n14473), .C2(n16422), .A(n14460), .B(n14459), .ZN(
        P1_U3119) );
  INV_X1 U18112 ( .A(n16390), .ZN(n21284) );
  OAI22_X1 U18113 ( .A1(n16295), .A2(n14468), .B1(n21287), .B2(n14467), .ZN(
        n14461) );
  AOI21_X1 U18114 ( .B1(n21753), .B2(n21284), .A(n14461), .ZN(n14463) );
  NAND2_X1 U18115 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14462) );
  OAI211_X1 U18116 ( .C1(n14473), .C2(n16394), .A(n14463), .B(n14462), .ZN(
        P1_U3113) );
  OAI22_X1 U18117 ( .A1(n16312), .A2(n14468), .B1(n21305), .B2(n14467), .ZN(
        n14464) );
  AOI21_X1 U18118 ( .B1(n21753), .B2(n21302), .A(n14464), .ZN(n14466) );
  NAND2_X1 U18119 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14465) );
  OAI211_X1 U18120 ( .C1(n14473), .C2(n16407), .A(n14466), .B(n14465), .ZN(
        P1_U3116) );
  OAI22_X1 U18121 ( .A1(n16304), .A2(n14468), .B1(n21293), .B2(n14467), .ZN(
        n14469) );
  AOI21_X1 U18122 ( .B1(n21753), .B2(n21290), .A(n14469), .ZN(n14472) );
  NAND2_X1 U18123 ( .A1(n14470), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14471) );
  OAI211_X1 U18124 ( .C1(n14473), .C2(n16399), .A(n14472), .B(n14471), .ZN(
        P1_U3114) );
  INV_X1 U18125 ( .A(n16757), .ZN(n14481) );
  AND2_X1 U18126 ( .A1(n14616), .A2(n14474), .ZN(n14480) );
  INV_X1 U18127 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14475) );
  NOR2_X1 U18128 ( .A1(n14476), .A2(n14475), .ZN(n14479) );
  AND2_X1 U18129 ( .A1(n14618), .A2(n14477), .ZN(n14478) );
  NAND4_X1 U18130 ( .A1(n14481), .A2(n14480), .A3(n14479), .A4(n14478), .ZN(
        n14496) );
  OR2_X1 U18131 ( .A1(n14578), .A2(n14496), .ZN(n16760) );
  NOR2_X1 U18132 ( .A1(n16760), .A2(n14583), .ZN(n14531) );
  NAND2_X1 U18133 ( .A1(n14531), .A2(n14530), .ZN(n14623) );
  NOR2_X1 U18134 ( .A1(n14623), .A2(n14622), .ZN(n14500) );
  AOI22_X1 U18135 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14485) );
  AOI22_X1 U18136 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14484) );
  AOI22_X1 U18137 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U18138 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14482) );
  NAND4_X1 U18139 ( .A1(n14485), .A2(n14484), .A3(n14483), .A4(n14482), .ZN(
        n14491) );
  AOI22_X1 U18140 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14489) );
  AOI22_X1 U18141 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U18142 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U18143 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14486) );
  NAND4_X1 U18144 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        n14490) );
  OR2_X1 U18145 ( .A1(n14491), .A2(n14490), .ZN(n14499) );
  AND2_X1 U18146 ( .A1(n14499), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14494) );
  NAND4_X1 U18147 ( .A1(n14494), .A2(n14493), .A3(n14530), .A4(n14492), .ZN(
        n14495) );
  NOR3_X1 U18148 ( .A1(n14496), .A2(n14897), .A3(n14495), .ZN(n14497) );
  OAI21_X1 U18149 ( .B1(n14500), .B2(n14499), .A(n14641), .ZN(n14650) );
  INV_X1 U18150 ( .A(n14501), .ZN(n14502) );
  AOI21_X1 U18151 ( .B1(n14503), .B2(n14279), .A(n14502), .ZN(n20176) );
  INV_X1 U18152 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U18153 ( .A1(n14507), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U18154 ( .A1(n16858), .A2(n14508), .B1(n20306), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14509) );
  OAI211_X1 U18155 ( .C1(n14511), .C2(n16859), .A(n14510), .B(n14509), .ZN(
        n14512) );
  AOI21_X1 U18156 ( .B1(n20176), .B2(n20307), .A(n14512), .ZN(n14513) );
  OAI21_X1 U18157 ( .B1(n20311), .B2(n14650), .A(n14513), .ZN(P2_U2903) );
  INV_X1 U18158 ( .A(n14514), .ZN(n14517) );
  INV_X1 U18159 ( .A(n14331), .ZN(n14516) );
  AOI21_X1 U18160 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14522) );
  INV_X1 U18161 ( .A(n14522), .ZN(n21138) );
  AOI22_X1 U18162 ( .A1(n21135), .A2(n15554), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n15553), .ZN(n14518) );
  OAI21_X1 U18163 ( .B1(n21138), .B2(n15530), .A(n14518), .ZN(P1_U2866) );
  AOI21_X1 U18164 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14519), .ZN(n14520) );
  OAI21_X1 U18165 ( .B1(n21136), .B2(n17665), .A(n14520), .ZN(n14521) );
  AOI21_X1 U18166 ( .B1(n14522), .B2(n17654), .A(n14521), .ZN(n14523) );
  OAI21_X1 U18167 ( .B1(n21094), .B2(n14524), .A(n14523), .ZN(P1_U2993) );
  AND2_X1 U18168 ( .A1(n14526), .A2(n14525), .ZN(n14625) );
  INV_X1 U18169 ( .A(n14526), .ZN(n16754) );
  NOR2_X1 U18170 ( .A1(n16754), .A2(n14527), .ZN(n14588) );
  NOR2_X1 U18171 ( .A1(n14588), .A2(n14528), .ZN(n14529) );
  OAI211_X1 U18172 ( .C1(n14531), .C2(n14530), .A(n14623), .B(n20288), .ZN(
        n14533) );
  NAND2_X1 U18173 ( .A1(n16764), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14532) );
  OAI211_X1 U18174 ( .C1(n20191), .C2(n16764), .A(n14533), .B(n14532), .ZN(
        P2_U2873) );
  OAI222_X1 U18175 ( .A1(n21138), .A2(n15643), .B1(n15646), .B2(n14534), .C1(
        n15644), .C2(n11229), .ZN(P1_U2898) );
  NAND2_X1 U18176 ( .A1(n16079), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16084) );
  INV_X1 U18177 ( .A(n16084), .ZN(n15023) );
  AOI21_X1 U18178 ( .B1(n14541), .B2(n15023), .A(n16385), .ZN(n14538) );
  INV_X1 U18179 ( .A(n16159), .ZN(n14536) );
  AOI21_X1 U18180 ( .B1(n14536), .B2(n16382), .A(n10457), .ZN(n14540) );
  NAND3_X1 U18181 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17600), .A3(
        n15029), .ZN(n16161) );
  AOI22_X1 U18182 ( .A1(n14538), .A2(n14540), .B1(n16385), .B2(n16161), .ZN(
        n14537) );
  NAND2_X1 U18183 ( .A1(n21281), .A2(n14537), .ZN(n14557) );
  INV_X1 U18184 ( .A(n14538), .ZN(n14539) );
  AOI22_X1 U18185 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n14557), .B1(
        n21278), .B2(n14556), .ZN(n14543) );
  AOI22_X1 U18186 ( .A1(n21279), .A2(n10457), .B1(n14558), .B2(n16297), .ZN(
        n14542) );
  OAI211_X1 U18187 ( .C1(n16390), .C2(n16237), .A(n14543), .B(n14542), .ZN(
        P1_U3057) );
  AOI22_X1 U18188 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14557), .B1(
        n21325), .B2(n14556), .ZN(n14545) );
  AOI22_X1 U18189 ( .A1(n21327), .A2(n10457), .B1(n14558), .B2(n16335), .ZN(
        n14544) );
  OAI211_X1 U18190 ( .C1(n16426), .C2(n16237), .A(n14545), .B(n14544), .ZN(
        P1_U3064) );
  AOI22_X1 U18191 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14557), .B1(
        n21318), .B2(n14556), .ZN(n14547) );
  AOI22_X1 U18192 ( .A1(n21319), .A2(n10457), .B1(n14558), .B2(n16329), .ZN(
        n14546) );
  OAI211_X1 U18193 ( .C1(n16418), .C2(n16237), .A(n14547), .B(n14546), .ZN(
        P1_U3063) );
  AOI22_X1 U18194 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14557), .B1(
        n21312), .B2(n14556), .ZN(n14549) );
  AOI22_X1 U18195 ( .A1(n21313), .A2(n10457), .B1(n14558), .B2(n16324), .ZN(
        n14548) );
  OAI211_X1 U18196 ( .C1(n16413), .C2(n16237), .A(n14549), .B(n14548), .ZN(
        P1_U3062) );
  AOI22_X1 U18197 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14557), .B1(
        n21300), .B2(n14556), .ZN(n14551) );
  AOI22_X1 U18198 ( .A1(n21301), .A2(n10457), .B1(n14558), .B2(n16314), .ZN(
        n14550) );
  OAI211_X1 U18199 ( .C1(n16403), .C2(n16237), .A(n14551), .B(n14550), .ZN(
        P1_U3060) );
  AOI22_X1 U18200 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14557), .B1(
        n21306), .B2(n14556), .ZN(n14553) );
  AOI22_X1 U18201 ( .A1(n21307), .A2(n10457), .B1(n14558), .B2(n16319), .ZN(
        n14552) );
  OAI211_X1 U18202 ( .C1(n16408), .C2(n16237), .A(n14553), .B(n14552), .ZN(
        P1_U3061) );
  AOI22_X1 U18203 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14557), .B1(
        n21288), .B2(n14556), .ZN(n14555) );
  AOI22_X1 U18204 ( .A1(n21289), .A2(n10457), .B1(n14558), .B2(n16306), .ZN(
        n14554) );
  OAI211_X1 U18205 ( .C1(n16395), .C2(n16237), .A(n14555), .B(n14554), .ZN(
        P1_U3058) );
  AOI22_X1 U18206 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14557), .B1(
        n21294), .B2(n14556), .ZN(n14560) );
  AOI22_X1 U18207 ( .A1(n21295), .A2(n10457), .B1(n14558), .B2(n21752), .ZN(
        n14559) );
  OAI211_X1 U18208 ( .C1(n21758), .C2(n16237), .A(n14560), .B(n14559), .ZN(
        P1_U3059) );
  XNOR2_X1 U18209 ( .A(n14562), .B(n14563), .ZN(n17373) );
  AOI21_X1 U18210 ( .B1(n21034), .B2(n21036), .A(n14564), .ZN(n20301) );
  NAND2_X1 U18211 ( .A1(n14567), .A2(n14566), .ZN(n14568) );
  NAND2_X1 U18212 ( .A1(n14565), .A2(n14568), .ZN(n16645) );
  XNOR2_X1 U18213 ( .A(n20422), .B(n16645), .ZN(n20300) );
  NOR2_X1 U18214 ( .A1(n20301), .A2(n20300), .ZN(n20299) );
  NOR2_X1 U18215 ( .A1(n21030), .A2(n21029), .ZN(n14571) );
  NAND2_X1 U18216 ( .A1(n14565), .A2(n14569), .ZN(n14570) );
  NAND2_X1 U18217 ( .A1(n14562), .A2(n14570), .ZN(n20292) );
  OAI21_X1 U18218 ( .B1(n20299), .B2(n14571), .A(n20292), .ZN(n20294) );
  INV_X1 U18219 ( .A(n14572), .ZN(n14573) );
  NAND2_X1 U18220 ( .A1(n14574), .A2(n14573), .ZN(n14575) );
  OR2_X1 U18221 ( .A1(n14576), .A2(n14575), .ZN(n14577) );
  NAND2_X1 U18222 ( .A1(n14578), .A2(n14577), .ZN(n20293) );
  INV_X1 U18223 ( .A(n20293), .ZN(n20289) );
  NAND3_X1 U18224 ( .A1(n20294), .A2(n20295), .A3(n20289), .ZN(n14581) );
  AOI22_X1 U18225 ( .A1(n14579), .A2(n20396), .B1(n20306), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n14580) );
  OAI211_X1 U18226 ( .C1(n17373), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        P2_U2914) );
  XNOR2_X1 U18227 ( .A(n16760), .B(n14583), .ZN(n14591) );
  INV_X1 U18228 ( .A(n16753), .ZN(n14585) );
  AND2_X1 U18229 ( .A1(n14619), .A2(n14585), .ZN(n14586) );
  NAND2_X1 U18230 ( .A1(n14584), .A2(n14586), .ZN(n16756) );
  AND2_X1 U18231 ( .A1(n16756), .A2(n14587), .ZN(n14589) );
  MUX2_X1 U18232 ( .A(n17281), .B(n12861), .S(n16764), .Z(n14590) );
  OAI21_X1 U18233 ( .B1(n14591), .B2(n20283), .A(n14590), .ZN(P2_U2874) );
  OAI21_X1 U18234 ( .B1(n20787), .B2(n20808), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14599) );
  INV_X1 U18235 ( .A(n20818), .ZN(n14593) );
  NAND2_X1 U18236 ( .A1(n14593), .A2(n14592), .ZN(n20511) );
  OR2_X1 U18237 ( .A1(n21494), .A2(n20511), .ZN(n14598) );
  AOI21_X1 U18238 ( .B1(n14594), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14596) );
  OAI21_X1 U18239 ( .B1(n14596), .B2(n20785), .A(n20874), .ZN(n14597) );
  INV_X1 U18240 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14607) );
  INV_X1 U18241 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17762) );
  INV_X1 U18242 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U18243 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20405), .ZN(n20897) );
  AOI22_X1 U18244 ( .A1(n20787), .A2(n20894), .B1(n20808), .B2(n20839), .ZN(
        n14606) );
  INV_X1 U18245 ( .A(n14600), .ZN(n14603) );
  OAI21_X1 U18246 ( .B1(n14601), .B2(n20785), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14602) );
  NOR2_X2 U18247 ( .A1(n20823), .A2(n20305), .ZN(n20893) );
  AOI22_X1 U18248 ( .A1(n20786), .A2(n20893), .B1(n20785), .B2(n20892), .ZN(
        n14605) );
  OAI211_X1 U18249 ( .C1(n20790), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        P2_U3147) );
  INV_X1 U18250 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14612) );
  INV_X1 U18251 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17831) );
  INV_X1 U18252 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17764) );
  AOI22_X1 U18253 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20405), .ZN(n20891) );
  AOI22_X1 U18254 ( .A1(n20787), .A2(n20888), .B1(n20808), .B2(n20835), .ZN(
        n14611) );
  NOR2_X2 U18255 ( .A1(n20823), .A2(n14608), .ZN(n20887) );
  AOI22_X1 U18256 ( .A1(n20786), .A2(n20887), .B1(n20785), .B2(n20886), .ZN(
        n14610) );
  OAI211_X1 U18257 ( .C1(n20790), .C2(n14612), .A(n14611), .B(n14610), .ZN(
        P2_U3146) );
  INV_X1 U18258 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14615) );
  AOI22_X1 U18259 ( .A1(n20787), .A2(n20876), .B1(n20808), .B2(n20828), .ZN(
        n14614) );
  AOI22_X1 U18260 ( .A1(n20786), .A2(n20867), .B1(n20866), .B2(n20785), .ZN(
        n14613) );
  OAI211_X1 U18261 ( .C1(n20790), .C2(n14615), .A(n14614), .B(n14613), .ZN(
        P2_U3144) );
  NAND2_X1 U18262 ( .A1(n14617), .A2(n14616), .ZN(n20284) );
  NOR2_X1 U18263 ( .A1(n20284), .A2(n20285), .ZN(n20282) );
  XNOR2_X1 U18264 ( .A(n20282), .B(n14618), .ZN(n14621) );
  OAI21_X1 U18265 ( .B1(n14584), .B2(n14619), .A(n16754), .ZN(n17040) );
  MUX2_X1 U18266 ( .A(n12906), .B(n17040), .S(n20291), .Z(n14620) );
  OAI21_X1 U18267 ( .B1(n14621), .B2(n20283), .A(n14620), .ZN(P2_U2876) );
  XNOR2_X1 U18268 ( .A(n14623), .B(n14622), .ZN(n14628) );
  OR2_X1 U18269 ( .A1(n14625), .A2(n14624), .ZN(n14626) );
  NAND2_X1 U18270 ( .A1(n14645), .A2(n14626), .ZN(n17247) );
  MUX2_X1 U18271 ( .A(n12913), .B(n17247), .S(n20291), .Z(n14627) );
  OAI21_X1 U18272 ( .B1(n14628), .B2(n20283), .A(n14627), .ZN(P2_U2872) );
  OAI21_X1 U18273 ( .B1(n9911), .B2(n9910), .A(n14630), .ZN(n16964) );
  AOI22_X1 U18274 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12352), .B1(
        n14803), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U18275 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14633) );
  AOI22_X1 U18276 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12349), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U18277 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12252), .B1(
        n12273), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14631) );
  NAND4_X1 U18278 ( .A1(n14634), .A2(n14633), .A3(n14632), .A4(n14631), .ZN(
        n14640) );
  AOI22_X1 U18279 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12278), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U18280 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12245), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U18281 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12232), .B1(
        n12231), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U18282 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12234), .B1(
        n12233), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14635) );
  NAND4_X1 U18283 ( .A1(n14638), .A2(n14637), .A3(n14636), .A4(n14635), .ZN(
        n14639) );
  NOR2_X1 U18284 ( .A1(n14640), .A2(n14639), .ZN(n14642) );
  AOI21_X1 U18285 ( .B1(n14642), .B2(n14641), .A(n14740), .ZN(n16866) );
  AOI22_X1 U18286 ( .A1(n16866), .A2(n20288), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16764), .ZN(n14643) );
  OAI21_X1 U18287 ( .B1(n16964), .B2(n16764), .A(n14643), .ZN(P2_U2870) );
  NAND2_X1 U18288 ( .A1(n14645), .A2(n14644), .ZN(n14646) );
  NAND2_X1 U18289 ( .A1(n14647), .A2(n14646), .ZN(n17235) );
  NOR2_X1 U18290 ( .A1(n17235), .A2(n16764), .ZN(n14648) );
  AOI21_X1 U18291 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16764), .A(n14648), .ZN(
        n14649) );
  OAI21_X1 U18292 ( .B1(n20283), .B2(n14650), .A(n14649), .ZN(P2_U2871) );
  OR2_X1 U18293 ( .A1(n14709), .A2(n14651), .ZN(n14652) );
  OAI211_X1 U18294 ( .C1(n14707), .C2(n17379), .A(n14652), .B(n17396), .ZN(
        n14655) );
  NOR2_X1 U18295 ( .A1(n14709), .A2(n17379), .ZN(n14654) );
  MUX2_X1 U18296 ( .A(n14655), .B(n14654), .S(n14653), .Z(n14666) );
  AOI22_X1 U18297 ( .A1(n17726), .A2(n14656), .B1(n20355), .B2(n16655), .ZN(
        n14664) );
  AOI21_X1 U18298 ( .B1(n20356), .B2(n16661), .A(n14657), .ZN(n14663) );
  NAND2_X1 U18299 ( .A1(n14659), .A2(n14658), .ZN(n14660) );
  OR2_X1 U18300 ( .A1(n20360), .A2(n14660), .ZN(n14661) );
  NAND4_X1 U18301 ( .A1(n14664), .A2(n14663), .A3(n14662), .A4(n14661), .ZN(
        n14665) );
  OR2_X1 U18302 ( .A1(n14666), .A2(n14665), .ZN(P2_U3044) );
  AOI21_X1 U18303 ( .B1(n14667), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17566) );
  NAND2_X1 U18304 ( .A1(n10611), .A2(n17566), .ZN(n19483) );
  NOR2_X1 U18305 ( .A1(n19483), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(n14668) );
  OAI21_X1 U18306 ( .B1(n14668), .B2(n20068), .A(n19565), .ZN(n19488) );
  INV_X1 U18307 ( .A(n19488), .ZN(n14669) );
  AOI22_X1 U18308 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n17560), .B2(n19105), .ZN(n17563) );
  NOR2_X1 U18309 ( .A1(n14669), .A2(n17563), .ZN(n14671) );
  NAND2_X1 U18310 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n10656), .ZN(n19566) );
  NAND2_X1 U18311 ( .A1(n19566), .A2(n19488), .ZN(n17561) );
  OR2_X1 U18312 ( .A1(n19837), .A2(n17561), .ZN(n14670) );
  MUX2_X1 U18313 ( .A(n14671), .B(n14670), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XNOR2_X1 U18314 ( .A(n9814), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15156) );
  OAI21_X1 U18315 ( .B1(n17723), .B2(n15175), .A(n14672), .ZN(n14673) );
  AOI21_X1 U18316 ( .B1(n15156), .B2(n17714), .A(n14673), .ZN(n14675) );
  OAI21_X1 U18317 ( .B1(n17116), .B2(n14677), .A(n14676), .ZN(P2_U2984) );
  INV_X1 U18318 ( .A(n14678), .ZN(n14706) );
  AND2_X1 U18319 ( .A1(n14680), .A2(n14679), .ZN(n14681) );
  NAND2_X1 U18320 ( .A1(n14682), .A2(n14681), .ZN(n15194) );
  NAND2_X1 U18321 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n17708), .ZN(n17616) );
  NAND2_X1 U18322 ( .A1(n14683), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14684) );
  MUX2_X1 U18323 ( .A(n17616), .B(n14684), .S(n21654), .Z(n14685) );
  NAND2_X1 U18324 ( .A1(n14685), .A2(n17669), .ZN(n14686) );
  INV_X1 U18325 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15498) );
  NOR2_X1 U18326 ( .A1(n13040), .A2(n15498), .ZN(n14700) );
  AND2_X1 U18327 ( .A1(n21434), .A2(n21428), .ZN(n17614) );
  INV_X1 U18328 ( .A(n17614), .ZN(n14688) );
  NAND2_X1 U18329 ( .A1(n14700), .A2(n14688), .ZN(n14689) );
  OAI21_X1 U18330 ( .B1(n14691), .B2(n14690), .A(n17614), .ZN(n14698) );
  INV_X1 U18331 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21665) );
  INV_X1 U18332 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21372) );
  NAND3_X1 U18333 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n21164) );
  NOR2_X1 U18334 ( .A1(n21363), .A2(n21164), .ZN(n15453) );
  NOR2_X1 U18335 ( .A1(n21584), .A2(n21367), .ZN(n21128) );
  AND3_X1 U18336 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n21128), .ZN(n15454) );
  NAND2_X1 U18337 ( .A1(n15453), .A2(n15454), .ZN(n21111) );
  NOR2_X1 U18338 ( .A1(n21372), .A2(n21111), .ZN(n17639) );
  NAND2_X1 U18339 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n17639), .ZN(n17629) );
  NOR2_X1 U18340 ( .A1(n21665), .A2(n17629), .ZN(n15441) );
  AND2_X1 U18341 ( .A1(n15441), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U18342 ( .A1(n17640), .A2(n14692), .ZN(n15432) );
  NAND2_X1 U18343 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14693) );
  INV_X1 U18344 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21382) );
  INV_X1 U18345 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21381) );
  NAND3_X1 U18346 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14694) );
  NAND2_X1 U18347 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15294) );
  INV_X1 U18348 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15712) );
  NOR2_X1 U18349 ( .A1(n15294), .A2(n15712), .ZN(n14695) );
  NAND2_X1 U18350 ( .A1(n15293), .A2(n14695), .ZN(n15281) );
  NAND3_X1 U18351 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n15244) );
  INV_X1 U18352 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21399) );
  NOR3_X1 U18353 ( .A1(n15281), .A2(n15244), .A3(n21399), .ZN(n15228) );
  NAND2_X1 U18354 ( .A1(n15228), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U18355 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14696) );
  NOR3_X1 U18356 ( .A1(n15219), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14696), 
        .ZN(n14704) );
  INV_X1 U18357 ( .A(n17628), .ZN(n15471) );
  NAND2_X1 U18358 ( .A1(n15471), .A2(n14692), .ZN(n15428) );
  NOR2_X1 U18359 ( .A1(n15428), .A2(n14693), .ZN(n15376) );
  NAND4_X1 U18360 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n15376), .ZN(n15341) );
  NOR2_X1 U18361 ( .A1(n14694), .A2(n15341), .ZN(n15305) );
  NAND2_X1 U18362 ( .A1(n15305), .A2(n14695), .ZN(n15268) );
  NOR2_X1 U18363 ( .A1(n15244), .A2(n15268), .ZN(n15242) );
  NAND3_X1 U18364 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n15242), .ZN(n15217) );
  NAND2_X1 U18365 ( .A1(n21173), .A2(n15471), .ZN(n15429) );
  OAI21_X1 U18366 ( .B1(n15217), .B2(n14696), .A(n15429), .ZN(n15206) );
  NAND2_X1 U18367 ( .A1(n14698), .A2(n14697), .ZN(n14699) );
  OR2_X1 U18368 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  AOI22_X1 U18369 ( .A1(n21182), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21174), .ZN(n14702) );
  OAI21_X1 U18370 ( .B1(n15206), .B2(n21409), .A(n14702), .ZN(n14703) );
  AOI211_X1 U18371 ( .C1(n15497), .C2(n21176), .A(n14704), .B(n14703), .ZN(
        n14705) );
  OAI21_X1 U18372 ( .B1(n14706), .B2(n21137), .A(n14705), .ZN(P1_U2809) );
  NAND2_X1 U18373 ( .A1(n20358), .A2(n14707), .ZN(n14708) );
  AND2_X1 U18374 ( .A1(n17246), .A2(n9836), .ZN(n14710) );
  AOI21_X1 U18375 ( .B1(n14714), .B2(n14501), .A(n9758), .ZN(n16856) );
  NAND2_X1 U18376 ( .A1(n16856), .A2(n20355), .ZN(n14715) );
  NAND2_X1 U18377 ( .A1(n20263), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16966) );
  OAI211_X1 U18378 ( .C1(n16964), .C2(n17352), .A(n14715), .B(n16966), .ZN(
        n14717) );
  INV_X1 U18379 ( .A(n16738), .ZN(n14725) );
  OR2_X1 U18380 ( .A1(n15135), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14721) );
  NAND2_X1 U18381 ( .A1(n14720), .A2(n14721), .ZN(n16547) );
  AOI21_X1 U18382 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14722), .ZN(n14723) );
  OAI21_X1 U18383 ( .B1(n16547), .B2(n17112), .A(n14723), .ZN(n14724) );
  AOI21_X1 U18384 ( .B1(n14725), .B2(n17716), .A(n14724), .ZN(n14728) );
  NAND3_X1 U18385 ( .A1(n13447), .A2(n17718), .A3(n14726), .ZN(n14727) );
  OAI211_X1 U18386 ( .C1(n14729), .C2(n17136), .A(n14728), .B(n14727), .ZN(
        P2_U2993) );
  AOI22_X1 U18387 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14733) );
  AOI22_X1 U18388 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U18389 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14731) );
  AOI22_X1 U18390 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14730) );
  NAND4_X1 U18391 ( .A1(n14733), .A2(n14732), .A3(n14731), .A4(n14730), .ZN(
        n14739) );
  AOI22_X1 U18392 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14737) );
  AOI22_X1 U18393 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U18394 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14735) );
  AOI22_X1 U18395 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14734) );
  NAND4_X1 U18396 ( .A1(n14737), .A2(n14736), .A3(n14735), .A4(n14734), .ZN(
        n14738) );
  AOI22_X1 U18397 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14803), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U18398 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14743) );
  AOI22_X1 U18399 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14742) );
  AOI22_X1 U18400 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12273), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14741) );
  NAND4_X1 U18401 ( .A1(n14744), .A2(n14743), .A3(n14742), .A4(n14741), .ZN(
        n14750) );
  AOI22_X1 U18402 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14748) );
  AOI22_X1 U18403 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12245), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U18404 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12231), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U18405 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12234), .B1(
        n12233), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14745) );
  NAND4_X1 U18406 ( .A1(n14748), .A2(n14747), .A3(n14746), .A4(n14745), .ZN(
        n14749) );
  NOR2_X1 U18407 ( .A1(n14750), .A2(n14749), .ZN(n16748) );
  INV_X1 U18408 ( .A(n16748), .ZN(n14751) );
  AOI22_X1 U18409 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U18410 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14754) );
  AOI22_X1 U18411 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14753) );
  AOI22_X1 U18412 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14752) );
  NAND4_X1 U18413 ( .A1(n14755), .A2(n14754), .A3(n14753), .A4(n14752), .ZN(
        n14761) );
  AOI22_X1 U18414 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14759) );
  AOI22_X1 U18415 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U18416 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14757) );
  AOI22_X1 U18417 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14756) );
  NAND4_X1 U18418 ( .A1(n14759), .A2(n14758), .A3(n14757), .A4(n14756), .ZN(
        n14760) );
  NOR2_X1 U18419 ( .A1(n14761), .A2(n14760), .ZN(n16740) );
  AOI22_X1 U18420 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U18421 ( .A1(n14802), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14764) );
  AOI22_X1 U18422 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U18423 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14762) );
  NAND4_X1 U18424 ( .A1(n14765), .A2(n14764), .A3(n14763), .A4(n14762), .ZN(
        n14771) );
  AOI22_X1 U18425 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14769) );
  AOI22_X1 U18426 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14768) );
  AOI22_X1 U18427 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14767) );
  AOI22_X1 U18428 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14766) );
  NAND4_X1 U18429 ( .A1(n14769), .A2(n14768), .A3(n14767), .A4(n14766), .ZN(
        n14770) );
  OR2_X1 U18430 ( .A1(n14771), .A2(n14770), .ZN(n16735) );
  AOI22_X1 U18431 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14776) );
  AOI22_X1 U18432 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14775) );
  AOI22_X1 U18433 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14774) );
  AOI22_X1 U18434 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14773) );
  NAND4_X1 U18435 ( .A1(n14776), .A2(n14775), .A3(n14774), .A4(n14773), .ZN(
        n14782) );
  AOI22_X1 U18436 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14780) );
  AOI22_X1 U18437 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U18438 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U18439 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14777) );
  NAND4_X1 U18440 ( .A1(n14780), .A2(n14779), .A3(n14778), .A4(n14777), .ZN(
        n14781) );
  NOR2_X1 U18441 ( .A1(n14782), .A2(n14781), .ZN(n16730) );
  AOI22_X1 U18442 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14952), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14793) );
  AND2_X1 U18443 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14785) );
  OR2_X1 U18444 ( .A1(n14785), .A2(n14784), .ZN(n14955) );
  INV_X1 U18445 ( .A(n14955), .ZN(n14931) );
  NAND2_X1 U18446 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14787) );
  NAND2_X1 U18447 ( .A1(n12001), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14786) );
  AND3_X1 U18448 ( .A1(n14931), .A2(n14787), .A3(n14786), .ZN(n14792) );
  AOI22_X1 U18449 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14791) );
  AOI22_X1 U18450 ( .A1(n14947), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14790) );
  NAND4_X1 U18451 ( .A1(n14793), .A2(n14792), .A3(n14791), .A4(n14790), .ZN(
        n14801) );
  AOI22_X1 U18452 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U18453 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14798) );
  AOI22_X1 U18454 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U18455 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14795) );
  NAND2_X1 U18456 ( .A1(n12001), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14794) );
  AND3_X1 U18457 ( .A1(n14795), .A2(n14794), .A3(n14955), .ZN(n14796) );
  NAND4_X1 U18458 ( .A1(n14799), .A2(n14798), .A3(n14797), .A4(n14796), .ZN(
        n14800) );
  NAND2_X1 U18459 ( .A1(n21078), .A2(n14836), .ZN(n14816) );
  AOI22_X1 U18460 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14802), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U18461 ( .A1(n12349), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12240), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U18462 ( .A1(n14803), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14807) );
  AOI22_X1 U18463 ( .A1(n12278), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14804), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14806) );
  NAND4_X1 U18464 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(
        n14815) );
  AOI22_X1 U18465 ( .A1(n12273), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12252), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U18466 ( .A1(n12257), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14812) );
  AOI22_X1 U18467 ( .A1(n12231), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12232), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U18468 ( .A1(n12233), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12234), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14810) );
  NAND4_X1 U18469 ( .A1(n14813), .A2(n14812), .A3(n14811), .A4(n14810), .ZN(
        n14814) );
  OR2_X1 U18470 ( .A1(n14815), .A2(n14814), .ZN(n14819) );
  XNOR2_X1 U18471 ( .A(n14816), .B(n14819), .ZN(n14839) );
  XNOR2_X1 U18472 ( .A(n14817), .B(n14839), .ZN(n16727) );
  NAND2_X1 U18473 ( .A1(n14904), .A2(n14836), .ZN(n16726) );
  NAND2_X1 U18474 ( .A1(n14819), .A2(n14836), .ZN(n14841) );
  AOI22_X1 U18475 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U18476 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U18477 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U18478 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14821) );
  NAND2_X1 U18479 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14820) );
  AND3_X1 U18480 ( .A1(n14821), .A2(n14820), .A3(n14955), .ZN(n14822) );
  NAND4_X1 U18481 ( .A1(n14825), .A2(n14824), .A3(n14823), .A4(n14822), .ZN(
        n14833) );
  AOI22_X1 U18482 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14831) );
  NAND2_X1 U18483 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14827) );
  NAND2_X1 U18484 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14826) );
  AND3_X1 U18485 ( .A1(n14931), .A2(n14827), .A3(n14826), .ZN(n14830) );
  AOI22_X1 U18486 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14829) );
  AOI22_X1 U18487 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14828) );
  NAND4_X1 U18488 ( .A1(n14831), .A2(n14830), .A3(n14829), .A4(n14828), .ZN(
        n14832) );
  NAND2_X1 U18489 ( .A1(n14833), .A2(n14832), .ZN(n14840) );
  XOR2_X1 U18490 ( .A(n14841), .B(n14840), .Z(n14834) );
  NAND2_X1 U18491 ( .A1(n14834), .A2(n14876), .ZN(n16719) );
  INV_X1 U18492 ( .A(n14840), .ZN(n14835) );
  NAND2_X1 U18493 ( .A1(n14904), .A2(n14835), .ZN(n16722) );
  INV_X1 U18494 ( .A(n14836), .ZN(n14837) );
  NOR2_X1 U18495 ( .A1(n16722), .A2(n14837), .ZN(n14838) );
  NOR2_X1 U18496 ( .A1(n14841), .A2(n14840), .ZN(n14856) );
  AOI22_X1 U18497 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14948), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14847) );
  AOI22_X1 U18498 ( .A1(n14947), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U18499 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14845) );
  INV_X1 U18500 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20491) );
  NAND2_X1 U18501 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14843) );
  NAND2_X1 U18502 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14842) );
  AND3_X1 U18503 ( .A1(n14843), .A2(n14842), .A3(n14955), .ZN(n14844) );
  NAND4_X1 U18504 ( .A1(n14847), .A2(n14846), .A3(n14845), .A4(n14844), .ZN(
        n14855) );
  AOI22_X1 U18505 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14952), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14853) );
  INV_X1 U18506 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U18507 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U18508 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14849) );
  NAND2_X1 U18509 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14848) );
  AND3_X1 U18510 ( .A1(n14931), .A2(n14849), .A3(n14848), .ZN(n14851) );
  AOI22_X1 U18511 ( .A1(n9749), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14850) );
  NAND4_X1 U18512 ( .A1(n14853), .A2(n14852), .A3(n14851), .A4(n14850), .ZN(
        n14854) );
  NAND2_X1 U18513 ( .A1(n14856), .A2(n14857), .ZN(n14896) );
  OAI211_X1 U18514 ( .C1(n14856), .C2(n14857), .A(n14876), .B(n14896), .ZN(
        n14874) );
  INV_X1 U18515 ( .A(n14857), .ZN(n14858) );
  NOR2_X1 U18516 ( .A1(n21078), .A2(n14858), .ZN(n16716) );
  AOI22_X1 U18517 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U18518 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14860) );
  NAND2_X1 U18519 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14859) );
  AND3_X1 U18520 ( .A1(n14931), .A2(n14860), .A3(n14859), .ZN(n14863) );
  AOI22_X1 U18521 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14862) );
  AOI22_X1 U18522 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14861) );
  NAND4_X1 U18523 ( .A1(n14864), .A2(n14863), .A3(n14862), .A4(n14861), .ZN(
        n14872) );
  AOI22_X1 U18524 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U18525 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U18526 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U18527 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14866) );
  NAND2_X1 U18528 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14865) );
  AND3_X1 U18529 ( .A1(n14866), .A2(n14865), .A3(n14955), .ZN(n14867) );
  NAND4_X1 U18530 ( .A1(n14870), .A2(n14869), .A3(n14868), .A4(n14867), .ZN(
        n14871) );
  NAND2_X1 U18531 ( .A1(n16706), .A2(n14873), .ZN(n14881) );
  INV_X1 U18532 ( .A(n16707), .ZN(n14879) );
  INV_X1 U18533 ( .A(n14875), .ZN(n16708) );
  XOR2_X1 U18534 ( .A(n14896), .B(n16708), .Z(n14877) );
  NAND2_X1 U18535 ( .A1(n14877), .A2(n14876), .ZN(n16710) );
  INV_X1 U18536 ( .A(n16710), .ZN(n14878) );
  NAND2_X1 U18537 ( .A1(n14881), .A2(n14880), .ZN(n14900) );
  AOI22_X1 U18538 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14887) );
  AOI22_X1 U18539 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U18540 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14885) );
  NAND2_X1 U18541 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14883) );
  NAND2_X1 U18542 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14882) );
  AND3_X1 U18543 ( .A1(n14883), .A2(n14882), .A3(n14955), .ZN(n14884) );
  NAND4_X1 U18544 ( .A1(n14887), .A2(n14886), .A3(n14885), .A4(n14884), .ZN(
        n14895) );
  AOI22_X1 U18545 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14893) );
  NAND2_X1 U18546 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14889) );
  NAND2_X1 U18547 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14888) );
  AND3_X1 U18548 ( .A1(n14931), .A2(n14889), .A3(n14888), .ZN(n14892) );
  AOI22_X1 U18549 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14891) );
  AOI22_X1 U18550 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14890) );
  NAND4_X1 U18551 ( .A1(n14893), .A2(n14892), .A3(n14891), .A4(n14890), .ZN(
        n14894) );
  NAND2_X1 U18552 ( .A1(n14895), .A2(n14894), .ZN(n14902) );
  OR2_X1 U18553 ( .A1(n14896), .A2(n16708), .ZN(n14898) );
  NOR2_X1 U18554 ( .A1(n14898), .A2(n14902), .ZN(n14921) );
  AOI211_X1 U18555 ( .C1(n14902), .C2(n14898), .A(n14897), .B(n14921), .ZN(
        n14899) );
  INV_X1 U18556 ( .A(n14902), .ZN(n14903) );
  NAND2_X1 U18557 ( .A1(n14904), .A2(n14903), .ZN(n16702) );
  INV_X1 U18558 ( .A(n14905), .ZN(n14920) );
  AOI22_X1 U18559 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U18560 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14907) );
  NAND2_X1 U18561 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14906) );
  AND3_X1 U18562 ( .A1(n14931), .A2(n14907), .A3(n14906), .ZN(n14910) );
  AOI22_X1 U18563 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14909) );
  AOI22_X1 U18564 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14908) );
  NAND4_X1 U18565 ( .A1(n14911), .A2(n14910), .A3(n14909), .A4(n14908), .ZN(
        n14919) );
  AOI22_X1 U18566 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14917) );
  AOI22_X1 U18567 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14916) );
  AOI22_X1 U18568 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U18569 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14913) );
  NAND2_X1 U18570 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14912) );
  AND3_X1 U18571 ( .A1(n14913), .A2(n14912), .A3(n14955), .ZN(n14914) );
  NAND4_X1 U18572 ( .A1(n14917), .A2(n14916), .A3(n14915), .A4(n14914), .ZN(
        n14918) );
  INV_X1 U18573 ( .A(n14921), .ZN(n16696) );
  NAND2_X1 U18574 ( .A1(n21078), .A2(n16697), .ZN(n14922) );
  NOR2_X1 U18575 ( .A1(n16696), .A2(n14922), .ZN(n14939) );
  AOI22_X1 U18576 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14948), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14928) );
  AOI22_X1 U18577 ( .A1(n14947), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U18578 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U18579 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14924) );
  NAND2_X1 U18580 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14923) );
  AND3_X1 U18581 ( .A1(n14924), .A2(n14923), .A3(n14955), .ZN(n14925) );
  NAND4_X1 U18582 ( .A1(n14928), .A2(n14927), .A3(n14926), .A4(n14925), .ZN(
        n14937) );
  AOI22_X1 U18583 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14935) );
  NAND2_X1 U18584 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14930) );
  NAND2_X1 U18585 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14929) );
  AND3_X1 U18586 ( .A1(n14931), .A2(n14930), .A3(n14929), .ZN(n14934) );
  AOI22_X1 U18587 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14933) );
  INV_X1 U18588 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U18589 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14932) );
  NAND4_X1 U18590 ( .A1(n14935), .A2(n14934), .A3(n14933), .A4(n14932), .ZN(
        n14936) );
  AND2_X1 U18591 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  NAND2_X1 U18592 ( .A1(n14939), .A2(n14938), .ZN(n14940) );
  OAI21_X1 U18593 ( .B1(n14939), .B2(n14938), .A(n14940), .ZN(n16691) );
  AOI22_X1 U18594 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14942) );
  AOI22_X1 U18595 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14941) );
  NAND2_X1 U18596 ( .A1(n14942), .A2(n14941), .ZN(n14962) );
  AOI22_X1 U18597 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14789), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14944) );
  AOI21_X1 U18598 ( .B1(n14953), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n14955), .ZN(n14943) );
  OAI211_X1 U18599 ( .C1(n14946), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        n14961) );
  AOI22_X1 U18600 ( .A1(n14948), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14947), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U18601 ( .A1(n14949), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9727), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14950) );
  NAND2_X1 U18602 ( .A1(n14951), .A2(n14950), .ZN(n14960) );
  AOI22_X1 U18603 ( .A1(n14952), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9749), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U18604 ( .A1(n14953), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14957) );
  NAND2_X1 U18605 ( .A1(n14954), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14956) );
  NAND4_X1 U18606 ( .A1(n14958), .A2(n14957), .A3(n14956), .A4(n14955), .ZN(
        n14959) );
  OAI22_X1 U18607 ( .A1(n14962), .A2(n14961), .B1(n14960), .B2(n14959), .ZN(
        n14963) );
  INV_X1 U18608 ( .A(n14964), .ZN(n15181) );
  INV_X1 U18609 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14968) );
  NAND2_X1 U18610 ( .A1(n14507), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U18611 ( .A1(n16858), .A2(n14965), .B1(n20306), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14966) );
  OAI211_X1 U18612 ( .C1(n16859), .C2(n14968), .A(n14967), .B(n14966), .ZN(
        n14969) );
  AOI21_X1 U18613 ( .B1(n15181), .B2(n20307), .A(n14969), .ZN(n14970) );
  OAI21_X1 U18614 ( .B1(n14973), .B2(n20311), .A(n14970), .ZN(P2_U2889) );
  MUX2_X1 U18615 ( .A(n14971), .B(n15182), .S(n20291), .Z(n14972) );
  OAI21_X1 U18616 ( .B1(n14973), .B2(n20283), .A(n14972), .ZN(P2_U2857) );
  NOR2_X1 U18617 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21335), .ZN(n15016) );
  NAND2_X1 U18618 ( .A1(n14975), .A2(n14974), .ZN(n14977) );
  OR2_X1 U18619 ( .A1(n14977), .A2(n14976), .ZN(n14978) );
  NOR2_X1 U18620 ( .A1(n14979), .A2(n14978), .ZN(n14980) );
  NAND3_X1 U18621 ( .A1(n14981), .A2(n14980), .A3(n15013), .ZN(n16097) );
  INV_X1 U18622 ( .A(n16097), .ZN(n15006) );
  OR2_X1 U18623 ( .A1(n16291), .A2(n15006), .ZN(n14991) );
  XNOR2_X1 U18624 ( .A(n16091), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16108) );
  INV_X1 U18625 ( .A(n16108), .ZN(n14982) );
  NAND2_X1 U18626 ( .A1(n10878), .A2(n14982), .ZN(n14988) );
  XNOR2_X1 U18627 ( .A(n14983), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14986) );
  NAND2_X1 U18628 ( .A1(n14985), .A2(n14984), .ZN(n14999) );
  AOI22_X1 U18629 ( .A1(n16090), .A2(n14986), .B1(n14999), .B2(n16108), .ZN(
        n14987) );
  OAI21_X1 U18630 ( .B1(n16097), .B2(n14988), .A(n14987), .ZN(n14989) );
  INV_X1 U18631 ( .A(n14989), .ZN(n14990) );
  AND2_X1 U18632 ( .A1(n14991), .A2(n14990), .ZN(n16105) );
  NAND2_X1 U18633 ( .A1(n16105), .A2(n15012), .ZN(n14994) );
  INV_X1 U18634 ( .A(n15012), .ZN(n17592) );
  NAND2_X1 U18635 ( .A1(n17592), .A2(n14992), .ZN(n14993) );
  AOI22_X1 U18636 ( .A1(n15016), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17596), .B2(n21335), .ZN(n15010) );
  NAND2_X1 U18637 ( .A1(n15024), .A2(n16097), .ZN(n15008) );
  NAND2_X1 U18638 ( .A1(n16091), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14995) );
  NAND2_X1 U18639 ( .A1(n14995), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14996) );
  NAND2_X1 U18640 ( .A1(n10723), .A2(n14996), .ZN(n16111) );
  AND2_X1 U18641 ( .A1(n10878), .A2(n16111), .ZN(n15005) );
  XNOR2_X1 U18642 ( .A(n14997), .B(n10695), .ZN(n14998) );
  NAND2_X1 U18643 ( .A1(n16090), .A2(n14998), .ZN(n15003) );
  OAI21_X1 U18644 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(n15002) );
  NAND2_X1 U18645 ( .A1(n15003), .A2(n15002), .ZN(n15004) );
  AOI21_X1 U18646 ( .B1(n15006), .B2(n15005), .A(n15004), .ZN(n15007) );
  NAND2_X1 U18647 ( .A1(n15008), .A2(n15007), .ZN(n16110) );
  MUX2_X1 U18648 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16110), .S(
        n15012), .Z(n17599) );
  AOI22_X1 U18649 ( .A1(n15016), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21335), .B2(n17599), .ZN(n15009) );
  NOR2_X1 U18650 ( .A1(n15010), .A2(n15009), .ZN(n17608) );
  INV_X1 U18651 ( .A(n15011), .ZN(n16093) );
  NAND2_X1 U18652 ( .A1(n17608), .A2(n16093), .ZN(n16075) );
  OAI21_X1 U18653 ( .B1(n15014), .B2(n15013), .A(n15012), .ZN(n15018) );
  AOI21_X1 U18654 ( .B1(n17592), .B2(n15015), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15017) );
  AOI22_X1 U18655 ( .A1(n15018), .A2(n15017), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15016), .ZN(n17610) );
  NAND3_X1 U18656 ( .A1(n16075), .A2(n17610), .A3(n21095), .ZN(n15021) );
  INV_X1 U18657 ( .A(n17709), .ZN(n15020) );
  AOI21_X1 U18658 ( .B1(n21280), .B2(n15023), .A(n16385), .ZN(n16387) );
  INV_X1 U18659 ( .A(n15024), .ZN(n21179) );
  NAND2_X1 U18660 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n17711), .ZN(n16076) );
  INV_X1 U18661 ( .A(n16076), .ZN(n16088) );
  NOR2_X1 U18662 ( .A1(n21179), .A2(n16088), .ZN(n15026) );
  AOI211_X1 U18663 ( .C1(n16387), .C2(n14024), .A(n15026), .B(n15025), .ZN(
        n15028) );
  NAND2_X1 U18664 ( .A1(n21258), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15027) );
  OAI21_X1 U18665 ( .B1(n21258), .B2(n15028), .A(n15027), .ZN(P1_U3475) );
  NAND3_X1 U18666 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15029), .A3(
        n16294), .ZN(n15052) );
  NOR2_X1 U18667 ( .A1(n21271), .A2(n15052), .ZN(n21265) );
  INV_X1 U18668 ( .A(n21265), .ZN(n15048) );
  OAI22_X1 U18669 ( .A1(n14687), .A2(n15052), .B1(n16385), .B2(n15048), .ZN(
        n15030) );
  AOI21_X1 U18670 ( .B1(n15053), .B2(n15031), .A(n15030), .ZN(n21259) );
  OAI22_X1 U18671 ( .A1(n16422), .A2(n21259), .B1(n16327), .B2(n15048), .ZN(
        n15032) );
  AOI21_X1 U18672 ( .B1(n21266), .B2(n21320), .A(n15032), .ZN(n15038) );
  INV_X1 U18673 ( .A(n14024), .ZN(n15034) );
  NOR2_X1 U18674 ( .A1(n15034), .A2(n15033), .ZN(n15036) );
  INV_X1 U18675 ( .A(n15052), .ZN(n15035) );
  NAND2_X1 U18676 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15037) );
  OAI211_X1 U18677 ( .C1(n21323), .C2(n21270), .A(n15038), .B(n15037), .ZN(
        P1_U3111) );
  OAI22_X1 U18678 ( .A1(n16412), .A2(n21259), .B1(n16317), .B2(n15048), .ZN(
        n15039) );
  AOI21_X1 U18679 ( .B1(n21266), .B2(n21308), .A(n15039), .ZN(n15041) );
  NAND2_X1 U18680 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n15040) );
  OAI211_X1 U18681 ( .C1(n21311), .C2(n21270), .A(n15041), .B(n15040), .ZN(
        P1_U3109) );
  OAI22_X1 U18682 ( .A1(n16407), .A2(n21259), .B1(n16312), .B2(n15048), .ZN(
        n15042) );
  AOI21_X1 U18683 ( .B1(n21266), .B2(n21302), .A(n15042), .ZN(n15044) );
  NAND2_X1 U18684 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15043) );
  OAI211_X1 U18685 ( .C1(n21305), .C2(n21270), .A(n15044), .B(n15043), .ZN(
        P1_U3108) );
  OAI22_X1 U18686 ( .A1(n16399), .A2(n21259), .B1(n16304), .B2(n15048), .ZN(
        n15045) );
  AOI21_X1 U18687 ( .B1(n21266), .B2(n21290), .A(n15045), .ZN(n15047) );
  NAND2_X1 U18688 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n15046) );
  OAI211_X1 U18689 ( .C1(n21293), .C2(n21270), .A(n15047), .B(n15046), .ZN(
        P1_U3106) );
  OAI22_X1 U18690 ( .A1(n16394), .A2(n21259), .B1(n16295), .B2(n15048), .ZN(
        n15049) );
  AOI21_X1 U18691 ( .B1(n21266), .B2(n21284), .A(n15049), .ZN(n15051) );
  NAND2_X1 U18692 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15050) );
  OAI211_X1 U18693 ( .C1(n21287), .C2(n21270), .A(n15051), .B(n15050), .ZN(
        P1_U3105) );
  NOR2_X1 U18694 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15052), .ZN(
        n15060) );
  AOI21_X1 U18695 ( .B1(n15053), .B2(n14436), .A(n15060), .ZN(n15058) );
  INV_X1 U18696 ( .A(n16121), .ZN(n15054) );
  NAND2_X1 U18697 ( .A1(n15054), .A2(n16164), .ZN(n16298) );
  INV_X1 U18698 ( .A(n16203), .ZN(n15055) );
  INV_X1 U18699 ( .A(n15060), .ZN(n15085) );
  INV_X1 U18700 ( .A(n21270), .ZN(n15056) );
  OAI21_X1 U18701 ( .B1(n15056), .B2(n15083), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15057) );
  NAND2_X1 U18702 ( .A1(n15058), .A2(n15057), .ZN(n15059) );
  OAI211_X1 U18703 ( .C1(n15060), .C2(n17711), .A(n16166), .B(n15059), .ZN(
        n15082) );
  AOI22_X1 U18704 ( .A1(n15083), .A2(n16335), .B1(
        P1_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n15082), .ZN(n15061) );
  OAI21_X1 U18705 ( .B1(n16333), .B2(n15085), .A(n15061), .ZN(n15062) );
  AOI21_X1 U18706 ( .B1(n21325), .B2(n15087), .A(n15062), .ZN(n15063) );
  OAI21_X1 U18707 ( .B1(n16426), .B2(n21270), .A(n15063), .ZN(P1_U3104) );
  AOI22_X1 U18708 ( .A1(n15083), .A2(n16329), .B1(
        P1_INSTQUEUE_REG_8__6__SCAN_IN), .B2(n15082), .ZN(n15064) );
  OAI21_X1 U18709 ( .B1(n16327), .B2(n15085), .A(n15064), .ZN(n15065) );
  AOI21_X1 U18710 ( .B1(n21318), .B2(n15087), .A(n15065), .ZN(n15066) );
  OAI21_X1 U18711 ( .B1(n16418), .B2(n21270), .A(n15066), .ZN(P1_U3103) );
  AOI22_X1 U18712 ( .A1(n15083), .A2(n16324), .B1(
        P1_INSTQUEUE_REG_8__5__SCAN_IN), .B2(n15082), .ZN(n15067) );
  OAI21_X1 U18713 ( .B1(n16322), .B2(n15085), .A(n15067), .ZN(n15068) );
  AOI21_X1 U18714 ( .B1(n21312), .B2(n15087), .A(n15068), .ZN(n15069) );
  OAI21_X1 U18715 ( .B1(n16413), .B2(n21270), .A(n15069), .ZN(P1_U3102) );
  AOI22_X1 U18716 ( .A1(n15083), .A2(n16319), .B1(
        P1_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n15082), .ZN(n15070) );
  OAI21_X1 U18717 ( .B1(n16317), .B2(n15085), .A(n15070), .ZN(n15071) );
  AOI21_X1 U18718 ( .B1(n21306), .B2(n15087), .A(n15071), .ZN(n15072) );
  OAI21_X1 U18719 ( .B1(n16408), .B2(n21270), .A(n15072), .ZN(P1_U3101) );
  AOI22_X1 U18720 ( .A1(n15083), .A2(n16314), .B1(
        P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n15082), .ZN(n15073) );
  OAI21_X1 U18721 ( .B1(n16312), .B2(n15085), .A(n15073), .ZN(n15074) );
  AOI21_X1 U18722 ( .B1(n21300), .B2(n15087), .A(n15074), .ZN(n15075) );
  OAI21_X1 U18723 ( .B1(n16403), .B2(n21270), .A(n15075), .ZN(P1_U3100) );
  AOI22_X1 U18724 ( .A1(n15083), .A2(n21752), .B1(
        P1_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n15082), .ZN(n15076) );
  OAI21_X1 U18725 ( .B1(n21748), .B2(n15085), .A(n15076), .ZN(n15077) );
  AOI21_X1 U18726 ( .B1(n21294), .B2(n15087), .A(n15077), .ZN(n15078) );
  OAI21_X1 U18727 ( .B1(n21758), .B2(n21270), .A(n15078), .ZN(P1_U3099) );
  AOI22_X1 U18728 ( .A1(n15083), .A2(n16306), .B1(
        P1_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n15082), .ZN(n15079) );
  OAI21_X1 U18729 ( .B1(n16304), .B2(n15085), .A(n15079), .ZN(n15080) );
  AOI21_X1 U18730 ( .B1(n21288), .B2(n15087), .A(n15080), .ZN(n15081) );
  OAI21_X1 U18731 ( .B1(n16395), .B2(n21270), .A(n15081), .ZN(P1_U3098) );
  AOI22_X1 U18732 ( .A1(n15083), .A2(n16297), .B1(
        P1_INSTQUEUE_REG_8__0__SCAN_IN), .B2(n15082), .ZN(n15084) );
  OAI21_X1 U18733 ( .B1(n16295), .B2(n15085), .A(n15084), .ZN(n15086) );
  AOI21_X1 U18734 ( .B1(n21278), .B2(n15087), .A(n15086), .ZN(n15088) );
  OAI21_X1 U18735 ( .B1(n16390), .B2(n21270), .A(n15088), .ZN(P1_U3097) );
  NOR2_X1 U18736 ( .A1(n16094), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15089) );
  INV_X1 U18737 ( .A(n15092), .ZN(n16114) );
  INV_X1 U18738 ( .A(n16112), .ZN(n16102) );
  AOI22_X1 U18739 ( .A1(n16102), .A2(n15095), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n15090), .ZN(n15091) );
  OAI21_X1 U18740 ( .B1(n17590), .B2(n16114), .A(n15091), .ZN(n15093) );
  AND2_X1 U18741 ( .A1(n16090), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17588) );
  AOI22_X1 U18742 ( .A1(n15093), .A2(n16116), .B1(n15092), .B2(n17588), .ZN(
        n15094) );
  OAI21_X1 U18743 ( .B1(n15095), .B2(n16116), .A(n15094), .ZN(P1_U3474) );
  NAND2_X1 U18744 ( .A1(n21073), .A2(n20814), .ZN(n15166) );
  MUX2_X2 U18745 ( .A(n15097), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15144) );
  MUX2_X1 U18746 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n17407) );
  NOR2_X1 U18747 ( .A1(n17407), .A2(n16665), .ZN(n16667) );
  OAI21_X1 U18749 ( .B1(n15099), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15100), .ZN(n17124) );
  NAND2_X1 U18750 ( .A1(n16637), .A2(n17124), .ZN(n20271) );
  AND2_X1 U18751 ( .A1(n15100), .A2(n20259), .ZN(n15102) );
  OR2_X1 U18752 ( .A1(n15102), .A2(n15101), .ZN(n17111) );
  INV_X1 U18753 ( .A(n17111), .ZN(n20273) );
  NOR2_X1 U18754 ( .A1(n20271), .A2(n20273), .ZN(n20274) );
  OR2_X1 U18755 ( .A1(n15101), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15104) );
  NAND2_X1 U18756 ( .A1(n15103), .A2(n15104), .ZN(n17712) );
  NAND2_X1 U18757 ( .A1(n15103), .A2(n17094), .ZN(n15105) );
  AND2_X1 U18758 ( .A1(n15106), .A2(n15105), .ZN(n17096) );
  AND2_X1 U18759 ( .A1(n15106), .A2(n17089), .ZN(n15108) );
  NOR2_X1 U18760 ( .A1(n15107), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15109) );
  OR2_X1 U18761 ( .A1(n15111), .A2(n15109), .ZN(n17080) );
  INV_X1 U18762 ( .A(n17080), .ZN(n20226) );
  OR2_X1 U18763 ( .A1(n15111), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15112) );
  NAND2_X1 U18764 ( .A1(n15110), .A2(n15112), .ZN(n17062) );
  AND2_X1 U18765 ( .A1(n20227), .A2(n17062), .ZN(n20212) );
  NAND2_X1 U18766 ( .A1(n15110), .A2(n15114), .ZN(n15115) );
  NAND2_X1 U18767 ( .A1(n15116), .A2(n15115), .ZN(n20211) );
  NAND2_X1 U18768 ( .A1(n15116), .A2(n17036), .ZN(n15117) );
  AND2_X1 U18769 ( .A1(n15118), .A2(n15117), .ZN(n17038) );
  AND2_X1 U18770 ( .A1(n15118), .A2(n20202), .ZN(n15120) );
  OR2_X1 U18771 ( .A1(n15119), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15122) );
  NAND2_X1 U18772 ( .A1(n15121), .A2(n15122), .ZN(n17012) );
  INV_X1 U18773 ( .A(n15123), .ZN(n15126) );
  NAND2_X1 U18774 ( .A1(n15121), .A2(n20187), .ZN(n15124) );
  NAND2_X1 U18775 ( .A1(n15126), .A2(n15124), .ZN(n20182) );
  NAND2_X1 U18776 ( .A1(n20180), .A2(n20182), .ZN(n16578) );
  AND2_X1 U18777 ( .A1(n15126), .A2(n16988), .ZN(n15127) );
  NOR2_X1 U18778 ( .A1(n15125), .A2(n15127), .ZN(n16990) );
  NOR2_X1 U18780 ( .A1(n15125), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15128) );
  OR2_X1 U18781 ( .A1(n15129), .A2(n15128), .ZN(n16978) );
  INV_X1 U18782 ( .A(n16978), .ZN(n20165) );
  NOR2_X1 U18783 ( .A1(n20163), .A2(n20165), .ZN(n20166) );
  OR2_X1 U18784 ( .A1(n15129), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15130) );
  NAND2_X1 U18785 ( .A1(n13320), .A2(n15130), .ZN(n16967) );
  AND2_X1 U18786 ( .A1(n15131), .A2(n20137), .ZN(n15132) );
  NOR2_X1 U18787 ( .A1(n15133), .A2(n15132), .ZN(n20130) );
  NOR2_X1 U18788 ( .A1(n15133), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15134) );
  OR2_X1 U18789 ( .A1(n15135), .A2(n15134), .ZN(n16946) );
  INV_X1 U18790 ( .A(n16946), .ZN(n16556) );
  NAND2_X1 U18791 ( .A1(n16546), .A2(n16547), .ZN(n16535) );
  NAND2_X1 U18792 ( .A1(n15144), .A2(n16535), .ZN(n15138) );
  NAND2_X1 U18793 ( .A1(n14720), .A2(n15136), .ZN(n15137) );
  NAND2_X1 U18794 ( .A1(n15139), .A2(n15137), .ZN(n16939) );
  NAND2_X1 U18795 ( .A1(n15138), .A2(n16939), .ZN(n16515) );
  NAND2_X1 U18796 ( .A1(n16515), .A2(n15144), .ZN(n15141) );
  NAND2_X1 U18797 ( .A1(n15139), .A2(n16926), .ZN(n15140) );
  NAND2_X1 U18798 ( .A1(n15142), .A2(n15140), .ZN(n16516) );
  NAND2_X1 U18799 ( .A1(n15141), .A2(n16516), .ZN(n16502) );
  AND2_X1 U18800 ( .A1(n15142), .A2(n16916), .ZN(n15143) );
  NOR2_X1 U18801 ( .A1(n15146), .A2(n15143), .ZN(n16914) );
  INV_X1 U18802 ( .A(n15144), .ZN(n10238) );
  OR2_X1 U18803 ( .A1(n15146), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15147) );
  NAND2_X1 U18804 ( .A1(n15145), .A2(n15147), .ZN(n16909) );
  NAND2_X1 U18805 ( .A1(n15145), .A2(n16895), .ZN(n15148) );
  AND2_X1 U18806 ( .A1(n9813), .A2(n15148), .ZN(n16897) );
  AND2_X1 U18807 ( .A1(n9813), .A2(n16889), .ZN(n15150) );
  OR2_X1 U18808 ( .A1(n15150), .A2(n15149), .ZN(n16888) );
  NOR2_X1 U18809 ( .A1(n15149), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15151) );
  OR2_X1 U18810 ( .A1(n15152), .A2(n15151), .ZN(n16877) );
  INV_X1 U18811 ( .A(n16877), .ZN(n15153) );
  AOI21_X1 U18812 ( .B1(n16435), .B2(n15144), .A(n15156), .ZN(n15185) );
  INV_X1 U18813 ( .A(n15185), .ZN(n15161) );
  OR2_X2 U18814 ( .A1(n15155), .A2(n15154), .ZN(n20933) );
  AOI21_X1 U18815 ( .B1(n16435), .B2(n15156), .A(n20933), .ZN(n15157) );
  INV_X1 U18816 ( .A(n15157), .ZN(n15159) );
  INV_X1 U18817 ( .A(n16678), .ZN(n15158) );
  INV_X1 U18818 ( .A(n15162), .ZN(n15178) );
  NAND2_X1 U18819 ( .A1(n15166), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15163) );
  INV_X1 U18820 ( .A(n15164), .ZN(n15165) );
  AND2_X1 U18821 ( .A1(n20350), .A2(n15165), .ZN(n15186) );
  INV_X1 U18822 ( .A(n15186), .ZN(n15170) );
  INV_X1 U18823 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15167) );
  NAND3_X1 U18824 ( .A1(n15168), .A2(n15167), .A3(n15166), .ZN(n15169) );
  NAND2_X1 U18825 ( .A1(n20169), .A2(n20933), .ZN(n15171) );
  NOR2_X1 U18826 ( .A1(n15172), .A2(n15171), .ZN(n15173) );
  OAI22_X1 U18827 ( .A1(n20258), .A2(n15175), .B1(n15174), .B2(n20249), .ZN(
        n15176) );
  AOI21_X1 U18828 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n20245), .A(n15176), .ZN(
        n15177) );
  NAND2_X1 U18829 ( .A1(n16764), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U18830 ( .B1(n15183), .B2(n16764), .A(n15184), .ZN(P2_U2856) );
  NAND2_X1 U18831 ( .A1(n15144), .A2(n20276), .ZN(n16688) );
  AOI22_X1 U18832 ( .A1(P2_REIP_REG_31__SCAN_IN), .A2(n20264), .B1(n15186), 
        .B2(P2_EBX_REG_31__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U18833 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15187) );
  OAI211_X1 U18834 ( .C1(n15189), .C2(n20260), .A(n15188), .B(n15187), .ZN(
        n15190) );
  AOI21_X1 U18835 ( .B1(n15185), .B2(n16651), .A(n15190), .ZN(n15193) );
  NAND2_X1 U18836 ( .A1(n15191), .A2(n20235), .ZN(n15192) );
  OAI211_X1 U18837 ( .C1(n15183), .C2(n20251), .A(n15193), .B(n15192), .ZN(
        P2_U2824) );
  NAND2_X1 U18838 ( .A1(n21274), .A2(n21335), .ZN(n15339) );
  NAND2_X1 U18839 ( .A1(n15194), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n15195)
         );
  NAND3_X1 U18840 ( .A1(n15196), .A2(n15339), .A3(n15195), .ZN(P1_U2801) );
  INV_X1 U18841 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21710) );
  NAND2_X1 U18842 ( .A1(n21710), .A2(n15339), .ZN(n15199) );
  INV_X1 U18843 ( .A(n15197), .ZN(n15198) );
  MUX2_X1 U18844 ( .A(n15199), .B(n15198), .S(n21432), .Z(P1_U3487) );
  NAND2_X1 U18845 ( .A1(n15200), .A2(n21130), .ZN(n15211) );
  INV_X1 U18846 ( .A(n15201), .ZN(n15202) );
  INV_X1 U18847 ( .A(n15219), .ZN(n15204) );
  AOI21_X1 U18848 ( .B1(n15204), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n15207) );
  AOI22_X1 U18849 ( .A1(n21182), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21174), .ZN(n15205) );
  OAI21_X1 U18850 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15208) );
  AOI21_X1 U18851 ( .B1(n15209), .B2(n21185), .A(n15208), .ZN(n15210) );
  OAI211_X1 U18852 ( .C1(n21161), .C2(n15212), .A(n15211), .B(n15210), .ZN(
        P1_U2810) );
  OAI21_X1 U18853 ( .B1(n15224), .B2(n15213), .A(n13404), .ZN(n15657) );
  AND2_X1 U18854 ( .A1(n9773), .A2(n15214), .ZN(n15215) );
  INV_X1 U18855 ( .A(n15870), .ZN(n15221) );
  AND2_X1 U18856 ( .A1(n15429), .A2(n15217), .ZN(n15229) );
  OAI22_X1 U18857 ( .A1(n21122), .A2(n15500), .B1(n15218), .B2(n21149), .ZN(
        n15220) );
  OAI21_X1 U18858 ( .B1(n15657), .B2(n21137), .A(n15222), .ZN(P1_U2811) );
  AOI21_X1 U18859 ( .B1(n15225), .B2(n15223), .A(n15224), .ZN(n15671) );
  INV_X1 U18860 ( .A(n15671), .ZN(n15573) );
  OAI21_X1 U18861 ( .B1(n15226), .B2(n15227), .A(n9773), .ZN(n15501) );
  INV_X1 U18862 ( .A(n15501), .ZN(n15876) );
  NOR2_X1 U18863 ( .A1(n21170), .A2(n15669), .ZN(n15234) );
  INV_X1 U18864 ( .A(n15228), .ZN(n15232) );
  AOI22_X1 U18865 ( .A1(n21182), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21174), .ZN(n15231) );
  NAND2_X1 U18866 ( .A1(n15229), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15230) );
  OAI211_X1 U18867 ( .C1(n15232), .C2(P1_REIP_REG_28__SCAN_IN), .A(n15231), 
        .B(n15230), .ZN(n15233) );
  AOI211_X1 U18868 ( .C1(n15876), .C2(n21176), .A(n15234), .B(n15233), .ZN(
        n15235) );
  OAI21_X1 U18869 ( .B1(n15573), .B2(n21137), .A(n15235), .ZN(P1_U2812) );
  INV_X1 U18870 ( .A(n15223), .ZN(n15237) );
  AOI21_X1 U18871 ( .B1(n15238), .B2(n15236), .A(n15237), .ZN(n15682) );
  INV_X1 U18872 ( .A(n15682), .ZN(n15578) );
  INV_X1 U18873 ( .A(n15226), .ZN(n15240) );
  OAI21_X1 U18874 ( .B1(n15241), .B2(n15239), .A(n15240), .ZN(n15503) );
  INV_X1 U18875 ( .A(n15503), .ZN(n15884) );
  NOR2_X1 U18876 ( .A1(n21129), .A2(n15242), .ZN(n15256) );
  INV_X1 U18877 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15504) );
  OAI22_X1 U18878 ( .A1(n21122), .A2(n15504), .B1(n15243), .B2(n21149), .ZN(
        n15246) );
  NOR3_X1 U18879 ( .A1(n15281), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15244), 
        .ZN(n15245) );
  AOI211_X1 U18880 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n15256), .A(n15246), 
        .B(n15245), .ZN(n15247) );
  OAI21_X1 U18881 ( .B1(n15680), .B2(n21170), .A(n15247), .ZN(n15248) );
  AOI21_X1 U18882 ( .B1(n15884), .B2(n21176), .A(n15248), .ZN(n15249) );
  OAI21_X1 U18883 ( .B1(n15578), .B2(n21137), .A(n15249), .ZN(P1_U2813) );
  OAI21_X1 U18884 ( .B1(n15250), .B2(n15251), .A(n15236), .ZN(n15694) );
  AND2_X1 U18885 ( .A1(n10469), .A2(n15252), .ZN(n15253) );
  OR2_X1 U18886 ( .A1(n15253), .A2(n15239), .ZN(n15897) );
  INV_X1 U18887 ( .A(n15897), .ZN(n15261) );
  OAI22_X1 U18888 ( .A1(n21122), .A2(n21681), .B1(n15254), .B2(n21149), .ZN(
        n15255) );
  AOI21_X1 U18889 ( .B1(n15256), .B2(P1_REIP_REG_26__SCAN_IN), .A(n15255), 
        .ZN(n15259) );
  INV_X1 U18890 ( .A(n15281), .ZN(n15257) );
  INV_X1 U18891 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15684) );
  NAND4_X1 U18892 ( .A1(n15257), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(n15684), .ZN(n15258) );
  OAI211_X1 U18893 ( .C1(n21170), .C2(n15685), .A(n15259), .B(n15258), .ZN(
        n15260) );
  AOI21_X1 U18894 ( .B1(n15261), .B2(n21176), .A(n15260), .ZN(n15262) );
  OAI21_X1 U18895 ( .B1(n15694), .B2(n21137), .A(n15262), .ZN(P1_U2814) );
  NAND2_X1 U18896 ( .A1(n15263), .A2(n15264), .ZN(n15276) );
  AOI21_X1 U18897 ( .B1(n15265), .B2(n15276), .A(n15250), .ZN(n15702) );
  INV_X1 U18898 ( .A(n15702), .ZN(n15583) );
  AOI21_X1 U18899 ( .B1(n15267), .B2(n15266), .A(n10264), .ZN(n15902) );
  NOR2_X1 U18900 ( .A1(n21170), .A2(n15700), .ZN(n15273) );
  XNOR2_X1 U18901 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n15271) );
  AOI22_X1 U18902 ( .A1(n21182), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21174), .ZN(n15270) );
  AND2_X1 U18903 ( .A1(n15429), .A2(n15268), .ZN(n15295) );
  NAND2_X1 U18904 ( .A1(n15295), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15269) );
  OAI211_X1 U18905 ( .C1(n15281), .C2(n15271), .A(n15270), .B(n15269), .ZN(
        n15272) );
  AOI211_X1 U18906 ( .C1(n15902), .C2(n21176), .A(n15273), .B(n15272), .ZN(
        n15274) );
  OAI21_X1 U18907 ( .B1(n15583), .B2(n21137), .A(n15274), .ZN(P1_U2815) );
  NAND2_X1 U18908 ( .A1(n15263), .A2(n15275), .ZN(n15287) );
  INV_X1 U18909 ( .A(n15276), .ZN(n15277) );
  AOI21_X1 U18910 ( .B1(n15278), .B2(n15287), .A(n15277), .ZN(n15710) );
  INV_X1 U18911 ( .A(n15710), .ZN(n15588) );
  INV_X1 U18912 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15506) );
  OAI22_X1 U18913 ( .A1(n21122), .A2(n15506), .B1(n21549), .B2(n21149), .ZN(
        n15279) );
  AOI21_X1 U18914 ( .B1(n15295), .B2(P1_REIP_REG_24__SCAN_IN), .A(n15279), 
        .ZN(n15280) );
  OAI21_X1 U18915 ( .B1(n15281), .B2(P1_REIP_REG_24__SCAN_IN), .A(n15280), 
        .ZN(n15285) );
  OR2_X1 U18916 ( .A1(n15291), .A2(n15282), .ZN(n15283) );
  NAND2_X1 U18917 ( .A1(n15266), .A2(n15283), .ZN(n15906) );
  NOR2_X1 U18918 ( .A1(n15906), .A2(n21161), .ZN(n15284) );
  AOI211_X1 U18919 ( .C1(n21185), .C2(n15707), .A(n15285), .B(n15284), .ZN(
        n15286) );
  OAI21_X1 U18920 ( .B1(n15588), .B2(n21137), .A(n15286), .ZN(P1_U2816) );
  AND2_X1 U18921 ( .A1(n15263), .A2(n15304), .ZN(n15302) );
  OAI21_X1 U18922 ( .B1(n15302), .B2(n15288), .A(n15287), .ZN(n15718) );
  AND2_X1 U18923 ( .A1(n15289), .A2(n15290), .ZN(n15292) );
  OR2_X1 U18924 ( .A1(n15292), .A2(n15291), .ZN(n15923) );
  INV_X1 U18925 ( .A(n15923), .ZN(n15300) );
  AOI22_X1 U18926 ( .A1(n21182), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21174), .ZN(n15298) );
  INV_X1 U18927 ( .A(n15293), .ZN(n15318) );
  NOR2_X1 U18928 ( .A1(n15318), .A2(n15294), .ZN(n15296) );
  OAI21_X1 U18929 ( .B1(n15296), .B2(P1_REIP_REG_23__SCAN_IN), .A(n15295), 
        .ZN(n15297) );
  OAI211_X1 U18930 ( .C1(n21170), .C2(n15713), .A(n15298), .B(n15297), .ZN(
        n15299) );
  AOI21_X1 U18931 ( .B1(n15300), .B2(n21176), .A(n15299), .ZN(n15301) );
  OAI21_X1 U18932 ( .B1(n15718), .B2(n21137), .A(n15301), .ZN(P1_U2817) );
  INV_X1 U18933 ( .A(n15302), .ZN(n15303) );
  OAI21_X1 U18934 ( .B1(n15304), .B2(n15263), .A(n15303), .ZN(n15727) );
  XNOR2_X1 U18935 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15308) );
  AOI22_X1 U18936 ( .A1(n21182), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21174), .ZN(n15307) );
  NOR2_X1 U18937 ( .A1(n21129), .A2(n15305), .ZN(n15327) );
  NAND2_X1 U18938 ( .A1(n15327), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15306) );
  OAI211_X1 U18939 ( .C1(n15318), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        n15309) );
  AOI21_X1 U18940 ( .B1(n15721), .B2(n21185), .A(n15309), .ZN(n15312) );
  AOI21_X1 U18941 ( .B1(n15310), .B2(n9756), .A(n10279), .ZN(n15924) );
  NAND2_X1 U18942 ( .A1(n15924), .A2(n21176), .ZN(n15311) );
  OAI211_X1 U18943 ( .C1(n15727), .C2(n21137), .A(n15312), .B(n15311), .ZN(
        P1_U2818) );
  OAI21_X1 U18944 ( .B1(n15324), .B2(n15313), .A(n9756), .ZN(n15932) );
  AOI21_X1 U18945 ( .B1(n15315), .B2(n15314), .A(n15263), .ZN(n15732) );
  NAND2_X1 U18946 ( .A1(n15732), .A2(n21130), .ZN(n15321) );
  AOI22_X1 U18947 ( .A1(n21182), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21174), .ZN(n15317) );
  NAND2_X1 U18948 ( .A1(n15327), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15316) );
  OAI211_X1 U18949 ( .C1(n15318), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15317), 
        .B(n15316), .ZN(n15319) );
  AOI21_X1 U18950 ( .B1(n15735), .B2(n21185), .A(n15319), .ZN(n15320) );
  OAI211_X1 U18951 ( .C1(n15932), .C2(n21161), .A(n15321), .B(n15320), .ZN(
        P1_U2819) );
  AOI21_X1 U18952 ( .B1(n15323), .B2(n15322), .A(n10428), .ZN(n15745) );
  INV_X1 U18953 ( .A(n15745), .ZN(n15602) );
  AOI21_X1 U18954 ( .B1(n15325), .B2(n15336), .A(n15324), .ZN(n15326) );
  INV_X1 U18955 ( .A(n15326), .ZN(n15952) );
  AOI22_X1 U18956 ( .A1(n21182), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21174), .ZN(n15330) );
  INV_X1 U18957 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15747) );
  INV_X1 U18958 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21386) );
  NOR3_X1 U18959 ( .A1(n15357), .A2(n15747), .A3(n21386), .ZN(n15328) );
  OAI21_X1 U18960 ( .B1(n15328), .B2(P1_REIP_REG_20__SCAN_IN), .A(n15327), 
        .ZN(n15329) );
  OAI211_X1 U18961 ( .C1(n15952), .C2(n21161), .A(n15330), .B(n15329), .ZN(
        n15331) );
  AOI21_X1 U18962 ( .B1(n15741), .B2(n21185), .A(n15331), .ZN(n15332) );
  OAI21_X1 U18963 ( .B1(n15602), .B2(n21137), .A(n15332), .ZN(P1_U2820) );
  OAI21_X1 U18964 ( .B1(n15333), .B2(n15334), .A(n15322), .ZN(n15756) );
  INV_X1 U18965 ( .A(n15336), .ZN(n15337) );
  AOI21_X1 U18966 ( .B1(n15338), .B2(n15351), .A(n15337), .ZN(n15956) );
  XNOR2_X1 U18967 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15345) );
  OR2_X1 U18968 ( .A1(n17628), .A2(n15339), .ZN(n21147) );
  OAI21_X1 U18969 ( .B1(n21149), .B2(n15340), .A(n21147), .ZN(n15343) );
  NAND2_X1 U18970 ( .A1(n15429), .A2(n15341), .ZN(n15366) );
  NOR2_X1 U18971 ( .A1(n15366), .A2(n15747), .ZN(n15342) );
  AOI211_X1 U18972 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n21182), .A(n15343), .B(
        n15342), .ZN(n15344) );
  OAI21_X1 U18973 ( .B1(n15357), .B2(n15345), .A(n15344), .ZN(n15347) );
  NOR2_X1 U18974 ( .A1(n21170), .A2(n15748), .ZN(n15346) );
  AOI211_X1 U18975 ( .C1(n15956), .C2(n21176), .A(n15347), .B(n15346), .ZN(
        n15348) );
  OAI21_X1 U18976 ( .B1(n15756), .B2(n21137), .A(n15348), .ZN(P1_U2821) );
  XNOR2_X1 U18977 ( .A(n9753), .B(n15349), .ZN(n15763) );
  INV_X1 U18978 ( .A(n15763), .ZN(n15609) );
  AOI21_X1 U18979 ( .B1(n15352), .B2(n15350), .A(n15335), .ZN(n15980) );
  NAND2_X1 U18980 ( .A1(n15980), .A2(n21176), .ZN(n15356) );
  OAI21_X1 U18981 ( .B1(n21149), .B2(n15761), .A(n21147), .ZN(n15354) );
  NOR2_X1 U18982 ( .A1(n15366), .A2(n21386), .ZN(n15353) );
  AOI211_X1 U18983 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n21182), .A(n15354), .B(
        n15353), .ZN(n15355) );
  OAI211_X1 U18984 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15357), .A(n15356), 
        .B(n15355), .ZN(n15358) );
  AOI21_X1 U18985 ( .B1(n15759), .B2(n21185), .A(n15358), .ZN(n15359) );
  OAI21_X1 U18986 ( .B1(n15609), .B2(n21137), .A(n15359), .ZN(P1_U2822) );
  AOI21_X1 U18987 ( .B1(n15361), .B2(n15360), .A(n9753), .ZN(n15778) );
  INV_X1 U18988 ( .A(n15778), .ZN(n15616) );
  INV_X1 U18989 ( .A(n15776), .ZN(n15371) );
  OAI21_X1 U18990 ( .B1(n15362), .B2(n15363), .A(n15350), .ZN(n15985) );
  OAI21_X1 U18991 ( .B1(n21149), .B2(n15364), .A(n21147), .ZN(n15365) );
  AOI21_X1 U18992 ( .B1(n21182), .B2(P1_EBX_REG_17__SCAN_IN), .A(n15365), .ZN(
        n15369) );
  INV_X1 U18993 ( .A(n15366), .ZN(n15367) );
  OAI21_X1 U18994 ( .B1(n9804), .B2(P1_REIP_REG_17__SCAN_IN), .A(n15367), .ZN(
        n15368) );
  OAI211_X1 U18995 ( .C1(n15985), .C2(n21161), .A(n15369), .B(n15368), .ZN(
        n15370) );
  AOI21_X1 U18996 ( .B1(n15371), .B2(n21185), .A(n15370), .ZN(n15372) );
  OAI21_X1 U18997 ( .B1(n15616), .B2(n21137), .A(n15372), .ZN(P1_U2823) );
  INV_X1 U18998 ( .A(n15360), .ZN(n15374) );
  AOI21_X1 U18999 ( .B1(n15375), .B2(n15373), .A(n15374), .ZN(n15789) );
  INV_X1 U19000 ( .A(n15789), .ZN(n15623) );
  NOR2_X1 U19001 ( .A1(n21129), .A2(n15376), .ZN(n15414) );
  NAND2_X1 U19002 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15377) );
  OAI21_X1 U19003 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15377), .ZN(n15382) );
  NOR2_X1 U19004 ( .A1(n15378), .A2(n15379), .ZN(n15380) );
  OR2_X1 U19005 ( .A1(n15362), .A2(n15380), .ZN(n15994) );
  OR2_X1 U19006 ( .A1(n21161), .A2(n15994), .ZN(n15381) );
  OAI21_X1 U19007 ( .B1(n15401), .B2(n15382), .A(n15381), .ZN(n15385) );
  AOI22_X1 U19008 ( .A1(n15785), .A2(n21185), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n21182), .ZN(n15383) );
  OAI211_X1 U19009 ( .C1(n21149), .C2(n15787), .A(n15383), .B(n21147), .ZN(
        n15384) );
  AOI211_X1 U19010 ( .C1(n15414), .C2(P1_REIP_REG_16__SCAN_IN), .A(n15385), 
        .B(n15384), .ZN(n15386) );
  OAI21_X1 U19011 ( .B1(n15623), .B2(n21137), .A(n15386), .ZN(P1_U2824) );
  INV_X1 U19012 ( .A(n15388), .ZN(n15390) );
  INV_X1 U19013 ( .A(n15389), .ZN(n15419) );
  NAND2_X1 U19014 ( .A1(n15388), .A2(n15419), .ZN(n15420) );
  OAI21_X1 U19015 ( .B1(n15390), .B2(n15525), .A(n15420), .ZN(n15391) );
  INV_X1 U19016 ( .A(n15392), .ZN(n15393) );
  OAI21_X1 U19017 ( .B1(n15406), .B2(n15393), .A(n15373), .ZN(n15800) );
  AND2_X1 U19018 ( .A1(n15411), .A2(n15395), .ZN(n15396) );
  NOR2_X1 U19019 ( .A1(n15378), .A2(n15396), .ZN(n16004) );
  NAND2_X1 U19020 ( .A1(n15414), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15400) );
  OAI21_X1 U19021 ( .B1(n21149), .B2(n15397), .A(n21147), .ZN(n15398) );
  AOI21_X1 U19022 ( .B1(n21182), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15398), .ZN(
        n15399) );
  OAI211_X1 U19023 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15401), .A(n15400), 
        .B(n15399), .ZN(n15403) );
  NOR2_X1 U19024 ( .A1(n21170), .A2(n15791), .ZN(n15402) );
  AOI211_X1 U19025 ( .C1(n16004), .C2(n21176), .A(n15403), .B(n15402), .ZN(
        n15404) );
  OAI21_X1 U19026 ( .B1(n15800), .B2(n21137), .A(n15404), .ZN(P1_U2825) );
  INV_X1 U19027 ( .A(n15405), .ZN(n15408) );
  INV_X1 U19028 ( .A(n15422), .ZN(n15407) );
  AOI21_X1 U19029 ( .B1(n15408), .B2(n15407), .A(n15406), .ZN(n15809) );
  NAND2_X1 U19030 ( .A1(n9840), .A2(n15409), .ZN(n15410) );
  NAND2_X1 U19031 ( .A1(n15411), .A2(n15410), .ZN(n16012) );
  OAI22_X1 U19032 ( .A1(n15518), .A2(n21122), .B1(n21161), .B2(n16012), .ZN(
        n15412) );
  AOI211_X1 U19033 ( .C1(n21174), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15412), .B(n21163), .ZN(n15416) );
  INV_X1 U19034 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21378) );
  INV_X1 U19035 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21379) );
  OAI21_X1 U19036 ( .B1(n15432), .B2(n21378), .A(n21379), .ZN(n15413) );
  NAND2_X1 U19037 ( .A1(n15414), .A2(n15413), .ZN(n15415) );
  OAI211_X1 U19038 ( .C1(n21170), .C2(n15807), .A(n15416), .B(n15415), .ZN(
        n15417) );
  AOI21_X1 U19039 ( .B1(n15809), .B2(n21130), .A(n15417), .ZN(n15418) );
  INV_X1 U19040 ( .A(n15418), .ZN(P1_U2826) );
  OAI21_X1 U19041 ( .B1(n15388), .B2(n15419), .A(n15420), .ZN(n15524) );
  OAI21_X1 U19042 ( .B1(n15524), .B2(n15525), .A(n15420), .ZN(n15439) );
  NAND2_X1 U19043 ( .A1(n15439), .A2(n15438), .ZN(n15437) );
  INV_X1 U19044 ( .A(n15421), .ZN(n15423) );
  AOI21_X1 U19045 ( .B1(n15437), .B2(n15423), .A(n15422), .ZN(n15820) );
  NAND2_X1 U19046 ( .A1(n15820), .A2(n21130), .ZN(n15436) );
  INV_X1 U19047 ( .A(n9840), .ZN(n15427) );
  AOI21_X1 U19048 ( .B1(n15424), .B2(n15440), .A(n15425), .ZN(n15426) );
  NOR2_X1 U19049 ( .A1(n15427), .A2(n15426), .ZN(n16018) );
  NAND2_X1 U19050 ( .A1(n15429), .A2(n15428), .ZN(n15445) );
  NOR2_X1 U19051 ( .A1(n15445), .A2(n21378), .ZN(n15434) );
  AOI21_X1 U19052 ( .B1(n21174), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21163), .ZN(n15431) );
  NAND2_X1 U19053 ( .A1(n21182), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n15430) );
  OAI211_X1 U19054 ( .C1(n15432), .C2(P1_REIP_REG_13__SCAN_IN), .A(n15431), 
        .B(n15430), .ZN(n15433) );
  AOI211_X1 U19055 ( .C1(n16018), .C2(n21176), .A(n15434), .B(n15433), .ZN(
        n15435) );
  OAI211_X1 U19056 ( .C1(n21170), .C2(n15818), .A(n15436), .B(n15435), .ZN(
        P1_U2827) );
  OAI21_X1 U19057 ( .B1(n15439), .B2(n15438), .A(n15437), .ZN(n15830) );
  XNOR2_X1 U19058 ( .A(n15424), .B(n15440), .ZN(n15523) );
  INV_X1 U19059 ( .A(n15523), .ZN(n16037) );
  AOI21_X1 U19060 ( .B1(n17640), .B2(n15441), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15446) );
  OAI21_X1 U19061 ( .B1(n21149), .B2(n15442), .A(n21147), .ZN(n15443) );
  AOI21_X1 U19062 ( .B1(n21182), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15443), .ZN(
        n15444) );
  OAI21_X1 U19063 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n15448) );
  NOR2_X1 U19064 ( .A1(n21170), .A2(n15826), .ZN(n15447) );
  AOI211_X1 U19065 ( .C1(n21176), .C2(n16037), .A(n15448), .B(n15447), .ZN(
        n15449) );
  OAI21_X1 U19066 ( .B1(n15830), .B2(n21137), .A(n15449), .ZN(P1_U2828) );
  INV_X1 U19067 ( .A(n15450), .ZN(n15452) );
  OAI21_X1 U19068 ( .B1(n15452), .B2(n10466), .A(n15451), .ZN(n15855) );
  INV_X1 U19069 ( .A(n15453), .ZN(n15455) );
  NOR2_X1 U19070 ( .A1(n17628), .A2(n15455), .ZN(n21127) );
  AOI21_X1 U19071 ( .B1(n15454), .B2(n21127), .A(n21129), .ZN(n21117) );
  INV_X1 U19072 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21369) );
  NOR2_X1 U19073 ( .A1(n21173), .A2(n15455), .ZN(n21151) );
  NAND2_X1 U19074 ( .A1(n21128), .A2(n21151), .ZN(n21134) );
  INV_X1 U19075 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21564) );
  OAI21_X1 U19076 ( .B1(n21369), .B2(n21134), .A(n21564), .ZN(n15464) );
  OR2_X1 U19077 ( .A1(n15551), .A2(n15458), .ZN(n15459) );
  NAND2_X1 U19078 ( .A1(n15457), .A2(n15459), .ZN(n17675) );
  OAI22_X1 U19079 ( .A1(n15460), .A2(n21149), .B1(n21161), .B2(n17675), .ZN(
        n15463) );
  AOI21_X1 U19080 ( .B1(n21182), .B2(P1_EBX_REG_8__SCAN_IN), .A(n21163), .ZN(
        n15461) );
  OAI21_X1 U19081 ( .B1(n21170), .B2(n15859), .A(n15461), .ZN(n15462) );
  AOI211_X1 U19082 ( .C1(n21117), .C2(n15464), .A(n15463), .B(n15462), .ZN(
        n15465) );
  OAI21_X1 U19083 ( .B1(n21137), .B2(n15855), .A(n15465), .ZN(P1_U2832) );
  NAND2_X1 U19084 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n21172) );
  NAND2_X1 U19085 ( .A1(n17640), .A2(n21172), .ZN(n15472) );
  INV_X1 U19086 ( .A(n15472), .ZN(n15475) );
  OR2_X1 U19087 ( .A1(n15476), .A2(n15466), .ZN(n21178) );
  INV_X1 U19088 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15468) );
  OAI22_X1 U19089 ( .A1(n15468), .A2(n21122), .B1(n21161), .B2(n15467), .ZN(
        n15469) );
  AOI21_X1 U19090 ( .B1(n21174), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15469), .ZN(n15470) );
  OAI21_X1 U19091 ( .B1(n16291), .B2(n21178), .A(n15470), .ZN(n15474) );
  AND2_X1 U19092 ( .A1(n15472), .A2(n15471), .ZN(n21190) );
  INV_X1 U19093 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21361) );
  NOR2_X1 U19094 ( .A1(n21190), .A2(n21361), .ZN(n15473) );
  AOI211_X1 U19095 ( .C1(n15475), .C2(P1_REIP_REG_1__SCAN_IN), .A(n15474), .B(
        n15473), .ZN(n15480) );
  OAI21_X1 U19096 ( .B1(n15477), .B2(n15476), .A(n21137), .ZN(n21187) );
  NAND2_X1 U19097 ( .A1(n21187), .A2(n15478), .ZN(n15479) );
  OAI211_X1 U19098 ( .C1(n21170), .C2(n15481), .A(n15480), .B(n15479), .ZN(
        P1_U2838) );
  INV_X1 U19099 ( .A(n21187), .ZN(n15496) );
  AOI22_X1 U19100 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n21182), .B1(n17628), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n15487) );
  OAI22_X1 U19101 ( .A1(n21178), .A2(n14436), .B1(n15485), .B2(n21149), .ZN(
        n15484) );
  INV_X1 U19102 ( .A(n13799), .ZN(n15482) );
  OAI22_X1 U19103 ( .A1(n15482), .A2(n21161), .B1(n21173), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n15483) );
  AOI211_X1 U19104 ( .C1(n21185), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15486) );
  OAI211_X1 U19105 ( .C1(n15496), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        P1_U2839) );
  OAI22_X1 U19106 ( .A1(n15490), .A2(n21122), .B1(n21178), .B2(n15489), .ZN(
        n15492) );
  NOR2_X1 U19107 ( .A1(n21129), .A2(n13791), .ZN(n15491) );
  AOI211_X1 U19108 ( .C1(n21176), .C2(n21249), .A(n15492), .B(n15491), .ZN(
        n15494) );
  OAI21_X1 U19109 ( .B1(n21185), .B2(n21174), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15493) );
  OAI211_X1 U19110 ( .C1(n15496), .C2(n15495), .A(n15494), .B(n15493), .ZN(
        P1_U2840) );
  INV_X1 U19111 ( .A(n15497), .ZN(n15499) );
  OAI22_X1 U19112 ( .A1(n15499), .A2(n15545), .B1(n15498), .B2(n15544), .ZN(
        P1_U2841) );
  OAI222_X1 U19113 ( .A1(n15500), .A2(n15544), .B1(n15545), .B2(n15870), .C1(
        n15657), .C2(n15530), .ZN(P1_U2843) );
  INV_X1 U19114 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15502) );
  OAI222_X1 U19115 ( .A1(n15502), .A2(n15544), .B1(n15545), .B2(n15501), .C1(
        n15573), .C2(n15530), .ZN(P1_U2844) );
  OAI222_X1 U19116 ( .A1(n15504), .A2(n15544), .B1(n15545), .B2(n15503), .C1(
        n15578), .C2(n15530), .ZN(P1_U2845) );
  OAI222_X1 U19117 ( .A1(n15897), .A2(n15545), .B1(n21681), .B2(n15544), .C1(
        n15694), .C2(n15530), .ZN(P1_U2846) );
  AOI22_X1 U19118 ( .A1(n15902), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n15505) );
  OAI21_X1 U19119 ( .B1(n15583), .B2(n15556), .A(n15505), .ZN(P1_U2847) );
  OAI222_X1 U19120 ( .A1(n15506), .A2(n15544), .B1(n15545), .B2(n15906), .C1(
        n15588), .C2(n15530), .ZN(P1_U2848) );
  INV_X1 U19121 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15507) );
  OAI222_X1 U19122 ( .A1(n15923), .A2(n15545), .B1(n15507), .B2(n15544), .C1(
        n15718), .C2(n15530), .ZN(P1_U2849) );
  AOI22_X1 U19123 ( .A1(n15924), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15508) );
  OAI21_X1 U19124 ( .B1(n15727), .B2(n15556), .A(n15508), .ZN(P1_U2850) );
  INV_X1 U19125 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15509) );
  INV_X1 U19126 ( .A(n15732), .ZN(n15598) );
  OAI222_X1 U19127 ( .A1(n15932), .A2(n15545), .B1(n15509), .B2(n15544), .C1(
        n15598), .C2(n15530), .ZN(P1_U2851) );
  OAI222_X1 U19128 ( .A1(n15952), .A2(n15545), .B1(n15510), .B2(n15544), .C1(
        n15602), .C2(n15530), .ZN(P1_U2852) );
  AOI22_X1 U19129 ( .A1(n15956), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n15511) );
  OAI21_X1 U19130 ( .B1(n15756), .B2(n15556), .A(n15511), .ZN(P1_U2853) );
  AOI22_X1 U19131 ( .A1(n15980), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15512) );
  OAI21_X1 U19132 ( .B1(n15609), .B2(n15556), .A(n15512), .ZN(P1_U2854) );
  INV_X1 U19133 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15513) );
  OAI222_X1 U19134 ( .A1(n15985), .A2(n15545), .B1(n15513), .B2(n15544), .C1(
        n15616), .C2(n15530), .ZN(P1_U2855) );
  INV_X1 U19135 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15514) );
  OAI22_X1 U19136 ( .A1(n15994), .A2(n15545), .B1(n15514), .B2(n15544), .ZN(
        n15515) );
  AOI21_X1 U19137 ( .B1(n15789), .B2(n15536), .A(n15515), .ZN(n15516) );
  INV_X1 U19138 ( .A(n15516), .ZN(P1_U2856) );
  AOI22_X1 U19139 ( .A1(n16004), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n15517) );
  OAI21_X1 U19140 ( .B1(n15800), .B2(n15556), .A(n15517), .ZN(P1_U2857) );
  OAI22_X1 U19141 ( .A1(n16012), .A2(n15545), .B1(n15518), .B2(n15544), .ZN(
        n15519) );
  AOI21_X1 U19142 ( .B1(n15809), .B2(n15536), .A(n15519), .ZN(n15520) );
  INV_X1 U19143 ( .A(n15520), .ZN(P1_U2858) );
  INV_X1 U19144 ( .A(n15820), .ZN(n15629) );
  AOI22_X1 U19145 ( .A1(n16018), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15521) );
  OAI21_X1 U19146 ( .B1(n15629), .B2(n15556), .A(n15521), .ZN(P1_U2859) );
  INV_X1 U19147 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15522) );
  OAI222_X1 U19148 ( .A1(n15830), .A2(n15530), .B1(n15545), .B2(n15523), .C1(
        n15544), .C2(n15522), .ZN(P1_U2860) );
  XOR2_X1 U19149 ( .A(n15525), .B(n15524), .Z(n17636) );
  INV_X1 U19150 ( .A(n17636), .ZN(n15633) );
  INV_X1 U19151 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15529) );
  NOR2_X1 U19152 ( .A1(n15526), .A2(n15527), .ZN(n15528) );
  OR2_X1 U19153 ( .A1(n15424), .A2(n15528), .ZN(n17631) );
  OAI222_X1 U19154 ( .A1(n15633), .A2(n15530), .B1(n15544), .B2(n15529), .C1(
        n17631), .C2(n15545), .ZN(P1_U2861) );
  AOI21_X1 U19155 ( .B1(n9848), .B2(n10122), .A(n15388), .ZN(n17646) );
  AND2_X1 U19156 ( .A1(n15532), .A2(n15533), .ZN(n15534) );
  OR2_X1 U19157 ( .A1(n15534), .A2(n15526), .ZN(n17641) );
  OAI22_X1 U19158 ( .A1(n17641), .A2(n15545), .B1(n17642), .B2(n15544), .ZN(
        n15535) );
  AOI21_X1 U19159 ( .B1(n17646), .B2(n15536), .A(n15535), .ZN(n15537) );
  INV_X1 U19160 ( .A(n15537), .ZN(P1_U2862) );
  AND2_X1 U19161 ( .A1(n15451), .A2(n15538), .ZN(n15539) );
  OR2_X1 U19162 ( .A1(n15539), .A2(n15531), .ZN(n21115) );
  NAND2_X1 U19163 ( .A1(n15457), .A2(n15540), .ZN(n15541) );
  AND2_X1 U19164 ( .A1(n15532), .A2(n15541), .ZN(n21110) );
  AOI22_X1 U19165 ( .A1(n21110), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n15542) );
  OAI21_X1 U19166 ( .B1(n21115), .B2(n15556), .A(n15542), .ZN(P1_U2863) );
  INV_X1 U19167 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15543) );
  OAI222_X1 U19168 ( .A1(n17675), .A2(n15545), .B1(n15544), .B2(n15543), .C1(
        n15556), .C2(n15855), .ZN(P1_U2864) );
  OR2_X1 U19169 ( .A1(n14515), .A2(n15546), .ZN(n15547) );
  INV_X1 U19170 ( .A(n21131), .ZN(n15647) );
  AOI21_X1 U19171 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15552) );
  NOR2_X1 U19172 ( .A1(n15552), .A2(n15551), .ZN(n21126) );
  AOI22_X1 U19173 ( .A1(n21126), .A2(n15554), .B1(n15553), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n15555) );
  OAI21_X1 U19174 ( .B1(n15647), .B2(n15556), .A(n15555), .ZN(P1_U2865) );
  AOI22_X1 U19175 ( .A1(n15617), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15637), .ZN(n15563) );
  NOR3_X1 U19176 ( .A1(n15637), .A2(n15558), .A3(n15557), .ZN(n15559) );
  INV_X1 U19177 ( .A(DATAI_14_), .ZN(n15561) );
  NAND2_X1 U19178 ( .A1(n15585), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15560) );
  OAI21_X1 U19179 ( .B1(n15585), .B2(n15561), .A(n15560), .ZN(n21230) );
  AOI22_X1 U19180 ( .A1(n15620), .A2(n21230), .B1(n15618), .B2(DATAI_30_), 
        .ZN(n15562) );
  OAI211_X1 U19181 ( .C1(n15564), .C2(n15643), .A(n15563), .B(n15562), .ZN(
        P1_U2874) );
  AOI22_X1 U19182 ( .A1(n15617), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15637), .ZN(n15568) );
  INV_X1 U19183 ( .A(DATAI_13_), .ZN(n15566) );
  NAND2_X1 U19184 ( .A1(n15585), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15565) );
  OAI21_X1 U19185 ( .B1(n15585), .B2(n15566), .A(n15565), .ZN(n21228) );
  AOI22_X1 U19186 ( .A1(n15620), .A2(n21228), .B1(n15618), .B2(DATAI_29_), 
        .ZN(n15567) );
  OAI211_X1 U19187 ( .C1(n15657), .C2(n15643), .A(n15568), .B(n15567), .ZN(
        P1_U2875) );
  AOI22_X1 U19188 ( .A1(n15617), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15637), .ZN(n15572) );
  INV_X1 U19189 ( .A(DATAI_12_), .ZN(n15570) );
  NAND2_X1 U19190 ( .A1(n15585), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15569) );
  OAI21_X1 U19191 ( .B1(n15585), .B2(n15570), .A(n15569), .ZN(n21226) );
  AOI22_X1 U19192 ( .A1(n15620), .A2(n21226), .B1(n15618), .B2(DATAI_28_), 
        .ZN(n15571) );
  OAI211_X1 U19193 ( .C1(n15573), .C2(n15643), .A(n15572), .B(n15571), .ZN(
        P1_U2876) );
  AOI22_X1 U19194 ( .A1(n15617), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15637), .ZN(n15577) );
  INV_X1 U19195 ( .A(DATAI_11_), .ZN(n15575) );
  NAND2_X1 U19196 ( .A1(n15585), .A2(BUF1_REG_11__SCAN_IN), .ZN(n15574) );
  OAI21_X1 U19197 ( .B1(n15585), .B2(n15575), .A(n15574), .ZN(n21224) );
  AOI22_X1 U19198 ( .A1(n15620), .A2(n21224), .B1(n15618), .B2(DATAI_27_), 
        .ZN(n15576) );
  OAI211_X1 U19199 ( .C1(n15578), .C2(n15643), .A(n15577), .B(n15576), .ZN(
        P1_U2877) );
  AOI22_X1 U19200 ( .A1(n15617), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15637), .ZN(n15580) );
  AOI22_X1 U19201 ( .A1(n15620), .A2(n15634), .B1(n15618), .B2(DATAI_26_), 
        .ZN(n15579) );
  OAI211_X1 U19202 ( .C1(n15694), .C2(n15643), .A(n15580), .B(n15579), .ZN(
        P1_U2878) );
  AOI22_X1 U19203 ( .A1(n15617), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15637), .ZN(n15582) );
  AOI22_X1 U19204 ( .A1(n15620), .A2(n15638), .B1(n15618), .B2(DATAI_25_), 
        .ZN(n15581) );
  OAI211_X1 U19205 ( .C1(n15583), .C2(n15643), .A(n15582), .B(n15581), .ZN(
        P1_U2879) );
  AOI22_X1 U19206 ( .A1(n15617), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15637), .ZN(n15587) );
  INV_X1 U19207 ( .A(DATAI_8_), .ZN(n21634) );
  NAND2_X1 U19208 ( .A1(n15585), .A2(BUF1_REG_8__SCAN_IN), .ZN(n15584) );
  OAI21_X1 U19209 ( .B1(n15585), .B2(n21634), .A(n15584), .ZN(n21222) );
  AOI22_X1 U19210 ( .A1(n15620), .A2(n21222), .B1(n15618), .B2(DATAI_24_), 
        .ZN(n15586) );
  OAI211_X1 U19211 ( .C1(n15588), .C2(n15643), .A(n15587), .B(n15586), .ZN(
        P1_U2880) );
  AOI22_X1 U19212 ( .A1(n15617), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15637), .ZN(n15591) );
  AOI22_X1 U19213 ( .A1(n15620), .A2(n15589), .B1(n15618), .B2(DATAI_23_), 
        .ZN(n15590) );
  OAI211_X1 U19214 ( .C1(n15718), .C2(n15643), .A(n15591), .B(n15590), .ZN(
        P1_U2881) );
  AOI22_X1 U19215 ( .A1(n15617), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15637), .ZN(n15594) );
  AOI22_X1 U19216 ( .A1(n15620), .A2(n15592), .B1(n15618), .B2(DATAI_22_), 
        .ZN(n15593) );
  OAI211_X1 U19217 ( .C1(n15727), .C2(n15643), .A(n15594), .B(n15593), .ZN(
        P1_U2882) );
  AOI22_X1 U19218 ( .A1(n15617), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15637), .ZN(n15597) );
  AOI22_X1 U19219 ( .A1(n15620), .A2(n15595), .B1(n15618), .B2(DATAI_21_), 
        .ZN(n15596) );
  OAI211_X1 U19220 ( .C1(n15598), .C2(n15643), .A(n15597), .B(n15596), .ZN(
        P1_U2883) );
  AOI22_X1 U19221 ( .A1(n15617), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n15637), .ZN(n15601) );
  AOI22_X1 U19222 ( .A1(n15620), .A2(n15599), .B1(n15618), .B2(DATAI_20_), 
        .ZN(n15600) );
  OAI211_X1 U19223 ( .C1(n15602), .C2(n15643), .A(n15601), .B(n15600), .ZN(
        P1_U2884) );
  AOI22_X1 U19224 ( .A1(n15617), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15637), .ZN(n15605) );
  AOI22_X1 U19225 ( .A1(n15620), .A2(n15603), .B1(n15618), .B2(DATAI_19_), 
        .ZN(n15604) );
  OAI211_X1 U19226 ( .C1(n15756), .C2(n15643), .A(n15605), .B(n15604), .ZN(
        P1_U2885) );
  AOI22_X1 U19227 ( .A1(n15617), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15637), .ZN(n15608) );
  AOI22_X1 U19228 ( .A1(n15620), .A2(n15606), .B1(n15618), .B2(DATAI_18_), 
        .ZN(n15607) );
  OAI211_X1 U19229 ( .C1(n15609), .C2(n15643), .A(n15608), .B(n15607), .ZN(
        P1_U2886) );
  INV_X1 U19230 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16863) );
  OAI22_X1 U19231 ( .A1(n15611), .A2(n16863), .B1(n15610), .B2(n15644), .ZN(
        n15612) );
  INV_X1 U19232 ( .A(n15612), .ZN(n15615) );
  AOI22_X1 U19233 ( .A1(n15620), .A2(n15613), .B1(n15618), .B2(DATAI_17_), 
        .ZN(n15614) );
  OAI211_X1 U19234 ( .C1(n15616), .C2(n15643), .A(n15615), .B(n15614), .ZN(
        P1_U2887) );
  AOI22_X1 U19235 ( .A1(n15617), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n15637), .ZN(n15622) );
  AOI22_X1 U19236 ( .A1(n15620), .A2(n15619), .B1(n15618), .B2(DATAI_16_), 
        .ZN(n15621) );
  OAI211_X1 U19237 ( .C1(n15623), .C2(n15643), .A(n15622), .B(n15621), .ZN(
        P1_U2888) );
  AOI22_X1 U19238 ( .A1(n15639), .A2(n15624), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n15637), .ZN(n15625) );
  OAI21_X1 U19239 ( .B1(n15800), .B2(n15643), .A(n15625), .ZN(P1_U2889) );
  INV_X1 U19240 ( .A(n15809), .ZN(n15627) );
  AOI22_X1 U19241 ( .A1(n15639), .A2(n21230), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15637), .ZN(n15626) );
  OAI21_X1 U19242 ( .B1(n15627), .B2(n15643), .A(n15626), .ZN(P1_U2890) );
  AOI22_X1 U19243 ( .A1(n15639), .A2(n21228), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15637), .ZN(n15628) );
  OAI21_X1 U19244 ( .B1(n15629), .B2(n15643), .A(n15628), .ZN(P1_U2891) );
  AOI22_X1 U19245 ( .A1(n15639), .A2(n21226), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15637), .ZN(n15630) );
  OAI21_X1 U19246 ( .B1(n15830), .B2(n15643), .A(n15630), .ZN(P1_U2892) );
  INV_X1 U19247 ( .A(n21224), .ZN(n15632) );
  OAI222_X1 U19248 ( .A1(n15633), .A2(n15643), .B1(n15646), .B2(n15632), .C1(
        n15631), .C2(n15644), .ZN(P1_U2893) );
  INV_X1 U19249 ( .A(n17646), .ZN(n15636) );
  AOI22_X1 U19250 ( .A1(n15639), .A2(n15634), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15637), .ZN(n15635) );
  OAI21_X1 U19251 ( .B1(n15636), .B2(n15643), .A(n15635), .ZN(P1_U2894) );
  AOI22_X1 U19252 ( .A1(n15639), .A2(n15638), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15637), .ZN(n15640) );
  OAI21_X1 U19253 ( .B1(n21115), .B2(n15643), .A(n15640), .ZN(P1_U2895) );
  INV_X1 U19254 ( .A(n21222), .ZN(n15642) );
  OAI222_X1 U19255 ( .A1(n15855), .A2(n15643), .B1(n15646), .B2(n15642), .C1(
        n15641), .C2(n15644), .ZN(P1_U2896) );
  OAI222_X1 U19256 ( .A1(n15647), .A2(n15643), .B1(n15646), .B2(n15645), .C1(
        n15644), .C2(n11237), .ZN(P1_U2897) );
  INV_X1 U19257 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21668) );
  NOR2_X1 U19258 ( .A1(n17669), .A2(n21668), .ZN(n15867) );
  NOR2_X1 U19259 ( .A1(n15648), .A2(n17665), .ZN(n15649) );
  AOI211_X1 U19260 ( .C1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n15857), .A(
        n15867), .B(n15649), .ZN(n15656) );
  XNOR2_X2 U19261 ( .A(n15654), .B(n15653), .ZN(n15864) );
  NAND2_X1 U19262 ( .A1(n15864), .A2(n17668), .ZN(n15655) );
  OAI211_X1 U19263 ( .C1(n15657), .C2(n17666), .A(n15656), .B(n15655), .ZN(
        P1_U2970) );
  NAND2_X1 U19264 ( .A1(n15729), .A2(n15891), .ZN(n15659) );
  NAND2_X1 U19265 ( .A1(n15658), .A2(n15659), .ZN(n15663) );
  NAND2_X1 U19266 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15660) );
  NOR2_X1 U19267 ( .A1(n15663), .A2(n15660), .ZN(n15666) );
  AND4_X1 U19268 ( .A1(n15661), .A2(n10347), .A3(n15690), .A4(n15677), .ZN(
        n15662) );
  AND2_X1 U19269 ( .A1(n15663), .A2(n15662), .ZN(n15665) );
  MUX2_X1 U19270 ( .A(n15666), .B(n15665), .S(n15840), .Z(n15667) );
  XNOR2_X1 U19271 ( .A(n15667), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15879) );
  INV_X1 U19272 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21401) );
  NOR2_X1 U19273 ( .A1(n17669), .A2(n21401), .ZN(n15875) );
  AOI21_X1 U19274 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15875), .ZN(n15668) );
  OAI21_X1 U19275 ( .B1(n15669), .B2(n17665), .A(n15668), .ZN(n15670) );
  AOI21_X1 U19276 ( .B1(n15671), .B2(n17654), .A(n15670), .ZN(n15672) );
  OAI21_X1 U19277 ( .B1(n21094), .B2(n15879), .A(n15672), .ZN(P1_U2971) );
  INV_X1 U19278 ( .A(n11169), .ZN(n15673) );
  NAND2_X1 U19279 ( .A1(n15674), .A2(n15673), .ZN(n15676) );
  MUX2_X1 U19280 ( .A(n15676), .B(n15675), .S(n15840), .Z(n15678) );
  XNOR2_X1 U19281 ( .A(n15678), .B(n15677), .ZN(n15887) );
  NOR2_X1 U19282 ( .A1(n17669), .A2(n21399), .ZN(n15882) );
  AOI21_X1 U19283 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15882), .ZN(n15679) );
  OAI21_X1 U19284 ( .B1(n15680), .B2(n17665), .A(n15679), .ZN(n15681) );
  AOI21_X1 U19285 ( .B1(n15682), .B2(n17654), .A(n15681), .ZN(n15683) );
  OAI21_X1 U19286 ( .B1(n21094), .B2(n15887), .A(n15683), .ZN(P1_U2972) );
  NOR2_X1 U19287 ( .A1(n17669), .A2(n15684), .ZN(n15893) );
  NOR2_X1 U19288 ( .A1(n15685), .A2(n17665), .ZN(n15686) );
  AOI211_X1 U19289 ( .C1(n15857), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15893), .B(n15686), .ZN(n15693) );
  AOI21_X1 U19290 ( .B1(n15658), .B2(n15687), .A(n15840), .ZN(n15688) );
  NOR2_X1 U19291 ( .A1(n15689), .A2(n15688), .ZN(n15691) );
  XNOR2_X1 U19292 ( .A(n15691), .B(n15690), .ZN(n15888) );
  NAND2_X1 U19293 ( .A1(n15888), .A2(n17668), .ZN(n15692) );
  OAI211_X1 U19294 ( .C1(n15694), .C2(n17666), .A(n15693), .B(n15692), .ZN(
        P1_U2973) );
  MUX2_X1 U19295 ( .A(n15696), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .S(
        n15729), .Z(n15697) );
  OAI21_X1 U19296 ( .B1(n15704), .B2(n21683), .A(n15697), .ZN(n15698) );
  XOR2_X1 U19297 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n15698), .Z(
        n15905) );
  NAND2_X1 U19298 ( .A1(n15856), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15898) );
  NAND2_X1 U19299 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15699) );
  OAI211_X1 U19300 ( .C1(n15700), .C2(n17665), .A(n15898), .B(n15699), .ZN(
        n15701) );
  AOI21_X1 U19301 ( .B1(n15702), .B2(n17654), .A(n15701), .ZN(n15703) );
  OAI21_X1 U19302 ( .B1(n21094), .B2(n15905), .A(n15703), .ZN(P1_U2974) );
  NOR2_X1 U19303 ( .A1(n15704), .A2(n15658), .ZN(n15705) );
  MUX2_X1 U19304 ( .A(n15705), .B(n15704), .S(n15729), .Z(n15706) );
  XNOR2_X1 U19305 ( .A(n15706), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15915) );
  NAND2_X1 U19306 ( .A1(n15707), .A2(n17655), .ZN(n15708) );
  NAND2_X1 U19307 ( .A1(n15856), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15910) );
  OAI211_X1 U19308 ( .C1(n17671), .C2(n21549), .A(n15708), .B(n15910), .ZN(
        n15709) );
  AOI21_X1 U19309 ( .B1(n15710), .B2(n17654), .A(n15709), .ZN(n15711) );
  OAI21_X1 U19310 ( .B1(n21094), .B2(n15915), .A(n15711), .ZN(P1_U2975) );
  NOR2_X1 U19311 ( .A1(n17669), .A2(n15712), .ZN(n15919) );
  NOR2_X1 U19312 ( .A1(n15713), .A2(n17665), .ZN(n15714) );
  AOI211_X1 U19313 ( .C1(n15857), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15919), .B(n15714), .ZN(n15717) );
  XNOR2_X1 U19314 ( .A(n15729), .B(n10347), .ZN(n15715) );
  XNOR2_X1 U19315 ( .A(n15658), .B(n15715), .ZN(n15916) );
  NAND2_X1 U19316 ( .A1(n15916), .A2(n17668), .ZN(n15716) );
  OAI211_X1 U19317 ( .C1(n15718), .C2(n17666), .A(n15717), .B(n15716), .ZN(
        P1_U2976) );
  INV_X1 U19318 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21393) );
  NOR2_X1 U19319 ( .A1(n17669), .A2(n21393), .ZN(n15928) );
  NOR2_X1 U19320 ( .A1(n17671), .A2(n15719), .ZN(n15720) );
  AOI211_X1 U19321 ( .C1(n15721), .C2(n17655), .A(n15928), .B(n15720), .ZN(
        n15726) );
  NAND2_X1 U19322 ( .A1(n15723), .A2(n15722), .ZN(n15724) );
  XNOR2_X1 U19323 ( .A(n15724), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15925) );
  NAND2_X1 U19324 ( .A1(n15925), .A2(n17668), .ZN(n15725) );
  OAI211_X1 U19325 ( .C1(n15727), .C2(n17666), .A(n15726), .B(n15725), .ZN(
        P1_U2977) );
  NOR2_X1 U19326 ( .A1(n15831), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15738) );
  OAI21_X1 U19327 ( .B1(n15729), .B2(n15977), .A(n15728), .ZN(n15752) );
  OAI22_X1 U19328 ( .A1(n15752), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15840), .B2(n15728), .ZN(n15730) );
  OAI21_X1 U19329 ( .B1(n15943), .B2(n15738), .A(n15730), .ZN(n15731) );
  XNOR2_X1 U19330 ( .A(n15731), .B(n15938), .ZN(n15942) );
  NAND2_X1 U19331 ( .A1(n15732), .A2(n17654), .ZN(n15737) );
  INV_X1 U19332 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21391) );
  NOR2_X1 U19333 ( .A1(n17669), .A2(n21391), .ZN(n15934) );
  NOR2_X1 U19334 ( .A1(n17671), .A2(n15733), .ZN(n15734) );
  AOI211_X1 U19335 ( .C1(n17655), .C2(n15735), .A(n15934), .B(n15734), .ZN(
        n15736) );
  OAI211_X1 U19336 ( .C1(n15942), .C2(n21094), .A(n15737), .B(n15736), .ZN(
        P1_U2978) );
  INV_X1 U19337 ( .A(n15738), .ZN(n15751) );
  NAND2_X1 U19338 ( .A1(n15831), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15750) );
  OAI22_X1 U19339 ( .A1(n15739), .A2(n15751), .B1(n15728), .B2(n15750), .ZN(
        n15740) );
  XNOR2_X1 U19340 ( .A(n15740), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15955) );
  NAND2_X1 U19341 ( .A1(n17655), .A2(n15741), .ZN(n15742) );
  NAND2_X1 U19342 ( .A1(n15856), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15951) );
  OAI211_X1 U19343 ( .C1(n17671), .C2(n15743), .A(n15742), .B(n15951), .ZN(
        n15744) );
  AOI21_X1 U19344 ( .B1(n15745), .B2(n17654), .A(n15744), .ZN(n15746) );
  OAI21_X1 U19345 ( .B1(n15955), .B2(n21094), .A(n15746), .ZN(P1_U2979) );
  NOR2_X1 U19346 ( .A1(n17669), .A2(n15747), .ZN(n15960) );
  NOR2_X1 U19347 ( .A1(n17665), .A2(n15748), .ZN(n15749) );
  AOI211_X1 U19348 ( .C1(n15857), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15960), .B(n15749), .ZN(n15755) );
  NAND2_X1 U19349 ( .A1(n15751), .A2(n15750), .ZN(n15753) );
  XOR2_X1 U19350 ( .A(n15753), .B(n15752), .Z(n15957) );
  NAND2_X1 U19351 ( .A1(n15957), .A2(n17668), .ZN(n15754) );
  OAI211_X1 U19352 ( .C1(n15756), .C2(n17666), .A(n15755), .B(n15754), .ZN(
        P1_U2980) );
  OAI21_X1 U19353 ( .B1(n15758), .B2(n15757), .A(n15728), .ZN(n15982) );
  NAND2_X1 U19354 ( .A1(n17655), .A2(n15759), .ZN(n15760) );
  NAND2_X1 U19355 ( .A1(n15856), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15976) );
  OAI211_X1 U19356 ( .C1(n17671), .C2(n15761), .A(n15760), .B(n15976), .ZN(
        n15762) );
  AOI21_X1 U19357 ( .B1(n15763), .B2(n17654), .A(n15762), .ZN(n15764) );
  OAI21_X1 U19358 ( .B1(n21094), .B2(n15982), .A(n15764), .ZN(P1_U2981) );
  INV_X1 U19359 ( .A(n15765), .ZN(n15767) );
  NAND2_X1 U19360 ( .A1(n15767), .A2(n15766), .ZN(n15839) );
  OAI21_X1 U19361 ( .B1(n15840), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15839), .ZN(n15838) );
  INV_X1 U19362 ( .A(n15768), .ZN(n15770) );
  OAI21_X1 U19363 ( .B1(n15803), .B2(n15770), .A(n15769), .ZN(n15773) );
  NAND2_X1 U19364 ( .A1(n15773), .A2(n15771), .ZN(n15772) );
  MUX2_X1 U19365 ( .A(n15773), .B(n15772), .S(n15840), .Z(n15774) );
  XNOR2_X1 U19366 ( .A(n15774), .B(n15983), .ZN(n15991) );
  INV_X1 U19367 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21383) );
  NOR2_X1 U19368 ( .A1(n17669), .A2(n21383), .ZN(n15987) );
  AOI21_X1 U19369 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15987), .ZN(n15775) );
  OAI21_X1 U19370 ( .B1(n15776), .B2(n17665), .A(n15775), .ZN(n15777) );
  AOI21_X1 U19371 ( .B1(n15778), .B2(n17654), .A(n15777), .ZN(n15779) );
  OAI21_X1 U19372 ( .B1(n15991), .B2(n21094), .A(n15779), .ZN(P1_U2982) );
  INV_X1 U19373 ( .A(n15780), .ZN(n15781) );
  OAI21_X1 U19374 ( .B1(n15838), .B2(n15782), .A(n15781), .ZN(n15797) );
  OAI21_X1 U19375 ( .B1(n15797), .B2(n15793), .A(n15794), .ZN(n15783) );
  XOR2_X1 U19376 ( .A(n15784), .B(n15783), .Z(n15999) );
  NAND2_X1 U19377 ( .A1(n17655), .A2(n15785), .ZN(n15786) );
  OR2_X1 U19378 ( .A1(n17669), .A2(n21382), .ZN(n15993) );
  OAI211_X1 U19379 ( .C1(n17671), .C2(n15787), .A(n15786), .B(n15993), .ZN(
        n15788) );
  AOI21_X1 U19380 ( .B1(n15789), .B2(n17654), .A(n15788), .ZN(n15790) );
  OAI21_X1 U19381 ( .B1(n15999), .B2(n21094), .A(n15790), .ZN(P1_U2983) );
  NOR2_X1 U19382 ( .A1(n17669), .A2(n21381), .ZN(n16003) );
  NOR2_X1 U19383 ( .A1(n17665), .A2(n15791), .ZN(n15792) );
  AOI211_X1 U19384 ( .C1(n15857), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16003), .B(n15792), .ZN(n15799) );
  INV_X1 U19385 ( .A(n15793), .ZN(n15795) );
  NAND2_X1 U19386 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  XNOR2_X1 U19387 ( .A(n15797), .B(n15796), .ZN(n16000) );
  NAND2_X1 U19388 ( .A1(n16000), .A2(n17668), .ZN(n15798) );
  OAI211_X1 U19389 ( .C1(n15800), .C2(n17666), .A(n15799), .B(n15798), .ZN(
        P1_U2984) );
  INV_X1 U19390 ( .A(n15801), .ZN(n15802) );
  XNOR2_X1 U19391 ( .A(n15729), .B(n15970), .ZN(n15804) );
  XNOR2_X1 U19392 ( .A(n15805), .B(n15804), .ZN(n16016) );
  NAND2_X1 U19393 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15806) );
  NAND2_X1 U19394 ( .A1(n15856), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16011) );
  OAI211_X1 U19395 ( .C1(n17665), .C2(n15807), .A(n15806), .B(n16011), .ZN(
        n15808) );
  AOI21_X1 U19396 ( .B1(n15809), .B2(n17654), .A(n15808), .ZN(n15810) );
  OAI21_X1 U19397 ( .B1(n16016), .B2(n21094), .A(n15810), .ZN(P1_U2985) );
  INV_X1 U19398 ( .A(n15811), .ZN(n15813) );
  OAI21_X1 U19399 ( .B1(n15838), .B2(n15813), .A(n15812), .ZN(n15825) );
  INV_X1 U19400 ( .A(n15823), .ZN(n15814) );
  OAI21_X1 U19401 ( .B1(n15825), .B2(n15814), .A(n15822), .ZN(n15815) );
  XNOR2_X1 U19402 ( .A(n15816), .B(n15815), .ZN(n16023) );
  NOR2_X1 U19403 ( .A1(n17669), .A2(n21378), .ZN(n16017) );
  AOI21_X1 U19404 ( .B1(n15857), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16017), .ZN(n15817) );
  OAI21_X1 U19405 ( .B1(n15818), .B2(n17665), .A(n15817), .ZN(n15819) );
  AOI21_X1 U19406 ( .B1(n15820), .B2(n17654), .A(n15819), .ZN(n15821) );
  OAI21_X1 U19407 ( .B1(n16023), .B2(n21094), .A(n15821), .ZN(P1_U2986) );
  NAND2_X1 U19408 ( .A1(n15823), .A2(n15822), .ZN(n15824) );
  XNOR2_X1 U19409 ( .A(n15825), .B(n15824), .ZN(n16032) );
  NAND2_X1 U19410 ( .A1(n16032), .A2(n17668), .ZN(n15829) );
  INV_X1 U19411 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21706) );
  NOR2_X1 U19412 ( .A1(n17669), .A2(n21706), .ZN(n16036) );
  NOR2_X1 U19413 ( .A1(n17665), .A2(n15826), .ZN(n15827) );
  AOI211_X1 U19414 ( .C1(n15857), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16036), .B(n15827), .ZN(n15828) );
  OAI211_X1 U19415 ( .C1(n15830), .C2(n17666), .A(n15829), .B(n15828), .ZN(
        P1_U2987) );
  NAND2_X1 U19416 ( .A1(n15831), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15833) );
  INV_X1 U19417 ( .A(n15839), .ZN(n15832) );
  NAND3_X1 U19418 ( .A1(n15832), .A2(n15840), .A3(n16059), .ZN(n15843) );
  OAI21_X1 U19419 ( .B1(n15838), .B2(n15833), .A(n15843), .ZN(n15834) );
  XNOR2_X1 U19420 ( .A(n15834), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16048) );
  NAND2_X1 U19421 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15835) );
  NAND2_X1 U19422 ( .A1(n15856), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n16043) );
  OAI211_X1 U19423 ( .C1(n17665), .C2(n17638), .A(n15835), .B(n16043), .ZN(
        n15836) );
  AOI21_X1 U19424 ( .B1(n17636), .B2(n17654), .A(n15836), .ZN(n15837) );
  OAI21_X1 U19425 ( .B1(n16048), .B2(n21094), .A(n15837), .ZN(P1_U2988) );
  XNOR2_X1 U19426 ( .A(n15838), .B(n16059), .ZN(n15842) );
  NAND2_X1 U19427 ( .A1(n15839), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15841) );
  MUX2_X1 U19428 ( .A(n15842), .B(n15841), .S(n15840), .Z(n15844) );
  NAND2_X1 U19429 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15845) );
  NAND2_X1 U19430 ( .A1(n15856), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16050) );
  OAI211_X1 U19431 ( .C1(n17665), .C2(n17644), .A(n15845), .B(n16050), .ZN(
        n15846) );
  AOI21_X1 U19432 ( .B1(n17646), .B2(n17654), .A(n15846), .ZN(n15847) );
  OAI21_X1 U19433 ( .B1(n16065), .B2(n21094), .A(n15847), .ZN(P1_U2989) );
  XNOR2_X1 U19434 ( .A(n15840), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15848) );
  XNOR2_X1 U19435 ( .A(n15765), .B(n15848), .ZN(n16072) );
  NAND2_X1 U19436 ( .A1(n16072), .A2(n17668), .ZN(n15852) );
  NOR2_X1 U19437 ( .A1(n17669), .A2(n21372), .ZN(n16066) );
  NOR2_X1 U19438 ( .A1(n17671), .A2(n15849), .ZN(n15850) );
  AOI211_X1 U19439 ( .C1(n17655), .C2(n21118), .A(n16066), .B(n15850), .ZN(
        n15851) );
  OAI211_X1 U19440 ( .C1(n17666), .C2(n21115), .A(n15852), .B(n15851), .ZN(
        P1_U2990) );
  XNOR2_X1 U19441 ( .A(n15854), .B(n15853), .ZN(n17680) );
  INV_X1 U19442 ( .A(n17680), .ZN(n15863) );
  INV_X1 U19443 ( .A(n15855), .ZN(n15861) );
  AOI22_X1 U19444 ( .A1(n15857), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n15856), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15858) );
  OAI21_X1 U19445 ( .B1(n15859), .B2(n17665), .A(n15858), .ZN(n15860) );
  AOI21_X1 U19446 ( .B1(n15861), .B2(n17654), .A(n15860), .ZN(n15862) );
  OAI21_X1 U19447 ( .B1(n15863), .B2(n21094), .A(n15862), .ZN(P1_U2991) );
  NAND2_X1 U19448 ( .A1(n15864), .A2(n21251), .ZN(n15869) );
  INV_X1 U19449 ( .A(n15873), .ZN(n15880) );
  NOR3_X1 U19450 ( .A1(n15880), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15871), .ZN(n15866) );
  AOI211_X1 U19451 ( .C1(n10214), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15867), .B(n15866), .ZN(n15868) );
  OAI211_X1 U19452 ( .C1(n15870), .C2(n16051), .A(n15869), .B(n15868), .ZN(
        P1_U3002) );
  AND3_X1 U19453 ( .A1(n15873), .A2(n15872), .A3(n15871), .ZN(n15874) );
  AOI211_X1 U19454 ( .C1(n15883), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15875), .B(n15874), .ZN(n15878) );
  NAND2_X1 U19455 ( .A1(n15876), .A2(n21250), .ZN(n15877) );
  OAI211_X1 U19456 ( .C1(n15879), .C2(n16064), .A(n15878), .B(n15877), .ZN(
        P1_U3003) );
  NOR2_X1 U19457 ( .A1(n15880), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15881) );
  AOI211_X1 U19458 ( .C1(n15883), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15882), .B(n15881), .ZN(n15886) );
  NAND2_X1 U19459 ( .A1(n15884), .A2(n21250), .ZN(n15885) );
  OAI211_X1 U19460 ( .C1(n15887), .C2(n16064), .A(n15886), .B(n15885), .ZN(
        P1_U3004) );
  NAND2_X1 U19461 ( .A1(n15888), .A2(n21251), .ZN(n15896) );
  NAND3_X1 U19462 ( .A1(n15889), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15890) );
  NOR2_X1 U19463 ( .A1(n15908), .A2(n15890), .ZN(n15899) );
  OR2_X1 U19464 ( .A1(n15901), .A2(n15899), .ZN(n15894) );
  NOR3_X1 U19465 ( .A1(n15908), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15891), .ZN(n15892) );
  AOI211_X1 U19466 ( .C1(n15894), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15893), .B(n15892), .ZN(n15895) );
  OAI211_X1 U19467 ( .C1(n16051), .C2(n15897), .A(n15896), .B(n15895), .ZN(
        P1_U3005) );
  INV_X1 U19468 ( .A(n15898), .ZN(n15900) );
  AOI211_X1 U19469 ( .C1(n15901), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15900), .B(n15899), .ZN(n15904) );
  NAND2_X1 U19470 ( .A1(n15902), .A2(n21250), .ZN(n15903) );
  OAI211_X1 U19471 ( .C1(n15905), .C2(n16064), .A(n15904), .B(n15903), .ZN(
        P1_U3006) );
  INV_X1 U19472 ( .A(n15906), .ZN(n15913) );
  AOI21_X1 U19473 ( .B1(n10347), .B2(n16031), .A(n15907), .ZN(n15911) );
  INV_X1 U19474 ( .A(n15908), .ZN(n15920) );
  NAND3_X1 U19475 ( .A1(n15920), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n21683), .ZN(n15909) );
  OAI211_X1 U19476 ( .C1(n15911), .C2(n21683), .A(n15910), .B(n15909), .ZN(
        n15912) );
  AOI21_X1 U19477 ( .B1(n15913), .B2(n21250), .A(n15912), .ZN(n15914) );
  OAI21_X1 U19478 ( .B1(n15915), .B2(n16064), .A(n15914), .ZN(P1_U3007) );
  NAND2_X1 U19479 ( .A1(n15916), .A2(n21251), .ZN(n15922) );
  NOR2_X1 U19480 ( .A1(n15917), .A2(n10347), .ZN(n15918) );
  AOI211_X1 U19481 ( .C1(n15920), .C2(n10347), .A(n15919), .B(n15918), .ZN(
        n15921) );
  OAI211_X1 U19482 ( .C1(n16051), .C2(n15923), .A(n15922), .B(n15921), .ZN(
        P1_U3008) );
  INV_X1 U19483 ( .A(n15924), .ZN(n15931) );
  NAND2_X1 U19484 ( .A1(n15925), .A2(n21251), .ZN(n15930) );
  XNOR2_X1 U19485 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15926) );
  NOR2_X1 U19486 ( .A1(n15933), .A2(n15926), .ZN(n15927) );
  AOI211_X1 U19487 ( .C1(n10224), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15928), .B(n15927), .ZN(n15929) );
  OAI211_X1 U19488 ( .C1(n16051), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        P1_U3009) );
  INV_X1 U19489 ( .A(n15932), .ZN(n15940) );
  INV_X1 U19490 ( .A(n15933), .ZN(n15935) );
  AOI21_X1 U19491 ( .B1(n15935), .B2(n15938), .A(n15934), .ZN(n15936) );
  OAI21_X1 U19492 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15939) );
  AOI21_X1 U19493 ( .B1(n15940), .B2(n21250), .A(n15939), .ZN(n15941) );
  OAI21_X1 U19494 ( .B1(n15942), .B2(n16064), .A(n15941), .ZN(P1_U3010) );
  INV_X1 U19495 ( .A(n16031), .ZN(n15945) );
  AOI21_X1 U19496 ( .B1(n15945), .B2(n15944), .A(n15943), .ZN(n15949) );
  OAI21_X1 U19497 ( .B1(n15958), .B2(n15947), .A(n15946), .ZN(n15948) );
  OAI21_X1 U19498 ( .B1(n15949), .B2(n15961), .A(n15948), .ZN(n15950) );
  OAI211_X1 U19499 ( .C1(n15952), .C2(n16051), .A(n15951), .B(n15950), .ZN(
        n15953) );
  INV_X1 U19500 ( .A(n15953), .ZN(n15954) );
  OAI21_X1 U19501 ( .B1(n15955), .B2(n16064), .A(n15954), .ZN(P1_U3011) );
  INV_X1 U19502 ( .A(n15956), .ZN(n15964) );
  NAND2_X1 U19503 ( .A1(n15957), .A2(n21251), .ZN(n15963) );
  NOR2_X1 U19504 ( .A1(n15958), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15959) );
  AOI211_X1 U19505 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15961), .A(
        n15960), .B(n15959), .ZN(n15962) );
  OAI211_X1 U19506 ( .C1(n16051), .C2(n15964), .A(n15963), .B(n15962), .ZN(
        P1_U3012) );
  OAI21_X1 U19507 ( .B1(n16010), .B2(n15966), .A(n15965), .ZN(n15967) );
  OAI211_X1 U19508 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15969), .A(
        n15968), .B(n15967), .ZN(n16019) );
  AOI21_X1 U19509 ( .B1(n15970), .B2(n17673), .A(n16019), .ZN(n16008) );
  OAI21_X1 U19510 ( .B1(n16030), .B2(n15973), .A(n16008), .ZN(n15989) );
  INV_X1 U19511 ( .A(n15989), .ZN(n15978) );
  INV_X1 U19512 ( .A(n15971), .ZN(n15972) );
  NAND2_X1 U19513 ( .A1(n16020), .A2(n15972), .ZN(n16001) );
  INV_X1 U19514 ( .A(n16001), .ZN(n15974) );
  NAND3_X1 U19515 ( .A1(n15974), .A2(n15973), .A3(n15977), .ZN(n15975) );
  OAI211_X1 U19516 ( .C1(n15978), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        n15979) );
  AOI21_X1 U19517 ( .B1(n15980), .B2(n21250), .A(n15979), .ZN(n15981) );
  OAI21_X1 U19518 ( .B1(n15982), .B2(n16064), .A(n15981), .ZN(P1_U3013) );
  NAND2_X1 U19519 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15984) );
  OAI21_X1 U19520 ( .B1(n16001), .B2(n15984), .A(n15983), .ZN(n15988) );
  NOR2_X1 U19521 ( .A1(n15985), .A2(n16051), .ZN(n15986) );
  AOI211_X1 U19522 ( .C1(n15989), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        n15990) );
  OAI21_X1 U19523 ( .B1(n15991), .B2(n16064), .A(n15990), .ZN(P1_U3014) );
  INV_X1 U19524 ( .A(n16008), .ZN(n15997) );
  XNOR2_X1 U19525 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15992) );
  NOR2_X1 U19526 ( .A1(n16001), .A2(n15992), .ZN(n15996) );
  OAI21_X1 U19527 ( .B1(n15994), .B2(n16051), .A(n15993), .ZN(n15995) );
  AOI211_X1 U19528 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15997), .A(
        n15996), .B(n15995), .ZN(n15998) );
  OAI21_X1 U19529 ( .B1(n15999), .B2(n16064), .A(n15998), .ZN(P1_U3015) );
  NAND2_X1 U19530 ( .A1(n16000), .A2(n21251), .ZN(n16006) );
  NOR2_X1 U19531 ( .A1(n16001), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16002) );
  AOI211_X1 U19532 ( .C1(n16004), .C2(n21250), .A(n16003), .B(n16002), .ZN(
        n16005) );
  OAI211_X1 U19533 ( .C1(n16008), .C2(n16007), .A(n16006), .B(n16005), .ZN(
        P1_U3016) );
  NOR4_X1 U19534 ( .A1(n16049), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16010), .A4(n16009), .ZN(n16014) );
  OAI21_X1 U19535 ( .B1(n16012), .B2(n16051), .A(n16011), .ZN(n16013) );
  AOI211_X1 U19536 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16019), .A(
        n16014), .B(n16013), .ZN(n16015) );
  OAI21_X1 U19537 ( .B1(n16016), .B2(n16064), .A(n16015), .ZN(P1_U3017) );
  AOI21_X1 U19538 ( .B1(n16018), .B2(n21250), .A(n16017), .ZN(n16022) );
  OAI21_X1 U19539 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16020), .A(
        n16019), .ZN(n16021) );
  OAI211_X1 U19540 ( .C1(n16023), .C2(n16064), .A(n16022), .B(n16021), .ZN(
        P1_U3018) );
  INV_X1 U19541 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16034) );
  INV_X1 U19542 ( .A(n16024), .ZN(n16029) );
  NAND2_X1 U19543 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16025), .ZN(
        n16026) );
  NAND2_X1 U19544 ( .A1(n16027), .A2(n16026), .ZN(n16028) );
  OAI211_X1 U19545 ( .C1(n16030), .C2(n16029), .A(n16055), .B(n16028), .ZN(
        n16046) );
  AOI21_X1 U19546 ( .B1(n16034), .B2(n16031), .A(n16046), .ZN(n16041) );
  NAND2_X1 U19547 ( .A1(n16032), .A2(n21251), .ZN(n16039) );
  INV_X1 U19548 ( .A(n16033), .ZN(n16042) );
  NOR4_X1 U19549 ( .A1(n16049), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n16034), .A4(n16042), .ZN(n16035) );
  AOI211_X1 U19550 ( .C1(n21250), .C2(n16037), .A(n16036), .B(n16035), .ZN(
        n16038) );
  OAI211_X1 U19551 ( .C1(n16041), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P1_U3019) );
  NOR3_X1 U19552 ( .A1(n16049), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16042), .ZN(n16045) );
  OAI21_X1 U19553 ( .B1(n17631), .B2(n16051), .A(n16043), .ZN(n16044) );
  AOI211_X1 U19554 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16046), .A(
        n16045), .B(n16044), .ZN(n16047) );
  OAI21_X1 U19555 ( .B1(n16048), .B2(n16064), .A(n16047), .ZN(P1_U3020) );
  NOR2_X1 U19556 ( .A1(n16049), .A2(n21461), .ZN(n17683) );
  NOR3_X1 U19557 ( .A1(n17674), .A2(n16069), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16062) );
  OAI21_X1 U19558 ( .B1(n17641), .B2(n16051), .A(n16050), .ZN(n16061) );
  INV_X1 U19559 ( .A(n16052), .ZN(n16053) );
  NAND3_X1 U19560 ( .A1(n16055), .A2(n16054), .A3(n16053), .ZN(n16057) );
  NAND2_X1 U19561 ( .A1(n16057), .A2(n16056), .ZN(n16070) );
  NOR2_X1 U19562 ( .A1(n17674), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16058) );
  NAND2_X1 U19563 ( .A1(n17683), .A2(n16058), .ZN(n16067) );
  AOI21_X1 U19564 ( .B1(n16070), .B2(n16067), .A(n16059), .ZN(n16060) );
  AOI211_X1 U19565 ( .C1(n17683), .C2(n16062), .A(n16061), .B(n16060), .ZN(
        n16063) );
  OAI21_X1 U19566 ( .B1(n16065), .B2(n16064), .A(n16063), .ZN(P1_U3021) );
  AOI21_X1 U19567 ( .B1(n21110), .B2(n21250), .A(n16066), .ZN(n16068) );
  OAI211_X1 U19568 ( .C1(n16070), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        n16071) );
  AOI21_X1 U19569 ( .B1(n16072), .B2(n21251), .A(n16071), .ZN(n16073) );
  INV_X1 U19570 ( .A(n16073), .ZN(P1_U3022) );
  NAND3_X1 U19571 ( .A1(n16075), .A2(n17610), .A3(n16074), .ZN(n17617) );
  OAI211_X1 U19572 ( .C1(n16385), .C2(n9720), .A(n17617), .B(n16077), .ZN(
        n16078) );
  MUX2_X1 U19573 ( .A(n16078), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n21258), .Z(P1_U3478) );
  NAND2_X1 U19574 ( .A1(n21274), .A2(n21428), .ZN(n16080) );
  MUX2_X1 U19575 ( .A(n16081), .B(n16080), .S(n16079), .Z(n16082) );
  OAI21_X1 U19576 ( .B1(n16088), .B2(n14436), .A(n16082), .ZN(n16083) );
  MUX2_X1 U19577 ( .A(n16083), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n21258), .Z(P1_U3477) );
  NAND2_X1 U19578 ( .A1(n16084), .A2(n21274), .ZN(n16086) );
  MUX2_X1 U19579 ( .A(n16086), .B(n16085), .S(n11176), .Z(n16087) );
  OAI21_X1 U19580 ( .B1(n16088), .B2(n16291), .A(n16087), .ZN(n16089) );
  MUX2_X1 U19581 ( .A(n16089), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n21258), .Z(P1_U3476) );
  INV_X1 U19582 ( .A(n16090), .ZN(n16095) );
  INV_X1 U19583 ( .A(n16091), .ZN(n16092) );
  NAND2_X1 U19584 ( .A1(n16093), .A2(n16092), .ZN(n16098) );
  OAI22_X1 U19585 ( .A1(n16095), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n16098), .B2(n16094), .ZN(n16096) );
  AOI21_X1 U19586 ( .B1(n16341), .B2(n16097), .A(n16096), .ZN(n17593) );
  INV_X1 U19587 ( .A(n16098), .ZN(n16101) );
  AOI22_X1 U19588 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16099), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13202), .ZN(n16106) );
  NAND2_X1 U19589 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16107) );
  INV_X1 U19590 ( .A(n16107), .ZN(n16100) );
  AOI22_X1 U19591 ( .A1(n16102), .A2(n16101), .B1(n16106), .B2(n16100), .ZN(
        n16103) );
  OAI21_X1 U19592 ( .B1(n17593), .B2(n16114), .A(n16103), .ZN(n16104) );
  MUX2_X1 U19593 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16104), .S(
        n16116), .Z(P1_U3473) );
  OAI222_X1 U19594 ( .A1(n16108), .A2(n16112), .B1(n16107), .B2(n16106), .C1(
        n16114), .C2(n16105), .ZN(n16109) );
  MUX2_X1 U19595 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16109), .S(
        n16116), .Z(P1_U3472) );
  INV_X1 U19596 ( .A(n16110), .ZN(n16115) );
  INV_X1 U19597 ( .A(n16111), .ZN(n16113) );
  OAI22_X1 U19598 ( .A1(n16115), .A2(n16114), .B1(n16113), .B2(n16112), .ZN(
        n16117) );
  MUX2_X1 U19599 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16117), .S(
        n16116), .Z(P1_U3469) );
  INV_X1 U19600 ( .A(n16155), .ZN(n16119) );
  NAND2_X1 U19601 ( .A1(n21280), .A2(n16118), .ZN(n16425) );
  NAND2_X1 U19602 ( .A1(n16119), .A2(n16425), .ZN(n16120) );
  AOI21_X1 U19603 ( .B1(n16120), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n16385), 
        .ZN(n16126) );
  NOR2_X1 U19604 ( .A1(n16159), .A2(n16341), .ZN(n16124) );
  NAND2_X1 U19605 ( .A1(n16164), .A2(n16121), .ZN(n16206) );
  INV_X1 U19606 ( .A(n16206), .ZN(n16122) );
  NOR2_X1 U19607 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16123), .ZN(
        n16128) );
  INV_X1 U19608 ( .A(n16128), .ZN(n16153) );
  INV_X1 U19609 ( .A(n16425), .ZN(n16151) );
  INV_X1 U19610 ( .A(n16124), .ZN(n16125) );
  AOI22_X1 U19611 ( .A1(n16126), .A2(n16125), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16206), .ZN(n16127) );
  OAI211_X1 U19612 ( .C1(n16128), .C2(n17711), .A(n16166), .B(n16127), .ZN(
        n16150) );
  AOI22_X1 U19613 ( .A1(n16151), .A2(n16297), .B1(
        P1_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n16150), .ZN(n16129) );
  OAI21_X1 U19614 ( .B1(n16295), .B2(n16153), .A(n16129), .ZN(n16130) );
  AOI21_X1 U19615 ( .B1(n16155), .B2(n21284), .A(n16130), .ZN(n16131) );
  OAI21_X1 U19616 ( .B1(n16157), .B2(n16394), .A(n16131), .ZN(P1_U3033) );
  AOI22_X1 U19617 ( .A1(n16151), .A2(n16306), .B1(
        P1_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n16150), .ZN(n16132) );
  OAI21_X1 U19618 ( .B1(n16304), .B2(n16153), .A(n16132), .ZN(n16133) );
  AOI21_X1 U19619 ( .B1(n16155), .B2(n21290), .A(n16133), .ZN(n16134) );
  OAI21_X1 U19620 ( .B1(n16157), .B2(n16399), .A(n16134), .ZN(P1_U3034) );
  AOI22_X1 U19621 ( .A1(n16151), .A2(n21752), .B1(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n16150), .ZN(n16135) );
  OAI21_X1 U19622 ( .B1(n21748), .B2(n16153), .A(n16135), .ZN(n16136) );
  AOI21_X1 U19623 ( .B1(n16155), .B2(n21296), .A(n16136), .ZN(n16137) );
  OAI21_X1 U19624 ( .B1(n16157), .B2(n21750), .A(n16137), .ZN(P1_U3035) );
  AOI22_X1 U19625 ( .A1(n16151), .A2(n16314), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n16150), .ZN(n16138) );
  OAI21_X1 U19626 ( .B1(n16312), .B2(n16153), .A(n16138), .ZN(n16139) );
  AOI21_X1 U19627 ( .B1(n16155), .B2(n21302), .A(n16139), .ZN(n16140) );
  OAI21_X1 U19628 ( .B1(n16157), .B2(n16407), .A(n16140), .ZN(P1_U3036) );
  AOI22_X1 U19629 ( .A1(n16151), .A2(n16319), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n16150), .ZN(n16141) );
  OAI21_X1 U19630 ( .B1(n16317), .B2(n16153), .A(n16141), .ZN(n16142) );
  AOI21_X1 U19631 ( .B1(n16155), .B2(n21308), .A(n16142), .ZN(n16143) );
  OAI21_X1 U19632 ( .B1(n16157), .B2(n16412), .A(n16143), .ZN(P1_U3037) );
  AOI22_X1 U19633 ( .A1(n16151), .A2(n16324), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n16150), .ZN(n16144) );
  OAI21_X1 U19634 ( .B1(n16322), .B2(n16153), .A(n16144), .ZN(n16145) );
  AOI21_X1 U19635 ( .B1(n16155), .B2(n21314), .A(n16145), .ZN(n16146) );
  OAI21_X1 U19636 ( .B1(n16157), .B2(n16417), .A(n16146), .ZN(P1_U3038) );
  AOI22_X1 U19637 ( .A1(n16151), .A2(n16329), .B1(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n16150), .ZN(n16147) );
  OAI21_X1 U19638 ( .B1(n16327), .B2(n16153), .A(n16147), .ZN(n16148) );
  AOI21_X1 U19639 ( .B1(n16155), .B2(n21320), .A(n16148), .ZN(n16149) );
  OAI21_X1 U19640 ( .B1(n16157), .B2(n16422), .A(n16149), .ZN(P1_U3039) );
  AOI22_X1 U19641 ( .A1(n16151), .A2(n16335), .B1(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n16150), .ZN(n16152) );
  OAI21_X1 U19642 ( .B1(n16333), .B2(n16153), .A(n16152), .ZN(n16154) );
  AOI21_X1 U19643 ( .B1(n16155), .B2(n21328), .A(n16154), .ZN(n16156) );
  OAI21_X1 U19644 ( .B1(n16157), .B2(n16431), .A(n16156), .ZN(P1_U3040) );
  NAND2_X1 U19645 ( .A1(n16190), .A2(n16167), .ZN(n16158) );
  AOI21_X1 U19646 ( .B1(n16158), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n16385), 
        .ZN(n16163) );
  NOR2_X1 U19647 ( .A1(n16159), .A2(n14436), .ZN(n16160) );
  NOR2_X1 U19648 ( .A1(n16164), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16249) );
  INV_X1 U19649 ( .A(n16160), .ZN(n16162) );
  AOI22_X1 U19650 ( .A1(n16163), .A2(n16162), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n16191), .ZN(n16165) );
  OAI21_X1 U19651 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16164), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16256) );
  NAND2_X1 U19652 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n16170) );
  OAI22_X1 U19653 ( .A1(n16295), .A2(n16191), .B1(n16390), .B2(n16190), .ZN(
        n16168) );
  AOI21_X1 U19654 ( .B1(n16193), .B2(n16297), .A(n16168), .ZN(n16169) );
  OAI211_X1 U19655 ( .C1(n16196), .C2(n16394), .A(n16170), .B(n16169), .ZN(
        P1_U3049) );
  NAND2_X1 U19656 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n16173) );
  OAI22_X1 U19657 ( .A1(n16304), .A2(n16191), .B1(n16395), .B2(n16190), .ZN(
        n16171) );
  AOI21_X1 U19658 ( .B1(n16193), .B2(n16306), .A(n16171), .ZN(n16172) );
  OAI211_X1 U19659 ( .C1(n16196), .C2(n16399), .A(n16173), .B(n16172), .ZN(
        P1_U3050) );
  NAND2_X1 U19660 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n16176) );
  OAI22_X1 U19661 ( .A1(n21748), .A2(n16191), .B1(n21758), .B2(n16190), .ZN(
        n16174) );
  AOI21_X1 U19662 ( .B1(n16193), .B2(n21752), .A(n16174), .ZN(n16175) );
  OAI211_X1 U19663 ( .C1(n16196), .C2(n21750), .A(n16176), .B(n16175), .ZN(
        P1_U3051) );
  NAND2_X1 U19664 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n16179) );
  OAI22_X1 U19665 ( .A1(n16312), .A2(n16191), .B1(n16403), .B2(n16190), .ZN(
        n16177) );
  AOI21_X1 U19666 ( .B1(n16193), .B2(n16314), .A(n16177), .ZN(n16178) );
  OAI211_X1 U19667 ( .C1(n16196), .C2(n16407), .A(n16179), .B(n16178), .ZN(
        P1_U3052) );
  NAND2_X1 U19668 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n16182) );
  OAI22_X1 U19669 ( .A1(n16317), .A2(n16191), .B1(n16408), .B2(n16190), .ZN(
        n16180) );
  AOI21_X1 U19670 ( .B1(n16193), .B2(n16319), .A(n16180), .ZN(n16181) );
  OAI211_X1 U19671 ( .C1(n16196), .C2(n16412), .A(n16182), .B(n16181), .ZN(
        P1_U3053) );
  NAND2_X1 U19672 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n16185) );
  OAI22_X1 U19673 ( .A1(n16322), .A2(n16191), .B1(n16413), .B2(n16190), .ZN(
        n16183) );
  AOI21_X1 U19674 ( .B1(n16193), .B2(n16324), .A(n16183), .ZN(n16184) );
  OAI211_X1 U19675 ( .C1(n16196), .C2(n16417), .A(n16185), .B(n16184), .ZN(
        P1_U3054) );
  NAND2_X1 U19676 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n16188) );
  OAI22_X1 U19677 ( .A1(n16327), .A2(n16191), .B1(n16418), .B2(n16190), .ZN(
        n16186) );
  AOI21_X1 U19678 ( .B1(n16193), .B2(n16329), .A(n16186), .ZN(n16187) );
  OAI211_X1 U19679 ( .C1(n16196), .C2(n16422), .A(n16188), .B(n16187), .ZN(
        P1_U3055) );
  NAND2_X1 U19680 ( .A1(n16189), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n16195) );
  OAI22_X1 U19681 ( .A1(n16333), .A2(n16191), .B1(n16426), .B2(n16190), .ZN(
        n16192) );
  AOI21_X1 U19682 ( .B1(n16193), .B2(n16335), .A(n16192), .ZN(n16194) );
  OAI211_X1 U19683 ( .C1(n16196), .C2(n16431), .A(n16195), .B(n16194), .ZN(
        P1_U3056) );
  INV_X1 U19684 ( .A(n16237), .ZN(n16198) );
  OAI21_X1 U19685 ( .B1(n16198), .B2(n16197), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n16199) );
  OAI21_X1 U19686 ( .B1(n16341), .B2(n16247), .A(n16199), .ZN(n16201) );
  NOR2_X1 U19687 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16200), .ZN(
        n16209) );
  AOI21_X1 U19688 ( .B1(n16201), .B2(n17711), .A(n16209), .ZN(n16205) );
  INV_X1 U19689 ( .A(n16351), .ZN(n16204) );
  NAND2_X1 U19690 ( .A1(n14436), .A2(n21274), .ZN(n16208) );
  OR2_X1 U19691 ( .A1(n16248), .A2(n16206), .ZN(n16207) );
  NOR2_X1 U19692 ( .A1(n16237), .A2(n21287), .ZN(n16211) );
  INV_X1 U19693 ( .A(n16209), .ZN(n16239) );
  OAI22_X1 U19694 ( .A1(n16295), .A2(n16239), .B1(n16390), .B2(n16238), .ZN(
        n16210) );
  AOI211_X1 U19695 ( .C1(n21278), .C2(n16242), .A(n16211), .B(n16210), .ZN(
        n16212) );
  OAI21_X1 U19696 ( .B1(n16245), .B2(n16213), .A(n16212), .ZN(P1_U3065) );
  INV_X1 U19697 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16217) );
  NOR2_X1 U19698 ( .A1(n16237), .A2(n21293), .ZN(n16215) );
  OAI22_X1 U19699 ( .A1(n16304), .A2(n16239), .B1(n16395), .B2(n16238), .ZN(
        n16214) );
  AOI211_X1 U19700 ( .C1(n21288), .C2(n16242), .A(n16215), .B(n16214), .ZN(
        n16216) );
  OAI21_X1 U19701 ( .B1(n16245), .B2(n16217), .A(n16216), .ZN(P1_U3066) );
  NOR2_X1 U19702 ( .A1(n16237), .A2(n21299), .ZN(n16219) );
  OAI22_X1 U19703 ( .A1(n21748), .A2(n16239), .B1(n21758), .B2(n16238), .ZN(
        n16218) );
  AOI211_X1 U19704 ( .C1(n21294), .C2(n16242), .A(n16219), .B(n16218), .ZN(
        n16220) );
  OAI21_X1 U19705 ( .B1(n16245), .B2(n16221), .A(n16220), .ZN(P1_U3067) );
  NOR2_X1 U19706 ( .A1(n16237), .A2(n21305), .ZN(n16223) );
  OAI22_X1 U19707 ( .A1(n16312), .A2(n16239), .B1(n16403), .B2(n16238), .ZN(
        n16222) );
  AOI211_X1 U19708 ( .C1(n21300), .C2(n16242), .A(n16223), .B(n16222), .ZN(
        n16224) );
  OAI21_X1 U19709 ( .B1(n16245), .B2(n21619), .A(n16224), .ZN(P1_U3068) );
  INV_X1 U19710 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16228) );
  NOR2_X1 U19711 ( .A1(n16237), .A2(n21311), .ZN(n16226) );
  OAI22_X1 U19712 ( .A1(n16317), .A2(n16239), .B1(n16408), .B2(n16238), .ZN(
        n16225) );
  AOI211_X1 U19713 ( .C1(n21306), .C2(n16242), .A(n16226), .B(n16225), .ZN(
        n16227) );
  OAI21_X1 U19714 ( .B1(n16245), .B2(n16228), .A(n16227), .ZN(P1_U3069) );
  NOR2_X1 U19715 ( .A1(n16237), .A2(n21317), .ZN(n16230) );
  OAI22_X1 U19716 ( .A1(n16322), .A2(n16239), .B1(n16413), .B2(n16238), .ZN(
        n16229) );
  AOI211_X1 U19717 ( .C1(n21312), .C2(n16242), .A(n16230), .B(n16229), .ZN(
        n16231) );
  OAI21_X1 U19718 ( .B1(n16245), .B2(n16232), .A(n16231), .ZN(P1_U3070) );
  NOR2_X1 U19719 ( .A1(n16237), .A2(n21323), .ZN(n16234) );
  OAI22_X1 U19720 ( .A1(n16327), .A2(n16239), .B1(n16418), .B2(n16238), .ZN(
        n16233) );
  AOI211_X1 U19721 ( .C1(n21318), .C2(n16242), .A(n16234), .B(n16233), .ZN(
        n16235) );
  OAI21_X1 U19722 ( .B1(n16245), .B2(n16236), .A(n16235), .ZN(P1_U3071) );
  NOR2_X1 U19723 ( .A1(n16237), .A2(n21334), .ZN(n16241) );
  OAI22_X1 U19724 ( .A1(n16333), .A2(n16239), .B1(n16426), .B2(n16238), .ZN(
        n16240) );
  AOI211_X1 U19725 ( .C1(n21325), .C2(n16242), .A(n16241), .B(n16240), .ZN(
        n16243) );
  OAI21_X1 U19726 ( .B1(n16245), .B2(n16244), .A(n16243), .ZN(P1_U3072) );
  NAND2_X1 U19727 ( .A1(n16281), .A2(n16280), .ZN(n16246) );
  AOI21_X1 U19728 ( .B1(n16246), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n16385), 
        .ZN(n16255) );
  NOR2_X1 U19729 ( .A1(n16247), .A2(n14436), .ZN(n16250) );
  INV_X1 U19730 ( .A(n16248), .ZN(n16342) );
  INV_X1 U19731 ( .A(n16250), .ZN(n16254) );
  INV_X1 U19732 ( .A(n16251), .ZN(n16252) );
  NOR2_X1 U19733 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16252), .ZN(
        n16283) );
  INV_X1 U19734 ( .A(n16283), .ZN(n16253) );
  AOI22_X1 U19735 ( .A1(n16255), .A2(n16254), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n16253), .ZN(n16257) );
  NAND3_X1 U19736 ( .A1(n16351), .A2(n16257), .A3(n16256), .ZN(n16279) );
  NAND2_X1 U19737 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n16260) );
  OAI22_X1 U19738 ( .A1(n16390), .A2(n16281), .B1(n16280), .B2(n21287), .ZN(
        n16258) );
  AOI21_X1 U19739 ( .B1(n21279), .B2(n16283), .A(n16258), .ZN(n16259) );
  OAI211_X1 U19740 ( .C1(n16286), .C2(n16394), .A(n16260), .B(n16259), .ZN(
        P1_U3081) );
  NAND2_X1 U19741 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n16263) );
  OAI22_X1 U19742 ( .A1(n16395), .A2(n16281), .B1(n16280), .B2(n21293), .ZN(
        n16261) );
  AOI21_X1 U19743 ( .B1(n21289), .B2(n16283), .A(n16261), .ZN(n16262) );
  OAI211_X1 U19744 ( .C1(n16286), .C2(n16399), .A(n16263), .B(n16262), .ZN(
        P1_U3082) );
  NAND2_X1 U19745 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n16266) );
  OAI22_X1 U19746 ( .A1(n21758), .A2(n16281), .B1(n16280), .B2(n21299), .ZN(
        n16264) );
  AOI21_X1 U19747 ( .B1(n21295), .B2(n16283), .A(n16264), .ZN(n16265) );
  OAI211_X1 U19748 ( .C1(n16286), .C2(n21750), .A(n16266), .B(n16265), .ZN(
        P1_U3083) );
  NAND2_X1 U19749 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n16269) );
  OAI22_X1 U19750 ( .A1(n16403), .A2(n16281), .B1(n16280), .B2(n21305), .ZN(
        n16267) );
  AOI21_X1 U19751 ( .B1(n21301), .B2(n16283), .A(n16267), .ZN(n16268) );
  OAI211_X1 U19752 ( .C1(n16286), .C2(n16407), .A(n16269), .B(n16268), .ZN(
        P1_U3084) );
  NAND2_X1 U19753 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n16272) );
  OAI22_X1 U19754 ( .A1(n16408), .A2(n16281), .B1(n16280), .B2(n21311), .ZN(
        n16270) );
  AOI21_X1 U19755 ( .B1(n21307), .B2(n16283), .A(n16270), .ZN(n16271) );
  OAI211_X1 U19756 ( .C1(n16286), .C2(n16412), .A(n16272), .B(n16271), .ZN(
        P1_U3085) );
  NAND2_X1 U19757 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n16275) );
  OAI22_X1 U19758 ( .A1(n16413), .A2(n16281), .B1(n16280), .B2(n21317), .ZN(
        n16273) );
  AOI21_X1 U19759 ( .B1(n21313), .B2(n16283), .A(n16273), .ZN(n16274) );
  OAI211_X1 U19760 ( .C1(n16286), .C2(n16417), .A(n16275), .B(n16274), .ZN(
        P1_U3086) );
  NAND2_X1 U19761 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n16278) );
  OAI22_X1 U19762 ( .A1(n16418), .A2(n16281), .B1(n16280), .B2(n21323), .ZN(
        n16276) );
  AOI21_X1 U19763 ( .B1(n21319), .B2(n16283), .A(n16276), .ZN(n16277) );
  OAI211_X1 U19764 ( .C1(n16286), .C2(n16422), .A(n16278), .B(n16277), .ZN(
        P1_U3087) );
  NAND2_X1 U19765 ( .A1(n16279), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n16285) );
  OAI22_X1 U19766 ( .A1(n16426), .A2(n16281), .B1(n16280), .B2(n21334), .ZN(
        n16282) );
  AOI21_X1 U19767 ( .B1(n21327), .B2(n16283), .A(n16282), .ZN(n16284) );
  OAI211_X1 U19768 ( .C1(n16286), .C2(n16431), .A(n16285), .B(n16284), .ZN(
        P1_U3088) );
  INV_X1 U19769 ( .A(n21333), .ZN(n16288) );
  OAI21_X1 U19770 ( .B1(n16336), .B2(n16288), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n16289) );
  NAND2_X1 U19771 ( .A1(n16289), .A2(n21274), .ZN(n16301) );
  INV_X1 U19772 ( .A(n16301), .ZN(n16293) );
  AND2_X1 U19773 ( .A1(n21272), .A2(n14436), .ZN(n16300) );
  INV_X1 U19774 ( .A(n16298), .ZN(n16292) );
  NAND3_X1 U19775 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n16294), .ZN(n21273) );
  OR2_X1 U19776 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21273), .ZN(
        n16332) );
  OAI22_X1 U19777 ( .A1(n16295), .A2(n16332), .B1(n16390), .B2(n21333), .ZN(
        n16296) );
  AOI21_X1 U19778 ( .B1(n16336), .B2(n16297), .A(n16296), .ZN(n16303) );
  AOI22_X1 U19779 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16298), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n16332), .ZN(n16299) );
  NAND2_X1 U19780 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n16302) );
  OAI211_X1 U19781 ( .C1(n16340), .C2(n16394), .A(n16303), .B(n16302), .ZN(
        P1_U3129) );
  OAI22_X1 U19782 ( .A1(n16304), .A2(n16332), .B1(n16395), .B2(n21333), .ZN(
        n16305) );
  AOI21_X1 U19783 ( .B1(n16336), .B2(n16306), .A(n16305), .ZN(n16308) );
  NAND2_X1 U19784 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n16307) );
  OAI211_X1 U19785 ( .C1(n16340), .C2(n16399), .A(n16308), .B(n16307), .ZN(
        P1_U3130) );
  OAI22_X1 U19786 ( .A1(n21748), .A2(n16332), .B1(n21758), .B2(n21333), .ZN(
        n16309) );
  AOI21_X1 U19787 ( .B1(n16336), .B2(n21752), .A(n16309), .ZN(n16311) );
  NAND2_X1 U19788 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n16310) );
  OAI211_X1 U19789 ( .C1(n16340), .C2(n21750), .A(n16311), .B(n16310), .ZN(
        P1_U3131) );
  OAI22_X1 U19790 ( .A1(n16312), .A2(n16332), .B1(n16403), .B2(n21333), .ZN(
        n16313) );
  AOI21_X1 U19791 ( .B1(n16336), .B2(n16314), .A(n16313), .ZN(n16316) );
  NAND2_X1 U19792 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n16315) );
  OAI211_X1 U19793 ( .C1(n16340), .C2(n16407), .A(n16316), .B(n16315), .ZN(
        P1_U3132) );
  OAI22_X1 U19794 ( .A1(n16317), .A2(n16332), .B1(n16408), .B2(n21333), .ZN(
        n16318) );
  AOI21_X1 U19795 ( .B1(n16336), .B2(n16319), .A(n16318), .ZN(n16321) );
  NAND2_X1 U19796 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n16320) );
  OAI211_X1 U19797 ( .C1(n16340), .C2(n16412), .A(n16321), .B(n16320), .ZN(
        P1_U3133) );
  OAI22_X1 U19798 ( .A1(n16322), .A2(n16332), .B1(n16413), .B2(n21333), .ZN(
        n16323) );
  AOI21_X1 U19799 ( .B1(n16336), .B2(n16324), .A(n16323), .ZN(n16326) );
  NAND2_X1 U19800 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n16325) );
  OAI211_X1 U19801 ( .C1(n16340), .C2(n16417), .A(n16326), .B(n16325), .ZN(
        P1_U3134) );
  OAI22_X1 U19802 ( .A1(n16327), .A2(n16332), .B1(n16418), .B2(n21333), .ZN(
        n16328) );
  AOI21_X1 U19803 ( .B1(n16336), .B2(n16329), .A(n16328), .ZN(n16331) );
  NAND2_X1 U19804 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n16330) );
  OAI211_X1 U19805 ( .C1(n16340), .C2(n16422), .A(n16331), .B(n16330), .ZN(
        P1_U3135) );
  OAI22_X1 U19806 ( .A1(n16333), .A2(n16332), .B1(n16426), .B2(n21333), .ZN(
        n16334) );
  AOI21_X1 U19807 ( .B1(n16336), .B2(n16335), .A(n16334), .ZN(n16339) );
  NAND2_X1 U19808 ( .A1(n16337), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n16338) );
  OAI211_X1 U19809 ( .C1(n16340), .C2(n16431), .A(n16339), .B(n16338), .ZN(
        P1_U3136) );
  NAND2_X1 U19810 ( .A1(n21272), .A2(n16341), .ZN(n16348) );
  INV_X1 U19811 ( .A(n16348), .ZN(n16344) );
  INV_X1 U19812 ( .A(n16424), .ZN(n16347) );
  OAI21_X1 U19813 ( .B1(n16347), .B2(n21329), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n16349) );
  AOI21_X1 U19814 ( .B1(n16349), .B2(n16348), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n16352) );
  NOR2_X1 U19815 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16386), .ZN(
        n16377) );
  NAND2_X1 U19816 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n16355) );
  OAI22_X1 U19817 ( .A1(n16390), .A2(n16424), .B1(n16375), .B2(n21287), .ZN(
        n16353) );
  AOI21_X1 U19818 ( .B1(n21279), .B2(n16377), .A(n16353), .ZN(n16354) );
  OAI211_X1 U19819 ( .C1(n16380), .C2(n16394), .A(n16355), .B(n16354), .ZN(
        P1_U3145) );
  NAND2_X1 U19820 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n16358) );
  OAI22_X1 U19821 ( .A1(n16375), .A2(n21293), .B1(n16395), .B2(n16424), .ZN(
        n16356) );
  AOI21_X1 U19822 ( .B1(n21289), .B2(n16377), .A(n16356), .ZN(n16357) );
  OAI211_X1 U19823 ( .C1(n16380), .C2(n16399), .A(n16358), .B(n16357), .ZN(
        P1_U3146) );
  NAND2_X1 U19824 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n16361) );
  OAI22_X1 U19825 ( .A1(n16375), .A2(n21299), .B1(n21758), .B2(n16424), .ZN(
        n16359) );
  AOI21_X1 U19826 ( .B1(n21295), .B2(n16377), .A(n16359), .ZN(n16360) );
  OAI211_X1 U19827 ( .C1(n16380), .C2(n21750), .A(n16361), .B(n16360), .ZN(
        P1_U3147) );
  NAND2_X1 U19828 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n16364) );
  OAI22_X1 U19829 ( .A1(n16375), .A2(n21305), .B1(n16403), .B2(n16424), .ZN(
        n16362) );
  AOI21_X1 U19830 ( .B1(n21301), .B2(n16377), .A(n16362), .ZN(n16363) );
  OAI211_X1 U19831 ( .C1(n16380), .C2(n16407), .A(n16364), .B(n16363), .ZN(
        P1_U3148) );
  NAND2_X1 U19832 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n16367) );
  OAI22_X1 U19833 ( .A1(n16375), .A2(n21311), .B1(n16408), .B2(n16424), .ZN(
        n16365) );
  AOI21_X1 U19834 ( .B1(n21307), .B2(n16377), .A(n16365), .ZN(n16366) );
  OAI211_X1 U19835 ( .C1(n16380), .C2(n16412), .A(n16367), .B(n16366), .ZN(
        P1_U3149) );
  NAND2_X1 U19836 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n16370) );
  OAI22_X1 U19837 ( .A1(n16375), .A2(n21317), .B1(n16413), .B2(n16424), .ZN(
        n16368) );
  AOI21_X1 U19838 ( .B1(n21313), .B2(n16377), .A(n16368), .ZN(n16369) );
  OAI211_X1 U19839 ( .C1(n16380), .C2(n16417), .A(n16370), .B(n16369), .ZN(
        P1_U3150) );
  NAND2_X1 U19840 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n16373) );
  OAI22_X1 U19841 ( .A1(n16375), .A2(n21323), .B1(n16418), .B2(n16424), .ZN(
        n16371) );
  AOI21_X1 U19842 ( .B1(n21319), .B2(n16377), .A(n16371), .ZN(n16372) );
  OAI211_X1 U19843 ( .C1(n16380), .C2(n16422), .A(n16373), .B(n16372), .ZN(
        P1_U3151) );
  NAND2_X1 U19844 ( .A1(n16374), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n16379) );
  OAI22_X1 U19845 ( .A1(n16375), .A2(n21334), .B1(n16426), .B2(n16424), .ZN(
        n16376) );
  AOI21_X1 U19846 ( .B1(n21327), .B2(n16377), .A(n16376), .ZN(n16378) );
  OAI211_X1 U19847 ( .C1(n16380), .C2(n16431), .A(n16379), .B(n16378), .ZN(
        P1_U3152) );
  INV_X1 U19848 ( .A(n16381), .ZN(n16428) );
  AOI21_X1 U19849 ( .B1(n21272), .B2(n16382), .A(n16428), .ZN(n16388) );
  INV_X1 U19850 ( .A(n16388), .ZN(n16384) );
  AOI22_X1 U19851 ( .A1(n16384), .A2(n21274), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16383), .ZN(n16432) );
  AOI22_X1 U19852 ( .A1(n16388), .A2(n16387), .B1(n16386), .B2(n16385), .ZN(
        n16389) );
  NAND2_X1 U19853 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n16393) );
  OAI22_X1 U19854 ( .A1(n16390), .A2(n16425), .B1(n16424), .B2(n21287), .ZN(
        n16391) );
  AOI21_X1 U19855 ( .B1(n21279), .B2(n16428), .A(n16391), .ZN(n16392) );
  OAI211_X1 U19856 ( .C1(n16432), .C2(n16394), .A(n16393), .B(n16392), .ZN(
        P1_U3153) );
  NAND2_X1 U19857 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n16398) );
  OAI22_X1 U19858 ( .A1(n16395), .A2(n16425), .B1(n16424), .B2(n21293), .ZN(
        n16396) );
  AOI21_X1 U19859 ( .B1(n21289), .B2(n16428), .A(n16396), .ZN(n16397) );
  OAI211_X1 U19860 ( .C1(n16432), .C2(n16399), .A(n16398), .B(n16397), .ZN(
        P1_U3154) );
  NAND2_X1 U19861 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n16402) );
  OAI22_X1 U19862 ( .A1(n21758), .A2(n16425), .B1(n16424), .B2(n21299), .ZN(
        n16400) );
  AOI21_X1 U19863 ( .B1(n21295), .B2(n16428), .A(n16400), .ZN(n16401) );
  OAI211_X1 U19864 ( .C1(n16432), .C2(n21750), .A(n16402), .B(n16401), .ZN(
        P1_U3155) );
  NAND2_X1 U19865 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n16406) );
  OAI22_X1 U19866 ( .A1(n16403), .A2(n16425), .B1(n16424), .B2(n21305), .ZN(
        n16404) );
  AOI21_X1 U19867 ( .B1(n21301), .B2(n16428), .A(n16404), .ZN(n16405) );
  OAI211_X1 U19868 ( .C1(n16432), .C2(n16407), .A(n16406), .B(n16405), .ZN(
        P1_U3156) );
  NAND2_X1 U19869 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n16411) );
  OAI22_X1 U19870 ( .A1(n16408), .A2(n16425), .B1(n16424), .B2(n21311), .ZN(
        n16409) );
  AOI21_X1 U19871 ( .B1(n21307), .B2(n16428), .A(n16409), .ZN(n16410) );
  OAI211_X1 U19872 ( .C1(n16432), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        P1_U3157) );
  NAND2_X1 U19873 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n16416) );
  OAI22_X1 U19874 ( .A1(n16413), .A2(n16425), .B1(n16424), .B2(n21317), .ZN(
        n16414) );
  AOI21_X1 U19875 ( .B1(n21313), .B2(n16428), .A(n16414), .ZN(n16415) );
  OAI211_X1 U19876 ( .C1(n16432), .C2(n16417), .A(n16416), .B(n16415), .ZN(
        P1_U3158) );
  NAND2_X1 U19877 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n16421) );
  OAI22_X1 U19878 ( .A1(n16418), .A2(n16425), .B1(n16424), .B2(n21323), .ZN(
        n16419) );
  AOI21_X1 U19879 ( .B1(n21319), .B2(n16428), .A(n16419), .ZN(n16420) );
  OAI211_X1 U19880 ( .C1(n16432), .C2(n16422), .A(n16421), .B(n16420), .ZN(
        P1_U3159) );
  NAND2_X1 U19881 ( .A1(n16423), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n16430) );
  OAI22_X1 U19882 ( .A1(n16426), .A2(n16425), .B1(n16424), .B2(n21334), .ZN(
        n16427) );
  AOI21_X1 U19883 ( .B1(n21327), .B2(n16428), .A(n16427), .ZN(n16429) );
  OAI211_X1 U19884 ( .C1(n16432), .C2(n16431), .A(n16430), .B(n16429), .ZN(
        P1_U3160) );
  OAI21_X1 U19885 ( .B1(n16433), .B2(n16434), .A(n20276), .ZN(n16437) );
  INV_X1 U19886 ( .A(n16435), .ZN(n16436) );
  AOI21_X1 U19887 ( .B1(n15158), .B2(n16437), .A(n16436), .ZN(n16442) );
  AOI22_X1 U19888 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_29__SCAN_IN), .ZN(n16439) );
  NAND2_X1 U19889 ( .A1(n20245), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16438) );
  OAI211_X1 U19890 ( .C1(n16440), .C2(n20260), .A(n16439), .B(n16438), .ZN(
        n16441) );
  OAI21_X1 U19892 ( .B1(n16772), .B2(n20267), .A(n16443), .ZN(P2_U2826) );
  AND2_X1 U19893 ( .A1(n16462), .A2(n16445), .ZN(n16446) );
  NOR2_X1 U19894 ( .A1(n10471), .A2(n16446), .ZN(n17145) );
  INV_X1 U19895 ( .A(n17145), .ZN(n16459) );
  OAI21_X1 U19896 ( .B1(n16447), .B2(n16449), .A(n16448), .ZN(n17142) );
  INV_X1 U19897 ( .A(n17142), .ZN(n16457) );
  INV_X1 U19898 ( .A(n16450), .ZN(n16466) );
  OAI21_X1 U19899 ( .B1(n16466), .B2(n16877), .A(n20276), .ZN(n16451) );
  AOI21_X1 U19900 ( .B1(n15158), .B2(n16451), .A(n16433), .ZN(n16456) );
  AOI22_X1 U19901 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n16453) );
  NAND2_X1 U19902 ( .A1(n20245), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16452) );
  OAI211_X1 U19903 ( .C1(n16454), .C2(n20260), .A(n16453), .B(n16452), .ZN(
        n16455) );
  AOI211_X1 U19904 ( .C1(n16457), .C2(n20269), .A(n16456), .B(n16455), .ZN(
        n16458) );
  OAI21_X1 U19905 ( .B1(n16459), .B2(n20267), .A(n16458), .ZN(P2_U2827) );
  NAND2_X1 U19906 ( .A1(n13263), .A2(n16460), .ZN(n16461) );
  NAND2_X1 U19907 ( .A1(n16462), .A2(n16461), .ZN(n17150) );
  NOR2_X1 U19908 ( .A1(n13256), .A2(n16463), .ZN(n16464) );
  INV_X1 U19909 ( .A(n17159), .ZN(n16472) );
  OAI21_X1 U19910 ( .B1(n16465), .B2(n16888), .A(n20276), .ZN(n16467) );
  AOI21_X1 U19911 ( .B1(n15158), .B2(n16467), .A(n16466), .ZN(n16471) );
  OAI22_X1 U19912 ( .A1(n20258), .A2(n16889), .B1(n21001), .B2(n20249), .ZN(
        n16468) );
  AOI21_X1 U19913 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n20245), .A(n16468), .ZN(
        n16469) );
  OAI21_X1 U19914 ( .B1(n16872), .B2(n20260), .A(n16469), .ZN(n16470) );
  AOI211_X1 U19915 ( .C1(n16472), .C2(n20269), .A(n16471), .B(n16470), .ZN(
        n16473) );
  OAI21_X1 U19916 ( .B1(n17150), .B2(n20267), .A(n16473), .ZN(P2_U2828) );
  INV_X1 U19917 ( .A(n16899), .ZN(n16480) );
  AOI21_X1 U19918 ( .B1(n16474), .B2(n16897), .A(n20933), .ZN(n16476) );
  INV_X1 U19919 ( .A(n16465), .ZN(n16475) );
  OAI22_X1 U19920 ( .A1(n20258), .A2(n16895), .B1(n20997), .B2(n20249), .ZN(
        n16477) );
  AOI21_X1 U19921 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n20245), .A(n16477), .ZN(
        n16478) );
  INV_X1 U19922 ( .A(n13264), .ZN(n16482) );
  OAI21_X1 U19923 ( .B1(n16481), .B2(n16483), .A(n16482), .ZN(n17170) );
  AOI21_X1 U19924 ( .B1(n16485), .B2(n16501), .A(n16484), .ZN(n17173) );
  OAI21_X1 U19925 ( .B1(n16486), .B2(n16909), .A(n20276), .ZN(n16488) );
  INV_X1 U19926 ( .A(n16474), .ZN(n16487) );
  AOI21_X1 U19927 ( .B1(n15158), .B2(n16488), .A(n16487), .ZN(n16494) );
  XNOR2_X1 U19928 ( .A(n16489), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n16492) );
  AOI22_X1 U19929 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_25__SCAN_IN), .ZN(n16491) );
  NAND2_X1 U19930 ( .A1(n20245), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16490) );
  OAI211_X1 U19931 ( .C1(n16492), .C2(n20260), .A(n16491), .B(n16490), .ZN(
        n16493) );
  AOI211_X1 U19932 ( .C1(n17173), .C2(n20269), .A(n16494), .B(n16493), .ZN(
        n16495) );
  OAI21_X1 U19933 ( .B1(n17170), .B2(n20267), .A(n16495), .ZN(P2_U2830) );
  AOI21_X1 U19934 ( .B1(n16497), .B2(n16496), .A(n16481), .ZN(n17186) );
  INV_X1 U19935 ( .A(n17186), .ZN(n16511) );
  NAND2_X1 U19936 ( .A1(n16498), .A2(n16499), .ZN(n16500) );
  AOI21_X1 U19937 ( .B1(n16502), .B2(n16914), .A(n20933), .ZN(n16504) );
  INV_X1 U19938 ( .A(n16486), .ZN(n16503) );
  OAI21_X1 U19939 ( .B1(n16678), .B2(n16504), .A(n16503), .ZN(n16507) );
  OAI22_X1 U19940 ( .A1(n20258), .A2(n16916), .B1(n20993), .B2(n20249), .ZN(
        n16505) );
  AOI21_X1 U19941 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n20245), .A(n16505), .ZN(
        n16506) );
  OAI211_X1 U19942 ( .C1(n20260), .C2(n16508), .A(n16507), .B(n16506), .ZN(
        n16509) );
  AOI21_X1 U19943 ( .B1(n16918), .B2(n20269), .A(n16509), .ZN(n16510) );
  OAI21_X1 U19944 ( .B1(n16511), .B2(n20267), .A(n16510), .ZN(P2_U2831) );
  NAND2_X1 U19945 ( .A1(n16512), .A2(n16513), .ZN(n16514) );
  INV_X1 U19946 ( .A(n17204), .ZN(n16528) );
  INV_X1 U19947 ( .A(n16516), .ZN(n16928) );
  AOI21_X1 U19948 ( .B1(n16515), .B2(n16928), .A(n20933), .ZN(n16517) );
  OAI21_X1 U19949 ( .B1(n16517), .B2(n16678), .A(n16502), .ZN(n16520) );
  AOI22_X1 U19950 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_23__SCAN_IN), .ZN(n16519) );
  NAND2_X1 U19951 ( .A1(n20245), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16518) );
  NAND3_X1 U19952 ( .A1(n16520), .A2(n16519), .A3(n16518), .ZN(n16525) );
  OR2_X1 U19953 ( .A1(n16521), .A2(n16522), .ZN(n16523) );
  NAND2_X1 U19954 ( .A1(n16498), .A2(n16523), .ZN(n17199) );
  NOR2_X1 U19955 ( .A1(n17199), .A2(n20251), .ZN(n16524) );
  AOI211_X1 U19956 ( .C1(n20246), .C2(n16526), .A(n16525), .B(n16524), .ZN(
        n16527) );
  OAI21_X1 U19957 ( .B1(n16528), .B2(n20267), .A(n16527), .ZN(P2_U2832) );
  OAI21_X1 U19958 ( .B1(n13458), .B2(n16529), .A(n16512), .ZN(n17209) );
  INV_X1 U19959 ( .A(n16530), .ZN(n16532) );
  INV_X1 U19960 ( .A(n13449), .ZN(n16531) );
  AOI21_X1 U19961 ( .B1(n16532), .B2(n16531), .A(n16521), .ZN(n17218) );
  NOR2_X1 U19962 ( .A1(n16533), .A2(n20260), .ZN(n16541) );
  INV_X1 U19963 ( .A(n16939), .ZN(n16534) );
  AOI21_X1 U19964 ( .B1(n16535), .B2(n16534), .A(n20933), .ZN(n16536) );
  OAI21_X1 U19965 ( .B1(n16678), .B2(n16536), .A(n16515), .ZN(n16539) );
  AOI22_X1 U19966 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_22__SCAN_IN), .ZN(n16538) );
  NAND2_X1 U19967 ( .A1(n20245), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16537) );
  NAND3_X1 U19968 ( .A1(n16539), .A2(n16538), .A3(n16537), .ZN(n16540) );
  AOI211_X1 U19969 ( .C1(n17218), .C2(n20269), .A(n16541), .B(n16540), .ZN(
        n16542) );
  OAI21_X1 U19970 ( .B1(n17209), .B2(n20267), .A(n16542), .ZN(P2_U2833) );
  AOI22_X1 U19971 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_21__SCAN_IN), .ZN(n16543) );
  OAI21_X1 U19972 ( .B1(n20266), .B2(n16544), .A(n16543), .ZN(n16550) );
  INV_X1 U19973 ( .A(n16546), .ZN(n16545) );
  OAI21_X1 U19974 ( .B1(n16545), .B2(n20933), .A(n15158), .ZN(n16548) );
  NOR2_X1 U19975 ( .A1(n16688), .A2(n16546), .ZN(n16555) );
  MUX2_X1 U19976 ( .A(n16548), .B(n16555), .S(n16547), .Z(n16549) );
  AOI211_X1 U19977 ( .C1(n20246), .C2(n16551), .A(n16550), .B(n16549), .ZN(
        n16553) );
  NAND2_X1 U19978 ( .A1(n16826), .A2(n20235), .ZN(n16552) );
  OAI211_X1 U19979 ( .C1(n16738), .C2(n20251), .A(n16553), .B(n16552), .ZN(
        P2_U2834) );
  NAND2_X1 U19980 ( .A1(n20132), .A2(n16556), .ZN(n16554) );
  NAND2_X1 U19981 ( .A1(n16555), .A2(n16554), .ZN(n16560) );
  AOI22_X1 U19982 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n20264), .B2(P2_REIP_REG_20__SCAN_IN), .ZN(n16559) );
  NAND2_X1 U19983 ( .A1(n16678), .A2(n16556), .ZN(n16558) );
  NAND2_X1 U19984 ( .A1(n20245), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16557) );
  NAND4_X1 U19985 ( .A1(n16560), .A2(n16559), .A3(n16558), .A4(n16557), .ZN(
        n16562) );
  INV_X1 U19986 ( .A(n16948), .ZN(n16742) );
  NOR2_X1 U19987 ( .A1(n16742), .A2(n20251), .ZN(n16561) );
  AOI211_X1 U19988 ( .C1(n20246), .C2(n16563), .A(n16562), .B(n16561), .ZN(
        n16564) );
  OAI21_X1 U19989 ( .B1(n16839), .B2(n20267), .A(n16564), .ZN(P2_U2835) );
  NOR2_X1 U19990 ( .A1(n10238), .A2(n20166), .ZN(n16565) );
  XNOR2_X1 U19991 ( .A(n16565), .B(n16967), .ZN(n16571) );
  NAND2_X1 U19992 ( .A1(n20255), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16566) );
  OAI211_X1 U19993 ( .C1(n20979), .C2(n20249), .A(n16566), .B(n20169), .ZN(
        n16567) );
  AOI21_X1 U19994 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n20245), .A(n16567), .ZN(
        n16568) );
  OAI21_X1 U19995 ( .B1(n16569), .B2(n20260), .A(n16568), .ZN(n16570) );
  AOI21_X1 U19996 ( .B1(n16571), .B2(n20276), .A(n16570), .ZN(n16573) );
  NAND2_X1 U19997 ( .A1(n16856), .A2(n20235), .ZN(n16572) );
  OAI211_X1 U19998 ( .C1(n20251), .C2(n16964), .A(n16573), .B(n16572), .ZN(
        P2_U2838) );
  INV_X1 U19999 ( .A(n17247), .ZN(n16583) );
  OAI21_X1 U20000 ( .B1(n20249), .B2(n20975), .A(n20169), .ZN(n16575) );
  NOR2_X1 U20001 ( .A1(n20266), .A2(n12913), .ZN(n16574) );
  AOI211_X1 U20002 ( .C1(n20255), .C2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16575), .B(n16574), .ZN(n16576) );
  OAI21_X1 U20003 ( .B1(n16577), .B2(n20260), .A(n16576), .ZN(n16582) );
  INV_X1 U20004 ( .A(n16578), .ZN(n20183) );
  NOR2_X1 U20005 ( .A1(n16688), .A2(n20183), .ZN(n16580) );
  OAI21_X1 U20006 ( .B1(n16578), .B2(n20933), .A(n15158), .ZN(n16579) );
  MUX2_X1 U20007 ( .A(n16580), .B(n16579), .S(n16990), .Z(n16581) );
  AOI211_X1 U20008 ( .C1(n20269), .C2(n16583), .A(n16582), .B(n16581), .ZN(
        n16584) );
  OAI21_X1 U20009 ( .B1(n17253), .B2(n20267), .A(n16584), .ZN(P2_U2840) );
  NOR2_X1 U20010 ( .A1(n10238), .A2(n20198), .ZN(n16585) );
  XOR2_X1 U20011 ( .A(n17012), .B(n16585), .Z(n16593) );
  OAI21_X1 U20012 ( .B1(n21471), .B2(n20249), .A(n12586), .ZN(n16586) );
  AOI21_X1 U20013 ( .B1(n20255), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16586), .ZN(n16587) );
  OAI21_X1 U20014 ( .B1(n20266), .B2(n12861), .A(n16587), .ZN(n16589) );
  NOR2_X1 U20015 ( .A1(n17281), .A2(n20251), .ZN(n16588) );
  AOI211_X1 U20016 ( .C1(n20246), .C2(n16590), .A(n16589), .B(n16588), .ZN(
        n16592) );
  NAND2_X1 U20017 ( .A1(n17284), .A2(n20235), .ZN(n16591) );
  OAI211_X1 U20018 ( .C1(n16593), .C2(n20933), .A(n16592), .B(n16591), .ZN(
        P2_U2842) );
  NAND2_X1 U20019 ( .A1(n16651), .A2(n20215), .ZN(n16596) );
  NOR2_X1 U20020 ( .A1(n20215), .A2(n20933), .ZN(n16594) );
  NOR2_X1 U20021 ( .A1(n16678), .A2(n16594), .ZN(n16595) );
  MUX2_X1 U20022 ( .A(n16596), .B(n16595), .S(n17038), .Z(n16603) );
  INV_X1 U20023 ( .A(n17040), .ZN(n17304) );
  AOI21_X1 U20024 ( .B1(n20264), .B2(P2_REIP_REG_11__SCAN_IN), .A(n20263), 
        .ZN(n16597) );
  OAI21_X1 U20025 ( .B1(n20258), .B2(n17036), .A(n16597), .ZN(n16598) );
  AOI21_X1 U20026 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n20245), .A(n16598), .ZN(
        n16599) );
  OAI21_X1 U20027 ( .B1(n16600), .B2(n20260), .A(n16599), .ZN(n16601) );
  AOI21_X1 U20028 ( .B1(n17304), .B2(n20269), .A(n16601), .ZN(n16602) );
  OAI211_X1 U20029 ( .C1(n20267), .C2(n17308), .A(n16603), .B(n16602), .ZN(
        P2_U2844) );
  NOR2_X1 U20030 ( .A1(n10238), .A2(n20227), .ZN(n16604) );
  XOR2_X1 U20031 ( .A(n17062), .B(n16604), .Z(n16612) );
  OAI21_X1 U20032 ( .B1(n20966), .B2(n20249), .A(n12586), .ZN(n16605) );
  AOI21_X1 U20033 ( .B1(n20255), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16605), .ZN(n16606) );
  OAI21_X1 U20034 ( .B1(n20266), .B2(n10375), .A(n16606), .ZN(n16607) );
  AOI21_X1 U20035 ( .B1(n16608), .B2(n20246), .A(n16607), .ZN(n16609) );
  OAI21_X1 U20036 ( .B1(n17324), .B2(n20251), .A(n16609), .ZN(n16610) );
  AOI21_X1 U20037 ( .B1(n20235), .B2(n17331), .A(n16610), .ZN(n16611) );
  OAI21_X1 U20038 ( .B1(n16612), .B2(n20933), .A(n16611), .ZN(P2_U2846) );
  NAND2_X1 U20039 ( .A1(n16651), .A2(n16613), .ZN(n16616) );
  NOR2_X1 U20040 ( .A1(n16613), .A2(n20933), .ZN(n16614) );
  NOR2_X1 U20041 ( .A1(n16678), .A2(n16614), .ZN(n16615) );
  MUX2_X1 U20042 ( .A(n16616), .B(n16615), .S(n17096), .Z(n16624) );
  OAI21_X1 U20043 ( .B1(n20961), .B2(n20249), .A(n12586), .ZN(n16618) );
  NOR2_X1 U20044 ( .A1(n20258), .A2(n17094), .ZN(n16617) );
  AOI211_X1 U20045 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n20245), .A(n16618), .B(
        n16617), .ZN(n16619) );
  OAI21_X1 U20046 ( .B1(n16620), .B2(n20260), .A(n16619), .ZN(n16621) );
  AOI21_X1 U20047 ( .B1(n16622), .B2(n20269), .A(n16621), .ZN(n16623) );
  OAI211_X1 U20048 ( .C1(n20267), .C2(n16625), .A(n16624), .B(n16623), .ZN(
        P2_U2849) );
  NOR2_X1 U20049 ( .A1(n10238), .A2(n20274), .ZN(n16627) );
  XOR2_X1 U20050 ( .A(n17712), .B(n16627), .Z(n16635) );
  OAI21_X1 U20051 ( .B1(n12494), .B2(n20249), .A(n12586), .ZN(n16629) );
  INV_X1 U20052 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17724) );
  NOR2_X1 U20053 ( .A1(n20258), .A2(n17724), .ZN(n16628) );
  AOI211_X1 U20054 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n20245), .A(n16629), .B(
        n16628), .ZN(n16630) );
  OAI21_X1 U20055 ( .B1(n16631), .B2(n20260), .A(n16630), .ZN(n16633) );
  NOR2_X1 U20056 ( .A1(n17373), .A2(n20267), .ZN(n16632) );
  AOI211_X1 U20057 ( .C1(n17715), .C2(n20269), .A(n16633), .B(n16632), .ZN(
        n16634) );
  OAI21_X1 U20058 ( .B1(n16635), .B2(n20933), .A(n16634), .ZN(P2_U2850) );
  AND2_X1 U20059 ( .A1(n16637), .A2(n20276), .ZN(n16636) );
  NOR2_X1 U20060 ( .A1(n16678), .A2(n16636), .ZN(n16640) );
  INV_X1 U20061 ( .A(n16637), .ZN(n16638) );
  NAND2_X1 U20062 ( .A1(n16651), .A2(n16638), .ZN(n16639) );
  MUX2_X1 U20063 ( .A(n16640), .B(n16639), .S(n17124), .Z(n16648) );
  NOR2_X1 U20064 ( .A1(n16641), .A2(n20260), .ZN(n16643) );
  INV_X1 U20065 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17128) );
  OAI22_X1 U20066 ( .A1(n20258), .A2(n17128), .B1(n12152), .B2(n20249), .ZN(
        n16642) );
  AOI211_X1 U20067 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n20245), .A(n16643), .B(
        n16642), .ZN(n16644) );
  OAI21_X1 U20068 ( .B1(n16645), .B2(n20267), .A(n16644), .ZN(n16646) );
  AOI21_X1 U20069 ( .B1(n13953), .B2(n20269), .A(n16646), .ZN(n16647) );
  OAI211_X1 U20070 ( .C1(n20422), .C2(n16664), .A(n16648), .B(n16647), .ZN(
        P2_U2852) );
  AND2_X1 U20071 ( .A1(n16667), .A2(n20276), .ZN(n16649) );
  NOR2_X1 U20072 ( .A1(n16678), .A2(n16649), .ZN(n16654) );
  INV_X1 U20073 ( .A(n16667), .ZN(n16650) );
  NAND2_X1 U20074 ( .A1(n16651), .A2(n16650), .ZN(n16653) );
  MUX2_X1 U20075 ( .A(n16654), .B(n16653), .S(n16652), .Z(n16663) );
  NAND2_X1 U20076 ( .A1(n16655), .A2(n20235), .ZN(n16658) );
  OAI22_X1 U20077 ( .A1(n13644), .A2(n20258), .B1(n20959), .B2(n20249), .ZN(
        n16656) );
  AOI21_X1 U20078 ( .B1(n20245), .B2(P2_EBX_REG_2__SCAN_IN), .A(n16656), .ZN(
        n16657) );
  OAI211_X1 U20079 ( .C1(n20260), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        n16660) );
  AOI21_X1 U20080 ( .B1(n16661), .B2(n20269), .A(n16660), .ZN(n16662) );
  OAI211_X1 U20081 ( .C1(n16664), .C2(n21036), .A(n16663), .B(n16662), .ZN(
        P2_U2853) );
  AND2_X1 U20082 ( .A1(n16665), .A2(n17407), .ZN(n16666) );
  NOR2_X1 U20083 ( .A1(n16667), .A2(n16666), .ZN(n16668) );
  NAND2_X1 U20084 ( .A1(n15144), .A2(n16668), .ZN(n17416) );
  NAND2_X1 U20085 ( .A1(n16678), .A2(n15098), .ZN(n16677) );
  NAND2_X1 U20086 ( .A1(n20245), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U20087 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20255), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n20264), .ZN(n16669) );
  OAI211_X1 U20088 ( .C1(n20260), .C2(n16671), .A(n16670), .B(n16669), .ZN(
        n16672) );
  AOI21_X1 U20089 ( .B1(n20235), .B2(n21047), .A(n16672), .ZN(n16673) );
  OAI21_X1 U20090 ( .B1(n16674), .B2(n20251), .A(n16673), .ZN(n16675) );
  AOI21_X1 U20091 ( .B1(n21043), .B2(n20270), .A(n16675), .ZN(n16676) );
  OAI211_X1 U20092 ( .C1(n17416), .C2(n20933), .A(n16677), .B(n16676), .ZN(
        P2_U2854) );
  INV_X1 U20093 ( .A(n17407), .ZN(n16689) );
  OAI21_X1 U20094 ( .B1(n16678), .B2(n20255), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16687) );
  INV_X1 U20095 ( .A(n16679), .ZN(n16680) );
  OAI22_X1 U20096 ( .A1(n20123), .A2(n20249), .B1(n20260), .B2(n16680), .ZN(
        n16682) );
  NOR2_X1 U20097 ( .A1(n20266), .A2(n13642), .ZN(n16681) );
  AOI211_X1 U20098 ( .C1(n17394), .C2(n20235), .A(n16682), .B(n16681), .ZN(
        n16683) );
  OAI21_X1 U20099 ( .B1(n16684), .B2(n20251), .A(n16683), .ZN(n16685) );
  AOI21_X1 U20100 ( .B1(n20421), .B2(n20270), .A(n16685), .ZN(n16686) );
  OAI211_X1 U20101 ( .C1(n16689), .C2(n16688), .A(n16687), .B(n16686), .ZN(
        P2_U2855) );
  INV_X1 U20102 ( .A(n16690), .ZN(n16695) );
  NAND2_X1 U20103 ( .A1(n16692), .A2(n16691), .ZN(n16768) );
  NAND3_X1 U20104 ( .A1(n9777), .A2(n20288), .A3(n16768), .ZN(n16694) );
  NAND2_X1 U20105 ( .A1(n16764), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16693) );
  OAI211_X1 U20106 ( .C1(n16695), .C2(n16764), .A(n16694), .B(n16693), .ZN(
        P2_U2858) );
  NAND2_X1 U20107 ( .A1(n14905), .A2(n16696), .ZN(n16698) );
  XNOR2_X1 U20108 ( .A(n16698), .B(n16697), .ZN(n16783) );
  NOR2_X1 U20109 ( .A1(n17142), .A2(n16764), .ZN(n16699) );
  AOI21_X1 U20110 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16764), .A(n16699), .ZN(
        n16700) );
  OAI21_X1 U20111 ( .B1(n16783), .B2(n20283), .A(n16700), .ZN(P2_U2859) );
  AOI21_X1 U20112 ( .B1(n16703), .B2(n16702), .A(n16701), .ZN(n16784) );
  NAND2_X1 U20113 ( .A1(n16784), .A2(n20288), .ZN(n16705) );
  NAND2_X1 U20114 ( .A1(n16764), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16704) );
  OAI211_X1 U20115 ( .C1(n17159), .C2(n16764), .A(n16705), .B(n16704), .ZN(
        P2_U2860) );
  NAND2_X1 U20116 ( .A1(n16706), .A2(n16716), .ZN(n16715) );
  NAND2_X1 U20117 ( .A1(n16715), .A2(n16707), .ZN(n16712) );
  NOR2_X1 U20118 ( .A1(n16708), .A2(n21078), .ZN(n16709) );
  XNOR2_X1 U20119 ( .A(n16710), .B(n16709), .ZN(n16711) );
  XNOR2_X1 U20120 ( .A(n16712), .B(n16711), .ZN(n16797) );
  NOR2_X1 U20121 ( .A1(n16899), .A2(n16764), .ZN(n16713) );
  AOI21_X1 U20122 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16764), .A(n16713), .ZN(
        n16714) );
  OAI21_X1 U20123 ( .B1(n16797), .B2(n20283), .A(n16714), .ZN(P2_U2861) );
  OAI21_X1 U20124 ( .B1(n16706), .B2(n16716), .A(n16715), .ZN(n16804) );
  NAND2_X1 U20125 ( .A1(n16764), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16718) );
  NAND2_X1 U20126 ( .A1(n17173), .A2(n20291), .ZN(n16717) );
  OAI211_X1 U20127 ( .C1(n16804), .C2(n20283), .A(n16718), .B(n16717), .ZN(
        P2_U2862) );
  AOI21_X1 U20128 ( .B1(n16720), .B2(n16719), .A(n9805), .ZN(n16721) );
  XOR2_X1 U20129 ( .A(n16722), .B(n16721), .Z(n16810) );
  INV_X1 U20130 ( .A(n16918), .ZN(n17183) );
  NOR2_X1 U20131 ( .A1(n17183), .A2(n16764), .ZN(n16723) );
  AOI21_X1 U20132 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16764), .A(n16723), .ZN(
        n16724) );
  OAI21_X1 U20133 ( .B1(n16810), .B2(n20283), .A(n16724), .ZN(P2_U2863) );
  AOI21_X1 U20134 ( .B1(n16727), .B2(n16726), .A(n16725), .ZN(n16811) );
  NAND2_X1 U20135 ( .A1(n16811), .A2(n20288), .ZN(n16729) );
  NAND2_X1 U20136 ( .A1(n16764), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16728) );
  OAI211_X1 U20137 ( .C1(n17199), .C2(n16764), .A(n16729), .B(n16728), .ZN(
        P2_U2864) );
  INV_X1 U20138 ( .A(n17218), .ZN(n16732) );
  AOI21_X1 U20139 ( .B1(n16730), .B2(n16734), .A(n14817), .ZN(n16824) );
  AOI22_X1 U20140 ( .A1(n16824), .A2(n20288), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16764), .ZN(n16731) );
  OAI21_X1 U20141 ( .B1(n16732), .B2(n16764), .A(n16731), .ZN(P2_U2865) );
  OAI21_X1 U20142 ( .B1(n16733), .B2(n16735), .A(n16734), .ZN(n16832) );
  INV_X1 U20143 ( .A(n16832), .ZN(n16736) );
  AOI22_X1 U20144 ( .A1(n16736), .A2(n20288), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16764), .ZN(n16737) );
  OAI21_X1 U20145 ( .B1(n16738), .B2(n16764), .A(n16737), .ZN(P2_U2866) );
  AOI21_X1 U20146 ( .B1(n16740), .B2(n16739), .A(n16733), .ZN(n16837) );
  AOI22_X1 U20147 ( .A1(n16837), .A2(n20288), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n16764), .ZN(n16741) );
  OAI21_X1 U20148 ( .B1(n16742), .B2(n16764), .A(n16741), .ZN(P2_U2867) );
  OR2_X1 U20149 ( .A1(n16744), .A2(n16743), .ZN(n16745) );
  NAND2_X1 U20150 ( .A1(n13291), .A2(n16745), .ZN(n20141) );
  INV_X1 U20151 ( .A(n16739), .ZN(n16747) );
  AOI21_X1 U20152 ( .B1(n16748), .B2(n16746), .A(n16747), .ZN(n16847) );
  AOI22_X1 U20153 ( .A1(n16847), .A2(n20288), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16764), .ZN(n16749) );
  OAI21_X1 U20154 ( .B1(n20141), .B2(n16764), .A(n16749), .ZN(P2_U2868) );
  OAI21_X1 U20155 ( .B1(n14740), .B2(n16750), .A(n16746), .ZN(n16751) );
  INV_X1 U20156 ( .A(n16751), .ZN(n16854) );
  AOI22_X1 U20157 ( .A1(n16854), .A2(n20288), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16764), .ZN(n16752) );
  OAI21_X1 U20158 ( .B1(n20156), .B2(n16764), .A(n16752), .ZN(P2_U2869) );
  NAND2_X1 U20159 ( .A1(n16754), .A2(n16753), .ZN(n16755) );
  NAND2_X1 U20160 ( .A1(n16756), .A2(n16755), .ZN(n20204) );
  INV_X1 U20161 ( .A(n20282), .ZN(n16759) );
  OAI21_X1 U20162 ( .B1(n16759), .B2(n16758), .A(n16757), .ZN(n16761) );
  NAND3_X1 U20163 ( .A1(n16761), .A2(n20288), .A3(n16760), .ZN(n16763) );
  NAND2_X1 U20164 ( .A1(n16764), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n16762) );
  OAI211_X1 U20165 ( .C1(n20204), .C2(n16764), .A(n16763), .B(n16762), .ZN(
        P2_U2875) );
  INV_X1 U20166 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U20167 ( .A1(n15191), .A2(n20307), .ZN(n16766) );
  AOI22_X1 U20168 ( .A1(n14507), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n20306), .ZN(n16765) );
  OAI211_X1 U20169 ( .C1(n16859), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        P2_U2888) );
  NAND3_X1 U20170 ( .A1(n9777), .A2(n20295), .A3(n16768), .ZN(n16776) );
  INV_X1 U20171 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16771) );
  AOI22_X1 U20172 ( .A1(n16858), .A2(n16769), .B1(n20306), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16770) );
  OAI21_X1 U20173 ( .B1(n16859), .B2(n16771), .A(n16770), .ZN(n16774) );
  NOR2_X1 U20174 ( .A1(n16772), .A2(n16868), .ZN(n16773) );
  AOI211_X1 U20175 ( .C1(n14507), .C2(BUF1_REG_29__SCAN_IN), .A(n16774), .B(
        n16773), .ZN(n16775) );
  NAND2_X1 U20176 ( .A1(n16776), .A2(n16775), .ZN(P2_U2890) );
  INV_X1 U20177 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16780) );
  NAND2_X1 U20178 ( .A1(n14507), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U20179 ( .A1(n16858), .A2(n16777), .B1(n20306), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16778) );
  OAI211_X1 U20180 ( .C1(n16780), .C2(n16859), .A(n16779), .B(n16778), .ZN(
        n16781) );
  AOI21_X1 U20181 ( .B1(n17145), .B2(n20307), .A(n16781), .ZN(n16782) );
  OAI21_X1 U20182 ( .B1(n16783), .B2(n20311), .A(n16782), .ZN(P2_U2891) );
  INV_X1 U20183 ( .A(n16784), .ZN(n16790) );
  AOI22_X1 U20184 ( .A1(n16858), .A2(n16785), .B1(n20306), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16786) );
  OAI21_X1 U20185 ( .B1(n16859), .B2(n17834), .A(n16786), .ZN(n16788) );
  NOR2_X1 U20186 ( .A1(n17150), .A2(n16868), .ZN(n16787) );
  AOI211_X1 U20187 ( .C1(n14507), .C2(BUF1_REG_27__SCAN_IN), .A(n16788), .B(
        n16787), .ZN(n16789) );
  OAI21_X1 U20188 ( .B1(n16790), .B2(n20311), .A(n16789), .ZN(P2_U2892) );
  AOI22_X1 U20189 ( .A1(n16858), .A2(n16791), .B1(n20306), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16792) );
  OAI21_X1 U20190 ( .B1(n16859), .B2(n17831), .A(n16792), .ZN(n16795) );
  NOR2_X1 U20191 ( .A1(n16793), .A2(n16868), .ZN(n16794) );
  AOI211_X1 U20192 ( .C1(n14507), .C2(BUF1_REG_26__SCAN_IN), .A(n16795), .B(
        n16794), .ZN(n16796) );
  OAI21_X1 U20193 ( .B1(n16797), .B2(n20311), .A(n16796), .ZN(P2_U2893) );
  INV_X1 U20194 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U20195 ( .A1(n16858), .A2(n16798), .B1(n20306), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16799) );
  OAI21_X1 U20196 ( .B1(n16859), .B2(n16800), .A(n16799), .ZN(n16802) );
  NOR2_X1 U20197 ( .A1(n17170), .A2(n16868), .ZN(n16801) );
  AOI211_X1 U20198 ( .C1(n14507), .C2(BUF1_REG_25__SCAN_IN), .A(n16802), .B(
        n16801), .ZN(n16803) );
  OAI21_X1 U20199 ( .B1(n16804), .B2(n20311), .A(n16803), .ZN(P2_U2894) );
  NAND2_X1 U20200 ( .A1(n14507), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16807) );
  AOI22_X1 U20201 ( .A1(n16858), .A2(n16805), .B1(n20306), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16806) );
  OAI211_X1 U20202 ( .C1(n16859), .C2(n17829), .A(n16807), .B(n16806), .ZN(
        n16808) );
  AOI21_X1 U20203 ( .B1(n17186), .B2(n20307), .A(n16808), .ZN(n16809) );
  OAI21_X1 U20204 ( .B1(n16810), .B2(n20311), .A(n16809), .ZN(P2_U2895) );
  INV_X1 U20205 ( .A(n16811), .ZN(n16818) );
  INV_X1 U20206 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U20207 ( .A1(n14507), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16814) );
  AOI22_X1 U20208 ( .A1(n16858), .A2(n16812), .B1(n20306), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16813) );
  OAI211_X1 U20209 ( .C1(n16815), .C2(n16859), .A(n16814), .B(n16813), .ZN(
        n16816) );
  AOI21_X1 U20210 ( .B1(n17204), .B2(n20307), .A(n16816), .ZN(n16817) );
  OAI21_X1 U20211 ( .B1(n20311), .B2(n16818), .A(n16817), .ZN(P2_U2896) );
  INV_X1 U20212 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U20213 ( .A1(n14507), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U20214 ( .A1(n16858), .A2(n16819), .B1(n20306), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16820) );
  OAI211_X1 U20215 ( .C1(n16859), .C2(n16822), .A(n16821), .B(n16820), .ZN(
        n16823) );
  AOI21_X1 U20216 ( .B1(n16824), .B2(n20295), .A(n16823), .ZN(n16825) );
  OAI21_X1 U20217 ( .B1(n17209), .B2(n16868), .A(n16825), .ZN(P2_U2897) );
  NAND2_X1 U20218 ( .A1(n16826), .A2(n20307), .ZN(n16831) );
  INV_X1 U20219 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20220 ( .A1(n16858), .A2(n20396), .B1(n20306), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16827) );
  OAI21_X1 U20221 ( .B1(n16859), .B2(n16828), .A(n16827), .ZN(n16829) );
  AOI21_X1 U20222 ( .B1(n14507), .B2(BUF1_REG_21__SCAN_IN), .A(n16829), .ZN(
        n16830) );
  OAI211_X1 U20223 ( .C1(n20311), .C2(n16832), .A(n16831), .B(n16830), .ZN(
        P2_U2898) );
  NAND2_X1 U20224 ( .A1(n14507), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20225 ( .A1(n16858), .A2(n16833), .B1(n20306), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16834) );
  OAI211_X1 U20226 ( .C1(n16859), .C2(n21470), .A(n16835), .B(n16834), .ZN(
        n16836) );
  AOI21_X1 U20227 ( .B1(n16837), .B2(n20295), .A(n16836), .ZN(n16838) );
  OAI21_X1 U20228 ( .B1(n16839), .B2(n16868), .A(n16838), .ZN(P2_U2899) );
  XNOR2_X1 U20229 ( .A(n16841), .B(n16840), .ZN(n20140) );
  INV_X1 U20230 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16845) );
  NAND2_X1 U20231 ( .A1(n14507), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20232 ( .A1(n16858), .A2(n16842), .B1(n20306), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16843) );
  OAI211_X1 U20233 ( .C1(n16859), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        n16846) );
  AOI21_X1 U20234 ( .B1(n16847), .B2(n20295), .A(n16846), .ZN(n16848) );
  OAI21_X1 U20235 ( .B1(n20140), .B2(n16868), .A(n16848), .ZN(P2_U2900) );
  INV_X1 U20236 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16852) );
  NAND2_X1 U20237 ( .A1(n14507), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U20238 ( .A1(n16858), .A2(n16849), .B1(n20306), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16850) );
  OAI211_X1 U20239 ( .C1(n16859), .C2(n16852), .A(n16851), .B(n16850), .ZN(
        n16853) );
  AOI21_X1 U20240 ( .B1(n16854), .B2(n20295), .A(n16853), .ZN(n16855) );
  OAI21_X1 U20241 ( .B1(n20157), .B2(n16868), .A(n16855), .ZN(P2_U2901) );
  INV_X1 U20242 ( .A(n16856), .ZN(n16869) );
  INV_X1 U20243 ( .A(n14507), .ZN(n16864) );
  AOI22_X1 U20244 ( .A1(n16858), .A2(n16857), .B1(n20306), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16862) );
  INV_X1 U20245 ( .A(n16859), .ZN(n16860) );
  NAND2_X1 U20246 ( .A1(n16860), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16861) );
  OAI211_X1 U20247 ( .C1(n16864), .C2(n16863), .A(n16862), .B(n16861), .ZN(
        n16865) );
  AOI21_X1 U20248 ( .B1(n16866), .B2(n20295), .A(n16865), .ZN(n16867) );
  OAI21_X1 U20249 ( .B1(n16869), .B2(n16868), .A(n16867), .ZN(P2_U2902) );
  XNOR2_X1 U20250 ( .A(n16870), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17149) );
  OAI21_X1 U20251 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n12822), .ZN(n16873) );
  XNOR2_X1 U20252 ( .A(n16874), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16875) );
  NAND2_X1 U20253 ( .A1(n20263), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n17139) );
  NAND2_X1 U20254 ( .A1(n17109), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16876) );
  OAI211_X1 U20255 ( .C1(n16877), .C2(n17112), .A(n17139), .B(n16876), .ZN(
        n16878) );
  INV_X1 U20256 ( .A(n16878), .ZN(n16879) );
  OAI21_X1 U20257 ( .B1(n17116), .B2(n17149), .A(n16881), .ZN(P2_U2986) );
  INV_X1 U20258 ( .A(n16882), .ZN(n16883) );
  NOR2_X1 U20259 ( .A1(n16884), .A2(n16883), .ZN(n16887) );
  XNOR2_X1 U20260 ( .A(n16885), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16886) );
  XNOR2_X1 U20261 ( .A(n16887), .B(n16886), .ZN(n17163) );
  INV_X1 U20262 ( .A(n16888), .ZN(n16891) );
  NAND2_X1 U20263 ( .A1(n20263), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20264 ( .B1(n17723), .B2(n16889), .A(n17155), .ZN(n16890) );
  AOI21_X1 U20265 ( .B1(n16891), .B2(n17714), .A(n16890), .ZN(n16892) );
  OAI21_X1 U20266 ( .B1(n17159), .B2(n17098), .A(n16892), .ZN(n16893) );
  OAI21_X1 U20267 ( .B1(n17723), .B2(n16895), .A(n16894), .ZN(n16896) );
  AOI21_X1 U20268 ( .B1(n16897), .B2(n17714), .A(n16896), .ZN(n16898) );
  OAI21_X1 U20269 ( .B1(n16899), .B2(n17098), .A(n16898), .ZN(n16900) );
  AOI21_X1 U20270 ( .B1(n16901), .B2(n17718), .A(n16900), .ZN(n16902) );
  OAI21_X1 U20271 ( .B1(n16903), .B2(n17136), .A(n16902), .ZN(P2_U2988) );
  NAND2_X1 U20272 ( .A1(n16905), .A2(n16904), .ZN(n16906) );
  XNOR2_X1 U20273 ( .A(n16907), .B(n16906), .ZN(n17178) );
  NOR2_X1 U20274 ( .A1(n12586), .A2(n20995), .ZN(n17165) );
  AOI21_X1 U20275 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17165), .ZN(n16908) );
  OAI21_X1 U20276 ( .B1(n16909), .B2(n17112), .A(n16908), .ZN(n16910) );
  AOI21_X1 U20277 ( .B1(n17173), .B2(n17716), .A(n16910), .ZN(n16912) );
  NAND3_X1 U20278 ( .A1(n17175), .A2(n17718), .A3(n17174), .ZN(n16911) );
  OAI211_X1 U20279 ( .C1(n17136), .C2(n17178), .A(n16912), .B(n16911), .ZN(
        P2_U2989) );
  NAND2_X1 U20280 ( .A1(n16914), .A2(n17714), .ZN(n16915) );
  NAND2_X1 U20281 ( .A1(n20263), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n17179) );
  OAI211_X1 U20282 ( .C1(n16916), .C2(n17723), .A(n16915), .B(n17179), .ZN(
        n16917) );
  AOI21_X1 U20283 ( .B1(n16918), .B2(n17716), .A(n16917), .ZN(n16925) );
  INV_X1 U20284 ( .A(n16919), .ZN(n16921) );
  NAND2_X1 U20285 ( .A1(n16921), .A2(n16920), .ZN(n16922) );
  XNOR2_X1 U20286 ( .A(n16923), .B(n16922), .ZN(n17187) );
  NAND2_X1 U20287 ( .A1(n17187), .A2(n17719), .ZN(n16924) );
  OAI211_X1 U20288 ( .C1(n17190), .C2(n17116), .A(n16925), .B(n16924), .ZN(
        P2_U2990) );
  NOR2_X1 U20289 ( .A1(n13447), .A2(n17214), .ZN(n16937) );
  OAI21_X1 U20290 ( .B1(n16937), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10131), .ZN(n17206) );
  NAND2_X1 U20291 ( .A1(n20263), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U20292 ( .B1(n17723), .B2(n16926), .A(n17195), .ZN(n16927) );
  AOI21_X1 U20293 ( .B1(n16928), .B2(n17714), .A(n16927), .ZN(n16932) );
  INV_X1 U20294 ( .A(n16929), .ZN(n17200) );
  NOR2_X1 U20295 ( .A1(n16931), .A2(n16930), .ZN(n17201) );
  NAND2_X1 U20296 ( .A1(n16934), .A2(n16933), .ZN(n16936) );
  XOR2_X1 U20297 ( .A(n16936), .B(n16935), .Z(n17221) );
  INV_X1 U20298 ( .A(n16937), .ZN(n17208) );
  NAND2_X1 U20299 ( .A1(n13447), .A2(n17214), .ZN(n17207) );
  NAND3_X1 U20300 ( .A1(n17208), .A2(n17718), .A3(n17207), .ZN(n16942) );
  NOR2_X1 U20301 ( .A1(n12586), .A2(n20989), .ZN(n17211) );
  AOI21_X1 U20302 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17211), .ZN(n16938) );
  OAI21_X1 U20303 ( .B1(n16939), .B2(n17112), .A(n16938), .ZN(n16940) );
  AOI21_X1 U20304 ( .B1(n17218), .B2(n17716), .A(n16940), .ZN(n16941) );
  OAI211_X1 U20305 ( .C1(n17221), .C2(n17136), .A(n16942), .B(n16941), .ZN(
        P2_U2992) );
  NAND2_X1 U20306 ( .A1(n16943), .A2(n17719), .ZN(n16950) );
  AOI21_X1 U20307 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16944), .ZN(n16945) );
  OAI21_X1 U20308 ( .B1(n16946), .B2(n17112), .A(n16945), .ZN(n16947) );
  AOI21_X1 U20309 ( .B1(n16948), .B2(n17716), .A(n16947), .ZN(n16949) );
  OAI211_X1 U20310 ( .C1(n17116), .C2(n16951), .A(n16950), .B(n16949), .ZN(
        P2_U2994) );
  XNOR2_X1 U20311 ( .A(n16953), .B(n16952), .ZN(n17232) );
  NAND2_X1 U20312 ( .A1(n16956), .A2(n16955), .ZN(n16957) );
  XNOR2_X1 U20313 ( .A(n16958), .B(n16957), .ZN(n17230) );
  NAND2_X1 U20314 ( .A1(n20263), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17223) );
  OAI21_X1 U20315 ( .B1(n17723), .B2(n20137), .A(n17223), .ZN(n16959) );
  AOI21_X1 U20316 ( .B1(n20130), .B2(n17714), .A(n16959), .ZN(n16960) );
  OAI21_X1 U20317 ( .B1(n20141), .B2(n17098), .A(n16960), .ZN(n16961) );
  AOI21_X1 U20318 ( .B1(n17230), .B2(n17719), .A(n16961), .ZN(n16962) );
  OAI21_X1 U20319 ( .B1(n17116), .B2(n17232), .A(n16962), .ZN(P2_U2995) );
  XNOR2_X1 U20320 ( .A(n16963), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16972) );
  NOR2_X1 U20321 ( .A1(n16964), .A2(n17098), .ZN(n16969) );
  NAND2_X1 U20322 ( .A1(n17109), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16965) );
  OAI211_X1 U20323 ( .C1(n16967), .C2(n17112), .A(n16966), .B(n16965), .ZN(
        n16968) );
  AOI211_X1 U20324 ( .C1(n16970), .C2(n17719), .A(n16969), .B(n16968), .ZN(
        n16971) );
  OAI21_X1 U20325 ( .B1(n17116), .B2(n16972), .A(n16971), .ZN(P2_U2997) );
  XOR2_X1 U20326 ( .A(n16973), .B(n16974), .Z(n17237) );
  INV_X1 U20327 ( .A(n17237), .ZN(n16982) );
  OAI21_X1 U20328 ( .B1(n17239), .B2(n17250), .A(n17243), .ZN(n16975) );
  NAND3_X1 U20329 ( .A1(n16976), .A2(n17718), .A3(n16975), .ZN(n16981) );
  INV_X1 U20330 ( .A(n17235), .ZN(n20175) );
  NAND2_X1 U20331 ( .A1(n20263), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U20332 ( .A1(n17109), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16977) );
  OAI211_X1 U20333 ( .C1(n17112), .C2(n16978), .A(n17233), .B(n16977), .ZN(
        n16979) );
  AOI21_X1 U20334 ( .B1(n20175), .B2(n17716), .A(n16979), .ZN(n16980) );
  OAI211_X1 U20335 ( .C1(n16982), .C2(n17136), .A(n16981), .B(n16980), .ZN(
        P2_U2998) );
  XNOR2_X1 U20336 ( .A(n17239), .B(n17250), .ZN(n17257) );
  NAND2_X1 U20337 ( .A1(n16984), .A2(n16983), .ZN(n16987) );
  INV_X1 U20338 ( .A(n16985), .ZN(n16996) );
  NOR2_X1 U20339 ( .A1(n9785), .A2(n16996), .ZN(n16986) );
  XOR2_X1 U20340 ( .A(n16987), .B(n16986), .Z(n17255) );
  NAND2_X1 U20341 ( .A1(n20263), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n17245) );
  OAI21_X1 U20342 ( .B1(n17723), .B2(n16988), .A(n17245), .ZN(n16989) );
  AOI21_X1 U20343 ( .B1(n17714), .B2(n16990), .A(n16989), .ZN(n16991) );
  OAI21_X1 U20344 ( .B1(n17247), .B2(n17098), .A(n16991), .ZN(n16992) );
  AOI21_X1 U20345 ( .B1(n17255), .B2(n17719), .A(n16992), .ZN(n16993) );
  OAI21_X1 U20346 ( .B1(n17257), .B2(n17116), .A(n16993), .ZN(P2_U2999) );
  OAI21_X1 U20347 ( .B1(n16994), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17239), .ZN(n17273) );
  NOR2_X1 U20348 ( .A1(n16997), .A2(n16996), .ZN(n16998) );
  XNOR2_X1 U20349 ( .A(n16995), .B(n16998), .ZN(n17271) );
  NOR2_X1 U20350 ( .A1(n12586), .A2(n20973), .ZN(n17265) );
  NOR2_X1 U20351 ( .A1(n17112), .A2(n20182), .ZN(n16999) );
  AOI211_X1 U20352 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17109), .A(
        n17265), .B(n16999), .ZN(n17000) );
  OAI21_X1 U20353 ( .B1(n20191), .B2(n17098), .A(n17000), .ZN(n17001) );
  AOI21_X1 U20354 ( .B1(n17271), .B2(n17719), .A(n17001), .ZN(n17002) );
  OAI21_X1 U20355 ( .B1(n17273), .B2(n17116), .A(n17002), .ZN(P2_U3000) );
  INV_X1 U20356 ( .A(n16994), .ZN(n17004) );
  NAND2_X1 U20357 ( .A1(n17004), .A2(n17003), .ZN(n17288) );
  AOI21_X1 U20358 ( .B1(n17005), .B2(n17007), .A(n17006), .ZN(n17011) );
  NAND2_X1 U20359 ( .A1(n17009), .A2(n17008), .ZN(n17010) );
  XNOR2_X1 U20360 ( .A(n17011), .B(n17010), .ZN(n17285) );
  NOR2_X1 U20361 ( .A1(n12586), .A2(n21471), .ZN(n17276) );
  NOR2_X1 U20362 ( .A1(n17112), .A2(n17012), .ZN(n17013) );
  AOI211_X1 U20363 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17109), .A(
        n17276), .B(n17013), .ZN(n17014) );
  OAI21_X1 U20364 ( .B1(n17281), .B2(n17098), .A(n17014), .ZN(n17015) );
  AOI21_X1 U20365 ( .B1(n17285), .B2(n17719), .A(n17015), .ZN(n17016) );
  OAI21_X1 U20366 ( .B1(n17288), .B2(n17116), .A(n17016), .ZN(P2_U3001) );
  XNOR2_X1 U20367 ( .A(n17026), .B(n17277), .ZN(n17300) );
  NAND2_X1 U20368 ( .A1(n17005), .A2(n17017), .ZN(n17021) );
  NAND2_X1 U20369 ( .A1(n17019), .A2(n17018), .ZN(n17020) );
  XNOR2_X1 U20370 ( .A(n17021), .B(n17020), .ZN(n17297) );
  NAND2_X1 U20371 ( .A1(n20263), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U20372 ( .B1(n17723), .B2(n20202), .A(n17289), .ZN(n17022) );
  AOI21_X1 U20373 ( .B1(n17714), .B2(n10462), .A(n17022), .ZN(n17023) );
  OAI21_X1 U20374 ( .B1(n20204), .B2(n17098), .A(n17023), .ZN(n17024) );
  AOI21_X1 U20375 ( .B1(n17297), .B2(n17719), .A(n17024), .ZN(n17025) );
  OAI21_X1 U20376 ( .B1(n17300), .B2(n17116), .A(n17025), .ZN(P2_U3002) );
  NOR2_X1 U20377 ( .A1(n17056), .A2(n17319), .ZN(n17049) );
  OAI21_X1 U20378 ( .B1(n17049), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17026), .ZN(n17312) );
  NAND2_X1 U20379 ( .A1(n17027), .A2(n17028), .ZN(n17061) );
  INV_X1 U20380 ( .A(n17029), .ZN(n17059) );
  NOR2_X1 U20381 ( .A1(n17061), .A2(n17059), .ZN(n17044) );
  AOI21_X1 U20382 ( .B1(n17044), .B2(n17045), .A(n17030), .ZN(n17035) );
  INV_X1 U20383 ( .A(n17031), .ZN(n17033) );
  NOR2_X1 U20384 ( .A1(n17033), .A2(n17032), .ZN(n17034) );
  XNOR2_X1 U20385 ( .A(n17035), .B(n17034), .ZN(n17310) );
  NAND2_X1 U20386 ( .A1(n20263), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17301) );
  OAI21_X1 U20387 ( .B1(n17723), .B2(n17036), .A(n17301), .ZN(n17037) );
  AOI21_X1 U20388 ( .B1(n17714), .B2(n17038), .A(n17037), .ZN(n17039) );
  OAI21_X1 U20389 ( .B1(n17040), .B2(n17098), .A(n17039), .ZN(n17041) );
  AOI21_X1 U20390 ( .B1(n17310), .B2(n17719), .A(n17041), .ZN(n17042) );
  OAI21_X1 U20391 ( .B1(n17312), .B2(n17116), .A(n17042), .ZN(P2_U3003) );
  INV_X1 U20392 ( .A(n17043), .ZN(n17058) );
  NOR2_X1 U20393 ( .A1(n17044), .A2(n17058), .ZN(n17048) );
  NAND2_X1 U20394 ( .A1(n17046), .A2(n17045), .ZN(n17047) );
  XNOR2_X1 U20395 ( .A(n17048), .B(n17047), .ZN(n17323) );
  AOI21_X1 U20396 ( .B1(n17319), .B2(n17056), .A(n17049), .ZN(n17313) );
  NAND2_X1 U20397 ( .A1(n17313), .A2(n17718), .ZN(n17055) );
  NOR2_X1 U20398 ( .A1(n14410), .A2(n17050), .ZN(n17051) );
  NOR2_X1 U20399 ( .A1(n12586), .A2(n20968), .ZN(n17314) );
  AOI21_X1 U20400 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17314), .ZN(n17052) );
  OAI21_X1 U20401 ( .B1(n17112), .B2(n20211), .A(n17052), .ZN(n17053) );
  AOI21_X1 U20402 ( .B1(n10444), .B2(n17716), .A(n17053), .ZN(n17054) );
  OAI211_X1 U20403 ( .C1(n17323), .C2(n17136), .A(n17055), .B(n17054), .ZN(
        P2_U3004) );
  OAI21_X1 U20404 ( .B1(n17057), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17056), .ZN(n17337) );
  NOR2_X1 U20405 ( .A1(n17059), .A2(n17058), .ZN(n17060) );
  XNOR2_X1 U20406 ( .A(n17061), .B(n17060), .ZN(n17335) );
  NOR2_X1 U20407 ( .A1(n12586), .A2(n20966), .ZN(n17325) );
  NOR2_X1 U20408 ( .A1(n17112), .A2(n17062), .ZN(n17063) );
  AOI211_X1 U20409 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17109), .A(
        n17325), .B(n17063), .ZN(n17064) );
  OAI21_X1 U20410 ( .B1(n17324), .B2(n17098), .A(n17064), .ZN(n17065) );
  AOI21_X1 U20411 ( .B1(n17335), .B2(n17719), .A(n17065), .ZN(n17066) );
  OAI21_X1 U20412 ( .B1(n17337), .B2(n17116), .A(n17066), .ZN(P2_U3005) );
  XNOR2_X1 U20413 ( .A(n17067), .B(n17068), .ZN(n17349) );
  AOI22_X1 U20414 ( .A1(n17071), .A2(n17070), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17069), .ZN(n17087) );
  INV_X1 U20415 ( .A(n17085), .ZN(n17072) );
  OAI21_X1 U20416 ( .B1(n17087), .B2(n17072), .A(n17086), .ZN(n17076) );
  NAND2_X1 U20417 ( .A1(n17074), .A2(n17073), .ZN(n17075) );
  XNOR2_X1 U20418 ( .A(n17076), .B(n17075), .ZN(n17347) );
  NAND2_X1 U20419 ( .A1(n20237), .A2(n17716), .ZN(n17079) );
  NOR2_X1 U20420 ( .A1(n12586), .A2(n17077), .ZN(n17339) );
  AOI21_X1 U20421 ( .B1(n17109), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17339), .ZN(n17078) );
  OAI211_X1 U20422 ( .C1(n17112), .C2(n17080), .A(n17079), .B(n17078), .ZN(
        n17081) );
  AOI21_X1 U20423 ( .B1(n17347), .B2(n17719), .A(n17081), .ZN(n17082) );
  OAI21_X1 U20424 ( .B1(n17349), .B2(n17116), .A(n17082), .ZN(P2_U3006) );
  XNOR2_X1 U20425 ( .A(n17083), .B(n17084), .ZN(n17361) );
  NAND2_X1 U20426 ( .A1(n17086), .A2(n17085), .ZN(n17088) );
  XOR2_X1 U20427 ( .A(n17088), .B(n17087), .Z(n17359) );
  NAND2_X1 U20428 ( .A1(n20263), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n17351) );
  OAI21_X1 U20429 ( .B1(n17723), .B2(n17089), .A(n17351), .ZN(n17090) );
  AOI21_X1 U20430 ( .B1(n17714), .B2(n9774), .A(n17090), .ZN(n17091) );
  OAI21_X1 U20431 ( .B1(n20252), .B2(n17098), .A(n17091), .ZN(n17092) );
  AOI21_X1 U20432 ( .B1(n17359), .B2(n17719), .A(n17092), .ZN(n17093) );
  OAI21_X1 U20433 ( .B1(n17116), .B2(n17361), .A(n17093), .ZN(P2_U3007) );
  OAI22_X1 U20434 ( .A1(n17723), .A2(n17094), .B1(n20961), .B2(n20169), .ZN(
        n17095) );
  AOI21_X1 U20435 ( .B1(n17714), .B2(n17096), .A(n17095), .ZN(n17097) );
  OAI21_X1 U20436 ( .B1(n17099), .B2(n17098), .A(n17097), .ZN(n17100) );
  AOI21_X1 U20437 ( .B1(n17101), .B2(n17719), .A(n17100), .ZN(n17102) );
  OAI21_X1 U20438 ( .B1(n17103), .B2(n17116), .A(n17102), .ZN(P2_U3008) );
  XNOR2_X1 U20439 ( .A(n17105), .B(n17104), .ZN(n20361) );
  NAND2_X1 U20440 ( .A1(n17107), .A2(n17106), .ZN(n17108) );
  AND2_X1 U20441 ( .A1(n14014), .A2(n17108), .ZN(n20357) );
  AOI22_X1 U20442 ( .A1(n17109), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n20263), .ZN(n17110) );
  OAI21_X1 U20443 ( .B1(n17112), .B2(n17111), .A(n17110), .ZN(n17118) );
  XNOR2_X1 U20444 ( .A(n17114), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17115) );
  XNOR2_X1 U20445 ( .A(n17113), .B(n17115), .ZN(n20359) );
  NOR2_X1 U20446 ( .A1(n20359), .A2(n17116), .ZN(n17117) );
  AOI211_X1 U20447 ( .C1(n17716), .C2(n20357), .A(n17118), .B(n17117), .ZN(
        n17119) );
  OAI21_X1 U20448 ( .B1(n17136), .B2(n20361), .A(n17119), .ZN(P2_U3010) );
  NAND2_X1 U20449 ( .A1(n17121), .A2(n17120), .ZN(n17123) );
  XNOR2_X1 U20450 ( .A(n17123), .B(n17122), .ZN(n17736) );
  INV_X1 U20451 ( .A(n17124), .ZN(n17125) );
  NAND2_X1 U20452 ( .A1(n17714), .A2(n17125), .ZN(n17127) );
  NAND2_X1 U20453 ( .A1(n20263), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U20454 ( .C1(n17723), .C2(n17128), .A(n17127), .B(n17126), .ZN(
        n17129) );
  AOI21_X1 U20455 ( .B1(n13953), .B2(n17716), .A(n17129), .ZN(n17135) );
  INV_X1 U20456 ( .A(n17131), .ZN(n17133) );
  NAND2_X1 U20457 ( .A1(n17133), .A2(n17132), .ZN(n17727) );
  NAND3_X1 U20458 ( .A1(n17130), .A2(n17727), .A3(n17718), .ZN(n17134) );
  OAI211_X1 U20459 ( .C1(n17736), .C2(n17136), .A(n17135), .B(n17134), .ZN(
        P2_U3011) );
  NAND2_X1 U20460 ( .A1(n17137), .A2(n17140), .ZN(n17138) );
  OAI211_X1 U20461 ( .C1(n17141), .C2(n17140), .A(n17139), .B(n17138), .ZN(
        n17144) );
  NOR2_X1 U20462 ( .A1(n17142), .A2(n17352), .ZN(n17143) );
  AOI211_X1 U20463 ( .C1(n17145), .C2(n20355), .A(n17144), .B(n17143), .ZN(
        n17148) );
  NAND2_X1 U20464 ( .A1(n17146), .A2(n17383), .ZN(n17147) );
  OAI211_X1 U20465 ( .C1(n17149), .C2(n20358), .A(n17148), .B(n17147), .ZN(
        P2_U3018) );
  NOR2_X1 U20466 ( .A1(n17150), .A2(n17372), .ZN(n17161) );
  INV_X1 U20467 ( .A(n17151), .ZN(n17153) );
  NAND3_X1 U20468 ( .A1(n17153), .A2(n17152), .A3(n17166), .ZN(n17154) );
  NAND2_X1 U20469 ( .A1(n17155), .A2(n17154), .ZN(n17156) );
  AOI21_X1 U20470 ( .B1(n17157), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17156), .ZN(n17158) );
  OAI21_X1 U20471 ( .B1(n17159), .B2(n17352), .A(n17158), .ZN(n17160) );
  INV_X1 U20472 ( .A(n17164), .ZN(n17169) );
  AOI21_X1 U20473 ( .B1(n17168), .B2(n17166), .A(n17165), .ZN(n17167) );
  OAI21_X1 U20474 ( .B1(n17169), .B2(n17168), .A(n17167), .ZN(n17172) );
  NOR2_X1 U20475 ( .A1(n17170), .A2(n17372), .ZN(n17171) );
  AOI211_X1 U20476 ( .C1(n17173), .C2(n20356), .A(n17172), .B(n17171), .ZN(
        n17177) );
  NAND3_X1 U20477 ( .A1(n17175), .A2(n17726), .A3(n17174), .ZN(n17176) );
  OAI211_X1 U20478 ( .C1(n17178), .C2(n20360), .A(n17177), .B(n17176), .ZN(
        P2_U3021) );
  OAI211_X1 U20479 ( .C1(n17182), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        n17185) );
  NOR2_X1 U20480 ( .A1(n17183), .A2(n17352), .ZN(n17184) );
  AOI211_X1 U20481 ( .C1(n17186), .C2(n20355), .A(n17185), .B(n17184), .ZN(
        n17189) );
  NAND2_X1 U20482 ( .A1(n17187), .A2(n17383), .ZN(n17188) );
  OAI211_X1 U20483 ( .C1(n17190), .C2(n20358), .A(n17189), .B(n17188), .ZN(
        P2_U3022) );
  INV_X1 U20484 ( .A(n17191), .ZN(n17192) );
  NAND2_X1 U20485 ( .A1(n17193), .A2(n17192), .ZN(n17210) );
  OAI211_X1 U20486 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17212), .B(n17194), .ZN(
        n17196) );
  NAND2_X1 U20487 ( .A1(n17196), .A2(n17195), .ZN(n17197) );
  AOI21_X1 U20488 ( .B1(n17210), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n17197), .ZN(n17198) );
  OAI21_X1 U20489 ( .B1(n17199), .B2(n17352), .A(n17198), .ZN(n17203) );
  NOR3_X1 U20490 ( .A1(n17201), .A2(n17200), .A3(n20360), .ZN(n17202) );
  AOI211_X1 U20491 ( .C1(n20355), .C2(n17204), .A(n17203), .B(n17202), .ZN(
        n17205) );
  OAI21_X1 U20492 ( .B1(n20358), .B2(n17206), .A(n17205), .ZN(P2_U3023) );
  NAND3_X1 U20493 ( .A1(n17208), .A2(n17726), .A3(n17207), .ZN(n17220) );
  NOR2_X1 U20494 ( .A1(n17209), .A2(n17372), .ZN(n17217) );
  INV_X1 U20495 ( .A(n17210), .ZN(n17215) );
  AOI21_X1 U20496 ( .B1(n17212), .B2(n17214), .A(n17211), .ZN(n17213) );
  OAI21_X1 U20497 ( .B1(n17215), .B2(n17214), .A(n17213), .ZN(n17216) );
  AOI211_X1 U20498 ( .C1(n17218), .C2(n20356), .A(n17217), .B(n17216), .ZN(
        n17219) );
  OAI211_X1 U20499 ( .C1(n17221), .C2(n20360), .A(n17220), .B(n17219), .ZN(
        P2_U3024) );
  INV_X1 U20500 ( .A(n20141), .ZN(n17227) );
  NAND3_X1 U20501 ( .A1(n17222), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n17259), .ZN(n17224) );
  NAND2_X1 U20502 ( .A1(n17224), .A2(n17223), .ZN(n17225) );
  AOI211_X1 U20503 ( .C1(n17227), .C2(n20356), .A(n17226), .B(n17225), .ZN(
        n17228) );
  OAI21_X1 U20504 ( .B1(n20140), .B2(n17372), .A(n17228), .ZN(n17229) );
  AOI21_X1 U20505 ( .B1(n17230), .B2(n17383), .A(n17229), .ZN(n17231) );
  OAI21_X1 U20506 ( .B1(n20358), .B2(n17232), .A(n17231), .ZN(P2_U3027) );
  NAND2_X1 U20507 ( .A1(n20176), .A2(n20355), .ZN(n17234) );
  OAI211_X1 U20508 ( .C1(n17352), .C2(n17235), .A(n17234), .B(n17233), .ZN(
        n17236) );
  AOI21_X1 U20509 ( .B1(n17237), .B2(n17383), .A(n17236), .ZN(n17242) );
  OAI21_X1 U20510 ( .B1(n17239), .B2(n20358), .A(n17238), .ZN(n17240) );
  NAND3_X1 U20511 ( .A1(n17240), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n17243), .ZN(n17241) );
  OAI211_X1 U20512 ( .C1(n17244), .C2(n17243), .A(n17242), .B(n17241), .ZN(
        P2_U3030) );
  OAI21_X1 U20513 ( .B1(n17246), .B2(n17250), .A(n17245), .ZN(n17249) );
  NOR2_X1 U20514 ( .A1(n17247), .A2(n17352), .ZN(n17248) );
  AOI211_X1 U20515 ( .C1(n17251), .C2(n17250), .A(n17249), .B(n17248), .ZN(
        n17252) );
  OAI21_X1 U20516 ( .B1(n17372), .B2(n17253), .A(n17252), .ZN(n17254) );
  AOI21_X1 U20517 ( .B1(n17255), .B2(n17383), .A(n17254), .ZN(n17256) );
  OAI21_X1 U20518 ( .B1(n17257), .B2(n20358), .A(n17256), .ZN(P2_U3031) );
  NOR2_X1 U20519 ( .A1(n20190), .A2(n17372), .ZN(n17270) );
  NOR2_X1 U20520 ( .A1(n17278), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17292) );
  OAI21_X1 U20521 ( .B1(n17258), .B2(n17329), .A(n17259), .ZN(n17317) );
  NAND2_X1 U20522 ( .A1(n17259), .A2(n17305), .ZN(n17260) );
  NAND2_X1 U20523 ( .A1(n17317), .A2(n17260), .ZN(n17291) );
  NOR2_X1 U20524 ( .A1(n17292), .A2(n17291), .ZN(n17275) );
  INV_X1 U20525 ( .A(n20191), .ZN(n17266) );
  NAND2_X1 U20526 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17261) );
  OAI21_X1 U20527 ( .B1(n17262), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17261), .ZN(n17263) );
  NOR2_X1 U20528 ( .A1(n17278), .A2(n17263), .ZN(n17264) );
  AOI211_X1 U20529 ( .C1(n17266), .C2(n20356), .A(n17265), .B(n17264), .ZN(
        n17267) );
  OAI21_X1 U20530 ( .B1(n17275), .B2(n17268), .A(n17267), .ZN(n17269) );
  AOI211_X1 U20531 ( .C1(n17271), .C2(n17383), .A(n17270), .B(n17269), .ZN(
        n17272) );
  OAI21_X1 U20532 ( .B1(n17273), .B2(n20358), .A(n17272), .ZN(P2_U3032) );
  NOR2_X1 U20533 ( .A1(n17275), .A2(n17274), .ZN(n17283) );
  INV_X1 U20534 ( .A(n17276), .ZN(n17280) );
  OR3_X1 U20535 ( .A1(n17278), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n17277), .ZN(n17279) );
  OAI211_X1 U20536 ( .C1(n17281), .C2(n17352), .A(n17280), .B(n17279), .ZN(
        n17282) );
  AOI211_X1 U20537 ( .C1(n20355), .C2(n17284), .A(n17283), .B(n17282), .ZN(
        n17287) );
  NAND2_X1 U20538 ( .A1(n17285), .A2(n17383), .ZN(n17286) );
  OAI211_X1 U20539 ( .C1(n17288), .C2(n20358), .A(n17287), .B(n17286), .ZN(
        P2_U3033) );
  INV_X1 U20540 ( .A(n17289), .ZN(n17290) );
  AOI21_X1 U20541 ( .B1(n17291), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17290), .ZN(n17294) );
  INV_X1 U20542 ( .A(n17292), .ZN(n17293) );
  OAI211_X1 U20543 ( .C1(n20204), .C2(n17352), .A(n17294), .B(n17293), .ZN(
        n17296) );
  NOR2_X1 U20544 ( .A1(n20205), .A2(n17372), .ZN(n17295) );
  NOR2_X1 U20545 ( .A1(n17296), .A2(n17295), .ZN(n17299) );
  NAND2_X1 U20546 ( .A1(n17297), .A2(n17383), .ZN(n17298) );
  OAI211_X1 U20547 ( .C1(n17300), .C2(n20358), .A(n17299), .B(n17298), .ZN(
        P2_U3034) );
  OAI21_X1 U20548 ( .B1(n17317), .B2(n17302), .A(n17301), .ZN(n17303) );
  AOI21_X1 U20549 ( .B1(n17304), .B2(n20356), .A(n17303), .ZN(n17307) );
  OAI211_X1 U20550 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17320), .B(n17305), .ZN(
        n17306) );
  OAI211_X1 U20551 ( .C1(n17308), .C2(n17372), .A(n17307), .B(n17306), .ZN(
        n17309) );
  AOI21_X1 U20552 ( .B1(n17310), .B2(n17383), .A(n17309), .ZN(n17311) );
  OAI21_X1 U20553 ( .B1(n17312), .B2(n20358), .A(n17311), .ZN(P2_U3035) );
  NAND2_X1 U20554 ( .A1(n17313), .A2(n17726), .ZN(n17322) );
  AOI21_X1 U20555 ( .B1(n10444), .B2(n20356), .A(n17314), .ZN(n17316) );
  NAND2_X1 U20556 ( .A1(n20221), .A2(n20355), .ZN(n17315) );
  OAI211_X1 U20557 ( .C1(n17317), .C2(n17319), .A(n17316), .B(n17315), .ZN(
        n17318) );
  AOI21_X1 U20558 ( .B1(n17320), .B2(n17319), .A(n17318), .ZN(n17321) );
  OAI211_X1 U20559 ( .C1(n17323), .C2(n20360), .A(n17322), .B(n17321), .ZN(
        P2_U3036) );
  INV_X1 U20560 ( .A(n17324), .ZN(n17326) );
  AOI21_X1 U20561 ( .B1(n17326), .B2(n20356), .A(n17325), .ZN(n17327) );
  OAI21_X1 U20562 ( .B1(n17329), .B2(n17328), .A(n17327), .ZN(n17330) );
  AOI21_X1 U20563 ( .B1(n20355), .B2(n17331), .A(n17330), .ZN(n17332) );
  OAI21_X1 U20564 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17333), .A(
        n17332), .ZN(n17334) );
  AOI21_X1 U20565 ( .B1(n17335), .B2(n17383), .A(n17334), .ZN(n17336) );
  OAI21_X1 U20566 ( .B1(n17337), .B2(n20358), .A(n17336), .ZN(P2_U3037) );
  NAND2_X1 U20567 ( .A1(n17357), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17338) );
  OR2_X1 U20568 ( .A1(n17340), .A2(n17338), .ZN(n17354) );
  AOI21_X1 U20569 ( .B1(n17354), .B2(n17356), .A(n17341), .ZN(n17346) );
  AOI21_X1 U20570 ( .B1(n20237), .B2(n20356), .A(n17339), .ZN(n17344) );
  INV_X1 U20571 ( .A(n17340), .ZN(n17342) );
  NAND4_X1 U20572 ( .A1(n17342), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n17341), .ZN(n17343) );
  OAI211_X1 U20573 ( .C1(n17372), .C2(n20234), .A(n17344), .B(n17343), .ZN(
        n17345) );
  AOI211_X1 U20574 ( .C1(n17347), .C2(n17383), .A(n17346), .B(n17345), .ZN(
        n17348) );
  OAI21_X1 U20575 ( .B1(n17349), .B2(n20358), .A(n17348), .ZN(P2_U3038) );
  OR2_X1 U20576 ( .A1(n20250), .A2(n17372), .ZN(n17350) );
  OAI211_X1 U20577 ( .C1(n20252), .C2(n17352), .A(n17351), .B(n17350), .ZN(
        n17353) );
  INV_X1 U20578 ( .A(n17353), .ZN(n17355) );
  OAI211_X1 U20579 ( .C1(n17357), .C2(n17356), .A(n17355), .B(n17354), .ZN(
        n17358) );
  AOI21_X1 U20580 ( .B1(n17359), .B2(n17383), .A(n17358), .ZN(n17360) );
  OAI21_X1 U20581 ( .B1(n20358), .B2(n17361), .A(n17360), .ZN(P2_U3039) );
  NAND2_X1 U20582 ( .A1(n17363), .A2(n17362), .ZN(n17364) );
  XNOR2_X1 U20583 ( .A(n9781), .B(n17364), .ZN(n17717) );
  INV_X1 U20584 ( .A(n17717), .ZN(n17378) );
  XOR2_X1 U20585 ( .A(n17365), .B(n9738), .Z(n17720) );
  NAND2_X1 U20586 ( .A1(n17720), .A2(n17383), .ZN(n17377) );
  AOI21_X1 U20587 ( .B1(n20363), .B2(n17368), .A(n17367), .ZN(n17375) );
  NAND2_X1 U20588 ( .A1(n17715), .A2(n20356), .ZN(n17371) );
  NOR2_X1 U20589 ( .A1(n17369), .A2(n17730), .ZN(n20365) );
  AOI22_X1 U20590 ( .A1(n20263), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n20365), .ZN(n17370) );
  OAI211_X1 U20591 ( .C1(n17373), .C2(n17372), .A(n17371), .B(n17370), .ZN(
        n17374) );
  AOI21_X1 U20592 ( .B1(n20364), .B2(n17375), .A(n17374), .ZN(n17376) );
  OAI211_X1 U20593 ( .C1(n17378), .C2(n20358), .A(n17377), .B(n17376), .ZN(
        P2_U3041) );
  OAI211_X1 U20594 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n17380), .B(n17379), .ZN(n17389) );
  AOI22_X1 U20595 ( .A1(n17383), .A2(n17382), .B1(n17726), .B2(n17381), .ZN(
        n17388) );
  INV_X1 U20596 ( .A(n17396), .ZN(n17384) );
  AOI22_X1 U20597 ( .A1(n17384), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20355), .B2(n21047), .ZN(n17387) );
  AOI21_X1 U20598 ( .B1(n20356), .B2(n13767), .A(n17385), .ZN(n17386) );
  NAND4_X1 U20599 ( .A1(n17389), .A2(n17388), .A3(n17387), .A4(n17386), .ZN(
        P2_U3045) );
  NOR2_X1 U20600 ( .A1(n20360), .A2(n17390), .ZN(n17391) );
  AOI211_X1 U20601 ( .C1(n20356), .C2(n17393), .A(n17392), .B(n17391), .ZN(
        n17400) );
  AOI22_X1 U20602 ( .A1(n17726), .A2(n17395), .B1(n20355), .B2(n17394), .ZN(
        n17399) );
  MUX2_X1 U20603 ( .A(n17397), .B(n17396), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n17398) );
  NAND3_X1 U20604 ( .A1(n17400), .A2(n17399), .A3(n17398), .ZN(P2_U3046) );
  NAND2_X1 U20605 ( .A1(n20421), .A2(n21040), .ZN(n17402) );
  OAI211_X1 U20606 ( .C1(n20864), .C2(n17403), .A(n17402), .B(n17401), .ZN(
        n17406) );
  AOI21_X1 U20607 ( .B1(n21061), .B2(n12457), .A(n17404), .ZN(n17405) );
  MUX2_X1 U20608 ( .A(n17406), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n21051), .Z(P2_U3605) );
  MUX2_X1 U20609 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n17407), .S(
        n15144), .Z(n17415) );
  OAI222_X1 U20610 ( .A1(n21021), .A2(n13771), .B1(n17409), .B2(n17415), .C1(
        n21025), .C2(n17408), .ZN(n17414) );
  NAND2_X1 U20611 ( .A1(n17410), .A2(n20929), .ZN(n17413) );
  AOI22_X1 U20612 ( .A1(n17411), .A2(P2_FLUSH_REG_SCAN_IN), .B1(n21075), .B2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n17412) );
  NAND2_X1 U20613 ( .A1(n17413), .A2(n17412), .ZN(n17574) );
  MUX2_X1 U20614 ( .A(n17414), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n21022), .Z(P2_U3601) );
  NAND2_X1 U20615 ( .A1(n17415), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n21020) );
  OAI21_X1 U20616 ( .B1(n15144), .B2(n21596), .A(n17416), .ZN(n21017) );
  INV_X1 U20617 ( .A(n21025), .ZN(n17572) );
  AOI22_X1 U20618 ( .A1(n21043), .A2(n17418), .B1(n17572), .B2(n17417), .ZN(
        n17419) );
  OAI21_X1 U20619 ( .B1(n21020), .B2(n21017), .A(n17419), .ZN(n17420) );
  MUX2_X1 U20620 ( .A(n17420), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n21022), .Z(P2_U3600) );
  OAI22_X1 U20621 ( .A1(n20422), .A2(n21021), .B1(n17421), .B2(n21025), .ZN(
        n17422) );
  MUX2_X1 U20622 ( .A(n17422), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n21022), .Z(P2_U3596) );
  INV_X1 U20623 ( .A(n17423), .ZN(n17424) );
  XNOR2_X1 U20624 ( .A(n19174), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17427) );
  OAI211_X1 U20625 ( .C1(n17424), .C2(n17497), .A(n17427), .B(n17426), .ZN(
        n17431) );
  NAND2_X1 U20626 ( .A1(n17435), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17434) );
  NAND3_X1 U20627 ( .A1(n17426), .A2(n17425), .A3(n17434), .ZN(n17429) );
  INV_X1 U20628 ( .A(n17427), .ZN(n17428) );
  OAI211_X1 U20629 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17435), .A(
        n17429), .B(n17428), .ZN(n17430) );
  NAND2_X1 U20630 ( .A1(n17431), .A2(n17430), .ZN(n17490) );
  NAND2_X1 U20631 ( .A1(n17739), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17432) );
  XNOR2_X1 U20632 ( .A(n17432), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17488) );
  INV_X1 U20633 ( .A(n17512), .ZN(n17433) );
  NOR2_X1 U20634 ( .A1(n17433), .A2(n17476), .ZN(n17737) );
  INV_X1 U20635 ( .A(n17434), .ZN(n17482) );
  AOI21_X1 U20636 ( .B1(n17737), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n17435), .ZN(n17436) );
  AOI21_X1 U20637 ( .B1(n17737), .B2(n17482), .A(n17436), .ZN(n17486) );
  NOR2_X1 U20638 ( .A1(n17486), .A2(n19177), .ZN(n17444) );
  XOR2_X1 U20639 ( .A(n17437), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17441) );
  AND2_X1 U20640 ( .A1(n19477), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n17478) );
  AOI21_X1 U20641 ( .B1(n19124), .B2(n18132), .A(n17478), .ZN(n17440) );
  OR2_X1 U20642 ( .A1(n17438), .A2(n17437), .ZN(n17439) );
  OAI211_X1 U20643 ( .C1(n17442), .C2(n17441), .A(n17440), .B(n17439), .ZN(
        n17443) );
  AOI211_X1 U20644 ( .C1(n17488), .C2(n19220), .A(n17444), .B(n17443), .ZN(
        n17445) );
  OAI21_X1 U20645 ( .B1(n17490), .B2(n19178), .A(n17445), .ZN(P3_U2799) );
  NOR2_X1 U20646 ( .A1(n19507), .A2(n17447), .ZN(n17448) );
  NAND2_X1 U20647 ( .A1(n17448), .A2(n19134), .ZN(n17449) );
  OAI211_X1 U20648 ( .C1(n19217), .C2(n17451), .A(n17450), .B(n17449), .ZN(
        n17454) );
  OR2_X2 U20649 ( .A1(n19124), .A2(n19004), .ZN(n19190) );
  NOR2_X1 U20650 ( .A1(n18177), .A2(n17447), .ZN(n18145) );
  NAND2_X1 U20651 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18145), .ZN(
        n18120) );
  OAI21_X1 U20652 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18145), .A(
        n18120), .ZN(n18136) );
  OAI21_X1 U20653 ( .B1(n17447), .B2(n19507), .A(n19151), .ZN(n19200) );
  OAI22_X1 U20654 ( .A1(n19223), .A2(n18136), .B1(n19134), .B2(n19200), .ZN(
        n17453) );
  AOI211_X1 U20655 ( .C1(n19220), .C2(n17455), .A(n17454), .B(n17453), .ZN(
        n17456) );
  INV_X1 U20656 ( .A(n17456), .ZN(P3_U2824) );
  AOI21_X1 U20657 ( .B1(n19449), .B2(n17458), .A(n17457), .ZN(n19446) );
  INV_X1 U20658 ( .A(n19446), .ZN(n17468) );
  OAI21_X1 U20659 ( .B1(n9730), .B2(n19105), .A(n19202), .ZN(n19206) );
  NAND2_X1 U20660 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9730), .ZN(
        n18179) );
  AND2_X1 U20661 ( .A1(n17461), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18147) );
  AOI21_X1 U20662 ( .B1(n17460), .B2(n18179), .A(n18147), .ZN(n18159) );
  AOI22_X1 U20663 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19206), .B1(
        n18159), .B2(n19190), .ZN(n17467) );
  INV_X1 U20664 ( .A(n17462), .ZN(n17463) );
  XNOR2_X1 U20665 ( .A(n17464), .B(n17463), .ZN(n19442) );
  NOR3_X1 U20666 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17459), .A3(
        n19507), .ZN(n17465) );
  INV_X1 U20667 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20008) );
  NOR2_X1 U20668 ( .A1(n19428), .A2(n20008), .ZN(n19445) );
  AOI211_X1 U20669 ( .C1(n17471), .C2(n19442), .A(n17465), .B(n19445), .ZN(
        n17466) );
  OAI211_X1 U20670 ( .C1(n19210), .C2(n17468), .A(n17467), .B(n17466), .ZN(
        P3_U2826) );
  AOI22_X1 U20671 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19151), .B1(
        n19190), .B2(n18177), .ZN(n17473) );
  AOI21_X1 U20672 ( .B1(n17471), .B2(n17470), .A(n17469), .ZN(n17472) );
  OAI211_X1 U20673 ( .C1(n19210), .C2(n17474), .A(n17473), .B(n17472), .ZN(
        P3_U2829) );
  NAND2_X1 U20674 ( .A1(n19443), .A2(n18769), .ZN(n19413) );
  AOI22_X1 U20675 ( .A1(n19421), .A2(n17476), .B1(n17475), .B2(n19470), .ZN(
        n17498) );
  OAI211_X1 U20676 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17477), .A(
        n17498), .B(n19466), .ZN(n17479) );
  AOI21_X1 U20677 ( .B1(n17479), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n17478), .ZN(n17485) );
  INV_X1 U20678 ( .A(n18942), .ZN(n18934) );
  NAND2_X1 U20679 ( .A1(n18934), .A2(n17480), .ZN(n19236) );
  NOR3_X1 U20680 ( .A1(n17481), .A2(n19459), .A3(n19236), .ZN(n17492) );
  NAND3_X1 U20681 ( .A1(n17492), .A2(n17483), .A3(n17482), .ZN(n17484) );
  OAI211_X1 U20682 ( .C1(n17486), .C2(n19413), .A(n17485), .B(n17484), .ZN(
        n17487) );
  AOI21_X1 U20683 ( .B1(n17488), .B2(n19476), .A(n17487), .ZN(n17489) );
  OAI21_X1 U20684 ( .B1(n17490), .B2(n19416), .A(n17489), .ZN(P3_U2831) );
  INV_X1 U20685 ( .A(n17491), .ZN(n17503) );
  INV_X1 U20686 ( .A(n19413), .ZN(n17493) );
  AOI21_X1 U20687 ( .B1(n17512), .B2(n17493), .A(n17492), .ZN(n17494) );
  OAI21_X1 U20688 ( .B1(n17515), .B2(n19430), .A(n17494), .ZN(n17583) );
  INV_X1 U20689 ( .A(n17495), .ZN(n17500) );
  OAI22_X1 U20690 ( .A1(n17737), .A2(n19413), .B1(n17739), .B2(n19430), .ZN(
        n17496) );
  NOR2_X1 U20691 ( .A1(n19468), .A2(n17496), .ZN(n17581) );
  AOI21_X1 U20692 ( .B1(n17498), .B2(n17581), .A(n17497), .ZN(n17499) );
  OAI21_X1 U20693 ( .B1(n17503), .B2(n19416), .A(n17502), .ZN(P3_U2832) );
  INV_X1 U20694 ( .A(n17504), .ZN(n17505) );
  AOI21_X1 U20695 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n9791), .A(
        n17505), .ZN(n18923) );
  INV_X1 U20696 ( .A(n18921), .ZN(n17507) );
  OAI22_X1 U20697 ( .A1(n17516), .A2(n19459), .B1(n17507), .B2(n17506), .ZN(
        n17519) );
  INV_X1 U20698 ( .A(n17508), .ZN(n17509) );
  OAI22_X1 U20699 ( .A1(n19346), .A2(n17509), .B1(n19253), .B2(n18921), .ZN(
        n17514) );
  AOI21_X1 U20700 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n19406), .A(
        n17510), .ZN(n19258) );
  NOR2_X1 U20701 ( .A1(n19258), .A2(n19297), .ZN(n17511) );
  AOI21_X1 U20702 ( .B1(n19252), .B2(n17511), .A(n19454), .ZN(n17528) );
  NOR2_X1 U20703 ( .A1(n17528), .A2(n17530), .ZN(n19232) );
  OAI21_X1 U20704 ( .B1(n17512), .B2(n19381), .A(n19232), .ZN(n17513) );
  AOI211_X1 U20705 ( .C1(n19948), .C2(n17515), .A(n17514), .B(n17513), .ZN(
        n19226) );
  NAND2_X1 U20706 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n19226), .ZN(
        n17518) );
  NAND2_X1 U20707 ( .A1(n19477), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18932) );
  OAI21_X1 U20708 ( .B1(n19466), .B2(n17516), .A(n18932), .ZN(n17517) );
  AOI21_X1 U20709 ( .B1(n17519), .B2(n17518), .A(n17517), .ZN(n17520) );
  OAI21_X1 U20710 ( .B1(n18923), .B2(n19416), .A(n17520), .ZN(P3_U2836) );
  INV_X1 U20711 ( .A(n17521), .ZN(n17523) );
  OAI21_X1 U20712 ( .B1(n17523), .B2(n18957), .A(n17522), .ZN(n18955) );
  INV_X1 U20713 ( .A(n19267), .ZN(n17524) );
  NAND2_X1 U20714 ( .A1(n17525), .A2(n18957), .ZN(n18962) );
  NAND2_X1 U20715 ( .A1(n19477), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18949) );
  OAI21_X1 U20716 ( .B1(n17524), .B2(n18962), .A(n18949), .ZN(n17533) );
  INV_X1 U20717 ( .A(n19381), .ZN(n19332) );
  NAND2_X1 U20718 ( .A1(n17525), .A2(n19080), .ZN(n18953) );
  INV_X1 U20719 ( .A(n18954), .ZN(n17526) );
  OAI21_X1 U20720 ( .B1(n17526), .B2(n19384), .A(n19466), .ZN(n17527) );
  AOI211_X1 U20721 ( .C1(n19332), .C2(n18953), .A(n17528), .B(n17527), .ZN(
        n17531) );
  NAND2_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17531), .ZN(
        n17529) );
  OAI21_X1 U20723 ( .B1(n17530), .B2(n17529), .A(n19428), .ZN(n19251) );
  AOI211_X1 U20724 ( .C1(n19323), .C2(n17531), .A(n18957), .B(n19251), .ZN(
        n17532) );
  AOI211_X1 U20725 ( .C1(n19377), .C2(n18955), .A(n17533), .B(n17532), .ZN(
        n17534) );
  INV_X1 U20726 ( .A(n17534), .ZN(P3_U2838) );
  INV_X1 U20727 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17538) );
  NAND2_X1 U20728 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18636) );
  NAND2_X1 U20729 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18625), .ZN(n18621) );
  NAND4_X1 U20730 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17537)
         );
  NOR4_X1 U20731 ( .A1(n17538), .A2(n17924), .A3(n18400), .A4(n17537), .ZN(
        n17539) );
  NAND4_X1 U20732 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_27__SCAN_IN), .A4(n17539), .ZN(n18227) );
  NOR2_X1 U20733 ( .A1(n18228), .A2(n18227), .ZN(n18355) );
  INV_X1 U20734 ( .A(n18644), .ZN(n18651) );
  NAND2_X1 U20735 ( .A1(n18642), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17541) );
  NAND2_X1 U20736 ( .A1(n18355), .A2(n19521), .ZN(n17540) );
  OAI22_X1 U20737 ( .A1(n18355), .A2(n17541), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17540), .ZN(P3_U2672) );
  INV_X1 U20738 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18408) );
  AOI22_X1 U20739 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17543) );
  NAND2_X1 U20740 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n17542) );
  OAI211_X1 U20741 ( .C1(n18408), .C2(n9726), .A(n17543), .B(n17542), .ZN(
        n17544) );
  INV_X1 U20742 ( .A(n17544), .ZN(n17548) );
  AOI22_X1 U20743 ( .A1(n17545), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17547) );
  AOI22_X1 U20744 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11836), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17546) );
  NAND3_X1 U20745 ( .A1(n17548), .A2(n17547), .A3(n17546), .ZN(n17556) );
  AOI22_X1 U20746 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U20747 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11802), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17553) );
  AOI22_X1 U20748 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U20749 ( .A1(n17550), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17551) );
  NAND4_X1 U20750 ( .A1(n17554), .A2(n17553), .A3(n17552), .A4(n17551), .ZN(
        n17555) );
  NOR2_X1 U20751 ( .A1(n17556), .A2(n17555), .ZN(n18746) );
  INV_X1 U20752 ( .A(n18547), .ZN(n17557) );
  OAI33_X1 U20753 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18697), .A3(n18547), 
        .B1(n18050), .B2(n18648), .B3(n17557), .ZN(n17558) );
  INV_X1 U20754 ( .A(n17558), .ZN(n17559) );
  OAI21_X1 U20755 ( .B1(n18746), .B2(n18642), .A(n17559), .ZN(P3_U2690) );
  NAND2_X1 U20756 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19707) );
  AND2_X1 U20757 ( .A1(n17560), .A2(n19105), .ZN(n17562) );
  AOI221_X1 U20758 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19707), .C1(n17562), 
        .C2(n19707), .A(n17561), .ZN(n19487) );
  NOR2_X1 U20759 ( .A1(n17563), .A2(n19755), .ZN(n17564) );
  OAI21_X1 U20760 ( .B1(n17564), .B2(n19837), .A(n19488), .ZN(n19485) );
  AOI22_X1 U20761 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19487), .B1(
        n19485), .B2(n19938), .ZN(P3_U2865) );
  INV_X1 U20762 ( .A(n17565), .ZN(n17567) );
  NOR2_X1 U20763 ( .A1(n17567), .A2(n17566), .ZN(n19956) );
  NAND3_X1 U20764 ( .A1(n17569), .A2(n20103), .A3(n19956), .ZN(n17568) );
  OAI21_X1 U20765 ( .B1(n17569), .B2(n19961), .A(n17568), .ZN(P3_U3284) );
  NAND4_X1 U20766 ( .A1(n17574), .A2(n17572), .A3(n17571), .A4(n17570), .ZN(
        n17573) );
  OAI21_X1 U20767 ( .B1(n17574), .B2(n12394), .A(n17573), .ZN(P2_U3595) );
  AOI22_X1 U20768 ( .A1(n13212), .A2(n17576), .B1(n19113), .B2(n17578), .ZN(
        n17577) );
  XNOR2_X1 U20769 ( .A(n17577), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17752) );
  AOI22_X1 U20770 ( .A1(n19470), .A2(n17579), .B1(n19421), .B2(n17578), .ZN(
        n17580) );
  INV_X1 U20771 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17741) );
  AOI21_X1 U20772 ( .B1(n17581), .B2(n17580), .A(n17741), .ZN(n17582) );
  AOI21_X1 U20773 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n19477), .A(n17582), 
        .ZN(n17586) );
  NAND3_X1 U20774 ( .A1(n17584), .A2(n17741), .A3(n17583), .ZN(n17585) );
  OAI211_X1 U20775 ( .C1(n17752), .C2(n19416), .A(n17586), .B(n17585), .ZN(
        P3_U2833) );
  NOR2_X1 U20776 ( .A1(n17587), .A2(n17616), .ZN(n17624) );
  NOR2_X1 U20777 ( .A1(n17588), .A2(n21271), .ZN(n17589) );
  AND2_X1 U20778 ( .A1(n17590), .A2(n17589), .ZN(n17591) );
  NAND2_X1 U20779 ( .A1(n17591), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17595) );
  OAI22_X1 U20780 ( .A1(n17593), .A2(n17592), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17591), .ZN(n17594) );
  NAND2_X1 U20781 ( .A1(n17595), .A2(n17594), .ZN(n17598) );
  INV_X1 U20782 ( .A(n17596), .ZN(n17597) );
  AOI222_X1 U20783 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17598), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17597), .C1(n17598), 
        .C2(n17597), .ZN(n17601) );
  AOI222_X1 U20784 ( .A1(n17601), .A2(n17600), .B1(n17601), .B2(n17599), .C1(
        n17600), .C2(n17599), .ZN(n17611) );
  INV_X1 U20785 ( .A(n17602), .ZN(n17607) );
  AOI21_X1 U20786 ( .B1(n21095), .B2(n17604), .A(n17603), .ZN(n17606) );
  NOR4_X1 U20787 ( .A1(n17608), .A2(n17607), .A3(n17606), .A4(n17605), .ZN(
        n17609) );
  OAI211_X1 U20788 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n17611), .A(
        n17610), .B(n17609), .ZN(n17619) );
  INV_X1 U20789 ( .A(n17619), .ZN(n17615) );
  AOI21_X1 U20790 ( .B1(n21429), .B2(n21340), .A(n17620), .ZN(n17612) );
  AOI21_X1 U20791 ( .B1(n17614), .B2(n17613), .A(n17612), .ZN(n17703) );
  OAI221_X1 U20792 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n17615), 
        .A(n17703), .ZN(n17710) );
  NAND2_X1 U20793 ( .A1(n17710), .A2(n21654), .ZN(n17623) );
  OAI211_X1 U20794 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21434), .A(n17617), 
        .B(n17616), .ZN(n17618) );
  AOI21_X1 U20795 ( .B1(n17620), .B2(n17619), .A(n17618), .ZN(n17621) );
  AND2_X1 U20796 ( .A1(n17710), .A2(n17621), .ZN(n17622) );
  OAI22_X1 U20797 ( .A1(n17624), .A2(n17623), .B1(n17622), .B2(n21654), .ZN(
        P1_U3161) );
  INV_X1 U20798 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21341) );
  NAND2_X1 U20799 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21342) );
  OAI21_X1 U20800 ( .B1(n21355), .B2(n21341), .A(n21342), .ZN(n17625) );
  OAI21_X1 U20801 ( .B1(n21355), .B2(n21357), .A(n17625), .ZN(n17627) );
  OAI211_X1 U20802 ( .C1(n21434), .C2(n21341), .A(n17627), .B(n17626), .ZN(
        P1_U3195) );
  NOR2_X1 U20803 ( .A1(n21698), .A2(n21221), .ZN(P1_U2905) );
  INV_X1 U20804 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21631) );
  INV_X1 U20805 ( .A(n21051), .ZN(n21048) );
  NOR2_X1 U20806 ( .A1(n21631), .A2(n21048), .ZN(P2_U3047) );
  AOI21_X1 U20807 ( .B1(n17640), .B2(n17629), .A(n17628), .ZN(n17650) );
  NOR3_X1 U20808 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21173), .A3(n17629), 
        .ZN(n17630) );
  AOI211_X1 U20809 ( .C1(n21174), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21163), .B(n17630), .ZN(n17634) );
  INV_X1 U20810 ( .A(n17631), .ZN(n17632) );
  AOI22_X1 U20811 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n21182), .B1(n21176), 
        .B2(n17632), .ZN(n17633) );
  OAI211_X1 U20812 ( .C1(n17650), .C2(n21665), .A(n17634), .B(n17633), .ZN(
        n17635) );
  AOI21_X1 U20813 ( .B1(n17636), .B2(n21130), .A(n17635), .ZN(n17637) );
  OAI21_X1 U20814 ( .B1(n17638), .B2(n21170), .A(n17637), .ZN(P1_U2829) );
  AOI21_X1 U20815 ( .B1(n17640), .B2(n17639), .A(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n17649) );
  OAI22_X1 U20816 ( .A1(n17642), .A2(n21122), .B1(n21161), .B2(n17641), .ZN(
        n17643) );
  AOI211_X1 U20817 ( .C1(n21174), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21163), .B(n17643), .ZN(n17648) );
  INV_X1 U20818 ( .A(n17644), .ZN(n17645) );
  AOI22_X1 U20819 ( .A1(n17646), .A2(n21130), .B1(n17645), .B2(n21185), .ZN(
        n17647) );
  OAI211_X1 U20820 ( .C1(n17650), .C2(n17649), .A(n17648), .B(n17647), .ZN(
        P1_U2830) );
  INV_X1 U20821 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21121) );
  OAI21_X1 U20822 ( .B1(n17653), .B2(n17652), .A(n17651), .ZN(n17688) );
  INV_X1 U20823 ( .A(n21123), .ZN(n17656) );
  AOI222_X1 U20824 ( .A1(n17688), .A2(n17668), .B1(n17656), .B2(n17655), .C1(
        n17654), .C2(n21131), .ZN(n17657) );
  OR2_X1 U20825 ( .A1(n17669), .A2(n21369), .ZN(n17685) );
  OAI211_X1 U20826 ( .C1(n21121), .C2(n17671), .A(n17657), .B(n17685), .ZN(
        P1_U2992) );
  OAI22_X1 U20827 ( .A1(n17661), .A2(n17660), .B1(n17659), .B2(n17658), .ZN(
        n17664) );
  XNOR2_X1 U20828 ( .A(n17662), .B(n17695), .ZN(n17663) );
  XNOR2_X1 U20829 ( .A(n17664), .B(n17663), .ZN(n17698) );
  OAI22_X1 U20830 ( .A1(n21152), .A2(n17666), .B1(n21156), .B2(n17665), .ZN(
        n17667) );
  AOI21_X1 U20831 ( .B1(n17698), .B2(n17668), .A(n17667), .ZN(n17670) );
  OR2_X1 U20832 ( .A1(n17669), .A2(n21584), .ZN(n17693) );
  OAI211_X1 U20833 ( .C1(n21695), .C2(n17671), .A(n17670), .B(n17693), .ZN(
        P1_U2994) );
  AOI21_X1 U20834 ( .B1(n21461), .B2(n17673), .A(n17672), .ZN(n17691) );
  OAI211_X1 U20835 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n17683), .B(n17674), .ZN(n17678) );
  INV_X1 U20836 ( .A(n17675), .ZN(n17676) );
  NAND2_X1 U20837 ( .A1(n17676), .A2(n21250), .ZN(n17677) );
  OAI211_X1 U20838 ( .C1(n21564), .C2(n17669), .A(n17678), .B(n17677), .ZN(
        n17679) );
  AOI21_X1 U20839 ( .B1(n17680), .B2(n21251), .A(n17679), .ZN(n17681) );
  OAI21_X1 U20840 ( .B1(n17691), .B2(n17682), .A(n17681), .ZN(P1_U3023) );
  INV_X1 U20841 ( .A(n17683), .ZN(n17686) );
  NAND2_X1 U20842 ( .A1(n21250), .A2(n21126), .ZN(n17684) );
  OAI211_X1 U20843 ( .C1(n17686), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17685), .B(n17684), .ZN(n17687) );
  AOI21_X1 U20844 ( .B1(n17688), .B2(n21251), .A(n17687), .ZN(n17689) );
  OAI21_X1 U20845 ( .B1(n17691), .B2(n17690), .A(n17689), .ZN(P1_U3024) );
  INV_X1 U20846 ( .A(n17692), .ZN(n17701) );
  NAND2_X1 U20847 ( .A1(n21250), .A2(n21146), .ZN(n17694) );
  OAI211_X1 U20848 ( .C1(n17696), .C2(n17695), .A(n17694), .B(n17693), .ZN(
        n17697) );
  AOI21_X1 U20849 ( .B1(n17698), .B2(n21251), .A(n17697), .ZN(n17699) );
  OAI21_X1 U20850 ( .B1(n17701), .B2(n17700), .A(n17699), .ZN(P1_U3026) );
  NAND2_X1 U20851 ( .A1(n17711), .A2(n21434), .ZN(n17707) );
  AOI21_X1 U20852 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n17710), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17706) );
  NOR2_X1 U20853 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21340), .ZN(n17702) );
  OAI221_X1 U20854 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n21654), .C2(n17702), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21336) );
  AOI21_X1 U20855 ( .B1(n21336), .B2(n17704), .A(n17703), .ZN(n17705) );
  AOI211_X1 U20856 ( .C1(n17708), .C2(n17707), .A(n17706), .B(n17705), .ZN(
        P1_U3162) );
  OAI221_X1 U20857 ( .B1(n17711), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n17711), 
        .C2(n17710), .A(n17709), .ZN(P1_U3466) );
  INV_X1 U20858 ( .A(n17712), .ZN(n17713) );
  AOI22_X1 U20859 ( .A1(n17714), .A2(n17713), .B1(P2_REIP_REG_5__SCAN_IN), 
        .B2(n20263), .ZN(n17722) );
  AOI222_X1 U20860 ( .A1(n17720), .A2(n17719), .B1(n17718), .B2(n17717), .C1(
        n17716), .C2(n17715), .ZN(n17721) );
  OAI211_X1 U20861 ( .C1(n17724), .C2(n17723), .A(n17722), .B(n17721), .ZN(
        P2_U3009) );
  NAND2_X1 U20862 ( .A1(n13953), .A2(n20356), .ZN(n17725) );
  OAI21_X1 U20863 ( .B1(n12152), .B2(n20169), .A(n17725), .ZN(n17729) );
  AND3_X1 U20864 ( .A1(n17130), .A2(n17727), .A3(n17726), .ZN(n17728) );
  AOI211_X1 U20865 ( .C1(n21029), .C2(n20355), .A(n17729), .B(n17728), .ZN(
        n17735) );
  AOI21_X1 U20866 ( .B1(n17732), .B2(n17731), .A(n17730), .ZN(n17733) );
  INV_X1 U20867 ( .A(n17733), .ZN(n17734) );
  OAI211_X1 U20868 ( .C1(n17736), .C2(n20360), .A(n17735), .B(n17734), .ZN(
        P2_U3043) );
  AOI211_X1 U20869 ( .C1(n17741), .C2(n17738), .A(n17737), .B(n19177), .ZN(
        n17750) );
  AOI211_X1 U20870 ( .C1(n17741), .C2(n17740), .A(n17739), .B(n19210), .ZN(
        n17749) );
  AOI22_X1 U20871 ( .A1(n19477), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17742), .ZN(n17745) );
  OAI21_X1 U20872 ( .B1(n17743), .B2(n19124), .A(n17871), .ZN(n17744) );
  OAI211_X1 U20873 ( .C1(n17747), .C2(n17746), .A(n17745), .B(n17744), .ZN(
        n17748) );
  NOR3_X1 U20874 ( .A1(n17750), .A2(n17749), .A3(n17748), .ZN(n17751) );
  OAI21_X1 U20875 ( .B1(n19178), .B2(n17752), .A(n17751), .ZN(P3_U2801) );
  NOR3_X1 U20876 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17754) );
  NOR4_X1 U20877 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17753) );
  INV_X2 U20878 ( .A(n17833), .ZN(U215) );
  NAND4_X1 U20879 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17754), .A3(n17753), .A4(
        U215), .ZN(U213) );
  INV_X1 U20880 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21709) );
  OAI222_X1 U20881 ( .A1(U212), .A2(n21709), .B1(n17800), .B2(n17756), .C1(
        U214), .C2(n21698), .ZN(U216) );
  INV_X1 U20882 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n17758) );
  INV_X2 U20883 ( .A(U212), .ZN(n17804) );
  AOI22_X1 U20884 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17804), .ZN(n17757) );
  OAI21_X1 U20885 ( .B1(n17758), .B2(n17800), .A(n17757), .ZN(U217) );
  INV_X1 U20886 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20392) );
  AOI22_X1 U20887 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17804), .ZN(n17759) );
  OAI21_X1 U20888 ( .B1(n20392), .B2(n17800), .A(n17759), .ZN(U218) );
  INV_X1 U20889 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20387) );
  AOI22_X1 U20890 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17804), .ZN(n17760) );
  OAI21_X1 U20891 ( .B1(n20387), .B2(n17800), .A(n17760), .ZN(U219) );
  AOI22_X1 U20892 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17804), .ZN(n17761) );
  OAI21_X1 U20893 ( .B1(n17762), .B2(n17800), .A(n17761), .ZN(U220) );
  AOI22_X1 U20894 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17804), .ZN(n17763) );
  OAI21_X1 U20895 ( .B1(n17764), .B2(n17800), .A(n17763), .ZN(U221) );
  AOI222_X1 U20896 ( .A1(n17798), .A2(P1_DATAO_REG_25__SCAN_IN), .B1(n17803), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n17804), .C2(P2_DATAO_REG_25__SCAN_IN), 
        .ZN(n17765) );
  INV_X1 U20897 ( .A(n17765), .ZN(U222) );
  AOI22_X1 U20898 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17804), .ZN(n17766) );
  OAI21_X1 U20899 ( .B1(n17767), .B2(n17800), .A(n17766), .ZN(U223) );
  INV_X1 U20900 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17769) );
  AOI22_X1 U20901 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17804), .ZN(n17768) );
  OAI21_X1 U20902 ( .B1(n17769), .B2(n17800), .A(n17768), .ZN(U224) );
  INV_X1 U20903 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17771) );
  AOI22_X1 U20904 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17804), .ZN(n17770) );
  OAI21_X1 U20905 ( .B1(n17771), .B2(n17800), .A(n17770), .ZN(U225) );
  INV_X1 U20906 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U20907 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17804), .ZN(n17772) );
  OAI21_X1 U20908 ( .B1(n17773), .B2(n17800), .A(n17772), .ZN(U226) );
  INV_X1 U20909 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U20910 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17804), .ZN(n17774) );
  OAI21_X1 U20911 ( .B1(n17775), .B2(n17800), .A(n17774), .ZN(U227) );
  INV_X1 U20912 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U20913 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17804), .ZN(n17776) );
  OAI21_X1 U20914 ( .B1(n17777), .B2(n17800), .A(n17776), .ZN(U228) );
  AOI222_X1 U20915 ( .A1(n17804), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n17803), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n17798), .C2(P1_DATAO_REG_18__SCAN_IN), 
        .ZN(n17778) );
  INV_X1 U20916 ( .A(n17778), .ZN(U229) );
  AOI22_X1 U20917 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17804), .ZN(n17779) );
  OAI21_X1 U20918 ( .B1(n16863), .B2(n17800), .A(n17779), .ZN(U230) );
  INV_X1 U20919 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U20920 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17804), .ZN(n17780) );
  OAI21_X1 U20921 ( .B1(n17781), .B2(n17800), .A(n17780), .ZN(U231) );
  INV_X1 U20922 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n17783) );
  AOI22_X1 U20923 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17804), .ZN(n17782) );
  OAI21_X1 U20924 ( .B1(n17783), .B2(n17800), .A(n17782), .ZN(U232) );
  AOI22_X1 U20925 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17804), .ZN(n17784) );
  OAI21_X1 U20926 ( .B1(n13543), .B2(n17800), .A(n17784), .ZN(U233) );
  AOI22_X1 U20927 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17804), .ZN(n17785) );
  OAI21_X1 U20928 ( .B1(n13571), .B2(n17800), .A(n17785), .ZN(U234) );
  AOI222_X1 U20929 ( .A1(n17798), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n17803), 
        .B2(BUF1_REG_12__SCAN_IN), .C1(n17804), .C2(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n17786) );
  INV_X1 U20930 ( .A(n17786), .ZN(U235) );
  AOI22_X1 U20931 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17804), .ZN(n17787) );
  OAI21_X1 U20932 ( .B1(n13607), .B2(n17800), .A(n17787), .ZN(U236) );
  AOI22_X1 U20933 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17804), .ZN(n17788) );
  OAI21_X1 U20934 ( .B1(n17789), .B2(n17800), .A(n17788), .ZN(U237) );
  INV_X1 U20935 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17815) );
  INV_X1 U20936 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n21572) );
  OAI222_X1 U20937 ( .A1(U212), .A2(n17815), .B1(n17800), .B2(n13611), .C1(
        U214), .C2(n21572), .ZN(U238) );
  AOI22_X1 U20938 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17804), .ZN(n17790) );
  OAI21_X1 U20939 ( .B1(n17791), .B2(n17800), .A(n17790), .ZN(U239) );
  AOI22_X1 U20940 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17804), .ZN(n17792) );
  OAI21_X1 U20941 ( .B1(n13600), .B2(n17800), .A(n17792), .ZN(U240) );
  INV_X1 U20942 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U20943 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17804), .ZN(n17793) );
  OAI21_X1 U20944 ( .B1(n17794), .B2(n17800), .A(n17793), .ZN(U241) );
  INV_X1 U20945 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n21661) );
  AOI22_X1 U20946 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17804), .ZN(n17795) );
  OAI21_X1 U20947 ( .B1(n21661), .B2(n17800), .A(n17795), .ZN(U242) );
  AOI22_X1 U20948 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17804), .ZN(n17796) );
  OAI21_X1 U20949 ( .B1(n13575), .B2(n17800), .A(n17796), .ZN(U243) );
  AOI22_X1 U20950 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17804), .ZN(n17797) );
  OAI21_X1 U20951 ( .B1(n13579), .B2(n17800), .A(n17797), .ZN(U244) );
  AOI22_X1 U20952 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17798), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17804), .ZN(n17799) );
  OAI21_X1 U20953 ( .B1(n17801), .B2(n17800), .A(n17799), .ZN(U245) );
  INV_X1 U20954 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n21216) );
  AOI22_X1 U20955 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17803), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17804), .ZN(n17802) );
  OAI21_X1 U20956 ( .B1(n21216), .B2(U214), .A(n17802), .ZN(U246) );
  AOI222_X1 U20957 ( .A1(n17804), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n17803), 
        .B2(BUF1_REG_0__SCAN_IN), .C1(n17798), .C2(P1_DATAO_REG_0__SCAN_IN), 
        .ZN(n17805) );
  INV_X1 U20958 ( .A(n17805), .ZN(U247) );
  OAI22_X1 U20959 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n17833), .ZN(n17806) );
  INV_X1 U20960 ( .A(n17806), .ZN(U251) );
  OAI22_X1 U20961 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17833), .ZN(n17807) );
  INV_X1 U20962 ( .A(n17807), .ZN(U252) );
  INV_X1 U20963 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17808) );
  AOI22_X1 U20964 ( .A1(n17833), .A2(n17808), .B1(n19499), .B2(U215), .ZN(U253) );
  OAI22_X1 U20965 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n17833), .ZN(n17809) );
  INV_X1 U20966 ( .A(n17809), .ZN(U254) );
  INV_X1 U20967 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17810) );
  INV_X1 U20968 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19506) );
  AOI22_X1 U20969 ( .A1(n17833), .A2(n17810), .B1(n19506), .B2(U215), .ZN(U255) );
  OAI22_X1 U20970 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17833), .ZN(n17811) );
  INV_X1 U20971 ( .A(n17811), .ZN(U256) );
  INV_X1 U20972 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17812) );
  INV_X1 U20973 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19514) );
  AOI22_X1 U20974 ( .A1(n17833), .A2(n17812), .B1(n19514), .B2(U215), .ZN(U257) );
  INV_X1 U20975 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17813) );
  AOI22_X1 U20976 ( .A1(n17833), .A2(n17813), .B1(n19518), .B2(U215), .ZN(U258) );
  INV_X1 U20977 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17814) );
  INV_X1 U20978 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18889) );
  AOI22_X1 U20979 ( .A1(n17833), .A2(n17814), .B1(n18889), .B2(U215), .ZN(U259) );
  INV_X1 U20980 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18891) );
  AOI22_X1 U20981 ( .A1(n17833), .A2(n17815), .B1(n18891), .B2(U215), .ZN(U260) );
  INV_X1 U20982 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17816) );
  INV_X1 U20983 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18893) );
  AOI22_X1 U20984 ( .A1(n17833), .A2(n17816), .B1(n18893), .B2(U215), .ZN(U261) );
  INV_X1 U20985 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17817) );
  INV_X1 U20986 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18895) );
  AOI22_X1 U20987 ( .A1(n17833), .A2(n17817), .B1(n18895), .B2(U215), .ZN(U262) );
  INV_X1 U20988 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n21660) );
  INV_X1 U20989 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21555) );
  AOI22_X1 U20990 ( .A1(n17833), .A2(n21660), .B1(n21555), .B2(U215), .ZN(U263) );
  INV_X1 U20991 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17818) );
  INV_X1 U20992 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n18901) );
  AOI22_X1 U20993 ( .A1(n17833), .A2(n17818), .B1(n18901), .B2(U215), .ZN(U264) );
  OAI22_X1 U20994 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17833), .ZN(n17819) );
  INV_X1 U20995 ( .A(n17819), .ZN(U265) );
  OAI22_X1 U20996 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17833), .ZN(n17820) );
  INV_X1 U20997 ( .A(n17820), .ZN(U266) );
  OAI22_X1 U20998 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17833), .ZN(n17821) );
  INV_X1 U20999 ( .A(n17821), .ZN(U267) );
  OAI22_X1 U21000 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17833), .ZN(n17822) );
  INV_X1 U21001 ( .A(n17822), .ZN(U268) );
  OAI22_X1 U21002 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17833), .ZN(n17823) );
  INV_X1 U21003 ( .A(n17823), .ZN(U269) );
  OAI22_X1 U21004 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17833), .ZN(n17824) );
  INV_X1 U21005 ( .A(n17824), .ZN(U270) );
  INV_X1 U21006 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U21007 ( .A1(n17833), .A2(n17825), .B1(n21470), .B2(U215), .ZN(U271) );
  OAI22_X1 U21008 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17833), .ZN(n17826) );
  INV_X1 U21009 ( .A(n17826), .ZN(U272) );
  INV_X1 U21010 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U21011 ( .A1(n17833), .A2(n17827), .B1(n16822), .B2(U215), .ZN(U273) );
  INV_X1 U21012 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17828) );
  AOI22_X1 U21013 ( .A1(n17833), .A2(n17828), .B1(n16815), .B2(U215), .ZN(U274) );
  INV_X1 U21014 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n17830) );
  AOI22_X1 U21015 ( .A1(n17833), .A2(n17830), .B1(n17829), .B2(U215), .ZN(U275) );
  INV_X1 U21016 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n21519) );
  AOI22_X1 U21017 ( .A1(n17833), .A2(n21519), .B1(n16800), .B2(U215), .ZN(U276) );
  INV_X1 U21018 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U21019 ( .A1(n17833), .A2(n17832), .B1(n17831), .B2(U215), .ZN(U277) );
  INV_X1 U21020 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U21021 ( .A1(n17833), .A2(n17835), .B1(n17834), .B2(U215), .ZN(U278) );
  INV_X1 U21022 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U21023 ( .A1(n17833), .A2(n17836), .B1(n16780), .B2(U215), .ZN(U279) );
  INV_X1 U21024 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U21025 ( .A1(n17833), .A2(n17838), .B1(n16771), .B2(U215), .ZN(U280) );
  OAI22_X1 U21026 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17833), .ZN(n17839) );
  INV_X1 U21027 ( .A(n17839), .ZN(U281) );
  OAI22_X1 U21028 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n17833), .ZN(n17840) );
  INV_X1 U21029 ( .A(n17840), .ZN(U282) );
  AOI222_X1 U21030 ( .A1(n18797), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n21698), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n21709), .C2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n17841) );
  INV_X1 U21031 ( .A(n17843), .ZN(n17842) );
  INV_X1 U21032 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20019) );
  INV_X1 U21033 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20969) );
  AOI22_X1 U21034 ( .A1(n17842), .A2(n20019), .B1(n20969), .B2(n17843), .ZN(
        U347) );
  INV_X1 U21035 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n21452) );
  INV_X1 U21036 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U21037 ( .A1(n17844), .A2(n21452), .B1(n20967), .B2(n17843), .ZN(
        U348) );
  INV_X1 U21038 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20015) );
  INV_X1 U21039 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20965) );
  AOI22_X1 U21040 ( .A1(n17842), .A2(n20015), .B1(n20965), .B2(n17843), .ZN(
        U349) );
  INV_X1 U21041 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20014) );
  INV_X1 U21042 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U21043 ( .A1(n17842), .A2(n20014), .B1(n20964), .B2(n17843), .ZN(
        U350) );
  INV_X1 U21044 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20012) );
  INV_X1 U21045 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20962) );
  AOI22_X1 U21046 ( .A1(n17842), .A2(n20012), .B1(n20962), .B2(n17843), .ZN(
        U351) );
  INV_X1 U21047 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U21048 ( .A1(n17842), .A2(n20010), .B1(n20960), .B2(n17843), .ZN(
        U352) );
  INV_X1 U21049 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n20009) );
  INV_X1 U21050 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21678) );
  AOI22_X1 U21051 ( .A1(n17844), .A2(n20009), .B1(n21678), .B2(n17843), .ZN(
        U353) );
  INV_X1 U21052 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n21496) );
  INV_X1 U21053 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n21453) );
  AOI22_X1 U21054 ( .A1(n17842), .A2(n21496), .B1(n21453), .B2(n17843), .ZN(
        U354) );
  INV_X1 U21055 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20060) );
  INV_X1 U21056 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n21716) );
  AOI22_X1 U21057 ( .A1(n17842), .A2(n20060), .B1(n21716), .B2(n17843), .ZN(
        U355) );
  INV_X1 U21058 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20057) );
  INV_X1 U21059 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n21005) );
  AOI22_X1 U21060 ( .A1(n17842), .A2(n20057), .B1(n21005), .B2(n17843), .ZN(
        U356) );
  INV_X1 U21061 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20054) );
  INV_X1 U21062 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21003) );
  AOI22_X1 U21063 ( .A1(n17842), .A2(n20054), .B1(n21003), .B2(n17843), .ZN(
        U357) );
  INV_X1 U21064 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20053) );
  INV_X1 U21065 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n21000) );
  AOI22_X1 U21066 ( .A1(n17842), .A2(n20053), .B1(n21000), .B2(n17843), .ZN(
        U358) );
  INV_X1 U21067 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20051) );
  INV_X1 U21068 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U21069 ( .A1(n17842), .A2(n20051), .B1(n20998), .B2(n17843), .ZN(
        U359) );
  INV_X1 U21070 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20049) );
  INV_X1 U21071 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20996) );
  AOI22_X1 U21072 ( .A1(n17842), .A2(n20049), .B1(n20996), .B2(n17843), .ZN(
        U360) );
  INV_X1 U21073 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20047) );
  INV_X1 U21074 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20994) );
  AOI22_X1 U21075 ( .A1(n17842), .A2(n20047), .B1(n20994), .B2(n17843), .ZN(
        U361) );
  INV_X1 U21076 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20045) );
  INV_X1 U21077 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U21078 ( .A1(n17842), .A2(n20045), .B1(n20992), .B2(n17843), .ZN(
        U362) );
  INV_X1 U21079 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20043) );
  INV_X1 U21080 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U21081 ( .A1(n17842), .A2(n20043), .B1(n20990), .B2(n17843), .ZN(
        U363) );
  INV_X1 U21082 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20041) );
  INV_X1 U21083 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20988) );
  AOI22_X1 U21084 ( .A1(n17842), .A2(n20041), .B1(n20988), .B2(n17843), .ZN(
        U364) );
  INV_X1 U21085 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n20005) );
  INV_X1 U21086 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20958) );
  AOI22_X1 U21087 ( .A1(n17842), .A2(n20005), .B1(n20958), .B2(n17843), .ZN(
        U365) );
  INV_X1 U21088 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20039) );
  INV_X1 U21089 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20986) );
  AOI22_X1 U21090 ( .A1(n17842), .A2(n20039), .B1(n20986), .B2(n17843), .ZN(
        U366) );
  INV_X1 U21091 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20037) );
  INV_X1 U21092 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20984) );
  AOI22_X1 U21093 ( .A1(n17842), .A2(n20037), .B1(n20984), .B2(n17843), .ZN(
        U367) );
  INV_X1 U21094 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20035) );
  INV_X1 U21095 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20982) );
  AOI22_X1 U21096 ( .A1(n17842), .A2(n20035), .B1(n20982), .B2(n17843), .ZN(
        U368) );
  INV_X1 U21097 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20032) );
  INV_X1 U21098 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20980) );
  AOI22_X1 U21099 ( .A1(n17842), .A2(n20032), .B1(n20980), .B2(n17843), .ZN(
        U369) );
  INV_X1 U21100 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20031) );
  INV_X1 U21101 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20978) );
  AOI22_X1 U21102 ( .A1(n17842), .A2(n20031), .B1(n20978), .B2(n17843), .ZN(
        U370) );
  INV_X1 U21103 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20029) );
  INV_X1 U21104 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U21105 ( .A1(n17844), .A2(n20029), .B1(n20976), .B2(n17843), .ZN(
        U371) );
  INV_X1 U21106 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20026) );
  INV_X1 U21107 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U21108 ( .A1(n17844), .A2(n20026), .B1(n20974), .B2(n17843), .ZN(
        U372) );
  INV_X1 U21109 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20025) );
  INV_X1 U21110 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U21111 ( .A1(n17844), .A2(n20025), .B1(n20972), .B2(n17843), .ZN(
        U373) );
  INV_X1 U21112 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20023) );
  INV_X1 U21113 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20971) );
  AOI22_X1 U21114 ( .A1(n17844), .A2(n20023), .B1(n20971), .B2(n17843), .ZN(
        U374) );
  INV_X1 U21115 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20021) );
  INV_X1 U21116 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U21117 ( .A1(n17844), .A2(n20021), .B1(n20970), .B2(n17843), .ZN(
        U375) );
  INV_X1 U21118 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20004) );
  INV_X1 U21119 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U21120 ( .A1(n17844), .A2(n20004), .B1(n20956), .B2(n17843), .ZN(
        U376) );
  INV_X1 U21121 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17845) );
  INV_X1 U21122 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U21123 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n20003), .ZN(n19994) );
  INV_X1 U21124 ( .A(n20067), .ZN(n20065) );
  OAI21_X1 U21125 ( .B1(n20001), .B2(n17845), .A(n20065), .ZN(P3_U2633) );
  AOI21_X1 U21126 ( .B1(n18858), .B2(n17852), .A(n18857), .ZN(n17847) );
  INV_X1 U21127 ( .A(P3_CODEFETCH_REG_SCAN_IN), .ZN(n21568) );
  OAI22_X1 U21128 ( .A1(n17847), .A2(n21568), .B1(n19980), .B2(n17846), .ZN(
        P3_U2634) );
  AOI21_X1 U21129 ( .B1(n20001), .B2(n20003), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17848) );
  AOI22_X1 U21130 ( .A1(n20101), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17848), 
        .B2(n20099), .ZN(P3_U2635) );
  NOR2_X1 U21131 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19986) );
  OAI21_X1 U21132 ( .B1(n19986), .B2(BS16), .A(n20067), .ZN(n20066) );
  OAI21_X1 U21133 ( .B1(n20067), .B2(n17849), .A(n20066), .ZN(P3_U2636) );
  AOI211_X1 U21134 ( .C1(n18858), .C2(n17852), .A(n17851), .B(n17850), .ZN(
        n19957) );
  NOR2_X1 U21135 ( .A1(n19957), .A2(n19976), .ZN(n20081) );
  OAI21_X1 U21136 ( .B1(n20081), .B2(n19482), .A(n17853), .ZN(P3_U2637) );
  NOR4_X1 U21137 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17863) );
  NOR4_X1 U21138 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n17862) );
  AOI211_X1 U21139 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_3__SCAN_IN), .B(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n17854) );
  INV_X1 U21140 ( .A(P3_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21455) );
  INV_X1 U21141 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21533) );
  NAND3_X1 U21142 ( .A1(n17854), .A2(n21455), .A3(n21533), .ZN(n17860) );
  NOR4_X1 U21143 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17858) );
  NOR4_X1 U21144 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n17857) );
  NOR4_X1 U21145 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17856) );
  NOR4_X1 U21146 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17855) );
  NAND4_X1 U21147 ( .A1(n17858), .A2(n17857), .A3(n17856), .A4(n17855), .ZN(
        n17859) );
  NOR4_X1 U21148 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(n17860), .A4(n17859), .ZN(n17861) );
  NAND3_X1 U21149 ( .A1(n17863), .A2(n17862), .A3(n17861), .ZN(n20077) );
  NOR2_X1 U21150 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20077), .ZN(n20079) );
  INV_X1 U21151 ( .A(n20077), .ZN(n17864) );
  NOR2_X1 U21152 ( .A1(n17864), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17865)
         );
  INV_X1 U21153 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20078) );
  INV_X1 U21154 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20071) );
  INV_X1 U21155 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20072) );
  NAND4_X1 U21156 ( .A1(n17864), .A2(n20078), .A3(n20071), .A4(n20072), .ZN(
        n17866) );
  OAI21_X1 U21157 ( .B1(n20079), .B2(n17865), .A(n17866), .ZN(P3_U2638) );
  AOI22_X1 U21158 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n20077), .B1(n20079), .B2(n20071), .ZN(n17867) );
  NAND2_X1 U21159 ( .A1(n17867), .A2(n17866), .ZN(P3_U2639) );
  NOR2_X1 U21160 ( .A1(n17881), .A2(n17868), .ZN(n17879) );
  AOI211_X1 U21161 ( .C1(n17871), .C2(n17870), .A(n17869), .B(n13366), .ZN(
        n17875) );
  INV_X1 U21162 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20056) );
  OAI22_X1 U21163 ( .A1(n17873), .A2(n20056), .B1(n17872), .B2(n18219), .ZN(
        n17874) );
  AOI211_X1 U21164 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n18217), .A(n17875), .B(
        n17874), .ZN(n17877) );
  NAND4_X1 U21165 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17880), .A4(n20056), .ZN(n17876) );
  OAI211_X1 U21166 ( .C1(n17879), .C2(n17878), .A(n17877), .B(n17876), .ZN(
        P3_U2642) );
  NAND2_X1 U21167 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17880), .ZN(n17889) );
  AOI22_X1 U21168 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17888) );
  INV_X1 U21169 ( .A(n17909), .ZN(n17894) );
  INV_X1 U21170 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20052) );
  NAND2_X1 U21171 ( .A1(n17880), .A2(n20052), .ZN(n17900) );
  NAND2_X1 U21172 ( .A1(n17894), .A2(n17900), .ZN(n17886) );
  AOI211_X1 U21173 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17897), .A(n17881), .B(
        n18226), .ZN(n17885) );
  AOI211_X1 U21174 ( .C1(n10510), .C2(n17883), .A(n17882), .B(n13366), .ZN(
        n17884) );
  AOI211_X1 U21175 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17886), .A(n17885), 
        .B(n17884), .ZN(n17887) );
  OAI211_X1 U21176 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17889), .A(n17888), 
        .B(n17887), .ZN(P3_U2643) );
  INV_X1 U21177 ( .A(n17890), .ZN(n17893) );
  INV_X1 U21178 ( .A(n17891), .ZN(n17892) );
  AOI211_X1 U21179 ( .C1(n18913), .C2(n17893), .A(n17892), .B(n13366), .ZN(
        n17896) );
  OAI22_X1 U21180 ( .A1(n18916), .A2(n18219), .B1(n20052), .B2(n17894), .ZN(
        n17895) );
  AOI211_X1 U21181 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n18217), .A(n17896), .B(
        n17895), .ZN(n17901) );
  OAI211_X1 U21182 ( .C1(n17902), .C2(n17898), .A(n18171), .B(n17897), .ZN(
        n17899) );
  NAND3_X1 U21183 ( .A1(n17901), .A2(n17900), .A3(n17899), .ZN(P3_U2644) );
  AOI22_X1 U21184 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17911) );
  AOI211_X1 U21185 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17903), .A(n17902), .B(
        n18226), .ZN(n17908) );
  CLKBUF_X1 U21186 ( .A(n17904), .Z(n17905) );
  AOI211_X1 U21187 ( .C1(n18928), .C2(n17906), .A(n17905), .B(n13366), .ZN(
        n17907) );
  AOI211_X1 U21188 ( .C1(n17909), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17908), 
        .B(n17907), .ZN(n17910) );
  OAI211_X1 U21189 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17912), .A(n17911), 
        .B(n17910), .ZN(P3_U2645) );
  OR2_X1 U21190 ( .A1(n18226), .A2(n17913), .ZN(n17926) );
  AOI21_X1 U21191 ( .B1(n18171), .B2(n17913), .A(n18217), .ZN(n17923) );
  AOI211_X1 U21192 ( .C1(n18940), .C2(n17915), .A(n17914), .B(n13366), .ZN(
        n17921) );
  NOR2_X1 U21193 ( .A1(n18205), .A2(n17916), .ZN(n17919) );
  INV_X1 U21194 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20046) );
  OAI21_X1 U21195 ( .B1(n17937), .B2(n18205), .A(n18212), .ZN(n17933) );
  AOI21_X1 U21196 ( .B1(n18169), .B2(n20046), .A(n17933), .ZN(n17917) );
  INV_X1 U21197 ( .A(n17917), .ZN(n17918) );
  MUX2_X1 U21198 ( .A(n17919), .B(n17918), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n17920) );
  AOI211_X1 U21199 ( .C1(n18193), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17921), .B(n17920), .ZN(n17922) );
  OAI221_X1 U21200 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17926), .C1(n17924), 
        .C2(n17923), .A(n17922), .ZN(P3_U2646) );
  NOR2_X1 U21201 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18205), .ZN(n17925) );
  AOI22_X1 U21202 ( .A1(n18217), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17937), 
        .B2(n17925), .ZN(n17932) );
  AOI21_X1 U21203 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17942), .A(n17926), .ZN(
        n17930) );
  AOI211_X1 U21204 ( .C1(n18960), .C2(n17928), .A(n17927), .B(n13366), .ZN(
        n17929) );
  AOI211_X1 U21205 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17933), .A(n17930), 
        .B(n17929), .ZN(n17931) );
  OAI211_X1 U21206 ( .C1(n18951), .C2(n18219), .A(n17932), .B(n17931), .ZN(
        P3_U2647) );
  INV_X1 U21207 ( .A(n17933), .ZN(n17946) );
  INV_X1 U21208 ( .A(n17934), .ZN(n17935) );
  AOI211_X1 U21209 ( .C1(n18968), .C2(n17936), .A(n17935), .B(n13366), .ZN(
        n17941) );
  OR2_X1 U21210 ( .A1(n18205), .A2(n17937), .ZN(n17938) );
  OAI22_X1 U21211 ( .A1(n18967), .A2(n18219), .B1(n17939), .B2(n17938), .ZN(
        n17940) );
  AOI211_X1 U21212 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n18217), .A(n17941), .B(
        n17940), .ZN(n17945) );
  OAI211_X1 U21213 ( .C1(n17951), .C2(n17943), .A(n18171), .B(n17942), .ZN(
        n17944) );
  OAI211_X1 U21214 ( .C1(n17946), .C2(n20044), .A(n17945), .B(n17944), .ZN(
        P3_U2648) );
  NAND2_X1 U21215 ( .A1(n18169), .A2(n17949), .ZN(n17984) );
  NOR2_X1 U21216 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17984), .ZN(n17947) );
  AOI22_X1 U21217 ( .A1(n18217), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n17948), 
        .B2(n17947), .ZN(n17958) );
  NAND2_X1 U21218 ( .A1(n17949), .A2(n18212), .ZN(n18029) );
  OAI21_X1 U21219 ( .B1(n17950), .B2(n18029), .A(n18156), .ZN(n17959) );
  OR3_X1 U21220 ( .A1(n17950), .A2(n17984), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n17965) );
  NAND2_X1 U21221 ( .A1(n17959), .A2(n17965), .ZN(n17956) );
  AOI211_X1 U21222 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17963), .A(n17951), .B(
        n18226), .ZN(n17955) );
  AOI211_X1 U21223 ( .C1(n18985), .C2(n17953), .A(n17952), .B(n13366), .ZN(
        n17954) );
  AOI211_X1 U21224 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17956), .A(n17955), 
        .B(n17954), .ZN(n17957) );
  OAI211_X1 U21225 ( .C1(n18987), .C2(n18219), .A(n17958), .B(n17957), .ZN(
        P3_U2649) );
  AOI22_X1 U21226 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17967) );
  INV_X1 U21227 ( .A(n17959), .ZN(n17973) );
  AOI211_X1 U21228 ( .C1(n18996), .C2(n17961), .A(n17960), .B(n13366), .ZN(
        n17962) );
  AOI21_X1 U21229 ( .B1(n17973), .B2(P3_REIP_REG_21__SCAN_IN), .A(n17962), 
        .ZN(n17966) );
  OAI211_X1 U21230 ( .C1(n17970), .C2(n18419), .A(n18171), .B(n17963), .ZN(
        n17964) );
  NAND4_X1 U21231 ( .A1(n17967), .A2(n17966), .A3(n17965), .A4(n17964), .ZN(
        P3_U2650) );
  AOI211_X1 U21232 ( .C1(n19005), .C2(n17969), .A(n17968), .B(n13366), .ZN(
        n17972) );
  AOI211_X1 U21233 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17979), .A(n17970), .B(
        n18226), .ZN(n17971) );
  AOI211_X1 U21234 ( .C1(n18193), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17972), .B(n17971), .ZN(n17976) );
  INV_X1 U21235 ( .A(n17984), .ZN(n18013) );
  OAI221_X1 U21236 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17974), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n18013), .A(n17973), .ZN(n17975) );
  OAI211_X1 U21237 ( .C1(n10142), .C2(n18158), .A(n17976), .B(n17975), .ZN(
        P3_U2651) );
  OAI21_X1 U21238 ( .B1(n17985), .B2(n18029), .A(n18156), .ZN(n18008) );
  INV_X1 U21239 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20036) );
  INV_X1 U21240 ( .A(n17977), .ZN(n17978) );
  AOI211_X1 U21241 ( .C1(n19024), .C2(n9847), .A(n17978), .B(n13366), .ZN(
        n17983) );
  OAI211_X1 U21242 ( .C1(n17989), .C2(n17981), .A(n18171), .B(n17979), .ZN(
        n17980) );
  OAI211_X1 U21243 ( .C1(n18158), .C2(n17981), .A(n19428), .B(n17980), .ZN(
        n17982) );
  AOI211_X1 U21244 ( .C1(n18193), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n17983), .B(n17982), .ZN(n17988) );
  NOR2_X1 U21245 ( .A1(n17985), .A2(n17984), .ZN(n17995) );
  OAI211_X1 U21246 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17995), .B(n17986), .ZN(n17987) );
  OAI211_X1 U21247 ( .C1(n18008), .C2(n20036), .A(n17988), .B(n17987), .ZN(
        P3_U2652) );
  AOI211_X1 U21248 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n18001), .A(n17989), .B(
        n18226), .ZN(n17990) );
  AOI211_X1 U21249 ( .C1(n18217), .C2(P3_EBX_REG_18__SCAN_IN), .A(n19477), .B(
        n17990), .ZN(n17998) );
  INV_X1 U21250 ( .A(n18008), .ZN(n17996) );
  INV_X1 U21251 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n20034) );
  INV_X1 U21252 ( .A(n17991), .ZN(n17992) );
  AOI211_X1 U21253 ( .C1(n19036), .C2(n17993), .A(n17992), .B(n13366), .ZN(
        n17994) );
  AOI221_X1 U21254 ( .B1(n17996), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n17995), 
        .C2(n20034), .A(n17994), .ZN(n17997) );
  OAI211_X1 U21255 ( .C1(n21731), .C2(n18219), .A(n17998), .B(n17997), .ZN(
        P3_U2653) );
  INV_X1 U21256 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20030) );
  NAND2_X1 U21257 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18013), .ZN(n18019) );
  INV_X1 U21258 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U21259 ( .B1(n20030), .B2(n18019), .A(n20033), .ZN(n17999) );
  INV_X1 U21260 ( .A(n17999), .ZN(n18009) );
  INV_X1 U21261 ( .A(n18014), .ZN(n18000) );
  AOI21_X1 U21262 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18000), .A(n18226), .ZN(
        n18002) );
  AOI22_X1 U21263 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18193), .B1(
        n18002), .B2(n18001), .ZN(n18007) );
  AOI211_X1 U21264 ( .C1(n19046), .C2(n18004), .A(n18003), .B(n13366), .ZN(
        n18005) );
  AOI211_X1 U21265 ( .C1(n18217), .C2(P3_EBX_REG_17__SCAN_IN), .A(n19477), .B(
        n18005), .ZN(n18006) );
  OAI211_X1 U21266 ( .C1(n18009), .C2(n18008), .A(n18007), .B(n18006), .ZN(
        P3_U2654) );
  AOI211_X1 U21267 ( .C1(n19060), .C2(n18011), .A(n18010), .B(n13366), .ZN(
        n18012) );
  AOI211_X1 U21268 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18193), .A(
        n19477), .B(n18012), .ZN(n18018) );
  NAND2_X1 U21269 ( .A1(n18156), .A2(n18029), .ZN(n18028) );
  INV_X1 U21270 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20028) );
  NAND2_X1 U21271 ( .A1(n18013), .A2(n20028), .ZN(n18024) );
  AOI21_X1 U21272 ( .B1(n18028), .B2(n18024), .A(n20030), .ZN(n18016) );
  AOI211_X1 U21273 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18022), .A(n18014), .B(
        n18226), .ZN(n18015) );
  AOI211_X1 U21274 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n18217), .A(n18016), .B(
        n18015), .ZN(n18017) );
  OAI211_X1 U21275 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n18019), .A(n18018), 
        .B(n18017), .ZN(P3_U2655) );
  NOR2_X1 U21276 ( .A1(n18059), .A2(n18120), .ZN(n19104) );
  NAND2_X1 U21277 ( .A1(n19102), .A2(n19104), .ZN(n18043) );
  NOR2_X1 U21278 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18043), .ZN(
        n18033) );
  AOI21_X1 U21279 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18033), .A(
        n9750), .ZN(n18035) );
  INV_X1 U21280 ( .A(n19058), .ZN(n18032) );
  OAI21_X1 U21281 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18032), .A(
        n18020), .ZN(n19075) );
  XOR2_X1 U21282 ( .A(n18035), .B(n19075), .Z(n18021) );
  OAI22_X1 U21283 ( .A1(n18158), .A2(n18514), .B1(n13366), .B2(n18021), .ZN(
        n18026) );
  OAI211_X1 U21284 ( .C1(n18031), .C2(n18514), .A(n18171), .B(n18022), .ZN(
        n18023) );
  OAI211_X1 U21285 ( .C1(n18219), .C2(n19078), .A(n18024), .B(n18023), .ZN(
        n18025) );
  NOR3_X1 U21286 ( .A1(n19477), .A2(n18026), .A3(n18025), .ZN(n18027) );
  OAI21_X1 U21287 ( .B1(n20028), .B2(n18028), .A(n18027), .ZN(P3_U2656) );
  INV_X1 U21288 ( .A(n18029), .ZN(n18042) );
  NOR2_X1 U21289 ( .A1(n18205), .A2(n18030), .ZN(n18046) );
  AOI22_X1 U21290 ( .A1(n18046), .A2(P3_REIP_REG_13__SCAN_IN), .B1(
        P3_REIP_REG_14__SCAN_IN), .B2(n18156), .ZN(n18041) );
  AOI211_X1 U21291 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18049), .A(n18031), .B(
        n18226), .ZN(n18039) );
  INV_X1 U21292 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n18037) );
  INV_X1 U21293 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19087) );
  AOI21_X1 U21294 ( .B1(n19087), .B2(n18043), .A(n18032), .ZN(n19089) );
  NOR2_X1 U21295 ( .A1(n18132), .A2(n13366), .ZN(n18163) );
  INV_X1 U21296 ( .A(n18033), .ZN(n18044) );
  AOI21_X1 U21297 ( .B1(n19089), .B2(n18044), .A(n13366), .ZN(n18034) );
  OAI22_X1 U21298 ( .A1(n19089), .A2(n18035), .B1(n18163), .B2(n18034), .ZN(
        n18036) );
  OAI211_X1 U21299 ( .C1(n18158), .C2(n18037), .A(n19428), .B(n18036), .ZN(
        n18038) );
  AOI211_X1 U21300 ( .C1(n18193), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n18039), .B(n18038), .ZN(n18040) );
  OAI21_X1 U21301 ( .B1(n18042), .B2(n18041), .A(n18040), .ZN(P3_U2657) );
  INV_X1 U21302 ( .A(n19104), .ZN(n18057) );
  NOR2_X1 U21303 ( .A1(n19120), .A2(n18057), .ZN(n18056) );
  OAI21_X1 U21304 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18056), .A(
        n18043), .ZN(n19108) );
  OAI21_X1 U21305 ( .B1(n9750), .B2(n18221), .A(n18189), .ZN(n18218) );
  AOI211_X1 U21306 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18132), .A(
        n19108), .B(n18218), .ZN(n18055) );
  NAND2_X1 U21307 ( .A1(n19108), .A2(n18044), .ZN(n18045) );
  OAI22_X1 U21308 ( .A1(n18158), .A2(n18050), .B1(n18220), .B2(n18045), .ZN(
        n18054) );
  INV_X1 U21309 ( .A(n18046), .ZN(n18048) );
  OAI21_X1 U21310 ( .B1(n18065), .B2(n18205), .A(n18212), .ZN(n18073) );
  NOR2_X1 U21311 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18205), .ZN(n18064) );
  NOR2_X1 U21312 ( .A1(n18073), .A2(n18064), .ZN(n18047) );
  MUX2_X1 U21313 ( .A(n18048), .B(n18047), .S(P3_REIP_REG_13__SCAN_IN), .Z(
        n18052) );
  OAI211_X1 U21314 ( .C1(n18061), .C2(n18050), .A(n18171), .B(n18049), .ZN(
        n18051) );
  OAI211_X1 U21315 ( .C1(n18219), .C2(n19110), .A(n18052), .B(n18051), .ZN(
        n18053) );
  OR4_X1 U21316 ( .A1(n19477), .A2(n18055), .A3(n18054), .A4(n18053), .ZN(
        P3_U2658) );
  AOI21_X1 U21317 ( .B1(n19120), .B2(n18057), .A(n18056), .ZN(n19123) );
  NOR2_X1 U21318 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18177), .ZN(
        n18197) );
  NAND2_X1 U21319 ( .A1(n18058), .A2(n18197), .ZN(n18121) );
  OAI21_X1 U21320 ( .B1(n18059), .B2(n18121), .A(n18132), .ZN(n18060) );
  XNOR2_X1 U21321 ( .A(n19123), .B(n18060), .ZN(n18063) );
  AOI211_X1 U21322 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n18074), .A(n18061), .B(
        n18226), .ZN(n18062) );
  AOI211_X1 U21323 ( .C1(n18189), .C2(n18063), .A(n19477), .B(n18062), .ZN(
        n18068) );
  AOI22_X1 U21324 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U21325 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18073), .B1(n18065), 
        .B2(n18064), .ZN(n18066) );
  NAND3_X1 U21326 ( .A1(n18068), .A2(n18067), .A3(n18066), .ZN(P3_U2659) );
  INV_X1 U21327 ( .A(n18069), .ZN(n18089) );
  NAND3_X1 U21328 ( .A1(n18169), .A2(P3_REIP_REG_4__SCAN_IN), .A3(n18168), 
        .ZN(n18144) );
  NAND2_X1 U21329 ( .A1(n18089), .A2(n18140), .ZN(n18106) );
  OAI21_X1 U21330 ( .B1(n18070), .B2(n18106), .A(n20020), .ZN(n18072) );
  INV_X1 U21331 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19135) );
  OAI22_X1 U21332 ( .A1(n19135), .A2(n18219), .B1(n18158), .B2(n21456), .ZN(
        n18071) );
  AOI21_X1 U21333 ( .B1(n18073), .B2(n18072), .A(n18071), .ZN(n18081) );
  OAI211_X1 U21334 ( .C1(n18086), .C2(n21456), .A(n18171), .B(n18074), .ZN(
        n18080) );
  NOR2_X1 U21335 ( .A1(n19133), .A2(n18120), .ZN(n18119) );
  NAND2_X1 U21336 ( .A1(n18075), .A2(n18119), .ZN(n18082) );
  AOI21_X1 U21337 ( .B1(n19135), .B2(n18082), .A(n19104), .ZN(n19138) );
  OAI21_X1 U21338 ( .B1(n18082), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18132), .ZN(n18076) );
  INV_X1 U21339 ( .A(n18076), .ZN(n18078) );
  AOI21_X1 U21340 ( .B1(n19138), .B2(n18078), .A(n13366), .ZN(n18077) );
  OAI21_X1 U21341 ( .B1(n19138), .B2(n18078), .A(n18077), .ZN(n18079) );
  NAND4_X1 U21342 ( .A1(n18081), .A2(n19216), .A3(n18080), .A4(n18079), .ZN(
        P3_U2660) );
  AND3_X1 U21343 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n18119), .ZN(n18098) );
  OAI21_X1 U21344 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18098), .A(
        n18082), .ZN(n18083) );
  INV_X1 U21345 ( .A(n18083), .ZN(n19149) );
  NAND2_X1 U21346 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18084) );
  NAND2_X1 U21347 ( .A1(n18119), .A2(n18221), .ZN(n18109) );
  OAI21_X1 U21348 ( .B1(n18084), .B2(n18109), .A(n18132), .ZN(n18099) );
  XNOR2_X1 U21349 ( .A(n19149), .B(n18099), .ZN(n18085) );
  AOI22_X1 U21350 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18193), .B1(
        n18189), .B2(n18085), .ZN(n18095) );
  AOI211_X1 U21351 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18096), .A(n18086), .B(
        n18226), .ZN(n18093) );
  INV_X1 U21352 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20017) );
  NOR2_X1 U21353 ( .A1(n20017), .A2(n18106), .ZN(n18091) );
  INV_X1 U21354 ( .A(n18212), .ZN(n18087) );
  AOI21_X1 U21355 ( .B1(n18169), .B2(n18088), .A(n18087), .ZN(n18143) );
  OAI21_X1 U21356 ( .B1(n18089), .B2(n18205), .A(n18143), .ZN(n18115) );
  AOI21_X1 U21357 ( .B1(n18156), .B2(n20017), .A(n18115), .ZN(n18107) );
  INV_X1 U21358 ( .A(n18107), .ZN(n18090) );
  MUX2_X1 U21359 ( .A(n18091), .B(n18090), .S(P3_REIP_REG_10__SCAN_IN), .Z(
        n18092) );
  AOI211_X1 U21360 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n18217), .A(n18093), .B(
        n18092), .ZN(n18094) );
  NAND3_X1 U21361 ( .A1(n18095), .A2(n18094), .A3(n19216), .ZN(P3_U2661) );
  AOI22_X1 U21362 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n18104) );
  OAI211_X1 U21363 ( .C1(n18108), .C2(n18097), .A(n18171), .B(n18096), .ZN(
        n18103) );
  NAND2_X1 U21364 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18119), .ZN(
        n18110) );
  AOI21_X1 U21365 ( .B1(n19159), .B2(n18110), .A(n18098), .ZN(n19163) );
  INV_X1 U21366 ( .A(n18099), .ZN(n18101) );
  AOI221_X1 U21367 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19163), .C1(
        n18110), .C2(n19163), .A(n13366), .ZN(n18100) );
  OAI22_X1 U21368 ( .A1(n19163), .A2(n18101), .B1(n18163), .B2(n18100), .ZN(
        n18102) );
  AND4_X1 U21369 ( .A1(n18104), .A2(n19428), .A3(n18103), .A4(n18102), .ZN(
        n18105) );
  OAI221_X1 U21370 ( .B1(n18107), .B2(n20017), .C1(n18107), .C2(n18106), .A(
        n18105), .ZN(P3_U2662) );
  NAND3_X1 U21371 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n18140), .ZN(n18118) );
  AOI22_X1 U21372 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_8__SCAN_IN), .ZN(n18117) );
  AOI211_X1 U21373 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18122), .A(n18108), .B(
        n18226), .ZN(n18114) );
  NAND2_X1 U21374 ( .A1(n18132), .A2(n18109), .ZN(n18111) );
  OAI21_X1 U21375 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18119), .A(
        n18110), .ZN(n19168) );
  XNOR2_X1 U21376 ( .A(n18111), .B(n19168), .ZN(n18112) );
  OAI21_X1 U21377 ( .B1(n18112), .B2(n13366), .A(n19428), .ZN(n18113) );
  AOI211_X1 U21378 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18115), .A(n18114), .B(
        n18113), .ZN(n18116) );
  OAI211_X1 U21379 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18118), .A(n18117), .B(
        n18116), .ZN(P3_U2663) );
  INV_X1 U21380 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20013) );
  OAI22_X1 U21381 ( .A1(n19133), .A2(n18219), .B1(n18158), .B2(n18123), .ZN(
        n18127) );
  AOI21_X1 U21382 ( .B1(n19133), .B2(n18120), .A(n18119), .ZN(n19191) );
  NAND2_X1 U21383 ( .A1(n18132), .A2(n18121), .ZN(n18131) );
  XOR2_X1 U21384 ( .A(n19191), .B(n18131), .Z(n18125) );
  OAI211_X1 U21385 ( .C1(n18133), .C2(n18123), .A(n18171), .B(n18122), .ZN(
        n18124) );
  OAI211_X1 U21386 ( .C1(n13366), .C2(n18125), .A(n19428), .B(n18124), .ZN(
        n18126) );
  NOR2_X1 U21387 ( .A1(n18127), .A2(n18126), .ZN(n18130) );
  NAND2_X1 U21388 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n18128) );
  OAI211_X1 U21389 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n18140), .B(n18128), .ZN(n18129) );
  OAI211_X1 U21390 ( .C1(n18143), .C2(n20013), .A(n18130), .B(n18129), .ZN(
        P3_U2664) );
  NOR2_X1 U21391 ( .A1(n13366), .A2(n18131), .ZN(n18137) );
  AOI211_X1 U21392 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18132), .A(
        n18136), .B(n18218), .ZN(n18135) );
  AOI211_X1 U21393 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18148), .A(n18133), .B(
        n18226), .ZN(n18134) );
  AOI211_X1 U21394 ( .C1(n18137), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        n18142) );
  INV_X1 U21395 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20011) );
  INV_X1 U21396 ( .A(n18143), .ZN(n18139) );
  OAI22_X1 U21397 ( .A1(n19134), .A2(n18219), .B1(n18158), .B2(n18629), .ZN(
        n18138) );
  AOI221_X1 U21398 ( .B1(n18140), .B2(n20011), .C1(n18139), .C2(
        P3_REIP_REG_6__SCAN_IN), .A(n18138), .ZN(n18141) );
  NAND3_X1 U21399 ( .A1(n18142), .A2(n18141), .A3(n19216), .ZN(P3_U2665) );
  AOI21_X1 U21400 ( .B1(n21460), .B2(n18144), .A(n18143), .ZN(n18153) );
  AOI21_X1 U21401 ( .B1(n18147), .B2(n18221), .A(n9750), .ZN(n18160) );
  INV_X1 U21402 ( .A(n18145), .ZN(n18146) );
  OAI21_X1 U21403 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18147), .A(
        n18146), .ZN(n19195) );
  XOR2_X1 U21404 ( .A(n18160), .B(n19195), .Z(n18151) );
  OAI211_X1 U21405 ( .C1(n18149), .C2(n18155), .A(n18171), .B(n18148), .ZN(
        n18150) );
  OAI211_X1 U21406 ( .C1(n13366), .C2(n18151), .A(n19428), .B(n18150), .ZN(
        n18152) );
  AOI211_X1 U21407 ( .C1(n18193), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n18153), .B(n18152), .ZN(n18154) );
  OAI21_X1 U21408 ( .B1(n18158), .B2(n18155), .A(n18154), .ZN(P3_U2666) );
  NAND2_X1 U21409 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18212), .ZN(n18206) );
  OAI21_X1 U21410 ( .B1(n18157), .B2(n18206), .A(n18156), .ZN(n18192) );
  OAI21_X1 U21411 ( .B1(n18226), .B2(n18170), .A(n18158), .ZN(n18175) );
  NOR2_X1 U21412 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17459), .ZN(
        n18161) );
  INV_X1 U21413 ( .A(n18159), .ZN(n18164) );
  AOI22_X1 U21414 ( .A1(n18197), .A2(n18161), .B1(n18160), .B2(n18164), .ZN(
        n18162) );
  OAI22_X1 U21415 ( .A1(n18162), .A2(n13366), .B1(n17460), .B2(n18219), .ZN(
        n18167) );
  INV_X1 U21416 ( .A(n18163), .ZN(n18199) );
  NOR2_X1 U21417 ( .A1(n18199), .A2(n18164), .ZN(n18166) );
  AOI21_X1 U21418 ( .B1(n19961), .B2(n18258), .A(n18214), .ZN(n18165) );
  OR4_X1 U21419 ( .A1(n18167), .A2(n19477), .A3(n18166), .A4(n18165), .ZN(
        n18174) );
  NAND2_X1 U21420 ( .A1(n18169), .A2(n18168), .ZN(n18172) );
  NAND2_X1 U21421 ( .A1(n18171), .A2(n18170), .ZN(n18184) );
  OAI22_X1 U21422 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18172), .B1(
        P3_EBX_REG_4__SCAN_IN), .B2(n18184), .ZN(n18173) );
  AOI211_X1 U21423 ( .C1(n18175), .C2(P3_EBX_REG_4__SCAN_IN), .A(n18174), .B(
        n18173), .ZN(n18176) );
  OAI21_X1 U21424 ( .B1(n20008), .B2(n18192), .A(n18176), .ZN(P3_U2667) );
  INV_X1 U21425 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U21426 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n18191) );
  INV_X1 U21427 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21725) );
  NOR2_X1 U21428 ( .A1(n18177), .A2(n21725), .ZN(n18196) );
  AOI21_X1 U21429 ( .B1(n18196), .B2(n18221), .A(n9750), .ZN(n18180) );
  OAI21_X1 U21430 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18196), .A(
        n18179), .ZN(n19204) );
  XNOR2_X1 U21431 ( .A(n18180), .B(n19204), .ZN(n18188) );
  NOR4_X1 U21432 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n20006), .A3(n18205), .A4(
        n13863), .ZN(n18187) );
  NOR2_X1 U21433 ( .A1(n18194), .A2(n18181), .ZN(n18185) );
  AOI21_X1 U21434 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18182), .A(
        n9723), .ZN(n18183) );
  OAI22_X1 U21435 ( .A1(n18185), .A2(n18184), .B1(n18183), .B2(n18214), .ZN(
        n18186) );
  AOI211_X1 U21436 ( .C1(n18189), .C2(n18188), .A(n18187), .B(n18186), .ZN(
        n18190) );
  OAI211_X1 U21437 ( .C1(n20007), .C2(n18192), .A(n18191), .B(n18190), .ZN(
        P3_U2668) );
  AOI22_X1 U21438 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18193), .B1(
        n18217), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n18210) );
  OR2_X1 U21439 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n18211) );
  AOI211_X1 U21440 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18211), .A(n18194), .B(
        n18226), .ZN(n18204) );
  AND2_X1 U21441 ( .A1(n20107), .A2(n18195), .ZN(n18202) );
  INV_X1 U21442 ( .A(n18196), .ZN(n18198) );
  OAI21_X1 U21443 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18198), .ZN(n19222) );
  OAI22_X1 U21444 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18198), .B1(
        n18197), .B2(n19222), .ZN(n18200) );
  OAI22_X1 U21445 ( .A1(n18220), .A2(n18200), .B1(n19222), .B2(n18199), .ZN(
        n18201) );
  OR2_X1 U21446 ( .A1(n18202), .A2(n18201), .ZN(n18203) );
  NOR2_X1 U21447 ( .A1(n18204), .A2(n18203), .ZN(n18209) );
  NOR2_X1 U21448 ( .A1(n18205), .A2(n13863), .ZN(n18207) );
  NOR2_X1 U21449 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18205), .ZN(n18216) );
  OAI22_X1 U21450 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18207), .B1(n18216), 
        .B2(n18206), .ZN(n18208) );
  NAND3_X1 U21451 ( .A1(n18210), .A2(n18209), .A3(n18208), .ZN(P3_U2669) );
  NAND2_X1 U21452 ( .A1(n18211), .A2(n18636), .ZN(n18643) );
  OAI22_X1 U21453 ( .A1(n18214), .A2(n18213), .B1(n13863), .B2(n18212), .ZN(
        n18215) );
  AOI211_X1 U21454 ( .C1(P3_EBX_REG_1__SCAN_IN), .C2(n18217), .A(n18216), .B(
        n18215), .ZN(n18225) );
  INV_X1 U21455 ( .A(n18218), .ZN(n18223) );
  OAI211_X1 U21456 ( .C1(n18221), .C2(n18220), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n18219), .ZN(n18222) );
  OAI21_X1 U21457 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18223), .A(
        n18222), .ZN(n18224) );
  OAI211_X1 U21458 ( .C1(n18226), .C2(n18643), .A(n18225), .B(n18224), .ZN(
        P3_U2670) );
  NAND2_X1 U21459 ( .A1(n18228), .A2(n18227), .ZN(n18229) );
  NAND2_X1 U21460 ( .A1(n18229), .A2(n18642), .ZN(n18354) );
  AOI22_X1 U21461 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18234) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18570), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11842), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U21464 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18231) );
  NAND4_X1 U21465 ( .A1(n18234), .A2(n18233), .A3(n18232), .A4(n18231), .ZN(
        n18243) );
  INV_X1 U21466 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U21467 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18236) );
  NAND2_X1 U21468 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n18235) );
  OAI211_X1 U21469 ( .C1(n9745), .C2(n18237), .A(n18236), .B(n18235), .ZN(
        n18238) );
  INV_X1 U21470 ( .A(n18238), .ZN(n18241) );
  AOI22_X1 U21471 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18240) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18613), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18239) );
  NAND3_X1 U21473 ( .A1(n18241), .A2(n18240), .A3(n18239), .ZN(n18242) );
  NOR2_X1 U21474 ( .A1(n18243), .A2(n18242), .ZN(n18365) );
  INV_X1 U21475 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U21476 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18245) );
  NAND2_X1 U21477 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n18244) );
  OAI211_X1 U21478 ( .C1(n18246), .C2(n9744), .A(n18245), .B(n18244), .ZN(
        n18247) );
  INV_X1 U21479 ( .A(n18247), .ZN(n18250) );
  AOI22_X1 U21480 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U21481 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18248) );
  NAND3_X1 U21482 ( .A1(n18250), .A2(n18249), .A3(n18248), .ZN(n18257) );
  AOI22_X1 U21483 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18255) );
  AOI22_X1 U21484 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18254) );
  AOI22_X1 U21485 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U21486 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18252) );
  NAND4_X1 U21487 ( .A1(n18255), .A2(n18254), .A3(n18253), .A4(n18252), .ZN(
        n18256) );
  NOR2_X1 U21488 ( .A1(n18257), .A2(n18256), .ZN(n18373) );
  INV_X1 U21489 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18262) );
  AOI22_X1 U21490 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18260) );
  NAND2_X1 U21491 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n18259) );
  OAI211_X1 U21492 ( .C1(n18262), .C2(n18261), .A(n18260), .B(n18259), .ZN(
        n18263) );
  INV_X1 U21493 ( .A(n18263), .ZN(n18266) );
  AOI22_X1 U21494 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18265) );
  AOI22_X1 U21495 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18264) );
  NAND3_X1 U21496 ( .A1(n18266), .A2(n18265), .A3(n18264), .ZN(n18272) );
  AOI22_X1 U21497 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9728), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U21498 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U21499 ( .A1(n10603), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18268) );
  AOI22_X1 U21500 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18267) );
  NAND4_X1 U21501 ( .A1(n18270), .A2(n18269), .A3(n18268), .A4(n18267), .ZN(
        n18271) );
  NOR2_X1 U21502 ( .A1(n18272), .A2(n18271), .ZN(n18383) );
  AOI22_X1 U21503 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U21504 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U21505 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U21506 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18273) );
  NAND4_X1 U21507 ( .A1(n18276), .A2(n18275), .A3(n18274), .A4(n18273), .ZN(
        n18285) );
  INV_X1 U21508 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U21509 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18517), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18278) );
  NAND2_X1 U21510 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n18277) );
  OAI211_X1 U21511 ( .C1(n18279), .C2(n9726), .A(n18278), .B(n18277), .ZN(
        n18280) );
  INV_X1 U21512 ( .A(n18280), .ZN(n18283) );
  AOI22_X1 U21513 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18282) );
  AOI22_X1 U21514 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18281) );
  NAND3_X1 U21515 ( .A1(n18283), .A2(n18282), .A3(n18281), .ZN(n18284) );
  NOR2_X1 U21516 ( .A1(n18285), .A2(n18284), .ZN(n18382) );
  NOR2_X1 U21517 ( .A1(n18383), .A2(n18382), .ZN(n18378) );
  INV_X1 U21518 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18288) );
  NAND2_X1 U21519 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n18287) );
  AOI22_X1 U21520 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18286) );
  OAI211_X1 U21521 ( .C1(n18288), .C2(n9726), .A(n18287), .B(n18286), .ZN(
        n18299) );
  AOI22_X1 U21522 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U21523 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10603), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U21524 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18290) );
  AOI22_X1 U21525 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18289) );
  NAND4_X1 U21526 ( .A1(n18292), .A2(n18291), .A3(n18290), .A4(n18289), .ZN(
        n18298) );
  INV_X1 U21527 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18294) );
  INV_X1 U21528 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18293) );
  OAI22_X1 U21529 ( .A1(n18410), .A2(n18294), .B1(n18505), .B2(n18293), .ZN(
        n18297) );
  INV_X1 U21530 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18591) );
  INV_X1 U21531 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18295) );
  OAI22_X1 U21532 ( .A1(n18440), .A2(n18591), .B1(n18261), .B2(n18295), .ZN(
        n18296) );
  OR4_X1 U21533 ( .A1(n18299), .A2(n18298), .A3(n18297), .A4(n18296), .ZN(
        n18377) );
  NAND2_X1 U21534 ( .A1(n18378), .A2(n18377), .ZN(n18376) );
  NOR2_X1 U21535 ( .A1(n18373), .A2(n18376), .ZN(n18370) );
  INV_X1 U21536 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18302) );
  NAND2_X1 U21537 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n18301) );
  AOI22_X1 U21538 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18300) );
  OAI211_X1 U21539 ( .C1(n18302), .C2(n9745), .A(n18301), .B(n18300), .ZN(
        n18313) );
  AOI22_X1 U21540 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U21541 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U21542 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18304) );
  AOI22_X1 U21543 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18303) );
  NAND4_X1 U21544 ( .A1(n18306), .A2(n18305), .A3(n18304), .A4(n18303), .ZN(
        n18312) );
  INV_X1 U21545 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18308) );
  INV_X1 U21546 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18307) );
  OAI22_X1 U21547 ( .A1(n18410), .A2(n18308), .B1(n18505), .B2(n18307), .ZN(
        n18311) );
  INV_X1 U21548 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18309) );
  INV_X1 U21549 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n21548) );
  OAI22_X1 U21550 ( .A1(n18440), .A2(n18309), .B1(n18261), .B2(n21548), .ZN(
        n18310) );
  OR4_X1 U21551 ( .A1(n18313), .A2(n18312), .A3(n18311), .A4(n18310), .ZN(
        n18369) );
  NAND2_X1 U21552 ( .A1(n18370), .A2(n18369), .ZN(n18368) );
  NOR2_X1 U21553 ( .A1(n18365), .A2(n18368), .ZN(n18362) );
  INV_X1 U21554 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18316) );
  NAND2_X1 U21555 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n18315) );
  AOI22_X1 U21556 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18314) );
  OAI211_X1 U21557 ( .C1(n18316), .C2(n9726), .A(n18315), .B(n18314), .ZN(
        n18326) );
  AOI22_X1 U21558 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U21559 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U21560 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U21561 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18318) );
  NAND4_X1 U21562 ( .A1(n18321), .A2(n18320), .A3(n18319), .A4(n18318), .ZN(
        n18325) );
  INV_X1 U21563 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18322) );
  INV_X1 U21564 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18403) );
  OAI22_X1 U21565 ( .A1(n18410), .A2(n18322), .B1(n18505), .B2(n18403), .ZN(
        n18324) );
  INV_X1 U21566 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18409) );
  INV_X1 U21567 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n21569) );
  OAI22_X1 U21568 ( .A1(n18440), .A2(n18409), .B1(n18261), .B2(n21569), .ZN(
        n18323) );
  OR4_X1 U21569 ( .A1(n18326), .A2(n18325), .A3(n18324), .A4(n18323), .ZN(
        n18361) );
  NAND2_X1 U21570 ( .A1(n18362), .A2(n18361), .ZN(n18360) );
  AOI22_X1 U21571 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U21572 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U21573 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U21574 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18327) );
  NAND4_X1 U21575 ( .A1(n18330), .A2(n18329), .A3(n18328), .A4(n18327), .ZN(
        n18339) );
  INV_X1 U21576 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U21577 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18332) );
  NAND2_X1 U21578 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n18331) );
  OAI211_X1 U21579 ( .C1(n18333), .C2(n9745), .A(n18332), .B(n18331), .ZN(
        n18334) );
  INV_X1 U21580 ( .A(n18334), .ZN(n18337) );
  AOI22_X1 U21581 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U21582 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18335) );
  NAND3_X1 U21583 ( .A1(n18337), .A2(n18336), .A3(n18335), .ZN(n18338) );
  NOR2_X1 U21584 ( .A1(n18339), .A2(n18338), .ZN(n18357) );
  NOR2_X1 U21585 ( .A1(n18360), .A2(n18357), .ZN(n18353) );
  AOI22_X1 U21586 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18343) );
  AOI22_X1 U21587 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18342) );
  AOI22_X1 U21588 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18341) );
  AOI22_X1 U21589 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18340) );
  NAND4_X1 U21590 ( .A1(n18343), .A2(n18342), .A3(n18341), .A4(n18340), .ZN(
        n18351) );
  INV_X1 U21591 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U21592 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18344) );
  OAI21_X1 U21593 ( .B1(n18261), .B2(n18345), .A(n18344), .ZN(n18346) );
  AOI21_X1 U21594 ( .B1(n9723), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n18346), .ZN(n18349) );
  AOI22_X1 U21595 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18348) );
  AOI22_X1 U21596 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18347) );
  NAND3_X1 U21597 ( .A1(n18349), .A2(n18348), .A3(n18347), .ZN(n18350) );
  NOR2_X1 U21598 ( .A1(n18351), .A2(n18350), .ZN(n18352) );
  XOR2_X1 U21599 ( .A(n18353), .B(n18352), .Z(n18664) );
  OAI22_X1 U21600 ( .A1(n18355), .A2(n18354), .B1(n18664), .B2(n18638), .ZN(
        P3_U2673) );
  INV_X1 U21601 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n18356) );
  NAND3_X1 U21602 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18372), .ZN(n18359) );
  XNOR2_X1 U21603 ( .A(n18357), .B(n18360), .ZN(n18668) );
  NAND3_X1 U21604 ( .A1(n18359), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18642), 
        .ZN(n18358) );
  OAI221_X1 U21605 ( .B1(n18359), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18642), 
        .C2(n18668), .A(n18358), .ZN(P3_U2674) );
  INV_X1 U21606 ( .A(n18359), .ZN(n18364) );
  AOI22_X1 U21607 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18642), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(n18372), .ZN(n18363) );
  OAI21_X1 U21608 ( .B1(n18362), .B2(n18361), .A(n18360), .ZN(n18672) );
  OAI22_X1 U21609 ( .A1(n18364), .A2(n18363), .B1(n18642), .B2(n18672), .ZN(
        P3_U2675) );
  XNOR2_X1 U21610 ( .A(n18365), .B(n18368), .ZN(n18676) );
  NAND3_X1 U21611 ( .A1(n18367), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18642), 
        .ZN(n18366) );
  OAI221_X1 U21612 ( .B1(n18367), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18638), 
        .C2(n18676), .A(n18366), .ZN(P3_U2676) );
  AOI21_X1 U21613 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18642), .A(n18375), .ZN(
        n18371) );
  OAI21_X1 U21614 ( .B1(n18370), .B2(n18369), .A(n18368), .ZN(n18681) );
  OAI22_X1 U21615 ( .A1(n18372), .A2(n18371), .B1(n18642), .B2(n18681), .ZN(
        P3_U2677) );
  AOI21_X1 U21616 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18642), .A(n18380), .ZN(
        n18374) );
  XNOR2_X1 U21617 ( .A(n18373), .B(n18376), .ZN(n18686) );
  OAI22_X1 U21618 ( .A1(n18375), .A2(n18374), .B1(n18642), .B2(n18686), .ZN(
        P3_U2678) );
  AOI21_X1 U21619 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18642), .A(n9775), .ZN(
        n18379) );
  OAI21_X1 U21620 ( .B1(n18378), .B2(n18377), .A(n18376), .ZN(n18691) );
  OAI22_X1 U21621 ( .A1(n18380), .A2(n18379), .B1(n18642), .B2(n18691), .ZN(
        P3_U2679) );
  AOI21_X1 U21622 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18642), .A(n18381), .ZN(
        n18384) );
  XNOR2_X1 U21623 ( .A(n18383), .B(n18382), .ZN(n18696) );
  OAI22_X1 U21624 ( .A1(n9775), .A2(n18384), .B1(n18642), .B2(n18696), .ZN(
        P3_U2680) );
  INV_X1 U21625 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18387) );
  AOI22_X1 U21626 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18386) );
  NAND2_X1 U21627 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n18385) );
  OAI211_X1 U21628 ( .C1(n18387), .C2(n9744), .A(n18386), .B(n18385), .ZN(
        n18388) );
  INV_X1 U21629 ( .A(n18388), .ZN(n18391) );
  AOI22_X1 U21630 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18390) );
  AOI22_X1 U21631 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18389) );
  NAND3_X1 U21632 ( .A1(n18391), .A2(n18390), .A3(n18389), .ZN(n18397) );
  AOI22_X1 U21633 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U21634 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U21635 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18393) );
  AOI22_X1 U21636 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18392) );
  NAND4_X1 U21637 ( .A1(n18395), .A2(n18394), .A3(n18393), .A4(n18392), .ZN(
        n18396) );
  NOR2_X1 U21638 ( .A1(n18397), .A2(n18396), .ZN(n18698) );
  NAND3_X1 U21639 ( .A1(n18399), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n18642), 
        .ZN(n18398) );
  OAI221_X1 U21640 ( .B1(n18399), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n18638), 
        .C2(n18698), .A(n18398), .ZN(P3_U2681) );
  NAND2_X1 U21641 ( .A1(n18642), .A2(n18400), .ZN(n18433) );
  NAND2_X1 U21642 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n18402) );
  AOI22_X1 U21643 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18401) );
  OAI211_X1 U21644 ( .C1(n18403), .C2(n9745), .A(n18402), .B(n18401), .ZN(
        n18416) );
  AOI22_X1 U21645 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18407) );
  AOI22_X1 U21646 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U21647 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U21648 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18404) );
  NAND4_X1 U21649 ( .A1(n18407), .A2(n18406), .A3(n18405), .A4(n18404), .ZN(
        n18415) );
  OAI22_X1 U21650 ( .A1(n18410), .A2(n18409), .B1(n18505), .B2(n18408), .ZN(
        n18414) );
  INV_X1 U21651 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18412) );
  INV_X1 U21652 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18411) );
  OAI22_X1 U21653 ( .A1(n18440), .A2(n18412), .B1(n18261), .B2(n18411), .ZN(
        n18413) );
  OR4_X1 U21654 ( .A1(n18416), .A2(n18415), .A3(n18414), .A4(n18413), .ZN(
        n18703) );
  AOI22_X1 U21655 ( .A1(n18648), .A2(n18703), .B1(n18417), .B2(n18419), .ZN(
        n18418) );
  OAI21_X1 U21656 ( .B1(n18419), .B2(n18433), .A(n18418), .ZN(P3_U2682) );
  NOR2_X1 U21657 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n9816), .ZN(n18434) );
  INV_X1 U21658 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18422) );
  AOI22_X1 U21659 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18421) );
  NAND2_X1 U21660 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n18420) );
  OAI211_X1 U21661 ( .C1(n9726), .C2(n18422), .A(n18421), .B(n18420), .ZN(
        n18423) );
  INV_X1 U21662 ( .A(n18423), .ZN(n18426) );
  AOI22_X1 U21663 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U21664 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18424) );
  NAND3_X1 U21665 ( .A1(n18426), .A2(n18425), .A3(n18424), .ZN(n18432) );
  AOI22_X1 U21666 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U21667 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11802), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18429) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18565), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18428) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9728), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18427) );
  NAND4_X1 U21670 ( .A1(n18430), .A2(n18429), .A3(n18428), .A4(n18427), .ZN(
        n18431) );
  NOR2_X1 U21671 ( .A1(n18432), .A2(n18431), .ZN(n18709) );
  OAI22_X1 U21672 ( .A1(n18434), .A2(n18433), .B1(n18709), .B2(n18638), .ZN(
        P3_U2683) );
  INV_X1 U21673 ( .A(n18465), .ZN(n18435) );
  OAI21_X1 U21674 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18435), .A(n18642), .ZN(
        n18450) );
  INV_X1 U21675 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18437) );
  AOI22_X1 U21676 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18436) );
  OAI21_X1 U21677 ( .B1(n18261), .B2(n18437), .A(n18436), .ZN(n18438) );
  AOI21_X1 U21678 ( .B1(n9729), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n18438), .ZN(n18443) );
  AOI22_X1 U21679 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U21680 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18441) );
  NAND3_X1 U21681 ( .A1(n18443), .A2(n18442), .A3(n18441), .ZN(n18449) );
  AOI22_X1 U21682 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18517), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18447) );
  AOI22_X1 U21683 ( .A1(n9743), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18446) );
  AOI22_X1 U21684 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18445) );
  AOI22_X1 U21685 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18444) );
  NAND4_X1 U21686 ( .A1(n18447), .A2(n18446), .A3(n18445), .A4(n18444), .ZN(
        n18448) );
  NOR2_X1 U21687 ( .A1(n18449), .A2(n18448), .ZN(n18718) );
  OAI22_X1 U21688 ( .A1(n9816), .A2(n18450), .B1(n18718), .B2(n18638), .ZN(
        P3_U2684) );
  AOI22_X1 U21689 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18454) );
  AOI22_X1 U21690 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18453) );
  AOI22_X1 U21691 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18452) );
  AOI22_X1 U21692 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18451) );
  NAND4_X1 U21693 ( .A1(n18454), .A2(n18453), .A3(n18452), .A4(n18451), .ZN(
        n18463) );
  INV_X1 U21694 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U21695 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18456) );
  NAND2_X1 U21696 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n18455) );
  OAI211_X1 U21697 ( .C1(n18457), .C2(n9744), .A(n18456), .B(n18455), .ZN(
        n18458) );
  INV_X1 U21698 ( .A(n18458), .ZN(n18461) );
  AOI22_X1 U21699 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18460) );
  AOI22_X1 U21700 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18459) );
  NAND3_X1 U21701 ( .A1(n18461), .A2(n18460), .A3(n18459), .ZN(n18462) );
  NOR2_X1 U21702 ( .A1(n18463), .A2(n18462), .ZN(n18722) );
  NAND2_X1 U21703 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .ZN(n21547) );
  NAND2_X1 U21704 ( .A1(n19521), .A2(n18464), .ZN(n18481) );
  NOR2_X1 U21705 ( .A1(n21547), .A2(n18481), .ZN(n18480) );
  OAI21_X1 U21706 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n18480), .A(n18465), .ZN(
        n18466) );
  AOI22_X1 U21707 ( .A1(n18648), .A2(n18722), .B1(n18466), .B2(n18642), .ZN(
        P3_U2685) );
  INV_X1 U21708 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n21504) );
  NOR2_X1 U21709 ( .A1(n21504), .A2(n18481), .ZN(n18496) );
  AOI21_X1 U21710 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18642), .A(n18496), .ZN(
        n18479) );
  INV_X1 U21711 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18468) );
  AOI22_X1 U21712 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18467) );
  OAI21_X1 U21713 ( .B1(n18261), .B2(n18468), .A(n18467), .ZN(n18469) );
  AOI21_X1 U21714 ( .B1(n9723), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n18469), .ZN(n18472) );
  AOI22_X1 U21715 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18471) );
  AOI22_X1 U21716 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18470) );
  NAND3_X1 U21717 ( .A1(n18472), .A2(n18471), .A3(n18470), .ZN(n18478) );
  AOI22_X1 U21718 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18476) );
  AOI22_X1 U21719 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18475) );
  AOI22_X1 U21720 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18474) );
  AOI22_X1 U21721 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18473) );
  NAND4_X1 U21722 ( .A1(n18476), .A2(n18475), .A3(n18474), .A4(n18473), .ZN(
        n18477) );
  NOR2_X1 U21723 ( .A1(n18478), .A2(n18477), .ZN(n18728) );
  OAI22_X1 U21724 ( .A1(n18480), .A2(n18479), .B1(n18728), .B2(n18638), .ZN(
        P3_U2686) );
  INV_X1 U21725 ( .A(n18481), .ZN(n18513) );
  AOI21_X1 U21726 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18642), .A(n18513), .ZN(
        n18495) );
  AOI22_X1 U21727 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18485) );
  AOI22_X1 U21728 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11842), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18484) );
  AOI22_X1 U21729 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18483) );
  AOI22_X1 U21730 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18482) );
  NAND4_X1 U21731 ( .A1(n18485), .A2(n18484), .A3(n18483), .A4(n18482), .ZN(
        n18494) );
  INV_X1 U21732 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U21733 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18487) );
  NAND2_X1 U21734 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n18486) );
  OAI211_X1 U21735 ( .C1(n18488), .C2(n9744), .A(n18487), .B(n18486), .ZN(
        n18489) );
  INV_X1 U21736 ( .A(n18489), .ZN(n18492) );
  AOI22_X1 U21737 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18491) );
  AOI22_X1 U21738 ( .A1(n11825), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18490) );
  NAND3_X1 U21739 ( .A1(n18492), .A2(n18491), .A3(n18490), .ZN(n18493) );
  NOR2_X1 U21740 ( .A1(n18494), .A2(n18493), .ZN(n18734) );
  OAI22_X1 U21741 ( .A1(n18496), .A2(n18495), .B1(n18734), .B2(n18638), .ZN(
        P3_U2687) );
  AOI22_X1 U21742 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U21743 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18501) );
  AOI22_X1 U21744 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18500) );
  AOI22_X1 U21745 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18499) );
  NAND4_X1 U21746 ( .A1(n18502), .A2(n18501), .A3(n18500), .A4(n18499), .ZN(
        n18512) );
  AOI22_X1 U21747 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18504) );
  NAND2_X1 U21748 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n18503) );
  OAI211_X1 U21749 ( .C1(n18506), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        n18507) );
  INV_X1 U21750 ( .A(n18507), .ZN(n18510) );
  AOI22_X1 U21751 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U21752 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18508) );
  NAND3_X1 U21753 ( .A1(n18510), .A2(n18509), .A3(n18508), .ZN(n18511) );
  NOR2_X1 U21754 ( .A1(n18512), .A2(n18511), .ZN(n18738) );
  AOI21_X1 U21755 ( .B1(n18514), .B2(n18531), .A(n18513), .ZN(n18515) );
  INV_X1 U21756 ( .A(n18515), .ZN(n18516) );
  AOI22_X1 U21757 ( .A1(n18648), .A2(n18738), .B1(n18516), .B2(n18642), .ZN(
        P3_U2688) );
  INV_X1 U21758 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18520) );
  AOI22_X1 U21759 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18517), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18519) );
  NAND2_X1 U21760 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n18518) );
  OAI211_X1 U21761 ( .C1(n18520), .C2(n9745), .A(n18519), .B(n18518), .ZN(
        n18521) );
  INV_X1 U21762 ( .A(n18521), .ZN(n18524) );
  AOI22_X1 U21763 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18523) );
  AOI22_X1 U21764 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18522) );
  NAND3_X1 U21765 ( .A1(n18524), .A2(n18523), .A3(n18522), .ZN(n18530) );
  AOI22_X1 U21766 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18606), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18528) );
  AOI22_X1 U21767 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18614), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U21768 ( .A1(n11802), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18526) );
  AOI22_X1 U21769 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18525) );
  NAND4_X1 U21770 ( .A1(n18528), .A2(n18527), .A3(n18526), .A4(n18525), .ZN(
        n18529) );
  NOR2_X1 U21771 ( .A1(n18530), .A2(n18529), .ZN(n18744) );
  OAI21_X1 U21772 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18532), .A(n18531), .ZN(
        n18533) );
  AOI22_X1 U21773 ( .A1(n18648), .A2(n18744), .B1(n18533), .B2(n18642), .ZN(
        P3_U2689) );
  INV_X1 U21774 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18536) );
  AOI22_X1 U21775 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18535) );
  NAND2_X1 U21776 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n18534) );
  OAI211_X1 U21777 ( .C1(n9726), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        n18537) );
  INV_X1 U21778 ( .A(n18537), .ZN(n18540) );
  AOI22_X1 U21779 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18539) );
  AOI22_X1 U21780 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18538) );
  NAND3_X1 U21781 ( .A1(n18540), .A2(n18539), .A3(n18538), .ZN(n18546) );
  AOI22_X1 U21782 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18544) );
  AOI22_X1 U21783 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U21784 ( .A1(n18517), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11802), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18542) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9728), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18541) );
  NAND4_X1 U21786 ( .A1(n18544), .A2(n18543), .A3(n18542), .A4(n18541), .ZN(
        n18545) );
  NOR2_X1 U21787 ( .A1(n18546), .A2(n18545), .ZN(n18749) );
  OAI211_X1 U21788 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n9817), .A(n18547), .B(
        n18642), .ZN(n18548) );
  OAI21_X1 U21789 ( .B1(n18749), .B2(n18642), .A(n18548), .ZN(P3_U2691) );
  INV_X1 U21790 ( .A(n18581), .ZN(n18549) );
  OAI21_X1 U21791 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18549), .A(n18638), .ZN(
        n18563) );
  INV_X1 U21792 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18552) );
  AOI22_X1 U21793 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18551) );
  NAND2_X1 U21794 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n18550) );
  OAI211_X1 U21795 ( .C1(n18552), .C2(n9744), .A(n18551), .B(n18550), .ZN(
        n18553) );
  INV_X1 U21796 ( .A(n18553), .ZN(n18556) );
  AOI22_X1 U21797 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18555) );
  AOI22_X1 U21798 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18554) );
  NAND3_X1 U21799 ( .A1(n18556), .A2(n18555), .A3(n18554), .ZN(n18562) );
  AOI22_X1 U21800 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18560) );
  AOI22_X1 U21801 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18559) );
  AOI22_X1 U21802 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18558) );
  AOI22_X1 U21803 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18557) );
  NAND4_X1 U21804 ( .A1(n18560), .A2(n18559), .A3(n18558), .A4(n18557), .ZN(
        n18561) );
  NOR2_X1 U21805 ( .A1(n18562), .A2(n18561), .ZN(n18753) );
  OAI22_X1 U21806 ( .A1(n9817), .A2(n18563), .B1(n18753), .B2(n18638), .ZN(
        P3_U2692) );
  AOI22_X1 U21807 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18569) );
  AOI22_X1 U21808 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18610), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18568) );
  AOI22_X1 U21809 ( .A1(n18564), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18439), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18567) );
  AOI22_X1 U21810 ( .A1(n18565), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11843), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18566) );
  NAND4_X1 U21811 ( .A1(n18569), .A2(n18568), .A3(n18567), .A4(n18566), .ZN(
        n18580) );
  INV_X1 U21812 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18573) );
  NAND2_X1 U21813 ( .A1(n18570), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n18572) );
  NAND2_X1 U21814 ( .A1(n18251), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n18571) );
  OAI211_X1 U21815 ( .C1(n18573), .C2(n9726), .A(n18572), .B(n18571), .ZN(
        n18574) );
  INV_X1 U21816 ( .A(n18574), .ZN(n18578) );
  INV_X1 U21817 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21715) );
  AOI22_X1 U21818 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18577) );
  AOI22_X1 U21819 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18576) );
  NAND2_X1 U21820 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n18575) );
  NAND4_X1 U21821 ( .A1(n18578), .A2(n18577), .A3(n18576), .A4(n18575), .ZN(
        n18579) );
  NOR2_X1 U21822 ( .A1(n18580), .A2(n18579), .ZN(n18756) );
  OAI21_X1 U21823 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18601), .A(n18581), .ZN(
        n18582) );
  AOI22_X1 U21824 ( .A1(n18648), .A2(n18756), .B1(n18582), .B2(n18638), .ZN(
        P3_U2693) );
  INV_X1 U21825 ( .A(n18621), .ZN(n18583) );
  OAI21_X1 U21826 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18583), .A(n18638), .ZN(
        n18600) );
  AOI22_X1 U21827 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18517), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18587) );
  AOI22_X1 U21828 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18586) );
  AOI22_X1 U21829 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17549), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U21830 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18584) );
  NAND4_X1 U21831 ( .A1(n18587), .A2(n18586), .A3(n18585), .A4(n18584), .ZN(
        n18599) );
  INV_X1 U21832 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18590) );
  AOI22_X1 U21833 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18589) );
  NAND2_X1 U21834 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n18588) );
  OAI211_X1 U21835 ( .C1(n18590), .C2(n9726), .A(n18589), .B(n18588), .ZN(
        n18597) );
  INV_X1 U21836 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n21570) );
  OAI22_X1 U21837 ( .A1(n18592), .A2(n18591), .B1(n10540), .B2(n21570), .ZN(
        n18596) );
  INV_X1 U21838 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18594) );
  INV_X1 U21839 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18593) );
  OAI22_X1 U21840 ( .A1(n18440), .A2(n18594), .B1(n10539), .B2(n18593), .ZN(
        n18595) );
  OR3_X1 U21841 ( .A1(n18597), .A2(n18596), .A3(n18595), .ZN(n18598) );
  NOR2_X1 U21842 ( .A1(n18599), .A2(n18598), .ZN(n18762) );
  OAI22_X1 U21843 ( .A1(n18601), .A2(n18600), .B1(n18762), .B2(n18638), .ZN(
        P3_U2694) );
  INV_X1 U21844 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18604) );
  AOI22_X1 U21845 ( .A1(n11842), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18570), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18603) );
  NAND2_X1 U21846 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n18602) );
  OAI211_X1 U21847 ( .C1(n18604), .C2(n9745), .A(n18603), .B(n18602), .ZN(
        n18605) );
  INV_X1 U21848 ( .A(n18605), .ZN(n18609) );
  AOI22_X1 U21849 ( .A1(n18606), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18608) );
  AOI22_X1 U21850 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18565), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18607) );
  NAND3_X1 U21851 ( .A1(n18609), .A2(n18608), .A3(n18607), .ZN(n18620) );
  AOI22_X1 U21852 ( .A1(n18610), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18618) );
  AOI22_X1 U21853 ( .A1(n11841), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18611), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18617) );
  AOI22_X1 U21854 ( .A1(n18613), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18612), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18616) );
  AOI22_X1 U21855 ( .A1(n18614), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18251), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18615) );
  NAND4_X1 U21856 ( .A1(n18618), .A2(n18617), .A3(n18616), .A4(n18615), .ZN(
        n18619) );
  NOR2_X1 U21857 ( .A1(n18620), .A2(n18619), .ZN(n18765) );
  NOR2_X1 U21858 ( .A1(n18629), .A2(n18626), .ZN(n18623) );
  OAI221_X1 U21859 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n18623), .A(n18621), .ZN(n18622) );
  AOI22_X1 U21860 ( .A1(n18648), .A2(n18765), .B1(n18622), .B2(n18638), .ZN(
        P3_U2695) );
  OAI21_X1 U21861 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18623), .A(n18642), .ZN(
        n18624) );
  OAI22_X1 U21862 ( .A1(n18625), .A2(n18624), .B1(n18345), .B2(n18638), .ZN(
        P3_U2696) );
  NAND2_X1 U21863 ( .A1(n18642), .A2(n18626), .ZN(n18630) );
  NOR2_X1 U21864 ( .A1(n18697), .A2(n18626), .ZN(n18627) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18648), .B1(
        n18627), .B2(n18629), .ZN(n18628) );
  OAI21_X1 U21866 ( .B1(n18629), .B2(n18630), .A(n18628), .ZN(P3_U2697) );
  NOR2_X1 U21867 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18635), .ZN(n18631) );
  OAI22_X1 U21868 ( .A1(n18631), .A2(n18630), .B1(n21569), .B2(n18638), .ZN(
        P3_U2698) );
  OAI21_X1 U21869 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18632), .A(n18638), .ZN(
        n18634) );
  INV_X1 U21870 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18633) );
  OAI22_X1 U21871 ( .A1(n18635), .A2(n18634), .B1(n18633), .B2(n18638), .ZN(
        P3_U2699) );
  NOR2_X1 U21872 ( .A1(n18697), .A2(n18644), .ZN(n18647) );
  NAND3_X1 U21873 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n10138), .A3(n18647), .ZN(
        n18639) );
  NAND3_X1 U21874 ( .A1(n18639), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n18642), .ZN(
        n18637) );
  OAI221_X1 U21875 ( .B1(n18639), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n18638), 
        .C2(n21548), .A(n18637), .ZN(P3_U2700) );
  INV_X1 U21876 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18641) );
  OAI211_X1 U21877 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n9851), .A(n18639), .B(
        n18642), .ZN(n18640) );
  OAI21_X1 U21878 ( .B1(n18642), .B2(n18641), .A(n18640), .ZN(P3_U2701) );
  INV_X1 U21879 ( .A(n18643), .ZN(n18645) );
  AOI222_X1 U21880 ( .A1(n18647), .A2(n18645), .B1(P3_EBX_REG_1__SCAN_IN), 
        .B2(n18644), .C1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .C2(n18648), .ZN(
        n18646) );
  INV_X1 U21881 ( .A(n18646), .ZN(P3_U2702) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18648), .B1(
        n18647), .B2(n18650), .ZN(n18649) );
  OAI21_X1 U21883 ( .B1(n18651), .B2(n18650), .A(n18649), .ZN(P3_U2703) );
  INV_X1 U21884 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18806) );
  INV_X1 U21885 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21622) );
  INV_X1 U21886 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n21565) );
  NAND2_X1 U21887 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n18768) );
  INV_X1 U21888 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18840) );
  NOR4_X1 U21889 ( .A1(n21565), .A2(n18652), .A3(n18768), .A4(n18840), .ZN(
        n18653) );
  NAND3_X1 U21890 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n18653), .ZN(n18740) );
  NAND4_X1 U21891 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n18654)
         );
  NAND4_X1 U21892 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n18656), .ZN(n18741) );
  NOR2_X2 U21893 ( .A1(n18741), .A2(n18908), .ZN(n18735) );
  INV_X1 U21894 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18816) );
  NOR2_X2 U21895 ( .A1(n18806), .A2(n18682), .ZN(n18677) );
  INV_X1 U21896 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18802) );
  NAND2_X1 U21897 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18661), .ZN(n18660) );
  NAND2_X1 U21898 ( .A1(n18660), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n18658) );
  NOR2_X2 U21899 ( .A1(n19515), .A2(n18784), .ZN(n18729) );
  NAND2_X1 U21900 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18729), .ZN(n18657) );
  OAI221_X1 U21901 ( .B1(n18660), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n18658), 
        .C2(n18777), .A(n18657), .ZN(P3_U2704) );
  NOR2_X2 U21902 ( .A1(n18659), .A2(n18784), .ZN(n18730) );
  AOI22_X1 U21903 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18729), .ZN(n18663) );
  OAI211_X1 U21904 ( .C1(n18661), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18784), .B(
        n18660), .ZN(n18662) );
  OAI211_X1 U21905 ( .C1(n18664), .C2(n18794), .A(n18663), .B(n18662), .ZN(
        P3_U2705) );
  AOI22_X1 U21906 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18729), .ZN(n18667) );
  OAI211_X1 U21907 ( .C1(n9789), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18784), .B(
        n18665), .ZN(n18666) );
  OAI211_X1 U21908 ( .C1(n18794), .C2(n18668), .A(n18667), .B(n18666), .ZN(
        P3_U2706) );
  AOI22_X1 U21909 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18729), .ZN(n18671) );
  AOI211_X1 U21910 ( .C1(n18802), .C2(n18673), .A(n9789), .B(n18777), .ZN(
        n18669) );
  INV_X1 U21911 ( .A(n18669), .ZN(n18670) );
  OAI211_X1 U21912 ( .C1(n18794), .C2(n18672), .A(n18671), .B(n18670), .ZN(
        P3_U2707) );
  AOI22_X1 U21913 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18729), .ZN(n18675) );
  OAI211_X1 U21914 ( .C1(n18677), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18784), .B(
        n18673), .ZN(n18674) );
  OAI211_X1 U21915 ( .C1(n18794), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        P3_U2708) );
  AOI22_X1 U21916 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18729), .ZN(n18680) );
  AOI211_X1 U21917 ( .C1(n18806), .C2(n18682), .A(n18677), .B(n18777), .ZN(
        n18678) );
  INV_X1 U21918 ( .A(n18678), .ZN(n18679) );
  OAI211_X1 U21919 ( .C1(n18794), .C2(n18681), .A(n18680), .B(n18679), .ZN(
        P3_U2709) );
  AOI22_X1 U21920 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18729), .ZN(n18685) );
  OAI211_X1 U21921 ( .C1(n18683), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18784), .B(
        n18682), .ZN(n18684) );
  OAI211_X1 U21922 ( .C1(n18794), .C2(n18686), .A(n18685), .B(n18684), .ZN(
        P3_U2710) );
  AOI22_X1 U21923 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18729), .ZN(n18690) );
  OAI211_X1 U21924 ( .C1(n18688), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18784), .B(
        n18687), .ZN(n18689) );
  OAI211_X1 U21925 ( .C1(n18794), .C2(n18691), .A(n18690), .B(n18689), .ZN(
        P3_U2711) );
  AOI22_X1 U21926 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18729), .ZN(n18695) );
  OAI211_X1 U21927 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n18693), .A(n18784), .B(
        n18692), .ZN(n18694) );
  OAI211_X1 U21928 ( .C1(n18794), .C2(n18696), .A(n18695), .B(n18694), .ZN(
        P3_U2712) );
  INV_X1 U21929 ( .A(n18730), .ZN(n18713) );
  INV_X1 U21930 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18864) );
  INV_X1 U21931 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18861) );
  NAND2_X1 U21932 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18723), .ZN(n18719) );
  NOR2_X2 U21933 ( .A1(n18864), .A2(n18719), .ZN(n18714) );
  NAND2_X1 U21934 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18714), .ZN(n18707) );
  NAND2_X1 U21935 ( .A1(n18784), .A2(n18707), .ZN(n18704) );
  OAI21_X1 U21936 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18739), .A(n18704), .ZN(
        n18701) );
  INV_X1 U21937 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18813) );
  AND4_X1 U21938 ( .A1(n18813), .A2(P3_EAX_REG_20__SCAN_IN), .A3(
        P3_EAX_REG_21__SCAN_IN), .A4(n18714), .ZN(n18700) );
  INV_X1 U21939 ( .A(n18729), .ZN(n18708) );
  OAI22_X1 U21940 ( .A1(n18698), .A2(n18794), .B1(n16822), .B2(n18708), .ZN(
        n18699) );
  AOI211_X1 U21941 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n18701), .A(n18700), .B(
        n18699), .ZN(n18702) );
  OAI21_X1 U21942 ( .B1(n19514), .B2(n18713), .A(n18702), .ZN(P3_U2713) );
  AOI22_X1 U21943 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18729), .B1(n18786), .B2(
        n18703), .ZN(n18706) );
  INV_X1 U21944 ( .A(n18704), .ZN(n18711) );
  AOI22_X1 U21945 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18730), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18711), .ZN(n18705) );
  OAI211_X1 U21946 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18707), .A(n18706), .B(
        n18705), .ZN(P3_U2714) );
  OAI22_X1 U21947 ( .A1(n18709), .A2(n18794), .B1(n21470), .B2(n18708), .ZN(
        n18710) );
  AOI221_X1 U21948 ( .B1(n18711), .B2(P3_EAX_REG_20__SCAN_IN), .C1(n18714), 
        .C2(n18816), .A(n18710), .ZN(n18712) );
  OAI21_X1 U21949 ( .B1(n19506), .B2(n18713), .A(n18712), .ZN(P3_U2715) );
  AOI22_X1 U21950 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18729), .ZN(n18717) );
  AOI211_X1 U21951 ( .C1(n18864), .C2(n18719), .A(n18714), .B(n18777), .ZN(
        n18715) );
  INV_X1 U21952 ( .A(n18715), .ZN(n18716) );
  OAI211_X1 U21953 ( .C1(n18718), .C2(n18794), .A(n18717), .B(n18716), .ZN(
        P3_U2716) );
  AOI22_X1 U21954 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18729), .ZN(n18721) );
  OAI211_X1 U21955 ( .C1(n18723), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18784), .B(
        n18719), .ZN(n18720) );
  OAI211_X1 U21956 ( .C1(n18722), .C2(n18794), .A(n18721), .B(n18720), .ZN(
        P3_U2717) );
  AOI22_X1 U21957 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18729), .ZN(n18727) );
  INV_X1 U21958 ( .A(n18731), .ZN(n18725) );
  INV_X1 U21959 ( .A(n18723), .ZN(n18724) );
  OAI211_X1 U21960 ( .C1(n18725), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18784), .B(
        n18724), .ZN(n18726) );
  OAI211_X1 U21961 ( .C1(n18728), .C2(n18794), .A(n18727), .B(n18726), .ZN(
        P3_U2718) );
  AOI22_X1 U21962 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18730), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18729), .ZN(n18733) );
  OAI211_X1 U21963 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18735), .A(n18784), .B(
        n18731), .ZN(n18732) );
  OAI211_X1 U21964 ( .C1(n18734), .C2(n18794), .A(n18733), .B(n18732), .ZN(
        P3_U2719) );
  AOI211_X1 U21965 ( .C1(n18908), .C2(n18741), .A(n18777), .B(n18735), .ZN(
        n18736) );
  AOI21_X1 U21966 ( .B1(n18787), .B2(BUF2_REG_15__SCAN_IN), .A(n18736), .ZN(
        n18737) );
  OAI21_X1 U21967 ( .B1(n18738), .B2(n18794), .A(n18737), .ZN(P3_U2720) );
  INV_X1 U21968 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18828) );
  INV_X1 U21969 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18832) );
  INV_X1 U21970 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18836) );
  NAND2_X1 U21971 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18771), .ZN(n18761) );
  NAND2_X1 U21972 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18764), .ZN(n18758) );
  NAND2_X1 U21973 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18755), .ZN(n18745) );
  NOR2_X1 U21974 ( .A1(n18828), .A2(n18745), .ZN(n18748) );
  INV_X1 U21975 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18903) );
  AOI22_X1 U21976 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18787), .B1(n18748), .B2(
        n18903), .ZN(n18743) );
  NAND3_X1 U21977 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18784), .A3(n18741), 
        .ZN(n18742) );
  OAI211_X1 U21978 ( .C1(n18744), .C2(n18794), .A(n18743), .B(n18742), .ZN(
        P3_U2721) );
  INV_X1 U21979 ( .A(n18745), .ZN(n18751) );
  AOI21_X1 U21980 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n18784), .A(n18751), .ZN(
        n18747) );
  OAI222_X1 U21981 ( .A1(n18795), .A2(n18901), .B1(n18748), .B2(n18747), .C1(
        n18794), .C2(n18746), .ZN(P3_U2722) );
  AOI21_X1 U21982 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18784), .A(n18755), .ZN(
        n18750) );
  OAI222_X1 U21983 ( .A1(n18795), .A2(n21555), .B1(n18751), .B2(n18750), .C1(
        n18794), .C2(n18749), .ZN(P3_U2723) );
  INV_X1 U21984 ( .A(n18758), .ZN(n18752) );
  AOI21_X1 U21985 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18784), .A(n18752), .ZN(
        n18754) );
  OAI222_X1 U21986 ( .A1(n18795), .A2(n18895), .B1(n18755), .B2(n18754), .C1(
        n18794), .C2(n18753), .ZN(P3_U2724) );
  INV_X1 U21987 ( .A(n18756), .ZN(n18757) );
  AOI22_X1 U21988 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18787), .B1(n18786), .B2(
        n18757), .ZN(n18760) );
  OAI211_X1 U21989 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n18764), .A(n18784), .B(
        n18758), .ZN(n18759) );
  NAND2_X1 U21990 ( .A1(n18760), .A2(n18759), .ZN(P3_U2725) );
  INV_X1 U21991 ( .A(n18761), .ZN(n18767) );
  AOI21_X1 U21992 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18784), .A(n18767), .ZN(
        n18763) );
  OAI222_X1 U21993 ( .A1(n18795), .A2(n18891), .B1(n18764), .B2(n18763), .C1(
        n18794), .C2(n18762), .ZN(P3_U2726) );
  AOI21_X1 U21994 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n18784), .A(n18771), .ZN(
        n18766) );
  OAI222_X1 U21995 ( .A1(n18795), .A2(n18889), .B1(n18767), .B2(n18766), .C1(
        n18794), .C2(n18765), .ZN(P3_U2727) );
  NAND3_X1 U21996 ( .A1(n19521), .A2(P3_EAX_REG_2__SCAN_IN), .A3(n18790), .ZN(
        n18789) );
  NOR2_X1 U21997 ( .A1(n21565), .A2(n18789), .ZN(n18780) );
  NAND2_X1 U21998 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18780), .ZN(n18779) );
  NOR2_X1 U21999 ( .A1(n18768), .A2(n18779), .ZN(n18774) );
  AOI21_X1 U22000 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18784), .A(n18774), .ZN(
        n18770) );
  OAI222_X1 U22001 ( .A1(n19518), .A2(n18795), .B1(n18771), .B2(n18770), .C1(
        n18794), .C2(n18769), .ZN(P3_U2728) );
  INV_X1 U22002 ( .A(n18779), .ZN(n18783) );
  AOI22_X1 U22003 ( .A1(n18783), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18784), .ZN(n18773) );
  OAI222_X1 U22004 ( .A1(n19514), .A2(n18795), .B1(n18774), .B2(n18773), .C1(
        n18794), .C2(n18772), .ZN(P3_U2729) );
  NAND2_X1 U22005 ( .A1(n18779), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n18778) );
  AOI22_X1 U22006 ( .A1(n18787), .A2(BUF2_REG_5__SCAN_IN), .B1(n18786), .B2(
        n18775), .ZN(n18776) );
  OAI221_X1 U22007 ( .B1(n18779), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n18778), 
        .C2(n18777), .A(n18776), .ZN(P3_U2730) );
  AOI21_X1 U22008 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18784), .A(n18780), .ZN(
        n18782) );
  OAI222_X1 U22009 ( .A1(n19506), .A2(n18795), .B1(n18783), .B2(n18782), .C1(
        n18794), .C2(n18781), .ZN(P3_U2731) );
  NAND2_X1 U22010 ( .A1(n18784), .A2(n18789), .ZN(n18792) );
  AOI22_X1 U22011 ( .A1(n18787), .A2(BUF2_REG_3__SCAN_IN), .B1(n18786), .B2(
        n18785), .ZN(n18788) );
  OAI221_X1 U22012 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18789), .C1(n21565), 
        .C2(n18792), .A(n18788), .ZN(P3_U2732) );
  NOR2_X1 U22013 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18790), .ZN(n18791) );
  OAI222_X1 U22014 ( .A1(n18795), .A2(n19499), .B1(n18794), .B2(n18793), .C1(
        n18792), .C2(n18791), .ZN(P3_U2733) );
  INV_X2 U22015 ( .A(n18843), .ZN(n20084) );
  NOR2_X1 U22016 ( .A1(n18821), .A2(n18797), .ZN(P3_U2736) );
  INV_X1 U22017 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18876) );
  INV_X2 U22018 ( .A(n18821), .ZN(n18850) );
  AOI22_X1 U22019 ( .A1(n20084), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18799) );
  OAI21_X1 U22020 ( .B1(n18876), .B2(n18823), .A(n18799), .ZN(P3_U2737) );
  AOI22_X1 U22021 ( .A1(n20084), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18800) );
  OAI21_X1 U22022 ( .B1(n10088), .B2(n18823), .A(n18800), .ZN(P3_U2738) );
  AOI22_X1 U22023 ( .A1(n20084), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18801) );
  OAI21_X1 U22024 ( .B1(n18802), .B2(n18823), .A(n18801), .ZN(P3_U2739) );
  INV_X1 U22025 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18804) );
  AOI22_X1 U22026 ( .A1(n20084), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18803) );
  OAI21_X1 U22027 ( .B1(n18804), .B2(n18823), .A(n18803), .ZN(P3_U2740) );
  AOI22_X1 U22028 ( .A1(n20084), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18805) );
  OAI21_X1 U22029 ( .B1(n18806), .B2(n18823), .A(n18805), .ZN(P3_U2741) );
  INV_X1 U22030 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18808) );
  AOI22_X1 U22031 ( .A1(n20084), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18807) );
  OAI21_X1 U22032 ( .B1(n18808), .B2(n18823), .A(n18807), .ZN(P3_U2742) );
  INV_X1 U22033 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n21506) );
  INV_X1 U22034 ( .A(n18823), .ZN(n18810) );
  AOI22_X1 U22035 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18810), .B1(n20084), 
        .B2(P3_UWORD_REG_8__SCAN_IN), .ZN(n18809) );
  OAI21_X1 U22036 ( .B1(n21506), .B2(n18821), .A(n18809), .ZN(P3_U2743) );
  INV_X1 U22037 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n21528) );
  AOI22_X1 U22038 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18810), .B1(n20084), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n18811) );
  OAI21_X1 U22039 ( .B1(n21528), .B2(n18821), .A(n18811), .ZN(P3_U2744) );
  AOI22_X1 U22040 ( .A1(n20084), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18812) );
  OAI21_X1 U22041 ( .B1(n18813), .B2(n18823), .A(n18812), .ZN(P3_U2745) );
  AOI22_X1 U22042 ( .A1(n20084), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18814) );
  OAI21_X1 U22043 ( .B1(n21622), .B2(n18823), .A(n18814), .ZN(P3_U2746) );
  AOI22_X1 U22044 ( .A1(n20084), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18815) );
  OAI21_X1 U22045 ( .B1(n18816), .B2(n18823), .A(n18815), .ZN(P3_U2747) );
  AOI22_X1 U22046 ( .A1(n20084), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18817) );
  OAI21_X1 U22047 ( .B1(n18864), .B2(n18823), .A(n18817), .ZN(P3_U2748) );
  INV_X1 U22048 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18819) );
  AOI22_X1 U22049 ( .A1(n20084), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18818) );
  OAI21_X1 U22050 ( .B1(n18819), .B2(n18823), .A(n18818), .ZN(P3_U2749) );
  AOI22_X1 U22051 ( .A1(n20084), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18820) );
  OAI21_X1 U22052 ( .B1(n18861), .B2(n18823), .A(n18820), .ZN(P3_U2750) );
  INV_X1 U22053 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18824) );
  AOI22_X1 U22054 ( .A1(n20084), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18822) );
  OAI21_X1 U22055 ( .B1(n18824), .B2(n18823), .A(n18822), .ZN(P3_U2751) );
  AOI22_X1 U22056 ( .A1(n20084), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18825) );
  OAI21_X1 U22057 ( .B1(n18908), .B2(n18853), .A(n18825), .ZN(P3_U2752) );
  AOI22_X1 U22058 ( .A1(n20084), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18826) );
  OAI21_X1 U22059 ( .B1(n18903), .B2(n18853), .A(n18826), .ZN(P3_U2753) );
  AOI22_X1 U22060 ( .A1(n20084), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18827) );
  OAI21_X1 U22061 ( .B1(n18828), .B2(n18853), .A(n18827), .ZN(P3_U2754) );
  INV_X1 U22062 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18830) );
  AOI22_X1 U22063 ( .A1(n20084), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18829) );
  OAI21_X1 U22064 ( .B1(n18830), .B2(n18853), .A(n18829), .ZN(P3_U2755) );
  AOI22_X1 U22065 ( .A1(n20084), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18831) );
  OAI21_X1 U22066 ( .B1(n18832), .B2(n18853), .A(n18831), .ZN(P3_U2756) );
  INV_X1 U22067 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18834) );
  AOI22_X1 U22068 ( .A1(n20084), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18833) );
  OAI21_X1 U22069 ( .B1(n18834), .B2(n18853), .A(n18833), .ZN(P3_U2757) );
  AOI22_X1 U22070 ( .A1(n20084), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18835) );
  OAI21_X1 U22071 ( .B1(n18836), .B2(n18853), .A(n18835), .ZN(P3_U2758) );
  INV_X1 U22072 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18838) );
  AOI22_X1 U22073 ( .A1(n20084), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18837) );
  OAI21_X1 U22074 ( .B1(n18838), .B2(n18853), .A(n18837), .ZN(P3_U2759) );
  AOI22_X1 U22075 ( .A1(n20084), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18839) );
  OAI21_X1 U22076 ( .B1(n18840), .B2(n18853), .A(n18839), .ZN(P3_U2760) );
  INV_X1 U22077 ( .A(P3_LWORD_REG_6__SCAN_IN), .ZN(n21532) );
  AOI22_X1 U22078 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18841), .B1(n18850), .B2(
        P3_DATAO_REG_6__SCAN_IN), .ZN(n18842) );
  OAI21_X1 U22079 ( .B1(n21532), .B2(n18843), .A(n18842), .ZN(P3_U2761) );
  INV_X1 U22080 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18885) );
  AOI22_X1 U22081 ( .A1(n20084), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18844) );
  OAI21_X1 U22082 ( .B1(n18885), .B2(n18853), .A(n18844), .ZN(P3_U2762) );
  INV_X1 U22083 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18846) );
  AOI22_X1 U22084 ( .A1(n20084), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18845) );
  OAI21_X1 U22085 ( .B1(n18846), .B2(n18853), .A(n18845), .ZN(P3_U2763) );
  AOI22_X1 U22086 ( .A1(n20084), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18847) );
  OAI21_X1 U22087 ( .B1(n21565), .B2(n18853), .A(n18847), .ZN(P3_U2764) );
  INV_X1 U22088 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18849) );
  AOI22_X1 U22089 ( .A1(n20084), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18848) );
  OAI21_X1 U22090 ( .B1(n18849), .B2(n18853), .A(n18848), .ZN(P3_U2765) );
  INV_X1 U22091 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18879) );
  AOI22_X1 U22092 ( .A1(n20084), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18851) );
  OAI21_X1 U22093 ( .B1(n18879), .B2(n18853), .A(n18851), .ZN(P3_U2766) );
  AOI22_X1 U22094 ( .A1(n20084), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18850), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18852) );
  OAI21_X1 U22095 ( .B1(n18854), .B2(n18853), .A(n18852), .ZN(P3_U2767) );
  INV_X1 U22096 ( .A(n18857), .ZN(n18855) );
  AOI22_X1 U22097 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18904), .ZN(n18859) );
  OAI21_X1 U22098 ( .B1(n19489), .B2(n18900), .A(n18859), .ZN(P3_U2768) );
  INV_X1 U22099 ( .A(n18898), .ZN(n18907) );
  AOI22_X1 U22100 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18905), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18882), .ZN(n18860) );
  OAI21_X1 U22101 ( .B1(n18861), .B2(n18907), .A(n18860), .ZN(P3_U2769) );
  AOI22_X1 U22102 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18904), .ZN(n18862) );
  OAI21_X1 U22103 ( .B1(n19499), .B2(n18900), .A(n18862), .ZN(P3_U2770) );
  AOI22_X1 U22104 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18905), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18882), .ZN(n18863) );
  OAI21_X1 U22105 ( .B1(n18864), .B2(n18907), .A(n18863), .ZN(P3_U2771) );
  AOI22_X1 U22106 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18904), .ZN(n18865) );
  OAI21_X1 U22107 ( .B1(n19506), .B2(n18900), .A(n18865), .ZN(P3_U2772) );
  AOI22_X1 U22108 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18905), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18882), .ZN(n18866) );
  OAI21_X1 U22109 ( .B1(n21622), .B2(n18907), .A(n18866), .ZN(P3_U2773) );
  AOI22_X1 U22110 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18898), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18904), .ZN(n18867) );
  OAI21_X1 U22111 ( .B1(n19514), .B2(n18900), .A(n18867), .ZN(P3_U2774) );
  AOI22_X1 U22112 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18882), .ZN(n18868) );
  OAI21_X1 U22113 ( .B1(n19518), .B2(n18900), .A(n18868), .ZN(P3_U2775) );
  AOI22_X1 U22114 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18904), .ZN(n18869) );
  OAI21_X1 U22115 ( .B1(n18889), .B2(n18900), .A(n18869), .ZN(P3_U2776) );
  AOI22_X1 U22116 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18882), .ZN(n18870) );
  OAI21_X1 U22117 ( .B1(n18891), .B2(n18900), .A(n18870), .ZN(P3_U2777) );
  AOI22_X1 U22118 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18898), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18882), .ZN(n18871) );
  OAI21_X1 U22119 ( .B1(n18893), .B2(n18900), .A(n18871), .ZN(P3_U2778) );
  AOI22_X1 U22120 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18904), .ZN(n18872) );
  OAI21_X1 U22121 ( .B1(n18895), .B2(n18900), .A(n18872), .ZN(P3_U2779) );
  AOI22_X1 U22122 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18882), .ZN(n18873) );
  OAI21_X1 U22123 ( .B1(n21555), .B2(n18900), .A(n18873), .ZN(P3_U2780) );
  AOI22_X1 U22124 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18896), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18882), .ZN(n18874) );
  OAI21_X1 U22125 ( .B1(n18901), .B2(n18900), .A(n18874), .ZN(P3_U2781) );
  AOI22_X1 U22126 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18905), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18904), .ZN(n18875) );
  OAI21_X1 U22127 ( .B1(n18876), .B2(n18907), .A(n18875), .ZN(P3_U2782) );
  AOI22_X1 U22128 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18898), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18904), .ZN(n18877) );
  OAI21_X1 U22129 ( .B1(n19489), .B2(n18900), .A(n18877), .ZN(P3_U2783) );
  AOI22_X1 U22130 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18905), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18904), .ZN(n18878) );
  OAI21_X1 U22131 ( .B1(n18879), .B2(n18907), .A(n18878), .ZN(P3_U2784) );
  AOI22_X1 U22132 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18904), .ZN(n18880) );
  OAI21_X1 U22133 ( .B1(n19499), .B2(n18900), .A(n18880), .ZN(P3_U2785) );
  AOI22_X1 U22134 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18905), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18904), .ZN(n18881) );
  OAI21_X1 U22135 ( .B1(n21565), .B2(n18907), .A(n18881), .ZN(P3_U2786) );
  AOI22_X1 U22136 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18882), .ZN(n18883) );
  OAI21_X1 U22137 ( .B1(n19506), .B2(n18900), .A(n18883), .ZN(P3_U2787) );
  AOI22_X1 U22138 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18905), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18904), .ZN(n18884) );
  OAI21_X1 U22139 ( .B1(n18885), .B2(n18907), .A(n18884), .ZN(P3_U2788) );
  AOI22_X1 U22140 ( .A1(P3_LWORD_REG_6__SCAN_IN), .A2(n18904), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18896), .ZN(n18886) );
  OAI21_X1 U22141 ( .B1(n19514), .B2(n18900), .A(n18886), .ZN(P3_U2789) );
  AOI22_X1 U22142 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18904), .ZN(n18887) );
  OAI21_X1 U22143 ( .B1(n19518), .B2(n18900), .A(n18887), .ZN(P3_U2790) );
  AOI22_X1 U22144 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18904), .ZN(n18888) );
  OAI21_X1 U22145 ( .B1(n18889), .B2(n18900), .A(n18888), .ZN(P3_U2791) );
  AOI22_X1 U22146 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18898), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18904), .ZN(n18890) );
  OAI21_X1 U22147 ( .B1(n18891), .B2(n18900), .A(n18890), .ZN(P3_U2792) );
  AOI22_X1 U22148 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18904), .ZN(n18892) );
  OAI21_X1 U22149 ( .B1(n18893), .B2(n18900), .A(n18892), .ZN(P3_U2793) );
  AOI22_X1 U22150 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18904), .ZN(n18894) );
  OAI21_X1 U22151 ( .B1(n18895), .B2(n18900), .A(n18894), .ZN(P3_U2794) );
  AOI22_X1 U22152 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18896), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18904), .ZN(n18897) );
  OAI21_X1 U22153 ( .B1(n21555), .B2(n18900), .A(n18897), .ZN(P3_U2795) );
  AOI22_X1 U22154 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18898), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18904), .ZN(n18899) );
  OAI21_X1 U22155 ( .B1(n18901), .B2(n18900), .A(n18899), .ZN(P3_U2796) );
  AOI22_X1 U22156 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18905), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18904), .ZN(n18902) );
  OAI21_X1 U22157 ( .B1(n18903), .B2(n18907), .A(n18902), .ZN(P3_U2797) );
  AOI22_X1 U22158 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18905), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18904), .ZN(n18906) );
  OAI21_X1 U22159 ( .B1(n18908), .B2(n18907), .A(n18906), .ZN(P3_U2798) );
  NAND2_X1 U22160 ( .A1(n10340), .A2(n18910), .ZN(n18911) );
  MUX2_X1 U22161 ( .A(n18911), .B(n10340), .S(n19113), .Z(n18912) );
  NAND2_X1 U22162 ( .A1(n18912), .A2(n13212), .ZN(n19231) );
  AOI22_X1 U22163 ( .A1(n19477), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n19124), 
        .B2(n18913), .ZN(n18914) );
  OAI221_X1 U22164 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18917), .C1(
        n18916), .C2(n18915), .A(n18914), .ZN(n18918) );
  AOI221_X1 U22165 ( .B1(n18919), .B2(n19225), .C1(n18925), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n18918), .ZN(n18920) );
  OAI21_X1 U22166 ( .B1(n19231), .B2(n19178), .A(n18920), .ZN(P3_U2803) );
  NAND2_X1 U22167 ( .A1(n18921), .A2(n17516), .ZN(n18922) );
  OAI22_X1 U22168 ( .A1(n18923), .A2(n19178), .B1(n18922), .B2(n18976), .ZN(
        n18924) );
  AOI21_X1 U22169 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18925), .A(
        n18924), .ZN(n18933) );
  AND3_X1 U22170 ( .A1(n19871), .A2(n13505), .A3(n18936), .ZN(n18927) );
  OAI21_X1 U22171 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18927), .A(
        n18926), .ZN(n18931) );
  OAI21_X1 U22172 ( .B1(n19124), .B2(n18929), .A(n18928), .ZN(n18930) );
  NAND4_X1 U22173 ( .A1(n18933), .A2(n18932), .A3(n18931), .A4(n18930), .ZN(
        P3_U2804) );
  NAND2_X1 U22174 ( .A1(n18934), .A2(n19080), .ZN(n18935) );
  XNOR2_X1 U22175 ( .A(n18935), .B(n19235), .ZN(n19244) );
  NAND2_X1 U22176 ( .A1(n13505), .A2(n19062), .ZN(n18952) );
  AOI211_X1 U22177 ( .C1(n21563), .C2(n18951), .A(n18936), .B(n18952), .ZN(
        n18939) );
  OR2_X1 U22178 ( .A1(n19507), .A2(n13505), .ZN(n18972) );
  OAI211_X1 U22179 ( .C1(n18937), .C2(n19103), .A(n19202), .B(n18972), .ZN(
        n18969) );
  AOI21_X1 U22180 ( .B1(n19004), .B2(n18967), .A(n18969), .ZN(n18950) );
  OAI22_X1 U22181 ( .A1(n18950), .A2(n21563), .B1(n19428), .B2(n20048), .ZN(
        n18938) );
  AOI211_X1 U22182 ( .C1(n18940), .C2(n19124), .A(n18939), .B(n18938), .ZN(
        n18948) );
  AOI221_X1 U22183 ( .B1(n19339), .B2(n19235), .C1(n18942), .C2(n19235), .A(
        n18941), .ZN(n19241) );
  INV_X1 U22184 ( .A(n18943), .ZN(n18944) );
  NAND2_X1 U22185 ( .A1(n18945), .A2(n18944), .ZN(n18946) );
  XNOR2_X1 U22186 ( .A(n18946), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n19240) );
  AOI22_X1 U22187 ( .A1(n19220), .A2(n19241), .B1(n19128), .B2(n19240), .ZN(
        n18947) );
  OAI211_X1 U22188 ( .C1(n19177), .C2(n19244), .A(n18948), .B(n18947), .ZN(
        P3_U2805) );
  OAI221_X1 U22189 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18952), .C1(
        n18951), .C2(n18950), .A(n18949), .ZN(n18959) );
  AOI22_X1 U22190 ( .A1(n18954), .A2(n19220), .B1(n18981), .B2(n18953), .ZN(
        n18975) );
  INV_X1 U22191 ( .A(n18955), .ZN(n18956) );
  OAI22_X1 U22192 ( .A1(n18975), .A2(n18957), .B1(n18956), .B2(n19178), .ZN(
        n18958) );
  AOI211_X1 U22193 ( .C1(n19124), .C2(n18960), .A(n18959), .B(n18958), .ZN(
        n18961) );
  OAI21_X1 U22194 ( .B1(n19067), .B2(n18962), .A(n18961), .ZN(P3_U2806) );
  NAND2_X1 U22195 ( .A1(n19174), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18964) );
  OAI211_X1 U22196 ( .C1(n18965), .C2(n18977), .A(n18964), .B(n18963), .ZN(
        n18966) );
  XNOR2_X1 U22197 ( .A(n18966), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19247) );
  NOR2_X1 U22198 ( .A1(n19428), .A2(n20044), .ZN(n19246) );
  NAND3_X1 U22199 ( .A1(n19004), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        n18967), .ZN(n18971) );
  AOI22_X1 U22200 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18969), .B1(
        n19124), .B2(n18968), .ZN(n18970) );
  OAI221_X1 U22201 ( .B1(n9853), .B2(n18972), .C1(n9853), .C2(n18971), .A(
        n18970), .ZN(n18973) );
  AOI211_X1 U22202 ( .C1(n19247), .C2(n19128), .A(n19246), .B(n18973), .ZN(
        n18974) );
  OAI221_X1 U22203 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18976), 
        .C1(n19250), .C2(n18975), .A(n18974), .ZN(P3_U2807) );
  INV_X1 U22204 ( .A(n18963), .ZN(n18979) );
  AOI21_X1 U22205 ( .B1(n19056), .B2(n19252), .A(n18977), .ZN(n18978) );
  NOR2_X1 U22206 ( .A1(n18979), .A2(n18978), .ZN(n18980) );
  XNOR2_X1 U22207 ( .A(n18980), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n19265) );
  INV_X1 U22208 ( .A(n19080), .ZN(n19331) );
  AOI22_X1 U22209 ( .A1(n19220), .A2(n19339), .B1(n18981), .B2(n19331), .ZN(
        n19066) );
  OAI21_X1 U22210 ( .B1(n19252), .B2(n19010), .A(n19066), .ZN(n18999) );
  NAND2_X1 U22211 ( .A1(n18982), .A2(n19062), .ZN(n18994) );
  AOI221_X1 U22212 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n18993), .C2(n18987), .A(
        n18994), .ZN(n18989) );
  NAND2_X1 U22213 ( .A1(n19059), .A2(n18983), .ZN(n18984) );
  OAI211_X1 U22214 ( .C1(n18982), .C2(n19105), .A(n19202), .B(n18984), .ZN(
        n19009) );
  AOI21_X1 U22215 ( .B1(n19004), .B2(n19002), .A(n19009), .ZN(n18992) );
  AOI22_X1 U22216 ( .A1(n19477), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n19124), 
        .B2(n18985), .ZN(n18986) );
  OAI21_X1 U22217 ( .B1(n18992), .B2(n18987), .A(n18986), .ZN(n18988) );
  AOI211_X1 U22218 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18999), .A(
        n18989), .B(n18988), .ZN(n18991) );
  NAND3_X1 U22219 ( .A1(n19252), .A2(n19048), .A3(n19261), .ZN(n18990) );
  OAI211_X1 U22220 ( .C1(n19178), .C2(n19265), .A(n18991), .B(n18990), .ZN(
        P3_U2808) );
  NAND2_X1 U22221 ( .A1(n19273), .A2(n19268), .ZN(n19279) );
  NOR2_X1 U22222 ( .A1(n19302), .A2(n19303), .ZN(n19266) );
  NAND2_X1 U22223 ( .A1(n19048), .A2(n19266), .ZN(n19032) );
  NAND2_X1 U22224 ( .A1(n19477), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19277) );
  OAI221_X1 U22225 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18994), .C1(
        n18993), .C2(n18992), .A(n19277), .ZN(n18995) );
  AOI21_X1 U22226 ( .B1(n19124), .B2(n18996), .A(n18995), .ZN(n19001) );
  INV_X1 U22227 ( .A(n19039), .ZN(n19026) );
  NAND4_X1 U22228 ( .A1(n19056), .A2(n19113), .A3(n19037), .A4(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19027) );
  INV_X1 U22229 ( .A(n19027), .ZN(n19013) );
  AOI22_X1 U22230 ( .A1(n19026), .A2(n18997), .B1(n19273), .B2(n19013), .ZN(
        n18998) );
  XNOR2_X1 U22231 ( .A(n18998), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n19276) );
  AOI22_X1 U22232 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18999), .B1(
        n19128), .B2(n19276), .ZN(n19000) );
  OAI211_X1 U22233 ( .C1(n19279), .C2(n19032), .A(n19001), .B(n19000), .ZN(
        P3_U2809) );
  NAND2_X1 U22234 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19257), .ZN(
        n19288) );
  NAND3_X1 U22235 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19003) );
  NAND2_X1 U22236 ( .A1(n19871), .A2(n19017), .ZN(n19049) );
  OAI21_X1 U22237 ( .B1(n19003), .B2(n19049), .A(n19002), .ZN(n19008) );
  INV_X1 U22238 ( .A(n19124), .ZN(n19109) );
  INV_X1 U22239 ( .A(n19005), .ZN(n19006) );
  AOI21_X1 U22240 ( .B1(n19109), .B2(n17452), .A(n19006), .ZN(n19007) );
  INV_X1 U22241 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20038) );
  NOR2_X1 U22242 ( .A1(n19428), .A2(n20038), .ZN(n19280) );
  AOI211_X1 U22243 ( .C1(n19009), .C2(n19008), .A(n19007), .B(n19280), .ZN(
        n19016) );
  INV_X1 U22244 ( .A(n19266), .ZN(n19269) );
  NOR2_X1 U22245 ( .A1(n19012), .A2(n19269), .ZN(n19284) );
  OAI21_X1 U22246 ( .B1(n19010), .B2(n19284), .A(n19066), .ZN(n19029) );
  INV_X1 U22247 ( .A(n19025), .ZN(n19038) );
  NAND2_X1 U22248 ( .A1(n19038), .A2(n19012), .ZN(n19011) );
  OAI211_X1 U22249 ( .C1(n19013), .C2(n19012), .A(n18963), .B(n19011), .ZN(
        n19014) );
  XNOR2_X1 U22250 ( .A(n19014), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n19281) );
  AOI22_X1 U22251 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19029), .B1(
        n19128), .B2(n19281), .ZN(n19015) );
  OAI211_X1 U22252 ( .C1(n19032), .C2(n19288), .A(n19016), .B(n19015), .ZN(
        P3_U2810) );
  NAND3_X1 U22253 ( .A1(n19017), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        n19062), .ZN(n19034) );
  AOI221_X1 U22254 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n21731), .C2(n19021), .A(
        n19034), .ZN(n19023) );
  NOR2_X1 U22255 ( .A1(n10482), .A2(n19018), .ZN(n19019) );
  OAI21_X1 U22256 ( .B1(n19019), .B2(n19105), .A(n19202), .ZN(n19050) );
  AOI21_X1 U22257 ( .B1(n19059), .B2(n19020), .A(n19050), .ZN(n19033) );
  OAI22_X1 U22258 ( .A1(n19033), .A2(n19021), .B1(n19428), .B2(n20036), .ZN(
        n19022) );
  AOI211_X1 U22259 ( .C1(n19024), .C2(n19124), .A(n19023), .B(n19022), .ZN(
        n19031) );
  NAND2_X1 U22260 ( .A1(n19026), .A2(n19025), .ZN(n19042) );
  NAND2_X1 U22261 ( .A1(n19042), .A2(n19027), .ZN(n19028) );
  XOR2_X1 U22262 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n19028), .Z(
        n19289) );
  AOI22_X1 U22263 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19029), .B1(
        n19128), .B2(n19289), .ZN(n19030) );
  OAI211_X1 U22264 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19032), .A(
        n19031), .B(n19030), .ZN(P3_U2811) );
  NAND2_X1 U22265 ( .A1(n19037), .A2(n19303), .ZN(n19309) );
  NAND2_X1 U22266 ( .A1(n19477), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n19307) );
  OAI221_X1 U22267 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19034), .C1(
        n21731), .C2(n19033), .A(n19307), .ZN(n19035) );
  AOI21_X1 U22268 ( .B1(n19124), .B2(n19036), .A(n19035), .ZN(n19045) );
  OAI21_X1 U22269 ( .B1(n19067), .B2(n19037), .A(n19066), .ZN(n19047) );
  NAND2_X1 U22270 ( .A1(n19113), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19041) );
  NAND2_X1 U22271 ( .A1(n19038), .A2(n19041), .ZN(n19040) );
  MUX2_X1 U22272 ( .A(n19041), .B(n19040), .S(n19039), .Z(n19043) );
  NAND2_X1 U22273 ( .A1(n19043), .A2(n19042), .ZN(n19304) );
  AOI22_X1 U22274 ( .A1(n19047), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19128), .B2(n19304), .ZN(n19044) );
  OAI211_X1 U22275 ( .C1(n19067), .C2(n19309), .A(n19045), .B(n19044), .ZN(
        P3_U2812) );
  XNOR2_X1 U22276 ( .A(n9834), .B(n19310), .ZN(n19312) );
  AOI22_X1 U22277 ( .A1(n19190), .A2(n19046), .B1(n19128), .B2(n19312), .ZN(
        n19054) );
  OAI221_X1 U22278 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n19048), .A(n19047), .ZN(
        n19053) );
  NAND2_X1 U22279 ( .A1(n19477), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n19314) );
  INV_X1 U22280 ( .A(n19049), .ZN(n19051) );
  OAI21_X1 U22281 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19051), .A(
        n19050), .ZN(n19052) );
  NAND4_X1 U22282 ( .A1(n19054), .A2(n19053), .A3(n19314), .A4(n19052), .ZN(
        P3_U2813) );
  NAND2_X1 U22283 ( .A1(n19382), .A2(n19113), .ZN(n19155) );
  OAI22_X1 U22284 ( .A1(n19056), .A2(n19113), .B1(n19155), .B2(n19055), .ZN(
        n19057) );
  XNOR2_X1 U22285 ( .A(n10181), .B(n19057), .ZN(n19325) );
  OAI21_X1 U22286 ( .B1(n10487), .B2(n19105), .A(n19202), .ZN(n19091) );
  AOI21_X1 U22287 ( .B1(n19059), .B2(n19058), .A(n19091), .ZN(n19076) );
  AOI22_X1 U22288 ( .A1(n19477), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19124), 
        .B2(n19060), .ZN(n19064) );
  NOR2_X1 U22289 ( .A1(n19063), .A2(n19121), .ZN(n19079) );
  NOR2_X1 U22290 ( .A1(n19093), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n19073) );
  INV_X1 U22291 ( .A(n19115), .ZN(n19071) );
  INV_X1 U22292 ( .A(n19068), .ZN(n19070) );
  AOI21_X1 U22293 ( .B1(n19071), .B2(n19070), .A(n19069), .ZN(n19072) );
  AOI211_X1 U22294 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19174), .A(
        n19073), .B(n19072), .ZN(n19074) );
  XNOR2_X1 U22295 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19074), .ZN(
        n19342) );
  NOR2_X1 U22296 ( .A1(n19428), .A2(n20028), .ZN(n19337) );
  OAI22_X1 U22297 ( .A1(n19076), .A2(n19078), .B1(n19109), .B2(n19075), .ZN(
        n19077) );
  AOI211_X1 U22298 ( .C1(n19079), .C2(n19078), .A(n19337), .B(n19077), .ZN(
        n19086) );
  NOR2_X1 U22299 ( .A1(n19080), .A2(n19177), .ZN(n19084) );
  INV_X1 U22300 ( .A(n19358), .ZN(n19372) );
  NOR2_X1 U22301 ( .A1(n19380), .A2(n19372), .ZN(n19343) );
  INV_X1 U22302 ( .A(n19343), .ZN(n19368) );
  NOR2_X1 U22303 ( .A1(n19081), .A2(n19368), .ZN(n19359) );
  NAND3_X1 U22304 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n19359), .ZN(n19097) );
  NAND2_X1 U22305 ( .A1(n11880), .A2(n19097), .ZN(n19330) );
  NOR2_X1 U22306 ( .A1(n19082), .A2(n19210), .ZN(n19083) );
  INV_X1 U22307 ( .A(n19095), .ZN(n19383) );
  NAND2_X1 U22308 ( .A1(n19329), .A2(n19383), .ZN(n19096) );
  NAND2_X1 U22309 ( .A1(n11880), .A2(n19096), .ZN(n19338) );
  AOI22_X1 U22310 ( .A1(n19084), .A2(n19330), .B1(n19083), .B2(n19338), .ZN(
        n19085) );
  OAI211_X1 U22311 ( .C1(n19178), .C2(n19342), .A(n19086), .B(n19085), .ZN(
        P3_U2815) );
  INV_X1 U22312 ( .A(n19102), .ZN(n19088) );
  NAND2_X1 U22313 ( .A1(n19871), .A2(n19061), .ZN(n19137) );
  OAI21_X1 U22314 ( .B1(n19088), .B2(n19137), .A(n19087), .ZN(n19090) );
  AOI22_X1 U22315 ( .A1(n19091), .A2(n19090), .B1(n19089), .B2(n19190), .ZN(
        n19100) );
  NAND2_X1 U22316 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19343), .ZN(
        n19347) );
  OAI21_X1 U22317 ( .B1(n19347), .B2(n19155), .A(n19092), .ZN(n19094) );
  XNOR2_X1 U22318 ( .A(n19094), .B(n19093), .ZN(n19353) );
  NOR2_X1 U22319 ( .A1(n19095), .A2(n19368), .ZN(n19360) );
  OAI221_X1 U22320 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n19360), .A(n19096), .ZN(
        n19357) );
  OAI221_X1 U22321 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n19359), .A(n19097), .ZN(
        n19352) );
  OAI22_X1 U22322 ( .A1(n19210), .A2(n19357), .B1(n19177), .B2(n19352), .ZN(
        n19098) );
  AOI21_X1 U22323 ( .B1(n19128), .B2(n19353), .A(n19098), .ZN(n19099) );
  OAI211_X1 U22324 ( .C1(n19216), .C2(n20027), .A(n19100), .B(n19099), .ZN(
        P3_U2816) );
  OAI22_X1 U22325 ( .A1(n19210), .A2(n19360), .B1(n19177), .B2(n19359), .ZN(
        n19101) );
  INV_X1 U22326 ( .A(n19101), .ZN(n19131) );
  AOI211_X1 U22327 ( .C1(n19120), .C2(n19110), .A(n19102), .B(n19121), .ZN(
        n19112) );
  OAI21_X1 U22328 ( .B1(n18058), .B2(n19105), .A(n19202), .ZN(n19183) );
  OAI22_X1 U22329 ( .A1(n19106), .A2(n19105), .B1(n19104), .B2(n19103), .ZN(
        n19107) );
  NOR2_X1 U22330 ( .A1(n19183), .A2(n19107), .ZN(n19119) );
  OAI22_X1 U22331 ( .A1(n19119), .A2(n19110), .B1(n19109), .B2(n19108), .ZN(
        n19111) );
  AOI211_X1 U22332 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n19477), .A(n19112), 
        .B(n19111), .ZN(n19118) );
  NAND2_X1 U22333 ( .A1(n19113), .A2(n19343), .ZN(n19114) );
  OAI22_X1 U22334 ( .A1(n19115), .A2(n19114), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n19125), .ZN(n19116) );
  XOR2_X1 U22335 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19116), .Z(
        n19365) );
  NOR2_X1 U22336 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n19368), .ZN(
        n19364) );
  AOI22_X1 U22337 ( .A1(n19128), .A2(n19365), .B1(n19364), .B2(n19164), .ZN(
        n19117) );
  OAI211_X1 U22338 ( .C1(n19131), .C2(n10343), .A(n19118), .B(n19117), .ZN(
        P3_U2817) );
  NAND2_X1 U22339 ( .A1(n19477), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19378) );
  OAI221_X1 U22340 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19121), .C1(
        n19120), .C2(n19119), .A(n19378), .ZN(n19122) );
  AOI21_X1 U22341 ( .B1(n19124), .B2(n19123), .A(n19122), .ZN(n19130) );
  OAI21_X1 U22342 ( .B1(n19155), .B2(n19372), .A(n19125), .ZN(n19126) );
  XNOR2_X1 U22343 ( .A(n19126), .B(n19380), .ZN(n19376) );
  NOR2_X1 U22344 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n19372), .ZN(
        n19127) );
  AOI22_X1 U22345 ( .A1(n19128), .A2(n19376), .B1(n19127), .B2(n19164), .ZN(
        n19129) );
  OAI211_X1 U22346 ( .C1(n19131), .C2(n19380), .A(n19130), .B(n19129), .ZN(
        P3_U2818) );
  OAI22_X1 U22347 ( .A1(n19177), .A2(n19382), .B1(n19383), .B2(n19210), .ZN(
        n19165) );
  AOI21_X1 U22348 ( .B1(n19386), .B2(n19164), .A(n19165), .ZN(n19145) );
  NOR2_X1 U22349 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19386), .ZN(
        n19392) );
  OAI22_X1 U22350 ( .A1(n19155), .A2(n19386), .B1(n19143), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19132) );
  XNOR2_X1 U22351 ( .A(n19132), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n19396) );
  INV_X1 U22352 ( .A(n19151), .ZN(n19158) );
  NOR4_X1 U22353 ( .A1(n19507), .A2(n17447), .A3(n19134), .A4(n19133), .ZN(
        n19170) );
  NAND2_X1 U22354 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19170), .ZN(
        n19160) );
  NOR2_X1 U22355 ( .A1(n19159), .A2(n19160), .ZN(n19157) );
  NAND2_X1 U22356 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19157), .ZN(
        n19150) );
  OAI21_X1 U22357 ( .B1(n19158), .B2(n19135), .A(n19150), .ZN(n19136) );
  AOI22_X1 U22358 ( .A1(n19138), .A2(n19190), .B1(n19137), .B2(n19136), .ZN(
        n19139) );
  NAND2_X1 U22359 ( .A1(n19477), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n19394) );
  OAI211_X1 U22360 ( .C1(n19178), .C2(n19396), .A(n19139), .B(n19394), .ZN(
        n19140) );
  AOI21_X1 U22361 ( .B1(n19392), .B2(n19164), .A(n19140), .ZN(n19141) );
  OAI21_X1 U22362 ( .B1(n19145), .B2(n19142), .A(n19141), .ZN(P3_U2819) );
  OAI21_X1 U22363 ( .B1(n19155), .B2(n10345), .A(n19143), .ZN(n19144) );
  XNOR2_X1 U22364 ( .A(n19144), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n19403) );
  INV_X1 U22365 ( .A(n19164), .ZN(n19146) );
  AOI221_X1 U22366 ( .B1(n19146), .B2(n19389), .C1(n10345), .C2(n19389), .A(
        n19145), .ZN(n19148) );
  INV_X1 U22367 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20018) );
  NOR2_X1 U22368 ( .A1(n19428), .A2(n20018), .ZN(n19147) );
  AOI211_X1 U22369 ( .C1(n19149), .C2(n19190), .A(n19148), .B(n19147), .ZN(
        n19153) );
  OAI211_X1 U22370 ( .C1(n19157), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19151), .B(n19150), .ZN(n19152) );
  OAI211_X1 U22371 ( .C1(n19403), .C2(n19178), .A(n19153), .B(n19152), .ZN(
        P3_U2820) );
  NAND2_X1 U22372 ( .A1(n19155), .A2(n19154), .ZN(n19156) );
  XNOR2_X1 U22373 ( .A(n19156), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n19412) );
  AOI211_X1 U22374 ( .C1(n19160), .C2(n19159), .A(n19158), .B(n19157), .ZN(
        n19162) );
  NOR2_X1 U22375 ( .A1(n19428), .A2(n20017), .ZN(n19161) );
  AOI211_X1 U22376 ( .C1(n19163), .C2(n19190), .A(n19162), .B(n19161), .ZN(
        n19167) );
  AOI22_X1 U22377 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n19165), .B1(
        n19164), .B2(n10345), .ZN(n19166) );
  OAI211_X1 U22378 ( .C1(n19412), .C2(n19178), .A(n19167), .B(n19166), .ZN(
        P3_U2821) );
  INV_X1 U22379 ( .A(n19168), .ZN(n19171) );
  INV_X1 U22380 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19169) );
  AOI22_X1 U22381 ( .A1(n19171), .A2(n19190), .B1(n19170), .B2(n19169), .ZN(
        n19182) );
  AOI21_X1 U22382 ( .B1(n19173), .B2(n9983), .A(n9731), .ZN(n19418) );
  NAND2_X1 U22383 ( .A1(n19414), .A2(n19174), .ZN(n19175) );
  AND2_X1 U22384 ( .A1(n19176), .A2(n19175), .ZN(n19415) );
  OAI22_X1 U22385 ( .A1(n19415), .A2(n19178), .B1(n19177), .B2(n19414), .ZN(
        n19179) );
  AOI21_X1 U22386 ( .B1(n19220), .B2(n19418), .A(n19179), .ZN(n19181) );
  NAND2_X1 U22387 ( .A1(n19477), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n19425) );
  NOR2_X1 U22388 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n19507), .ZN(
        n19184) );
  OAI21_X1 U22389 ( .B1(n19183), .B2(n19184), .A(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19180) );
  NAND4_X1 U22390 ( .A1(n19182), .A2(n19181), .A3(n19425), .A4(n19180), .ZN(
        P3_U2822) );
  AOI22_X1 U22391 ( .A1(n18058), .A2(n19184), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19183), .ZN(n19193) );
  NAND2_X1 U22392 ( .A1(n19186), .A2(n19185), .ZN(n19187) );
  XOR2_X1 U22393 ( .A(n19187), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n19431) );
  XNOR2_X1 U22394 ( .A(n19188), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19429) );
  OAI22_X1 U22395 ( .A1(n19431), .A2(n19210), .B1(n19429), .B2(n19217), .ZN(
        n19189) );
  AOI21_X1 U22396 ( .B1(n19191), .B2(n19190), .A(n19189), .ZN(n19192) );
  OAI211_X1 U22397 ( .C1(n19216), .C2(n20013), .A(n19193), .B(n19192), .ZN(
        P3_U2823) );
  AOI21_X1 U22398 ( .B1(n17461), .B2(n19202), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19201) );
  OAI22_X1 U22399 ( .A1(n19223), .A2(n19195), .B1(n19217), .B2(n19194), .ZN(
        n19196) );
  AOI211_X1 U22400 ( .C1(n19220), .C2(n19198), .A(n19197), .B(n19196), .ZN(
        n19199) );
  OAI21_X1 U22401 ( .B1(n19201), .B2(n19200), .A(n19199), .ZN(P3_U2825) );
  AND2_X1 U22402 ( .A1(n19202), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19213) );
  OAI22_X1 U22403 ( .A1(n19223), .A2(n19204), .B1(n19217), .B2(n19203), .ZN(
        n19205) );
  AOI221_X1 U22404 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19206), .C1(
        n19213), .C2(n19206), .A(n19205), .ZN(n19208) );
  OAI211_X1 U22405 ( .C1(n19210), .C2(n19209), .A(n19208), .B(n19207), .ZN(
        P3_U2827) );
  XNOR2_X1 U22406 ( .A(n19212), .B(n19211), .ZN(n19462) );
  AOI21_X1 U22407 ( .B1(n19507), .B2(n21725), .A(n19213), .ZN(n19219) );
  XNOR2_X1 U22408 ( .A(n19215), .B(n19214), .ZN(n19458) );
  OAI22_X1 U22409 ( .A1(n19217), .A2(n19458), .B1(n20006), .B2(n19216), .ZN(
        n19218) );
  AOI211_X1 U22410 ( .C1(n19220), .C2(n19462), .A(n19219), .B(n19218), .ZN(
        n19221) );
  OAI21_X1 U22411 ( .B1(n19223), .B2(n19222), .A(n19221), .ZN(P3_U2828) );
  AOI221_X1 U22412 ( .B1(n19262), .B2(n19225), .C1(n19224), .C2(n19225), .A(
        n19459), .ZN(n19228) );
  OAI211_X1 U22413 ( .C1(n19253), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n19226), .ZN(n19227) );
  AOI22_X1 U22414 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n19468), .B1(
        n19228), .B2(n19227), .ZN(n19230) );
  NAND2_X1 U22415 ( .A1(n19477), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n19229) );
  OAI211_X1 U22416 ( .C1(n19231), .C2(n19416), .A(n19230), .B(n19229), .ZN(
        P3_U2835) );
  NOR2_X1 U22417 ( .A1(n19428), .A2(n20048), .ZN(n19239) );
  NAND2_X1 U22418 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19234) );
  INV_X1 U22419 ( .A(n19232), .ZN(n19233) );
  AOI21_X1 U22420 ( .B1(n19440), .B2(n19234), .A(n19233), .ZN(n19237) );
  AOI221_X1 U22421 ( .B1(n19237), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n19236), .C2(n19235), .A(n19459), .ZN(n19238) );
  AOI211_X1 U22422 ( .C1(n19468), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n19239), .B(n19238), .ZN(n19243) );
  AOI22_X1 U22423 ( .A1(n19476), .A2(n19241), .B1(n19377), .B2(n19240), .ZN(
        n19242) );
  OAI211_X1 U22424 ( .C1(n19413), .C2(n19244), .A(n19243), .B(n19242), .ZN(
        P3_U2837) );
  OR3_X1 U22425 ( .A1(n19245), .A2(n19468), .A3(n19262), .ZN(n19249) );
  AOI21_X1 U22426 ( .B1(n19247), .B2(n19377), .A(n19246), .ZN(n19248) );
  OAI221_X1 U22427 ( .B1(n19251), .B2(n19250), .C1(n19251), .C2(n19249), .A(
        n19248), .ZN(P3_U2839) );
  INV_X1 U22428 ( .A(n19252), .ZN(n19260) );
  INV_X1 U22429 ( .A(n19273), .ZN(n19259) );
  AOI21_X1 U22430 ( .B1(n19254), .B2(n19284), .A(n19253), .ZN(n19256) );
  NAND2_X1 U22431 ( .A1(n19322), .A2(n19255), .ZN(n19300) );
  NAND2_X1 U22432 ( .A1(n19384), .A2(n19381), .ZN(n19385) );
  AOI22_X1 U22433 ( .A1(n19469), .A2(n19257), .B1(n19260), .B2(n19385), .ZN(
        n19272) );
  NAND2_X1 U22434 ( .A1(n19477), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19263) );
  OAI211_X1 U22435 ( .C1(n19265), .C2(n19416), .A(n19264), .B(n19263), .ZN(
        P3_U2840) );
  NAND2_X1 U22436 ( .A1(n19267), .A2(n19266), .ZN(n19293) );
  NOR2_X1 U22437 ( .A1(n19477), .A2(n19268), .ZN(n19275) );
  OAI21_X1 U22438 ( .B1(n19321), .B2(n19269), .A(n19390), .ZN(n19270) );
  AND3_X1 U22439 ( .A1(n19271), .A2(n19470), .A3(n19270), .ZN(n19283) );
  OAI211_X1 U22440 ( .C1(n19346), .C2(n19273), .A(n19283), .B(n19272), .ZN(
        n19274) );
  AOI22_X1 U22441 ( .A1(n19377), .A2(n19276), .B1(n19275), .B2(n19274), .ZN(
        n19278) );
  OAI211_X1 U22442 ( .C1(n19279), .C2(n19293), .A(n19278), .B(n19277), .ZN(
        P3_U2841) );
  AOI21_X1 U22443 ( .B1(n19281), .B2(n19377), .A(n19280), .ZN(n19287) );
  INV_X1 U22444 ( .A(n19385), .ZN(n19282) );
  AOI221_X1 U22445 ( .B1(n19284), .B2(n19283), .C1(n19282), .C2(n19283), .A(
        n19477), .ZN(n19290) );
  NOR3_X1 U22446 ( .A1(n19346), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n20102), .ZN(n19285) );
  OAI21_X1 U22447 ( .B1(n19290), .B2(n19285), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19286) );
  OAI211_X1 U22448 ( .C1(n19293), .C2(n19288), .A(n19287), .B(n19286), .ZN(
        P3_U2842) );
  AOI22_X1 U22449 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19290), .B1(
        n19377), .B2(n19289), .ZN(n19292) );
  NAND2_X1 U22450 ( .A1(n19477), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19291) );
  OAI211_X1 U22451 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n19293), .A(
        n19292), .B(n19291), .ZN(P3_U2843) );
  NOR2_X1 U22452 ( .A1(n19438), .A2(n19294), .ZN(n19349) );
  NOR2_X1 U22453 ( .A1(n19349), .A2(n19295), .ZN(n19373) );
  NAND2_X1 U22454 ( .A1(n19296), .A2(n19404), .ZN(n19328) );
  NOR3_X1 U22455 ( .A1(n19298), .A2(n19297), .A3(n10181), .ZN(n19299) );
  NOR2_X1 U22456 ( .A1(n19299), .A2(n19454), .ZN(n19301) );
  AOI211_X1 U22457 ( .C1(n19302), .C2(n19385), .A(n19301), .B(n19300), .ZN(
        n19311) );
  OAI211_X1 U22458 ( .C1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n19454), .A(
        n19311), .B(n19470), .ZN(n19306) );
  NOR2_X1 U22459 ( .A1(n19477), .A2(n19303), .ZN(n19305) );
  AOI22_X1 U22460 ( .A1(n19306), .A2(n19305), .B1(n19377), .B2(n19304), .ZN(
        n19308) );
  OAI211_X1 U22461 ( .C1(n19309), .C2(n19328), .A(n19308), .B(n19307), .ZN(
        P3_U2844) );
  NAND2_X1 U22462 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19310), .ZN(
        n19316) );
  OAI21_X1 U22463 ( .B1(n19311), .B2(n19459), .A(n19466), .ZN(n19313) );
  AOI22_X1 U22464 ( .A1(n19313), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19377), .B2(n19312), .ZN(n19315) );
  OAI211_X1 U22465 ( .C1(n19328), .C2(n19316), .A(n19315), .B(n19314), .ZN(
        P3_U2845) );
  INV_X1 U22466 ( .A(n19317), .ZN(n19319) );
  AOI22_X1 U22467 ( .A1(n19949), .A2(n19319), .B1(n19469), .B2(n19318), .ZN(
        n19405) );
  OAI21_X1 U22468 ( .B1(n19329), .B2(n19398), .A(n19405), .ZN(n19320) );
  AOI211_X1 U22469 ( .C1(n19321), .C2(n19390), .A(n19320), .B(n11880), .ZN(
        n19333) );
  OAI211_X1 U22470 ( .C1(n19323), .C2(n19333), .A(n19470), .B(n19322), .ZN(
        n19324) );
  NAND2_X1 U22471 ( .A1(n19428), .A2(n19324), .ZN(n19327) );
  AOI22_X1 U22472 ( .A1(n19477), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n19377), 
        .B2(n19325), .ZN(n19326) );
  OAI221_X1 U22473 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19328), 
        .C1(n10181), .C2(n19327), .A(n19326), .ZN(P3_U2846) );
  AOI21_X1 U22474 ( .B1(n19329), .B2(n19349), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19335) );
  NAND3_X1 U22475 ( .A1(n19332), .A2(n19331), .A3(n19330), .ZN(n19334) );
  AOI221_X1 U22476 ( .B1(n19335), .B2(n19334), .C1(n19333), .C2(n19334), .A(
        n19459), .ZN(n19336) );
  AOI211_X1 U22477 ( .C1(n19468), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n19337), .B(n19336), .ZN(n19341) );
  NAND3_X1 U22478 ( .A1(n19476), .A2(n19339), .A3(n19338), .ZN(n19340) );
  OAI211_X1 U22479 ( .C1(n19342), .C2(n19416), .A(n19341), .B(n19340), .ZN(
        P3_U2847) );
  AOI22_X1 U22480 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19468), .B1(
        n19477), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n19356) );
  INV_X1 U22481 ( .A(n19398), .ZN(n19344) );
  AOI21_X1 U22482 ( .B1(n19407), .B2(n19343), .A(n19406), .ZN(n19363) );
  AOI21_X1 U22483 ( .B1(n19344), .B2(n19347), .A(n19363), .ZN(n19345) );
  OAI211_X1 U22484 ( .C1(n19346), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n19405), .B(n19345), .ZN(n19350) );
  NOR2_X1 U22485 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19347), .ZN(
        n19348) );
  AOI22_X1 U22486 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n19350), .B1(
        n19349), .B2(n19348), .ZN(n19351) );
  OAI21_X1 U22487 ( .B1(n19381), .B2(n19352), .A(n19351), .ZN(n19354) );
  AOI22_X1 U22488 ( .A1(n19470), .A2(n19354), .B1(n19377), .B2(n19353), .ZN(
        n19355) );
  OAI211_X1 U22489 ( .C1(n19430), .C2(n19357), .A(n19356), .B(n19355), .ZN(
        P3_U2848) );
  AOI21_X1 U22490 ( .B1(n19358), .B2(n19405), .A(n19398), .ZN(n19388) );
  OAI22_X1 U22491 ( .A1(n19360), .A2(n19384), .B1(n19359), .B2(n19381), .ZN(
        n19361) );
  NOR2_X1 U22492 ( .A1(n19388), .A2(n19361), .ZN(n19371) );
  OAI211_X1 U22493 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n19398), .A(
        n19470), .B(n19371), .ZN(n19362) );
  OAI21_X1 U22494 ( .B1(n19363), .B2(n19362), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U22495 ( .A1(n19377), .A2(n19365), .B1(n19404), .B2(n19364), .ZN(
        n19366) );
  OAI221_X1 U22496 ( .B1(n19477), .B2(n19367), .C1(n19428), .C2(n20024), .A(
        n19366), .ZN(P3_U2849) );
  INV_X1 U22497 ( .A(n19407), .ZN(n19369) );
  OAI22_X1 U22498 ( .A1(n19390), .A2(n19380), .B1(n19369), .B2(n19368), .ZN(
        n19370) );
  AOI21_X1 U22499 ( .B1(n19371), .B2(n19370), .A(n19459), .ZN(n19375) );
  OAI21_X1 U22500 ( .B1(n19373), .B2(n19372), .A(n19380), .ZN(n19374) );
  AOI22_X1 U22501 ( .A1(n19377), .A2(n19376), .B1(n19375), .B2(n19374), .ZN(
        n19379) );
  OAI211_X1 U22502 ( .C1(n19466), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P3_U2850) );
  OAI22_X1 U22503 ( .A1(n19384), .A2(n19383), .B1(n19382), .B2(n19381), .ZN(
        n19409) );
  AOI21_X1 U22504 ( .B1(n19386), .B2(n19385), .A(n19409), .ZN(n19387) );
  OAI221_X1 U22505 ( .B1(n19406), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n19406), .C2(n19407), .A(n19387), .ZN(n19400) );
  AOI211_X1 U22506 ( .C1(n19390), .C2(n19389), .A(n19388), .B(n19400), .ZN(
        n19391) );
  OAI21_X1 U22507 ( .B1(n19391), .B2(n19459), .A(n19466), .ZN(n19393) );
  AOI22_X1 U22508 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n19393), .B1(
        n19404), .B2(n19392), .ZN(n19395) );
  OAI211_X1 U22509 ( .C1(n19416), .C2(n19396), .A(n19395), .B(n19394), .ZN(
        P3_U2851) );
  NOR2_X1 U22510 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10345), .ZN(
        n19397) );
  AOI22_X1 U22511 ( .A1(n19477), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n19404), 
        .B2(n19397), .ZN(n19402) );
  OAI211_X1 U22512 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n19398), .A(
        n19405), .B(n19466), .ZN(n19399) );
  OAI211_X1 U22513 ( .C1(n19400), .C2(n19399), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19428), .ZN(n19401) );
  OAI211_X1 U22514 ( .C1(n19403), .C2(n19416), .A(n19402), .B(n19401), .ZN(
        P3_U2852) );
  AOI22_X1 U22515 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n19477), .B1(n19404), 
        .B2(n10345), .ZN(n19411) );
  OAI211_X1 U22516 ( .C1(n19407), .C2(n19406), .A(n19405), .B(n19470), .ZN(
        n19408) );
  OAI211_X1 U22517 ( .C1(n19409), .C2(n19408), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n19428), .ZN(n19410) );
  OAI211_X1 U22518 ( .C1(n19412), .C2(n19416), .A(n19411), .B(n19410), .ZN(
        P3_U2853) );
  OAI22_X1 U22519 ( .A1(n19416), .A2(n19415), .B1(n19414), .B2(n19413), .ZN(
        n19417) );
  AOI21_X1 U22520 ( .B1(n19476), .B2(n19418), .A(n19417), .ZN(n19426) );
  AND2_X1 U22521 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n19419), .ZN(
        n19437) );
  AOI21_X1 U22522 ( .B1(n19421), .B2(n19420), .A(n19468), .ZN(n19422) );
  OAI21_X1 U22523 ( .B1(n19437), .B2(n19459), .A(n19422), .ZN(n19434) );
  OAI211_X1 U22524 ( .C1(n19468), .C2(n19440), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n19434), .ZN(n19424) );
  NAND4_X1 U22525 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n19427), .A4(n9983), .ZN(
        n19423) );
  NAND4_X1 U22526 ( .A1(n19426), .A2(n19425), .A3(n19424), .A4(n19423), .ZN(
        P3_U2854) );
  NAND2_X1 U22527 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19427), .ZN(
        n19436) );
  NOR2_X1 U22528 ( .A1(n19428), .A2(n20013), .ZN(n19433) );
  OAI22_X1 U22529 ( .A1(n19431), .A2(n19430), .B1(n19429), .B2(n19471), .ZN(
        n19432) );
  AOI211_X1 U22530 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n19434), .A(
        n19433), .B(n19432), .ZN(n19435) );
  OAI21_X1 U22531 ( .B1(n19437), .B2(n19436), .A(n19435), .ZN(P3_U2855) );
  NOR2_X1 U22532 ( .A1(n19438), .A2(n19459), .ZN(n19439) );
  NAND2_X1 U22533 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n19439), .ZN(
        n19450) );
  AOI21_X1 U22534 ( .B1(n19441), .B2(n19440), .A(n19468), .ZN(n19448) );
  AND2_X1 U22535 ( .A1(n19443), .A2(n19442), .ZN(n19444) );
  AOI211_X1 U22536 ( .C1(n19476), .C2(n19446), .A(n19445), .B(n19444), .ZN(
        n19447) );
  OAI221_X1 U22537 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19450), .C1(
        n19449), .C2(n19448), .A(n19447), .ZN(P3_U2858) );
  NOR2_X1 U22538 ( .A1(n11932), .A2(n19451), .ZN(n19457) );
  NAND3_X1 U22539 ( .A1(n19949), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19453) );
  OAI211_X1 U22540 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n19454), .A(
        n19453), .B(n19452), .ZN(n19456) );
  AOI221_X1 U22541 ( .B1(n19457), .B2(n19465), .C1(n19456), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n19455), .ZN(n19460) );
  OAI22_X1 U22542 ( .A1(n19460), .A2(n19459), .B1(n19458), .B2(n19471), .ZN(
        n19461) );
  AOI21_X1 U22543 ( .B1(n19476), .B2(n19462), .A(n19461), .ZN(n19464) );
  NAND2_X1 U22544 ( .A1(n19477), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19463) );
  OAI211_X1 U22545 ( .C1(n19466), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P3_U2860) );
  INV_X1 U22546 ( .A(n19467), .ZN(n19475) );
  AOI21_X1 U22547 ( .B1(n19470), .B2(n19469), .A(n19468), .ZN(n19473) );
  OAI22_X1 U22548 ( .A1(n19473), .A2(n19472), .B1(n19471), .B2(n19475), .ZN(
        n19474) );
  AOI21_X1 U22549 ( .B1(n19476), .B2(n19475), .A(n19474), .ZN(n19480) );
  NAND2_X1 U22550 ( .A1(n19477), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n19479) );
  NAND3_X1 U22551 ( .A1(n19480), .A2(n19479), .A3(n19478), .ZN(P3_U2862) );
  AOI211_X1 U22552 ( .C1(n19483), .C2(n19482), .A(n19481), .B(n20102), .ZN(
        n19970) );
  INV_X1 U22553 ( .A(n19566), .ZN(n19525) );
  OAI21_X1 U22554 ( .B1(n19970), .B2(n19525), .A(n19488), .ZN(n19484) );
  OAI221_X1 U22555 ( .B1(n10656), .B2(n20086), .C1(n10656), .C2(n19488), .A(
        n19484), .ZN(P3_U2863) );
  INV_X1 U22556 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19942) );
  NOR2_X1 U22557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19938), .ZN(
        n19657) );
  NOR2_X1 U22558 ( .A1(n19779), .A2(n19657), .ZN(n19486) );
  OAI22_X1 U22559 ( .A1(n19487), .A2(n19942), .B1(n19486), .B2(n19485), .ZN(
        P3_U2866) );
  NOR2_X1 U22560 ( .A1(n19943), .A2(n19488), .ZN(P3_U2867) );
  NAND2_X1 U22561 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19490) );
  NOR2_X1 U22562 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19490), .ZN(
        n19870) );
  NAND2_X1 U22563 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19870), .ZN(
        n19914) );
  NAND2_X1 U22564 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19871), .ZN(n19875) );
  NOR2_X2 U22565 ( .A1(n19565), .A2(n19489), .ZN(n19866) );
  NOR2_X1 U22566 ( .A1(n19755), .A2(n10656), .ZN(n19932) );
  INV_X1 U22567 ( .A(n19932), .ZN(n19757) );
  NOR2_X2 U22568 ( .A1(n19757), .A2(n19490), .ZN(n19920) );
  INV_X1 U22569 ( .A(n19920), .ZN(n19882) );
  NAND2_X1 U22570 ( .A1(n19755), .A2(n10656), .ZN(n19934) );
  NAND2_X1 U22571 ( .A1(n19938), .A2(n19942), .ZN(n19610) );
  NOR2_X1 U22572 ( .A1(n19934), .A2(n19610), .ZN(n19556) );
  INV_X1 U22573 ( .A(n19556), .ZN(n19587) );
  NAND2_X1 U22574 ( .A1(n19882), .A2(n19587), .ZN(n19544) );
  AND2_X1 U22575 ( .A1(n19865), .A2(n19544), .ZN(n19519) );
  AND2_X1 U22576 ( .A1(n19871), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19867) );
  NAND2_X1 U22577 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n10656), .ZN(
        n19633) );
  NOR2_X2 U22578 ( .A1(n19490), .A2(n19633), .ZN(n19860) );
  AOI22_X1 U22579 ( .A1(n19866), .A2(n19519), .B1(n19867), .B2(n19860), .ZN(
        n19495) );
  INV_X1 U22580 ( .A(n19633), .ZN(n19731) );
  NOR2_X1 U22581 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n10656), .ZN(
        n19705) );
  NOR2_X1 U22582 ( .A1(n19731), .A2(n19705), .ZN(n19781) );
  NOR2_X1 U22583 ( .A1(n19781), .A2(n19490), .ZN(n19838) );
  AOI21_X1 U22584 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n19565), .ZN(n19835) );
  AOI22_X1 U22585 ( .A1(n19871), .A2(n19838), .B1(n19835), .B2(n19544), .ZN(
        n19522) );
  NAND2_X1 U22586 ( .A1(n19492), .A2(n19491), .ZN(n19520) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19872), .ZN(n19494) );
  OAI211_X1 U22588 ( .C1(n19914), .C2(n19875), .A(n19495), .B(n19494), .ZN(
        P3_U2868) );
  INV_X1 U22589 ( .A(n19860), .ZN(n19850) );
  NAND2_X1 U22590 ( .A1(n19871), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19811) );
  INV_X1 U22591 ( .A(n19914), .ZN(n19918) );
  NOR2_X2 U22592 ( .A1(n16800), .A2(n19507), .ZN(n19878) );
  AND2_X1 U22593 ( .A1(n19783), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U22594 ( .A1(n19918), .A2(n19878), .B1(n19519), .B2(n19876), .ZN(
        n19498) );
  NOR2_X1 U22595 ( .A1(n19496), .A2(n19520), .ZN(n19808) );
  AOI22_X1 U22596 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19808), .ZN(n19497) );
  OAI211_X1 U22597 ( .C1(n19850), .C2(n19811), .A(n19498), .B(n19497), .ZN(
        P3_U2869) );
  NOR2_X2 U22598 ( .A1(n19565), .A2(n19499), .ZN(n19883) );
  AND2_X1 U22599 ( .A1(n19871), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U22600 ( .A1(n19519), .A2(n19883), .B1(n19860), .B2(n19884), .ZN(
        n19502) );
  AOI22_X1 U22601 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19885), .ZN(n19501) );
  OAI211_X1 U22602 ( .C1(n19914), .C2(n19888), .A(n19502), .B(n19501), .ZN(
        P3_U2870) );
  NAND2_X1 U22603 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19871), .ZN(n19894) );
  AND2_X1 U22604 ( .A1(n19871), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U22605 ( .A1(n19519), .A2(n19889), .B1(n19860), .B2(n19890), .ZN(
        n19505) );
  AOI22_X1 U22606 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19891), .ZN(n19504) );
  OAI211_X1 U22607 ( .C1(n19914), .C2(n19894), .A(n19505), .B(n19504), .ZN(
        P3_U2871) );
  NAND2_X1 U22608 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19871), .ZN(n19695) );
  NOR2_X2 U22609 ( .A1(n19565), .A2(n19506), .ZN(n19895) );
  NOR2_X1 U22610 ( .A1(n19507), .A2(n21470), .ZN(n19692) );
  AOI22_X1 U22611 ( .A1(n19519), .A2(n19895), .B1(n19860), .B2(n19692), .ZN(
        n19510) );
  NOR2_X2 U22612 ( .A1(n19508), .A2(n19520), .ZN(n19897) );
  AOI22_X1 U22613 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19897), .ZN(n19509) );
  OAI211_X1 U22614 ( .C1(n19914), .C2(n19695), .A(n19510), .B(n19509), .ZN(
        P3_U2872) );
  NAND2_X1 U22615 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19871), .ZN(n19824) );
  AND2_X1 U22616 ( .A1(n19783), .A2(BUF2_REG_5__SCAN_IN), .ZN(n19901) );
  NAND2_X1 U22617 ( .A1(n19871), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19906) );
  INV_X1 U22618 ( .A(n19906), .ZN(n19821) );
  AOI22_X1 U22619 ( .A1(n19519), .A2(n19901), .B1(n19860), .B2(n19821), .ZN(
        n19513) );
  NOR2_X2 U22620 ( .A1(n19511), .A2(n19520), .ZN(n19903) );
  AOI22_X1 U22621 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19903), .ZN(n19512) );
  OAI211_X1 U22622 ( .C1(n19914), .C2(n19824), .A(n19513), .B(n19512), .ZN(
        P3_U2873) );
  NAND2_X1 U22623 ( .A1(n19871), .A2(BUF2_REG_22__SCAN_IN), .ZN(n19913) );
  NAND2_X1 U22624 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19871), .ZN(n19828) );
  INV_X1 U22625 ( .A(n19828), .ZN(n19908) );
  NOR2_X2 U22626 ( .A1(n19565), .A2(n19514), .ZN(n19909) );
  AOI22_X1 U22627 ( .A1(n19918), .A2(n19908), .B1(n19519), .B2(n19909), .ZN(
        n19517) );
  NOR2_X2 U22628 ( .A1(n19515), .A2(n19520), .ZN(n19910) );
  AOI22_X1 U22629 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19910), .ZN(n19516) );
  OAI211_X1 U22630 ( .C1(n19850), .C2(n19913), .A(n19517), .B(n19516), .ZN(
        P3_U2874) );
  NAND2_X1 U22631 ( .A1(n19871), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19925) );
  INV_X1 U22632 ( .A(n19925), .ZN(n19858) );
  NOR2_X2 U22633 ( .A1(n19565), .A2(n19518), .ZN(n19916) );
  AOI22_X1 U22634 ( .A1(n19918), .A2(n19858), .B1(n19519), .B2(n19916), .ZN(
        n19524) );
  NOR2_X2 U22635 ( .A1(n19521), .A2(n19520), .ZN(n19919) );
  AOI22_X1 U22636 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19522), .B1(
        n19580), .B2(n19919), .ZN(n19523) );
  OAI211_X1 U22637 ( .C1(n19850), .C2(n19864), .A(n19524), .B(n19523), .ZN(
        P3_U2875) );
  INV_X1 U22638 ( .A(n19610), .ZN(n19567) );
  NAND2_X1 U22639 ( .A1(n19567), .A2(n19705), .ZN(n19609) );
  INV_X1 U22640 ( .A(n19875), .ZN(n19778) );
  NAND2_X1 U22641 ( .A1(n19755), .A2(n19865), .ZN(n19706) );
  NOR2_X1 U22642 ( .A1(n19610), .A2(n19706), .ZN(n19540) );
  AOI22_X1 U22643 ( .A1(n19778), .A2(n19860), .B1(n19866), .B2(n19540), .ZN(
        n19527) );
  NOR2_X1 U22644 ( .A1(n19942), .A2(n19707), .ZN(n19869) );
  NOR2_X1 U22645 ( .A1(n19565), .A2(n19525), .ZN(n19868) );
  AND2_X1 U22646 ( .A1(n19755), .A2(n19868), .ZN(n19611) );
  AOI22_X1 U22647 ( .A1(n19871), .A2(n19869), .B1(n19567), .B2(n19611), .ZN(
        n19541) );
  AOI22_X1 U22648 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19541), .B1(
        n19920), .B2(n19867), .ZN(n19526) );
  OAI211_X1 U22649 ( .C1(n19786), .C2(n19609), .A(n19527), .B(n19526), .ZN(
        P3_U2876) );
  INV_X1 U22650 ( .A(n19808), .ZN(n19881) );
  INV_X1 U22651 ( .A(n19811), .ZN(n19877) );
  AOI22_X1 U22652 ( .A1(n19920), .A2(n19877), .B1(n19876), .B2(n19540), .ZN(
        n19529) );
  AOI22_X1 U22653 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19541), .B1(
        n19860), .B2(n19878), .ZN(n19528) );
  OAI211_X1 U22654 ( .C1(n19881), .C2(n19609), .A(n19529), .B(n19528), .ZN(
        P3_U2877) );
  AOI22_X1 U22655 ( .A1(n19920), .A2(n19884), .B1(n19883), .B2(n19540), .ZN(
        n19531) );
  AOI22_X1 U22656 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19541), .B1(
        n19885), .B2(n19600), .ZN(n19530) );
  OAI211_X1 U22657 ( .C1(n19850), .C2(n19888), .A(n19531), .B(n19530), .ZN(
        P3_U2878) );
  INV_X1 U22658 ( .A(n19894), .ZN(n19846) );
  AOI22_X1 U22659 ( .A1(n19860), .A2(n19846), .B1(n19889), .B2(n19540), .ZN(
        n19533) );
  AOI22_X1 U22660 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19541), .B1(
        n19920), .B2(n19890), .ZN(n19532) );
  OAI211_X1 U22661 ( .C1(n19849), .C2(n19609), .A(n19533), .B(n19532), .ZN(
        P3_U2879) );
  AOI22_X1 U22662 ( .A1(n19920), .A2(n19692), .B1(n19895), .B2(n19540), .ZN(
        n19535) );
  AOI22_X1 U22663 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19541), .B1(
        n19897), .B2(n19600), .ZN(n19534) );
  OAI211_X1 U22664 ( .C1(n19850), .C2(n19695), .A(n19535), .B(n19534), .ZN(
        P3_U2880) );
  AOI22_X1 U22665 ( .A1(n19920), .A2(n19821), .B1(n19901), .B2(n19540), .ZN(
        n19537) );
  AOI22_X1 U22666 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19541), .B1(
        n19903), .B2(n19600), .ZN(n19536) );
  OAI211_X1 U22667 ( .C1(n19850), .C2(n19824), .A(n19537), .B(n19536), .ZN(
        P3_U2881) );
  INV_X1 U22668 ( .A(n19913), .ZN(n19825) );
  AOI22_X1 U22669 ( .A1(n19920), .A2(n19825), .B1(n19909), .B2(n19540), .ZN(
        n19539) );
  AOI22_X1 U22670 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19541), .B1(
        n19910), .B2(n19600), .ZN(n19538) );
  OAI211_X1 U22671 ( .C1(n19850), .C2(n19828), .A(n19539), .B(n19538), .ZN(
        P3_U2882) );
  INV_X1 U22672 ( .A(n19864), .ZN(n19917) );
  AOI22_X1 U22673 ( .A1(n19920), .A2(n19917), .B1(n19916), .B2(n19540), .ZN(
        n19543) );
  AOI22_X1 U22674 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19541), .B1(
        n19919), .B2(n19600), .ZN(n19542) );
  OAI211_X1 U22675 ( .C1(n19850), .C2(n19925), .A(n19543), .B(n19542), .ZN(
        P3_U2883) );
  NAND2_X1 U22676 ( .A1(n19567), .A2(n19731), .ZN(n19627) );
  NOR2_X1 U22677 ( .A1(n19600), .A2(n19628), .ZN(n19588) );
  NOR2_X1 U22678 ( .A1(n19978), .A2(n19588), .ZN(n19561) );
  AOI22_X1 U22679 ( .A1(n19778), .A2(n19920), .B1(n19866), .B2(n19561), .ZN(
        n19547) );
  INV_X1 U22680 ( .A(n19588), .ZN(n19545) );
  OAI221_X1 U22681 ( .B1(n19545), .B2(n19837), .C1(n19545), .C2(n19544), .A(
        n19835), .ZN(n19562) );
  AOI22_X1 U22682 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19562), .B1(
        n19580), .B2(n19867), .ZN(n19546) );
  OAI211_X1 U22683 ( .C1(n19786), .C2(n19627), .A(n19547), .B(n19546), .ZN(
        P3_U2884) );
  AOI22_X1 U22684 ( .A1(n19920), .A2(n19878), .B1(n19876), .B2(n19561), .ZN(
        n19549) );
  AOI22_X1 U22685 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19562), .B1(
        n19580), .B2(n19877), .ZN(n19548) );
  OAI211_X1 U22686 ( .C1(n19881), .C2(n19627), .A(n19549), .B(n19548), .ZN(
        P3_U2885) );
  AOI22_X1 U22687 ( .A1(n19920), .A2(n19812), .B1(n19883), .B2(n19561), .ZN(
        n19551) );
  AOI22_X1 U22688 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19562), .B1(
        n19580), .B2(n19884), .ZN(n19550) );
  OAI211_X1 U22689 ( .C1(n19815), .C2(n19627), .A(n19551), .B(n19550), .ZN(
        P3_U2886) );
  AOI22_X1 U22690 ( .A1(n19920), .A2(n19846), .B1(n19889), .B2(n19561), .ZN(
        n19553) );
  AOI22_X1 U22691 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19562), .B1(
        n19580), .B2(n19890), .ZN(n19552) );
  OAI211_X1 U22692 ( .C1(n19849), .C2(n19627), .A(n19553), .B(n19552), .ZN(
        P3_U2887) );
  AOI22_X1 U22693 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19562), .B1(
        n19895), .B2(n19561), .ZN(n19555) );
  AOI22_X1 U22694 ( .A1(n19580), .A2(n19692), .B1(n19897), .B2(n19628), .ZN(
        n19554) );
  OAI211_X1 U22695 ( .C1(n19882), .C2(n19695), .A(n19555), .B(n19554), .ZN(
        P3_U2888) );
  AOI22_X1 U22696 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19562), .B1(
        n19901), .B2(n19561), .ZN(n19558) );
  AOI22_X1 U22697 ( .A1(n19556), .A2(n19821), .B1(n19903), .B2(n19628), .ZN(
        n19557) );
  OAI211_X1 U22698 ( .C1(n19882), .C2(n19824), .A(n19558), .B(n19557), .ZN(
        P3_U2889) );
  AOI22_X1 U22699 ( .A1(n19580), .A2(n19825), .B1(n19909), .B2(n19561), .ZN(
        n19560) );
  AOI22_X1 U22700 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19562), .B1(
        n19910), .B2(n19628), .ZN(n19559) );
  OAI211_X1 U22701 ( .C1(n19882), .C2(n19828), .A(n19560), .B(n19559), .ZN(
        P3_U2890) );
  AOI22_X1 U22702 ( .A1(n19580), .A2(n19917), .B1(n19916), .B2(n19561), .ZN(
        n19564) );
  AOI22_X1 U22703 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19562), .B1(
        n19919), .B2(n19628), .ZN(n19563) );
  OAI211_X1 U22704 ( .C1(n19882), .C2(n19925), .A(n19564), .B(n19563), .ZN(
        P3_U2891) );
  NAND2_X1 U22705 ( .A1(n19932), .A2(n19567), .ZN(n19650) );
  INV_X1 U22706 ( .A(n19837), .ZN(n19732) );
  AOI21_X1 U22707 ( .B1(n19755), .B2(n19732), .A(n19565), .ZN(n19656) );
  NAND3_X1 U22708 ( .A1(n19567), .A2(n19656), .A3(n19566), .ZN(n19584) );
  AOI22_X1 U22709 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19584), .B1(
        n19866), .B2(n19583), .ZN(n19569) );
  AOI22_X1 U22710 ( .A1(n19778), .A2(n19580), .B1(n19867), .B2(n19600), .ZN(
        n19568) );
  OAI211_X1 U22711 ( .C1(n19786), .C2(n19650), .A(n19569), .B(n19568), .ZN(
        P3_U2892) );
  AOI22_X1 U22712 ( .A1(n19877), .A2(n19600), .B1(n19876), .B2(n19583), .ZN(
        n19571) );
  AOI22_X1 U22713 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19584), .B1(
        n19580), .B2(n19878), .ZN(n19570) );
  OAI211_X1 U22714 ( .C1(n19881), .C2(n19650), .A(n19571), .B(n19570), .ZN(
        P3_U2893) );
  AOI22_X1 U22715 ( .A1(n19580), .A2(n19812), .B1(n19883), .B2(n19583), .ZN(
        n19573) );
  AOI22_X1 U22716 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19584), .B1(
        n19884), .B2(n19600), .ZN(n19572) );
  OAI211_X1 U22717 ( .C1(n19815), .C2(n19650), .A(n19573), .B(n19572), .ZN(
        P3_U2894) );
  AOI22_X1 U22718 ( .A1(n19580), .A2(n19846), .B1(n19889), .B2(n19583), .ZN(
        n19575) );
  AOI22_X1 U22719 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19584), .B1(
        n19890), .B2(n19600), .ZN(n19574) );
  OAI211_X1 U22720 ( .C1(n19849), .C2(n19650), .A(n19575), .B(n19574), .ZN(
        P3_U2895) );
  AOI22_X1 U22721 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19584), .B1(
        n19895), .B2(n19583), .ZN(n19577) );
  AOI22_X1 U22722 ( .A1(n19897), .A2(n19651), .B1(n19692), .B2(n19600), .ZN(
        n19576) );
  OAI211_X1 U22723 ( .C1(n19587), .C2(n19695), .A(n19577), .B(n19576), .ZN(
        P3_U2896) );
  INV_X1 U22724 ( .A(n19824), .ZN(n19902) );
  AOI22_X1 U22725 ( .A1(n19580), .A2(n19902), .B1(n19901), .B2(n19583), .ZN(
        n19579) );
  AOI22_X1 U22726 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19584), .B1(
        n19903), .B2(n19651), .ZN(n19578) );
  OAI211_X1 U22727 ( .C1(n19906), .C2(n19609), .A(n19579), .B(n19578), .ZN(
        P3_U2897) );
  AOI22_X1 U22728 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19584), .B1(
        n19909), .B2(n19583), .ZN(n19582) );
  AOI22_X1 U22729 ( .A1(n19580), .A2(n19908), .B1(n19910), .B2(n19651), .ZN(
        n19581) );
  OAI211_X1 U22730 ( .C1(n19913), .C2(n19609), .A(n19582), .B(n19581), .ZN(
        P3_U2898) );
  AOI22_X1 U22731 ( .A1(n19917), .A2(n19600), .B1(n19916), .B2(n19583), .ZN(
        n19586) );
  AOI22_X1 U22732 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19584), .B1(
        n19919), .B2(n19651), .ZN(n19585) );
  OAI211_X1 U22733 ( .C1(n19587), .C2(n19925), .A(n19586), .B(n19585), .ZN(
        P3_U2899) );
  INV_X1 U22734 ( .A(n19934), .ZN(n19679) );
  NAND2_X1 U22735 ( .A1(n19679), .A2(n19657), .ZN(n19661) );
  AOI21_X1 U22736 ( .B1(n19650), .B2(n19661), .A(n19978), .ZN(n19605) );
  AOI22_X1 U22737 ( .A1(n19778), .A2(n19600), .B1(n19866), .B2(n19605), .ZN(
        n19591) );
  INV_X1 U22738 ( .A(n19661), .ZN(n19676) );
  AOI221_X1 U22739 ( .B1(n19588), .B2(n19650), .C1(n19732), .C2(n19650), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19589) );
  OAI21_X1 U22740 ( .B1(n19676), .B2(n19589), .A(n19783), .ZN(n19606) );
  AOI22_X1 U22741 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19606), .B1(
        n19867), .B2(n19628), .ZN(n19590) );
  OAI211_X1 U22742 ( .C1(n19786), .C2(n19661), .A(n19591), .B(n19590), .ZN(
        P3_U2900) );
  AOI22_X1 U22743 ( .A1(n19877), .A2(n19628), .B1(n19876), .B2(n19605), .ZN(
        n19593) );
  AOI22_X1 U22744 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19606), .B1(
        n19878), .B2(n19600), .ZN(n19592) );
  OAI211_X1 U22745 ( .C1(n19881), .C2(n19661), .A(n19593), .B(n19592), .ZN(
        P3_U2901) );
  AOI22_X1 U22746 ( .A1(n19884), .A2(n19628), .B1(n19883), .B2(n19605), .ZN(
        n19595) );
  AOI22_X1 U22747 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19606), .B1(
        n19885), .B2(n19676), .ZN(n19594) );
  OAI211_X1 U22748 ( .C1(n19888), .C2(n19609), .A(n19595), .B(n19594), .ZN(
        P3_U2902) );
  AOI22_X1 U22749 ( .A1(n19890), .A2(n19628), .B1(n19889), .B2(n19605), .ZN(
        n19597) );
  AOI22_X1 U22750 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19606), .B1(
        n19891), .B2(n19676), .ZN(n19596) );
  OAI211_X1 U22751 ( .C1(n19894), .C2(n19609), .A(n19597), .B(n19596), .ZN(
        P3_U2903) );
  AOI22_X1 U22752 ( .A1(n19692), .A2(n19628), .B1(n19895), .B2(n19605), .ZN(
        n19599) );
  AOI22_X1 U22753 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19606), .B1(
        n19897), .B2(n19676), .ZN(n19598) );
  OAI211_X1 U22754 ( .C1(n19695), .C2(n19609), .A(n19599), .B(n19598), .ZN(
        P3_U2904) );
  AOI22_X1 U22755 ( .A1(n19902), .A2(n19600), .B1(n19901), .B2(n19605), .ZN(
        n19602) );
  AOI22_X1 U22756 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19606), .B1(
        n19903), .B2(n19676), .ZN(n19601) );
  OAI211_X1 U22757 ( .C1(n19906), .C2(n19627), .A(n19602), .B(n19601), .ZN(
        P3_U2905) );
  AOI22_X1 U22758 ( .A1(n19825), .A2(n19628), .B1(n19909), .B2(n19605), .ZN(
        n19604) );
  AOI22_X1 U22759 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19606), .B1(
        n19910), .B2(n19676), .ZN(n19603) );
  OAI211_X1 U22760 ( .C1(n19828), .C2(n19609), .A(n19604), .B(n19603), .ZN(
        P3_U2906) );
  AOI22_X1 U22761 ( .A1(n19917), .A2(n19628), .B1(n19916), .B2(n19605), .ZN(
        n19608) );
  AOI22_X1 U22762 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19606), .B1(
        n19919), .B2(n19676), .ZN(n19607) );
  OAI211_X1 U22763 ( .C1(n19925), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        P3_U2907) );
  NOR2_X1 U22764 ( .A1(n19658), .A2(n19706), .ZN(n19629) );
  AOI22_X1 U22765 ( .A1(n19866), .A2(n19629), .B1(n19867), .B2(n19651), .ZN(
        n19614) );
  NOR2_X1 U22766 ( .A1(n19755), .A2(n19610), .ZN(n19612) );
  AOI22_X1 U22767 ( .A1(n19871), .A2(n19612), .B1(n19657), .B2(n19611), .ZN(
        n19630) );
  AOI22_X1 U22768 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19630), .B1(
        n19778), .B2(n19628), .ZN(n19613) );
  OAI211_X1 U22769 ( .C1(n19786), .C2(n19704), .A(n19614), .B(n19613), .ZN(
        P3_U2908) );
  AOI22_X1 U22770 ( .A1(n19878), .A2(n19628), .B1(n19876), .B2(n19629), .ZN(
        n19616) );
  AOI22_X1 U22771 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19630), .B1(
        n19877), .B2(n19651), .ZN(n19615) );
  OAI211_X1 U22772 ( .C1(n19881), .C2(n19704), .A(n19616), .B(n19615), .ZN(
        P3_U2909) );
  AOI22_X1 U22773 ( .A1(n19812), .A2(n19628), .B1(n19883), .B2(n19629), .ZN(
        n19618) );
  AOI22_X1 U22774 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19630), .B1(
        n19884), .B2(n19651), .ZN(n19617) );
  OAI211_X1 U22775 ( .C1(n19815), .C2(n19704), .A(n19618), .B(n19617), .ZN(
        P3_U2910) );
  AOI22_X1 U22776 ( .A1(n19890), .A2(n19651), .B1(n19889), .B2(n19629), .ZN(
        n19620) );
  AOI22_X1 U22777 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19630), .B1(
        n19846), .B2(n19628), .ZN(n19619) );
  OAI211_X1 U22778 ( .C1(n19849), .C2(n19704), .A(n19620), .B(n19619), .ZN(
        P3_U2911) );
  AOI22_X1 U22779 ( .A1(n19692), .A2(n19651), .B1(n19895), .B2(n19629), .ZN(
        n19622) );
  AOI22_X1 U22780 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19630), .B1(
        n19897), .B2(n19685), .ZN(n19621) );
  OAI211_X1 U22781 ( .C1(n19695), .C2(n19627), .A(n19622), .B(n19621), .ZN(
        P3_U2912) );
  AOI22_X1 U22782 ( .A1(n19821), .A2(n19651), .B1(n19901), .B2(n19629), .ZN(
        n19624) );
  AOI22_X1 U22783 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19630), .B1(
        n19903), .B2(n19685), .ZN(n19623) );
  OAI211_X1 U22784 ( .C1(n19824), .C2(n19627), .A(n19624), .B(n19623), .ZN(
        P3_U2913) );
  AOI22_X1 U22785 ( .A1(n19825), .A2(n19651), .B1(n19909), .B2(n19629), .ZN(
        n19626) );
  AOI22_X1 U22786 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19630), .B1(
        n19910), .B2(n19685), .ZN(n19625) );
  OAI211_X1 U22787 ( .C1(n19828), .C2(n19627), .A(n19626), .B(n19625), .ZN(
        P3_U2914) );
  AOI22_X1 U22788 ( .A1(n19916), .A2(n19629), .B1(n19858), .B2(n19628), .ZN(
        n19632) );
  AOI22_X1 U22789 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19630), .B1(
        n19919), .B2(n19685), .ZN(n19631) );
  OAI211_X1 U22790 ( .C1(n19864), .C2(n19650), .A(n19632), .B(n19631), .ZN(
        P3_U2915) );
  NOR2_X1 U22791 ( .A1(n19658), .A2(n19633), .ZN(n19726) );
  INV_X1 U22792 ( .A(n19726), .ZN(n19723) );
  NOR2_X1 U22793 ( .A1(n19651), .A2(n19676), .ZN(n19634) );
  NOR2_X1 U22794 ( .A1(n19685), .A2(n19718), .ZN(n19681) );
  OAI21_X1 U22795 ( .B1(n19634), .B2(n19732), .A(n19681), .ZN(n19635) );
  OAI211_X1 U22796 ( .C1(n19718), .C2(n20070), .A(n19783), .B(n19635), .ZN(
        n19653) );
  NOR2_X1 U22797 ( .A1(n19978), .A2(n19681), .ZN(n19652) );
  AOI22_X1 U22798 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19653), .B1(
        n19866), .B2(n19652), .ZN(n19637) );
  AOI22_X1 U22799 ( .A1(n19872), .A2(n19718), .B1(n19867), .B2(n19676), .ZN(
        n19636) );
  OAI211_X1 U22800 ( .C1(n19875), .C2(n19650), .A(n19637), .B(n19636), .ZN(
        P3_U2916) );
  AOI22_X1 U22801 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19653), .B1(
        n19876), .B2(n19652), .ZN(n19639) );
  AOI22_X1 U22802 ( .A1(n19808), .A2(n19718), .B1(n19878), .B2(n19651), .ZN(
        n19638) );
  OAI211_X1 U22803 ( .C1(n19811), .C2(n19661), .A(n19639), .B(n19638), .ZN(
        P3_U2917) );
  AOI22_X1 U22804 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19653), .B1(
        n19883), .B2(n19652), .ZN(n19641) );
  AOI22_X1 U22805 ( .A1(n19885), .A2(n19718), .B1(n19884), .B2(n19676), .ZN(
        n19640) );
  OAI211_X1 U22806 ( .C1(n19888), .C2(n19650), .A(n19641), .B(n19640), .ZN(
        P3_U2918) );
  AOI22_X1 U22807 ( .A1(n19890), .A2(n19676), .B1(n19889), .B2(n19652), .ZN(
        n19643) );
  AOI22_X1 U22808 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19653), .B1(
        n19891), .B2(n19718), .ZN(n19642) );
  OAI211_X1 U22809 ( .C1(n19894), .C2(n19650), .A(n19643), .B(n19642), .ZN(
        P3_U2919) );
  INV_X1 U22810 ( .A(n19692), .ZN(n19900) );
  INV_X1 U22811 ( .A(n19695), .ZN(n19896) );
  AOI22_X1 U22812 ( .A1(n19896), .A2(n19651), .B1(n19895), .B2(n19652), .ZN(
        n19645) );
  AOI22_X1 U22813 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19653), .B1(
        n19897), .B2(n19718), .ZN(n19644) );
  OAI211_X1 U22814 ( .C1(n19900), .C2(n19661), .A(n19645), .B(n19644), .ZN(
        P3_U2920) );
  AOI22_X1 U22815 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19653), .B1(
        n19901), .B2(n19652), .ZN(n19647) );
  AOI22_X1 U22816 ( .A1(n19902), .A2(n19651), .B1(n19903), .B2(n19726), .ZN(
        n19646) );
  OAI211_X1 U22817 ( .C1(n19906), .C2(n19661), .A(n19647), .B(n19646), .ZN(
        P3_U2921) );
  AOI22_X1 U22818 ( .A1(n19825), .A2(n19676), .B1(n19909), .B2(n19652), .ZN(
        n19649) );
  AOI22_X1 U22819 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19653), .B1(
        n19910), .B2(n19726), .ZN(n19648) );
  OAI211_X1 U22820 ( .C1(n19828), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P3_U2922) );
  AOI22_X1 U22821 ( .A1(n19916), .A2(n19652), .B1(n19858), .B2(n19651), .ZN(
        n19655) );
  AOI22_X1 U22822 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19653), .B1(
        n19919), .B2(n19726), .ZN(n19654) );
  OAI211_X1 U22823 ( .C1(n19864), .C2(n19661), .A(n19655), .B(n19654), .ZN(
        P3_U2923) );
  AOI22_X1 U22824 ( .A1(n19866), .A2(n19674), .B1(n19867), .B2(n19685), .ZN(
        n19660) );
  OAI211_X1 U22825 ( .C1(n19932), .C2(n20070), .A(n19657), .B(n19656), .ZN(
        n19675) );
  NOR2_X2 U22826 ( .A1(n19757), .A2(n19658), .ZN(n19750) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19675), .B1(
        n19872), .B2(n19750), .ZN(n19659) );
  OAI211_X1 U22828 ( .C1(n19875), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P3_U2924) );
  AOI22_X1 U22829 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19675), .B1(
        n19876), .B2(n19674), .ZN(n19663) );
  AOI22_X1 U22830 ( .A1(n19808), .A2(n19750), .B1(n19878), .B2(n19676), .ZN(
        n19662) );
  OAI211_X1 U22831 ( .C1(n19811), .C2(n19704), .A(n19663), .B(n19662), .ZN(
        P3_U2925) );
  AOI22_X1 U22832 ( .A1(n19812), .A2(n19676), .B1(n19883), .B2(n19674), .ZN(
        n19665) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19675), .B1(
        n19884), .B2(n19685), .ZN(n19664) );
  OAI211_X1 U22834 ( .C1(n19815), .C2(n19749), .A(n19665), .B(n19664), .ZN(
        P3_U2926) );
  AOI22_X1 U22835 ( .A1(n19846), .A2(n19676), .B1(n19889), .B2(n19674), .ZN(
        n19667) );
  AOI22_X1 U22836 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19675), .B1(
        n19890), .B2(n19685), .ZN(n19666) );
  OAI211_X1 U22837 ( .C1(n19849), .C2(n19749), .A(n19667), .B(n19666), .ZN(
        P3_U2927) );
  AOI22_X1 U22838 ( .A1(n19896), .A2(n19676), .B1(n19895), .B2(n19674), .ZN(
        n19669) );
  AOI22_X1 U22839 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19675), .B1(
        n19897), .B2(n19750), .ZN(n19668) );
  OAI211_X1 U22840 ( .C1(n19900), .C2(n19704), .A(n19669), .B(n19668), .ZN(
        P3_U2928) );
  AOI22_X1 U22841 ( .A1(n19902), .A2(n19676), .B1(n19901), .B2(n19674), .ZN(
        n19671) );
  AOI22_X1 U22842 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19675), .B1(
        n19903), .B2(n19750), .ZN(n19670) );
  OAI211_X1 U22843 ( .C1(n19906), .C2(n19704), .A(n19671), .B(n19670), .ZN(
        P3_U2929) );
  AOI22_X1 U22844 ( .A1(n19909), .A2(n19674), .B1(n19908), .B2(n19676), .ZN(
        n19673) );
  AOI22_X1 U22845 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19675), .B1(
        n19910), .B2(n19750), .ZN(n19672) );
  OAI211_X1 U22846 ( .C1(n19913), .C2(n19704), .A(n19673), .B(n19672), .ZN(
        P3_U2930) );
  AOI22_X1 U22847 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19675), .B1(
        n19916), .B2(n19674), .ZN(n19678) );
  AOI22_X1 U22848 ( .A1(n19919), .A2(n19750), .B1(n19858), .B2(n19676), .ZN(
        n19677) );
  OAI211_X1 U22849 ( .C1(n19864), .C2(n19704), .A(n19678), .B(n19677), .ZN(
        P3_U2931) );
  NAND2_X1 U22850 ( .A1(n19679), .A2(n19779), .ZN(n19772) );
  NOR2_X1 U22851 ( .A1(n19750), .A2(n19773), .ZN(n19733) );
  NOR2_X1 U22852 ( .A1(n19978), .A2(n19733), .ZN(n19700) );
  AOI22_X1 U22853 ( .A1(n19866), .A2(n19700), .B1(n19867), .B2(n19726), .ZN(
        n19684) );
  INV_X1 U22854 ( .A(n19835), .ZN(n19680) );
  AOI221_X1 U22855 ( .B1(n19733), .B2(n19732), .C1(n19733), .C2(n19681), .A(
        n19680), .ZN(n19682) );
  INV_X1 U22856 ( .A(n19682), .ZN(n19701) );
  AOI22_X1 U22857 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19701), .B1(
        n19778), .B2(n19685), .ZN(n19683) );
  OAI211_X1 U22858 ( .C1(n19786), .C2(n19772), .A(n19684), .B(n19683), .ZN(
        P3_U2932) );
  AOI22_X1 U22859 ( .A1(n19877), .A2(n19718), .B1(n19876), .B2(n19700), .ZN(
        n19687) );
  AOI22_X1 U22860 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19701), .B1(
        n19878), .B2(n19685), .ZN(n19686) );
  OAI211_X1 U22861 ( .C1(n19881), .C2(n19772), .A(n19687), .B(n19686), .ZN(
        P3_U2933) );
  AOI22_X1 U22862 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19701), .B1(
        n19883), .B2(n19700), .ZN(n19689) );
  AOI22_X1 U22863 ( .A1(n19885), .A2(n19773), .B1(n19884), .B2(n19726), .ZN(
        n19688) );
  OAI211_X1 U22864 ( .C1(n19888), .C2(n19704), .A(n19689), .B(n19688), .ZN(
        P3_U2934) );
  AOI22_X1 U22865 ( .A1(n19890), .A2(n19718), .B1(n19889), .B2(n19700), .ZN(
        n19691) );
  AOI22_X1 U22866 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19701), .B1(
        n19891), .B2(n19773), .ZN(n19690) );
  OAI211_X1 U22867 ( .C1(n19894), .C2(n19704), .A(n19691), .B(n19690), .ZN(
        P3_U2935) );
  AOI22_X1 U22868 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19701), .B1(
        n19895), .B2(n19700), .ZN(n19694) );
  AOI22_X1 U22869 ( .A1(n19897), .A2(n19773), .B1(n19692), .B2(n19726), .ZN(
        n19693) );
  OAI211_X1 U22870 ( .C1(n19695), .C2(n19704), .A(n19694), .B(n19693), .ZN(
        P3_U2936) );
  AOI22_X1 U22871 ( .A1(n19821), .A2(n19718), .B1(n19901), .B2(n19700), .ZN(
        n19697) );
  AOI22_X1 U22872 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19701), .B1(
        n19903), .B2(n19773), .ZN(n19696) );
  OAI211_X1 U22873 ( .C1(n19824), .C2(n19704), .A(n19697), .B(n19696), .ZN(
        P3_U2937) );
  AOI22_X1 U22874 ( .A1(n19825), .A2(n19718), .B1(n19909), .B2(n19700), .ZN(
        n19699) );
  AOI22_X1 U22875 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19701), .B1(
        n19910), .B2(n19773), .ZN(n19698) );
  OAI211_X1 U22876 ( .C1(n19828), .C2(n19704), .A(n19699), .B(n19698), .ZN(
        P3_U2938) );
  AOI22_X1 U22877 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19701), .B1(
        n19916), .B2(n19700), .ZN(n19703) );
  AOI22_X1 U22878 ( .A1(n19917), .A2(n19718), .B1(n19919), .B2(n19773), .ZN(
        n19702) );
  OAI211_X1 U22879 ( .C1(n19925), .C2(n19704), .A(n19703), .B(n19702), .ZN(
        P3_U2939) );
  NAND2_X1 U22880 ( .A1(n19779), .A2(n19705), .ZN(n19797) );
  INV_X1 U22881 ( .A(n19779), .ZN(n19756) );
  NOR2_X1 U22882 ( .A1(n19756), .A2(n19706), .ZN(n19727) );
  AOI22_X1 U22883 ( .A1(n19866), .A2(n19727), .B1(n19867), .B2(n19750), .ZN(
        n19711) );
  NOR2_X1 U22884 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19707), .ZN(
        n19709) );
  NOR2_X1 U22885 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19756), .ZN(
        n19708) );
  AOI22_X1 U22886 ( .A1(n19871), .A2(n19709), .B1(n19868), .B2(n19708), .ZN(
        n19728) );
  AOI22_X1 U22887 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19728), .B1(
        n19778), .B2(n19726), .ZN(n19710) );
  OAI211_X1 U22888 ( .C1(n19786), .C2(n19797), .A(n19711), .B(n19710), .ZN(
        P3_U2940) );
  AOI22_X1 U22889 ( .A1(n19878), .A2(n19718), .B1(n19876), .B2(n19727), .ZN(
        n19713) );
  AOI22_X1 U22890 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19728), .B1(
        n19877), .B2(n19750), .ZN(n19712) );
  OAI211_X1 U22891 ( .C1(n19881), .C2(n19797), .A(n19713), .B(n19712), .ZN(
        P3_U2941) );
  AOI22_X1 U22892 ( .A1(n19812), .A2(n19718), .B1(n19883), .B2(n19727), .ZN(
        n19715) );
  AOI22_X1 U22893 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19728), .B1(
        n19884), .B2(n19750), .ZN(n19714) );
  OAI211_X1 U22894 ( .C1(n19815), .C2(n19797), .A(n19715), .B(n19714), .ZN(
        P3_U2942) );
  AOI22_X1 U22895 ( .A1(n19890), .A2(n19750), .B1(n19889), .B2(n19727), .ZN(
        n19717) );
  AOI22_X1 U22896 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19728), .B1(
        n19846), .B2(n19726), .ZN(n19716) );
  OAI211_X1 U22897 ( .C1(n19849), .C2(n19797), .A(n19717), .B(n19716), .ZN(
        P3_U2943) );
  AOI22_X1 U22898 ( .A1(n19896), .A2(n19718), .B1(n19895), .B2(n19727), .ZN(
        n19720) );
  INV_X1 U22899 ( .A(n19797), .ZN(n19802) );
  AOI22_X1 U22900 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19728), .B1(
        n19897), .B2(n19802), .ZN(n19719) );
  OAI211_X1 U22901 ( .C1(n19900), .C2(n19749), .A(n19720), .B(n19719), .ZN(
        P3_U2944) );
  AOI22_X1 U22902 ( .A1(n19821), .A2(n19750), .B1(n19901), .B2(n19727), .ZN(
        n19722) );
  AOI22_X1 U22903 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19728), .B1(
        n19903), .B2(n19802), .ZN(n19721) );
  OAI211_X1 U22904 ( .C1(n19824), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P3_U2945) );
  AOI22_X1 U22905 ( .A1(n19909), .A2(n19727), .B1(n19908), .B2(n19726), .ZN(
        n19725) );
  AOI22_X1 U22906 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19728), .B1(
        n19910), .B2(n19802), .ZN(n19724) );
  OAI211_X1 U22907 ( .C1(n19913), .C2(n19749), .A(n19725), .B(n19724), .ZN(
        P3_U2946) );
  AOI22_X1 U22908 ( .A1(n19916), .A2(n19727), .B1(n19858), .B2(n19726), .ZN(
        n19730) );
  AOI22_X1 U22909 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19728), .B1(
        n19919), .B2(n19802), .ZN(n19729) );
  OAI211_X1 U22910 ( .C1(n19864), .C2(n19749), .A(n19730), .B(n19729), .ZN(
        P3_U2947) );
  NAND2_X1 U22911 ( .A1(n19779), .A2(n19731), .ZN(n19833) );
  AOI21_X1 U22912 ( .B1(n19797), .B2(n19833), .A(n19978), .ZN(n19751) );
  AOI22_X1 U22913 ( .A1(n19866), .A2(n19751), .B1(n19867), .B2(n19773), .ZN(
        n19736) );
  INV_X1 U22914 ( .A(n19833), .ZN(n19818) );
  OAI211_X1 U22915 ( .C1(n19733), .C2(n19732), .A(n19797), .B(n19833), .ZN(
        n19734) );
  OAI211_X1 U22916 ( .C1(n19818), .C2(n20070), .A(n19783), .B(n19734), .ZN(
        n19752) );
  AOI22_X1 U22917 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19752), .B1(
        n19872), .B2(n19818), .ZN(n19735) );
  OAI211_X1 U22918 ( .C1(n19875), .C2(n19749), .A(n19736), .B(n19735), .ZN(
        P3_U2948) );
  AOI22_X1 U22919 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19752), .B1(
        n19876), .B2(n19751), .ZN(n19738) );
  AOI22_X1 U22920 ( .A1(n19808), .A2(n19818), .B1(n19878), .B2(n19750), .ZN(
        n19737) );
  OAI211_X1 U22921 ( .C1(n19811), .C2(n19772), .A(n19738), .B(n19737), .ZN(
        P3_U2949) );
  AOI22_X1 U22922 ( .A1(n19884), .A2(n19773), .B1(n19883), .B2(n19751), .ZN(
        n19740) );
  AOI22_X1 U22923 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19752), .B1(
        n19885), .B2(n19818), .ZN(n19739) );
  OAI211_X1 U22924 ( .C1(n19888), .C2(n19749), .A(n19740), .B(n19739), .ZN(
        P3_U2950) );
  AOI22_X1 U22925 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19752), .B1(
        n19889), .B2(n19751), .ZN(n19742) );
  AOI22_X1 U22926 ( .A1(n19891), .A2(n19818), .B1(n19890), .B2(n19773), .ZN(
        n19741) );
  OAI211_X1 U22927 ( .C1(n19894), .C2(n19749), .A(n19742), .B(n19741), .ZN(
        P3_U2951) );
  AOI22_X1 U22928 ( .A1(n19896), .A2(n19750), .B1(n19895), .B2(n19751), .ZN(
        n19744) );
  AOI22_X1 U22929 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19752), .B1(
        n19897), .B2(n19818), .ZN(n19743) );
  OAI211_X1 U22930 ( .C1(n19900), .C2(n19772), .A(n19744), .B(n19743), .ZN(
        P3_U2952) );
  AOI22_X1 U22931 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19752), .B1(
        n19901), .B2(n19751), .ZN(n19746) );
  AOI22_X1 U22932 ( .A1(n19903), .A2(n19818), .B1(n19821), .B2(n19773), .ZN(
        n19745) );
  OAI211_X1 U22933 ( .C1(n19824), .C2(n19749), .A(n19746), .B(n19745), .ZN(
        P3_U2953) );
  AOI22_X1 U22934 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19752), .B1(
        n19909), .B2(n19751), .ZN(n19748) );
  AOI22_X1 U22935 ( .A1(n19825), .A2(n19773), .B1(n19910), .B2(n19818), .ZN(
        n19747) );
  OAI211_X1 U22936 ( .C1(n19828), .C2(n19749), .A(n19748), .B(n19747), .ZN(
        P3_U2954) );
  AOI22_X1 U22937 ( .A1(n19916), .A2(n19751), .B1(n19858), .B2(n19750), .ZN(
        n19754) );
  AOI22_X1 U22938 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19752), .B1(
        n19919), .B2(n19818), .ZN(n19753) );
  OAI211_X1 U22939 ( .C1(n19864), .C2(n19772), .A(n19754), .B(n19753), .ZN(
        P3_U2955) );
  NOR2_X1 U22940 ( .A1(n19755), .A2(n19756), .ZN(n19805) );
  AND2_X1 U22941 ( .A1(n19865), .A2(n19805), .ZN(n19774) );
  AOI22_X1 U22942 ( .A1(n19866), .A2(n19774), .B1(n19867), .B2(n19802), .ZN(
        n19759) );
  OAI211_X1 U22943 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19871), .A(
        n19868), .B(n19779), .ZN(n19775) );
  NOR2_X2 U22944 ( .A1(n19757), .A2(n19756), .ZN(n19857) );
  AOI22_X1 U22945 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19775), .B1(
        n19872), .B2(n19857), .ZN(n19758) );
  OAI211_X1 U22946 ( .C1(n19875), .C2(n19772), .A(n19759), .B(n19758), .ZN(
        P3_U2956) );
  INV_X1 U22947 ( .A(n19857), .ZN(n19845) );
  AOI22_X1 U22948 ( .A1(n19877), .A2(n19802), .B1(n19876), .B2(n19774), .ZN(
        n19761) );
  AOI22_X1 U22949 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19775), .B1(
        n19878), .B2(n19773), .ZN(n19760) );
  OAI211_X1 U22950 ( .C1(n19881), .C2(n19845), .A(n19761), .B(n19760), .ZN(
        P3_U2957) );
  AOI22_X1 U22951 ( .A1(n19884), .A2(n19802), .B1(n19883), .B2(n19774), .ZN(
        n19763) );
  AOI22_X1 U22952 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19775), .B1(
        n19885), .B2(n19857), .ZN(n19762) );
  OAI211_X1 U22953 ( .C1(n19888), .C2(n19772), .A(n19763), .B(n19762), .ZN(
        P3_U2958) );
  AOI22_X1 U22954 ( .A1(n19846), .A2(n19773), .B1(n19889), .B2(n19774), .ZN(
        n19765) );
  AOI22_X1 U22955 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19775), .B1(
        n19890), .B2(n19802), .ZN(n19764) );
  OAI211_X1 U22956 ( .C1(n19849), .C2(n19845), .A(n19765), .B(n19764), .ZN(
        P3_U2959) );
  AOI22_X1 U22957 ( .A1(n19896), .A2(n19773), .B1(n19895), .B2(n19774), .ZN(
        n19767) );
  AOI22_X1 U22958 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19775), .B1(
        n19897), .B2(n19857), .ZN(n19766) );
  OAI211_X1 U22959 ( .C1(n19900), .C2(n19797), .A(n19767), .B(n19766), .ZN(
        P3_U2960) );
  AOI22_X1 U22960 ( .A1(n19902), .A2(n19773), .B1(n19901), .B2(n19774), .ZN(
        n19769) );
  AOI22_X1 U22961 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19775), .B1(
        n19903), .B2(n19857), .ZN(n19768) );
  OAI211_X1 U22962 ( .C1(n19906), .C2(n19797), .A(n19769), .B(n19768), .ZN(
        P3_U2961) );
  AOI22_X1 U22963 ( .A1(n19825), .A2(n19802), .B1(n19909), .B2(n19774), .ZN(
        n19771) );
  AOI22_X1 U22964 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19775), .B1(
        n19910), .B2(n19857), .ZN(n19770) );
  OAI211_X1 U22965 ( .C1(n19828), .C2(n19772), .A(n19771), .B(n19770), .ZN(
        P3_U2962) );
  AOI22_X1 U22966 ( .A1(n19916), .A2(n19774), .B1(n19858), .B2(n19773), .ZN(
        n19777) );
  AOI22_X1 U22967 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19775), .B1(
        n19919), .B2(n19857), .ZN(n19776) );
  OAI211_X1 U22968 ( .C1(n19864), .C2(n19797), .A(n19777), .B(n19776), .ZN(
        P3_U2963) );
  NAND2_X1 U22969 ( .A1(n19870), .A2(n10656), .ZN(n19924) );
  INV_X1 U22970 ( .A(n19924), .ZN(n19907) );
  NOR2_X1 U22971 ( .A1(n19857), .A2(n19907), .ZN(n19834) );
  NOR2_X1 U22972 ( .A1(n19978), .A2(n19834), .ZN(n19800) );
  AOI22_X1 U22973 ( .A1(n19778), .A2(n19802), .B1(n19866), .B2(n19800), .ZN(
        n19785) );
  NAND2_X1 U22974 ( .A1(n19837), .A2(n19779), .ZN(n19780) );
  OAI21_X1 U22975 ( .B1(n19781), .B2(n19780), .A(n19834), .ZN(n19782) );
  OAI211_X1 U22976 ( .C1(n19907), .C2(n20070), .A(n19783), .B(n19782), .ZN(
        n19801) );
  AOI22_X1 U22977 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19801), .B1(
        n19867), .B2(n19818), .ZN(n19784) );
  OAI211_X1 U22978 ( .C1(n19786), .C2(n19924), .A(n19785), .B(n19784), .ZN(
        P3_U2964) );
  AOI22_X1 U22979 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19801), .B1(
        n19876), .B2(n19800), .ZN(n19788) );
  AOI22_X1 U22980 ( .A1(n19808), .A2(n19907), .B1(n19878), .B2(n19802), .ZN(
        n19787) );
  OAI211_X1 U22981 ( .C1(n19811), .C2(n19833), .A(n19788), .B(n19787), .ZN(
        P3_U2965) );
  AOI22_X1 U22982 ( .A1(n19812), .A2(n19802), .B1(n19883), .B2(n19800), .ZN(
        n19790) );
  AOI22_X1 U22983 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19801), .B1(
        n19884), .B2(n19818), .ZN(n19789) );
  OAI211_X1 U22984 ( .C1(n19815), .C2(n19924), .A(n19790), .B(n19789), .ZN(
        P3_U2966) );
  AOI22_X1 U22985 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19801), .B1(
        n19889), .B2(n19800), .ZN(n19792) );
  AOI22_X1 U22986 ( .A1(n19891), .A2(n19907), .B1(n19890), .B2(n19818), .ZN(
        n19791) );
  OAI211_X1 U22987 ( .C1(n19894), .C2(n19797), .A(n19792), .B(n19791), .ZN(
        P3_U2967) );
  AOI22_X1 U22988 ( .A1(n19896), .A2(n19802), .B1(n19895), .B2(n19800), .ZN(
        n19794) );
  AOI22_X1 U22989 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19801), .B1(
        n19897), .B2(n19907), .ZN(n19793) );
  OAI211_X1 U22990 ( .C1(n19900), .C2(n19833), .A(n19794), .B(n19793), .ZN(
        P3_U2968) );
  AOI22_X1 U22991 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19801), .B1(
        n19901), .B2(n19800), .ZN(n19796) );
  AOI22_X1 U22992 ( .A1(n19903), .A2(n19907), .B1(n19821), .B2(n19818), .ZN(
        n19795) );
  OAI211_X1 U22993 ( .C1(n19824), .C2(n19797), .A(n19796), .B(n19795), .ZN(
        P3_U2969) );
  AOI22_X1 U22994 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19801), .B1(
        n19909), .B2(n19800), .ZN(n19799) );
  AOI22_X1 U22995 ( .A1(n19910), .A2(n19907), .B1(n19908), .B2(n19802), .ZN(
        n19798) );
  OAI211_X1 U22996 ( .C1(n19913), .C2(n19833), .A(n19799), .B(n19798), .ZN(
        P3_U2970) );
  AOI22_X1 U22997 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19801), .B1(
        n19916), .B2(n19800), .ZN(n19804) );
  AOI22_X1 U22998 ( .A1(n19919), .A2(n19907), .B1(n19858), .B2(n19802), .ZN(
        n19803) );
  OAI211_X1 U22999 ( .C1(n19864), .C2(n19833), .A(n19804), .B(n19803), .ZN(
        P3_U2971) );
  AND2_X1 U23000 ( .A1(n19865), .A2(n19870), .ZN(n19829) );
  AOI22_X1 U23001 ( .A1(n19866), .A2(n19829), .B1(n19867), .B2(n19857), .ZN(
        n19807) );
  AOI22_X1 U23002 ( .A1(n19871), .A2(n19805), .B1(n19870), .B2(n19868), .ZN(
        n19830) );
  AOI22_X1 U23003 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19872), .ZN(n19806) );
  OAI211_X1 U23004 ( .C1(n19875), .C2(n19833), .A(n19807), .B(n19806), .ZN(
        P3_U2972) );
  AOI22_X1 U23005 ( .A1(n19878), .A2(n19818), .B1(n19876), .B2(n19829), .ZN(
        n19810) );
  AOI22_X1 U23006 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19808), .ZN(n19809) );
  OAI211_X1 U23007 ( .C1(n19811), .C2(n19845), .A(n19810), .B(n19809), .ZN(
        P3_U2973) );
  AOI22_X1 U23008 ( .A1(n19812), .A2(n19818), .B1(n19883), .B2(n19829), .ZN(
        n19814) );
  AOI22_X1 U23009 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19830), .B1(
        n19884), .B2(n19857), .ZN(n19813) );
  OAI211_X1 U23010 ( .C1(n19914), .C2(n19815), .A(n19814), .B(n19813), .ZN(
        P3_U2974) );
  AOI22_X1 U23011 ( .A1(n19890), .A2(n19857), .B1(n19889), .B2(n19829), .ZN(
        n19817) );
  AOI22_X1 U23012 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19891), .ZN(n19816) );
  OAI211_X1 U23013 ( .C1(n19894), .C2(n19833), .A(n19817), .B(n19816), .ZN(
        P3_U2975) );
  AOI22_X1 U23014 ( .A1(n19896), .A2(n19818), .B1(n19895), .B2(n19829), .ZN(
        n19820) );
  AOI22_X1 U23015 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19897), .ZN(n19819) );
  OAI211_X1 U23016 ( .C1(n19900), .C2(n19845), .A(n19820), .B(n19819), .ZN(
        P3_U2976) );
  AOI22_X1 U23017 ( .A1(n19821), .A2(n19857), .B1(n19901), .B2(n19829), .ZN(
        n19823) );
  AOI22_X1 U23018 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19903), .ZN(n19822) );
  OAI211_X1 U23019 ( .C1(n19824), .C2(n19833), .A(n19823), .B(n19822), .ZN(
        P3_U2977) );
  AOI22_X1 U23020 ( .A1(n19825), .A2(n19857), .B1(n19909), .B2(n19829), .ZN(
        n19827) );
  AOI22_X1 U23021 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19910), .ZN(n19826) );
  OAI211_X1 U23022 ( .C1(n19828), .C2(n19833), .A(n19827), .B(n19826), .ZN(
        P3_U2978) );
  AOI22_X1 U23023 ( .A1(n19917), .A2(n19857), .B1(n19916), .B2(n19829), .ZN(
        n19832) );
  AOI22_X1 U23024 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19830), .B1(
        n19918), .B2(n19919), .ZN(n19831) );
  OAI211_X1 U23025 ( .C1(n19925), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        P3_U2979) );
  AND2_X1 U23026 ( .A1(n19865), .A2(n19838), .ZN(n19859) );
  AOI22_X1 U23027 ( .A1(n19866), .A2(n19859), .B1(n19867), .B2(n19907), .ZN(
        n19840) );
  INV_X1 U23028 ( .A(n19834), .ZN(n19836) );
  OAI221_X1 U23029 ( .B1(n19838), .B2(n19837), .C1(n19838), .C2(n19836), .A(
        n19835), .ZN(n19861) );
  AOI22_X1 U23030 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19861), .B1(
        n19872), .B2(n19860), .ZN(n19839) );
  OAI211_X1 U23031 ( .C1(n19875), .C2(n19845), .A(n19840), .B(n19839), .ZN(
        P3_U2980) );
  AOI22_X1 U23032 ( .A1(n19877), .A2(n19907), .B1(n19876), .B2(n19859), .ZN(
        n19842) );
  AOI22_X1 U23033 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19861), .B1(
        n19878), .B2(n19857), .ZN(n19841) );
  OAI211_X1 U23034 ( .C1(n19850), .C2(n19881), .A(n19842), .B(n19841), .ZN(
        P3_U2981) );
  AOI22_X1 U23035 ( .A1(n19884), .A2(n19907), .B1(n19883), .B2(n19859), .ZN(
        n19844) );
  AOI22_X1 U23036 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19885), .ZN(n19843) );
  OAI211_X1 U23037 ( .C1(n19888), .C2(n19845), .A(n19844), .B(n19843), .ZN(
        P3_U2982) );
  AOI22_X1 U23038 ( .A1(n19846), .A2(n19857), .B1(n19889), .B2(n19859), .ZN(
        n19848) );
  AOI22_X1 U23039 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19861), .B1(
        n19890), .B2(n19907), .ZN(n19847) );
  OAI211_X1 U23040 ( .C1(n19850), .C2(n19849), .A(n19848), .B(n19847), .ZN(
        P3_U2983) );
  AOI22_X1 U23041 ( .A1(n19896), .A2(n19857), .B1(n19895), .B2(n19859), .ZN(
        n19852) );
  AOI22_X1 U23042 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19897), .ZN(n19851) );
  OAI211_X1 U23043 ( .C1(n19900), .C2(n19924), .A(n19852), .B(n19851), .ZN(
        P3_U2984) );
  AOI22_X1 U23044 ( .A1(n19902), .A2(n19857), .B1(n19901), .B2(n19859), .ZN(
        n19854) );
  AOI22_X1 U23045 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19903), .ZN(n19853) );
  OAI211_X1 U23046 ( .C1(n19906), .C2(n19924), .A(n19854), .B(n19853), .ZN(
        P3_U2985) );
  AOI22_X1 U23047 ( .A1(n19909), .A2(n19859), .B1(n19908), .B2(n19857), .ZN(
        n19856) );
  AOI22_X1 U23048 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19910), .ZN(n19855) );
  OAI211_X1 U23049 ( .C1(n19913), .C2(n19924), .A(n19856), .B(n19855), .ZN(
        P3_U2986) );
  AOI22_X1 U23050 ( .A1(n19916), .A2(n19859), .B1(n19858), .B2(n19857), .ZN(
        n19863) );
  AOI22_X1 U23051 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19861), .B1(
        n19860), .B2(n19919), .ZN(n19862) );
  OAI211_X1 U23052 ( .C1(n19864), .C2(n19924), .A(n19863), .B(n19862), .ZN(
        P3_U2987) );
  AND2_X1 U23053 ( .A1(n19865), .A2(n19869), .ZN(n19915) );
  AOI22_X1 U23054 ( .A1(n19918), .A2(n19867), .B1(n19866), .B2(n19915), .ZN(
        n19874) );
  AOI22_X1 U23055 ( .A1(n19871), .A2(n19870), .B1(n19869), .B2(n19868), .ZN(
        n19921) );
  AOI22_X1 U23056 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19872), .ZN(n19873) );
  OAI211_X1 U23057 ( .C1(n19875), .C2(n19924), .A(n19874), .B(n19873), .ZN(
        P3_U2988) );
  AOI22_X1 U23058 ( .A1(n19918), .A2(n19877), .B1(n19876), .B2(n19915), .ZN(
        n19880) );
  AOI22_X1 U23059 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19921), .B1(
        n19878), .B2(n19907), .ZN(n19879) );
  OAI211_X1 U23060 ( .C1(n19882), .C2(n19881), .A(n19880), .B(n19879), .ZN(
        P3_U2989) );
  AOI22_X1 U23061 ( .A1(n19918), .A2(n19884), .B1(n19883), .B2(n19915), .ZN(
        n19887) );
  AOI22_X1 U23062 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19885), .ZN(n19886) );
  OAI211_X1 U23063 ( .C1(n19888), .C2(n19924), .A(n19887), .B(n19886), .ZN(
        P3_U2990) );
  AOI22_X1 U23064 ( .A1(n19918), .A2(n19890), .B1(n19889), .B2(n19915), .ZN(
        n19893) );
  AOI22_X1 U23065 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19891), .ZN(n19892) );
  OAI211_X1 U23066 ( .C1(n19894), .C2(n19924), .A(n19893), .B(n19892), .ZN(
        P3_U2991) );
  AOI22_X1 U23067 ( .A1(n19896), .A2(n19907), .B1(n19895), .B2(n19915), .ZN(
        n19899) );
  AOI22_X1 U23068 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19897), .ZN(n19898) );
  OAI211_X1 U23069 ( .C1(n19914), .C2(n19900), .A(n19899), .B(n19898), .ZN(
        P3_U2992) );
  AOI22_X1 U23070 ( .A1(n19902), .A2(n19907), .B1(n19901), .B2(n19915), .ZN(
        n19905) );
  AOI22_X1 U23071 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19903), .ZN(n19904) );
  OAI211_X1 U23072 ( .C1(n19914), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P3_U2993) );
  AOI22_X1 U23073 ( .A1(n19909), .A2(n19915), .B1(n19908), .B2(n19907), .ZN(
        n19912) );
  AOI22_X1 U23074 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19910), .ZN(n19911) );
  OAI211_X1 U23075 ( .C1(n19914), .C2(n19913), .A(n19912), .B(n19911), .ZN(
        P3_U2994) );
  AOI22_X1 U23076 ( .A1(n19918), .A2(n19917), .B1(n19916), .B2(n19915), .ZN(
        n19923) );
  AOI22_X1 U23077 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19921), .B1(
        n19920), .B2(n19919), .ZN(n19922) );
  OAI211_X1 U23078 ( .C1(n19925), .C2(n19924), .A(n19923), .B(n19922), .ZN(
        P3_U2995) );
  AOI21_X1 U23079 ( .B1(n19960), .B2(n19927), .A(n19926), .ZN(n19929) );
  OAI22_X1 U23080 ( .A1(n19929), .A2(n19928), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19960), .ZN(n19944) );
  NOR2_X1 U23081 ( .A1(n19933), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19931) );
  OAI21_X1 U23082 ( .B1(n19931), .B2(n19930), .A(n19960), .ZN(n19935) );
  AOI22_X1 U23083 ( .A1(n19935), .A2(n19934), .B1(n19933), .B2(n19932), .ZN(
        n19939) );
  MUX2_X1 U23084 ( .A(n19937), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19936), .Z(n19941) );
  AOI222_X1 U23085 ( .A1(n19939), .A2(n19941), .B1(n19939), .B2(n19938), .C1(
        n19941), .C2(n19938), .ZN(n19940) );
  AOI211_X1 U23086 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n19944), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n19940), .ZN(n19964) );
  INV_X1 U23087 ( .A(n19941), .ZN(n19946) );
  NAND2_X1 U23088 ( .A1(n19943), .A2(n19942), .ZN(n19945) );
  AOI21_X1 U23089 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(n19963) );
  INV_X1 U23090 ( .A(n19947), .ZN(n19954) );
  NOR2_X1 U23091 ( .A1(n19949), .A2(n19948), .ZN(n19951) );
  OAI222_X1 U23092 ( .A1(n19955), .A2(n19954), .B1(n19953), .B2(n19952), .C1(
        n19951), .C2(n19950), .ZN(n20082) );
  AOI221_X1 U23093 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n19957), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n19957), .A(n19956), .ZN(n19958) );
  OAI211_X1 U23094 ( .C1(n19961), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        n19962) );
  NOR4_X1 U23095 ( .A1(n19964), .A2(n19963), .A3(n20082), .A4(n19962), .ZN(
        n19977) );
  NOR2_X1 U23096 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20095) );
  AOI22_X1 U23097 ( .A1(n19965), .A2(n20095), .B1(n20090), .B2(n20084), .ZN(
        n19966) );
  INV_X1 U23098 ( .A(n19966), .ZN(n19972) );
  INV_X1 U23099 ( .A(n19967), .ZN(n19969) );
  OAI211_X1 U23100 ( .C1(n19969), .C2(n19968), .A(n20087), .B(n19977), .ZN(
        n20069) );
  OAI21_X1 U23101 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n20083), .A(n20069), 
        .ZN(n19979) );
  NOR2_X1 U23102 ( .A1(n19970), .A2(n19979), .ZN(n19971) );
  MUX2_X1 U23103 ( .A(n19972), .B(n19971), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19975) );
  INV_X1 U23104 ( .A(n19973), .ZN(n19974) );
  OAI211_X1 U23105 ( .C1(n19977), .C2(n19976), .A(n19975), .B(n19974), .ZN(
        P3_U2996) );
  NAND2_X1 U23106 ( .A1(n20090), .A2(n20084), .ZN(n19982) );
  NAND4_X1 U23107 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n20090), .A4(n20102), .ZN(n19983) );
  OR3_X1 U23108 ( .A1(n19980), .A2(n19979), .A3(n19978), .ZN(n19981) );
  NAND4_X1 U23109 ( .A1(n13366), .A2(n19982), .A3(n19983), .A4(n19981), .ZN(
        P3_U2997) );
  INV_X1 U23110 ( .A(n20095), .ZN(n19985) );
  AND4_X1 U23111 ( .A1(n19985), .A2(n19984), .A3(n19983), .A4(n20068), .ZN(
        P3_U2998) );
  AND2_X1 U23112 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n20065), .ZN(
        P3_U2999) );
  AND2_X1 U23113 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n20065), .ZN(
        P3_U3000) );
  AND2_X1 U23114 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n20065), .ZN(
        P3_U3001) );
  AND2_X1 U23115 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n20065), .ZN(
        P3_U3002) );
  AND2_X1 U23116 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n20065), .ZN(
        P3_U3003) );
  AND2_X1 U23117 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n20065), .ZN(
        P3_U3004) );
  AND2_X1 U23118 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n20065), .ZN(
        P3_U3005) );
  NOR2_X1 U23119 ( .A1(n21455), .A2(n20067), .ZN(P3_U3006) );
  AND2_X1 U23120 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n20065), .ZN(
        P3_U3007) );
  AND2_X1 U23121 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n20065), .ZN(
        P3_U3008) );
  INV_X1 U23122 ( .A(P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21694) );
  NOR2_X1 U23123 ( .A1(n21694), .A2(n20067), .ZN(P3_U3009) );
  AND2_X1 U23124 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n20065), .ZN(
        P3_U3010) );
  AND2_X1 U23125 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n20065), .ZN(
        P3_U3011) );
  AND2_X1 U23126 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n20065), .ZN(
        P3_U3012) );
  AND2_X1 U23127 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n20065), .ZN(
        P3_U3013) );
  AND2_X1 U23128 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n20065), .ZN(
        P3_U3014) );
  AND2_X1 U23129 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n20065), .ZN(
        P3_U3015) );
  AND2_X1 U23130 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n20065), .ZN(
        P3_U3016) );
  AND2_X1 U23131 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n20065), .ZN(
        P3_U3017) );
  AND2_X1 U23132 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n20065), .ZN(
        P3_U3018) );
  AND2_X1 U23133 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n20065), .ZN(
        P3_U3019) );
  NOR2_X1 U23134 ( .A1(n21533), .A2(n20067), .ZN(P3_U3020) );
  AND2_X1 U23135 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n20065), .ZN(P3_U3021) );
  AND2_X1 U23136 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n20065), .ZN(P3_U3022) );
  AND2_X1 U23137 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n20065), .ZN(P3_U3023) );
  AND2_X1 U23138 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n20065), .ZN(P3_U3024) );
  AND2_X1 U23139 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n20065), .ZN(P3_U3025) );
  AND2_X1 U23140 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n20065), .ZN(P3_U3026) );
  AND2_X1 U23141 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n20065), .ZN(P3_U3027) );
  AND2_X1 U23142 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n20065), .ZN(P3_U3028) );
  OAI21_X1 U23143 ( .B1(n21355), .B2(n19986), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19987) );
  INV_X1 U23144 ( .A(n19987), .ZN(n19990) );
  NAND2_X1 U23145 ( .A1(n20090), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19997) );
  INV_X1 U23146 ( .A(n19997), .ZN(n19995) );
  OAI21_X1 U23147 ( .B1(n19995), .B2(n20001), .A(n20003), .ZN(n19989) );
  NAND3_X1 U23148 ( .A1(NA), .A2(n20001), .A3(n19988), .ZN(n19996) );
  OAI211_X1 U23149 ( .C1(n20101), .C2(n19990), .A(n19989), .B(n19996), .ZN(
        P3_U3029) );
  NOR2_X1 U23150 ( .A1(n20003), .A2(n21355), .ZN(n19999) );
  INV_X1 U23151 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20097) );
  NOR3_X1 U23152 ( .A1(n19999), .A2(n20097), .A3(n20001), .ZN(n19991) );
  NOR2_X1 U23153 ( .A1(n19991), .A2(n19995), .ZN(n19993) );
  OAI211_X1 U23154 ( .C1(n21355), .C2(n19994), .A(n19993), .B(n19992), .ZN(
        P3_U3030) );
  AOI21_X1 U23155 ( .B1(n20001), .B2(n19996), .A(n19995), .ZN(n20002) );
  OAI22_X1 U23156 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19997), .ZN(n19998) );
  OAI22_X1 U23157 ( .A1(n19999), .A2(n19998), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n20000) );
  OAI22_X1 U23158 ( .A1(n20002), .A2(n20003), .B1(n20001), .B2(n20000), .ZN(
        P3_U3031) );
  NAND2_X2 U23159 ( .A1(n20101), .A2(n20003), .ZN(n20058) );
  OAI222_X1 U23160 ( .A1(n20058), .A2(n20006), .B1(n20004), .B2(n20101), .C1(
        n13863), .C2(n20062), .ZN(P3_U3032) );
  OAI222_X1 U23161 ( .A1(n20006), .A2(n20062), .B1(n20005), .B2(n20101), .C1(
        n20007), .C2(n20058), .ZN(P3_U3033) );
  OAI222_X1 U23162 ( .A1(n20058), .A2(n20008), .B1(n21496), .B2(n20101), .C1(
        n20007), .C2(n20062), .ZN(P3_U3034) );
  OAI222_X1 U23163 ( .A1(n20058), .A2(n21460), .B1(n20009), .B2(n20101), .C1(
        n20008), .C2(n20062), .ZN(P3_U3035) );
  OAI222_X1 U23164 ( .A1(n21460), .A2(n20062), .B1(n20010), .B2(n20101), .C1(
        n20011), .C2(n20058), .ZN(P3_U3036) );
  OAI222_X1 U23165 ( .A1(n20058), .A2(n20013), .B1(n20012), .B2(n20101), .C1(
        n20011), .C2(n20062), .ZN(P3_U3037) );
  INV_X1 U23166 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20016) );
  OAI222_X1 U23167 ( .A1(n20058), .A2(n20016), .B1(n20014), .B2(n20101), .C1(
        n20013), .C2(n20062), .ZN(P3_U3038) );
  OAI222_X1 U23168 ( .A1(n20016), .A2(n20062), .B1(n20015), .B2(n20101), .C1(
        n20017), .C2(n20058), .ZN(P3_U3039) );
  OAI222_X1 U23169 ( .A1(n20058), .A2(n20018), .B1(n21452), .B2(n20101), .C1(
        n20017), .C2(n20062), .ZN(P3_U3040) );
  OAI222_X1 U23170 ( .A1(n20058), .A2(n20020), .B1(n20019), .B2(n20101), .C1(
        n20018), .C2(n20062), .ZN(P3_U3041) );
  INV_X1 U23171 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20022) );
  OAI222_X1 U23172 ( .A1(n20058), .A2(n20022), .B1(n20021), .B2(n20101), .C1(
        n20020), .C2(n20062), .ZN(P3_U3042) );
  OAI222_X1 U23173 ( .A1(n20058), .A2(n20024), .B1(n20023), .B2(n20101), .C1(
        n20022), .C2(n20062), .ZN(P3_U3043) );
  OAI222_X1 U23174 ( .A1(n20058), .A2(n20027), .B1(n20025), .B2(n20101), .C1(
        n20024), .C2(n20062), .ZN(P3_U3044) );
  OAI222_X1 U23175 ( .A1(n20027), .A2(n20062), .B1(n20026), .B2(n20101), .C1(
        n20028), .C2(n20058), .ZN(P3_U3045) );
  OAI222_X1 U23176 ( .A1(n20058), .A2(n20030), .B1(n20029), .B2(n20101), .C1(
        n20028), .C2(n20062), .ZN(P3_U3046) );
  OAI222_X1 U23177 ( .A1(n20058), .A2(n20033), .B1(n20031), .B2(n20101), .C1(
        n20030), .C2(n20062), .ZN(P3_U3047) );
  OAI222_X1 U23178 ( .A1(n20033), .A2(n20062), .B1(n20032), .B2(n20101), .C1(
        n20034), .C2(n20058), .ZN(P3_U3048) );
  OAI222_X1 U23179 ( .A1(n20058), .A2(n20036), .B1(n20035), .B2(n20101), .C1(
        n20034), .C2(n20062), .ZN(P3_U3049) );
  OAI222_X1 U23180 ( .A1(n20058), .A2(n20038), .B1(n20037), .B2(n20101), .C1(
        n20036), .C2(n20062), .ZN(P3_U3050) );
  OAI222_X1 U23181 ( .A1(n20058), .A2(n20040), .B1(n20039), .B2(n20101), .C1(
        n20038), .C2(n20062), .ZN(P3_U3051) );
  INV_X1 U23182 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U23183 ( .A1(n20058), .A2(n20042), .B1(n20041), .B2(n20101), .C1(
        n20040), .C2(n20062), .ZN(P3_U3052) );
  OAI222_X1 U23184 ( .A1(n20058), .A2(n20044), .B1(n20043), .B2(n20101), .C1(
        n20042), .C2(n20062), .ZN(P3_U3053) );
  OAI222_X1 U23185 ( .A1(n20058), .A2(n20046), .B1(n20045), .B2(n20101), .C1(
        n20044), .C2(n20062), .ZN(P3_U3054) );
  OAI222_X1 U23186 ( .A1(n20058), .A2(n20048), .B1(n20047), .B2(n20101), .C1(
        n20046), .C2(n20062), .ZN(P3_U3055) );
  OAI222_X1 U23187 ( .A1(n20058), .A2(n20050), .B1(n20049), .B2(n20101), .C1(
        n20048), .C2(n20062), .ZN(P3_U3056) );
  OAI222_X1 U23188 ( .A1(n20058), .A2(n20052), .B1(n20051), .B2(n20101), .C1(
        n20050), .C2(n20062), .ZN(P3_U3057) );
  INV_X1 U23189 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20055) );
  OAI222_X1 U23190 ( .A1(n20058), .A2(n20055), .B1(n20053), .B2(n20101), .C1(
        n20052), .C2(n20062), .ZN(P3_U3058) );
  OAI222_X1 U23191 ( .A1(n20055), .A2(n20062), .B1(n20054), .B2(n20101), .C1(
        n20056), .C2(n20058), .ZN(P3_U3059) );
  OAI222_X1 U23192 ( .A1(n20058), .A2(n20061), .B1(n20057), .B2(n20101), .C1(
        n20056), .C2(n20062), .ZN(P3_U3060) );
  OAI222_X1 U23193 ( .A1(n20062), .A2(n20061), .B1(n20060), .B2(n20101), .C1(
        n20059), .C2(n20058), .ZN(P3_U3061) );
  MUX2_X1 U23194 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n20101), .Z(P3_U3274) );
  MUX2_X1 U23195 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n20101), .Z(P3_U3275) );
  MUX2_X1 U23196 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n20101), .Z(P3_U3276) );
  INV_X1 U23197 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20076) );
  INV_X1 U23198 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n20063) );
  AOI22_X1 U23199 ( .A1(n20101), .A2(n20076), .B1(n20063), .B2(n20099), .ZN(
        P3_U3277) );
  INV_X1 U23200 ( .A(n20066), .ZN(n20064) );
  AOI21_X1 U23201 ( .B1(n20065), .B2(n20072), .A(n20064), .ZN(P3_U3280) );
  OAI21_X1 U23202 ( .B1(n20067), .B2(n20071), .A(n20066), .ZN(P3_U3281) );
  OAI221_X1 U23203 ( .B1(n20070), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n20070), 
        .C2(n20069), .A(n20068), .ZN(P3_U3282) );
  OAI211_X1 U23204 ( .C1(n20072), .C2(n20078), .A(n20071), .B(n20079), .ZN(
        n20075) );
  NOR2_X1 U23205 ( .A1(n20077), .A2(n20078), .ZN(n20073) );
  AOI22_X1 U23206 ( .A1(P3_BYTEENABLE_REG_2__SCAN_IN), .A2(n20077), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n20073), .ZN(n20074) );
  NAND2_X1 U23207 ( .A1(n20075), .A2(n20074), .ZN(P3_U3292) );
  AOI22_X1 U23208 ( .A1(n20079), .A2(n20078), .B1(n20077), .B2(n20076), .ZN(
        P3_U3293) );
  INV_X1 U23209 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20080) );
  AOI22_X1 U23210 ( .A1(n20101), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20080), 
        .B2(n20099), .ZN(P3_U3294) );
  MUX2_X1 U23211 ( .A(P3_MORE_REG_SCAN_IN), .B(n20082), .S(n20081), .Z(
        P3_U3295) );
  AOI21_X1 U23212 ( .B1(n20084), .B2(n20083), .A(n20105), .ZN(n20085) );
  OAI21_X1 U23213 ( .B1(n20087), .B2(n20086), .A(n20085), .ZN(n20098) );
  OAI21_X1 U23214 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20089), .A(n20088), 
        .ZN(n20091) );
  AOI211_X1 U23215 ( .C1(n20106), .C2(n20091), .A(n20090), .B(n20102), .ZN(
        n20093) );
  NOR2_X1 U23216 ( .A1(n20093), .A2(n20092), .ZN(n20094) );
  OAI21_X1 U23217 ( .B1(n20095), .B2(n20094), .A(n20098), .ZN(n20096) );
  OAI21_X1 U23218 ( .B1(n20098), .B2(n20097), .A(n20096), .ZN(P3_U3296) );
  INV_X1 U23219 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n20108) );
  INV_X1 U23220 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n20100) );
  AOI22_X1 U23221 ( .A1(n20101), .A2(n20108), .B1(n20100), .B2(n20099), .ZN(
        P3_U3297) );
  AOI21_X1 U23222 ( .B1(n20103), .B2(n20102), .A(n20105), .ZN(n20109) );
  INV_X1 U23223 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20104) );
  AOI22_X1 U23224 ( .A1(n20106), .A2(n20105), .B1(n20109), .B2(n20104), .ZN(
        P3_U3298) );
  AOI21_X1 U23225 ( .B1(n20109), .B2(n20108), .A(n20107), .ZN(P3_U3299) );
  INV_X1 U23226 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n20110) );
  NAND2_X1 U23227 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20955), .ZN(n20945) );
  NAND2_X1 U23228 ( .A1(n20937), .A2(n20936), .ZN(n20941) );
  OAI21_X1 U23229 ( .B1(n20937), .B2(n20945), .A(n20941), .ZN(n21016) );
  OAI21_X1 U23230 ( .B1(n20937), .B2(n20110), .A(n20935), .ZN(P2_U2815) );
  AOI21_X1 U23231 ( .B1(n20937), .B2(n20955), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n20111) );
  AOI22_X1 U23232 ( .A1(n20999), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n20111), 
        .B2(n21085), .ZN(P2_U2817) );
  OAI21_X1 U23233 ( .B1(n20949), .B2(BS16), .A(n21016), .ZN(n21014) );
  OAI21_X1 U23234 ( .B1(n21016), .B2(n20814), .A(n21014), .ZN(P2_U2818) );
  NOR4_X1 U23235 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20121) );
  NOR4_X1 U23236 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20120) );
  NOR4_X1 U23237 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20112) );
  INV_X1 U23238 ( .A(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21497) );
  INV_X1 U23239 ( .A(P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21623) );
  NAND3_X1 U23240 ( .A1(n20112), .A2(n21497), .A3(n21623), .ZN(n20118) );
  NOR4_X1 U23241 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20116) );
  NOR4_X1 U23242 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n20115) );
  NOR4_X1 U23243 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20114) );
  NOR4_X1 U23244 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20113) );
  NAND4_X1 U23245 ( .A1(n20116), .A2(n20115), .A3(n20114), .A4(n20113), .ZN(
        n20117) );
  AOI211_X1 U23246 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20118), .B(n20117), .ZN(n20119) );
  NAND3_X1 U23247 ( .A1(n20121), .A2(n20120), .A3(n20119), .ZN(n20128) );
  NOR2_X1 U23248 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n20128), .ZN(n20122) );
  INV_X1 U23249 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U23250 ( .A1(n20122), .A2(n20123), .B1(n20128), .B2(n21012), .ZN(
        P2_U2820) );
  OR3_X1 U23251 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20127) );
  INV_X1 U23252 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21632) );
  AOI22_X1 U23253 ( .A1(n20122), .A2(n20127), .B1(n21632), .B2(n20128), .ZN(
        P2_U2821) );
  INV_X1 U23254 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21015) );
  NAND2_X1 U23255 ( .A1(n20122), .A2(n21015), .ZN(n20126) );
  INV_X1 U23256 ( .A(n20128), .ZN(n20129) );
  OAI21_X1 U23257 ( .B1(n20123), .B2(n20957), .A(n20129), .ZN(n20124) );
  OAI21_X1 U23258 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n20129), .A(n20124), 
        .ZN(n20125) );
  OAI221_X1 U23259 ( .B1(n20126), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n20126), .C2(P2_REIP_REG_0__SCAN_IN), .A(n20125), .ZN(P2_U2822) );
  INV_X1 U23260 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21009) );
  OAI221_X1 U23261 ( .B1(n20129), .B2(n21009), .C1(n20128), .C2(n20127), .A(
        n20126), .ZN(P2_U2823) );
  NAND2_X1 U23262 ( .A1(n15144), .A2(n20149), .ZN(n20131) );
  MUX2_X1 U23263 ( .A(n15144), .B(n20131), .S(n20130), .Z(n20133) );
  NAND2_X1 U23264 ( .A1(n20133), .A2(n20132), .ZN(n20145) );
  NAND2_X1 U23265 ( .A1(n20245), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U23266 ( .B1(n20249), .B2(n20983), .A(n20169), .ZN(n20134) );
  INV_X1 U23267 ( .A(n20134), .ZN(n20135) );
  OAI211_X1 U23268 ( .C1(n20258), .C2(n20137), .A(n20136), .B(n20135), .ZN(
        n20138) );
  AOI21_X1 U23269 ( .B1(n20139), .B2(n20246), .A(n20138), .ZN(n20144) );
  OAI22_X1 U23270 ( .A1(n20141), .A2(n20251), .B1(n20140), .B2(n20267), .ZN(
        n20142) );
  INV_X1 U23271 ( .A(n20142), .ZN(n20143) );
  OAI211_X1 U23272 ( .C1(n20933), .C2(n20145), .A(n20144), .B(n20143), .ZN(
        P2_U2836) );
  NAND2_X1 U23273 ( .A1(n20146), .A2(n20148), .ZN(n20147) );
  MUX2_X1 U23274 ( .A(n20148), .B(n20147), .S(n15144), .Z(n20150) );
  NAND2_X1 U23275 ( .A1(n20150), .A2(n20149), .ZN(n20162) );
  OAI21_X1 U23276 ( .B1(n20249), .B2(n20981), .A(n20169), .ZN(n20151) );
  AOI21_X1 U23277 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20255), .A(
        n20151), .ZN(n20153) );
  NAND2_X1 U23278 ( .A1(n20245), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n20152) );
  OAI211_X1 U23279 ( .C1(n20154), .C2(n20260), .A(n20153), .B(n20152), .ZN(
        n20155) );
  INV_X1 U23280 ( .A(n20155), .ZN(n20161) );
  INV_X1 U23281 ( .A(n20156), .ZN(n20159) );
  INV_X1 U23282 ( .A(n20157), .ZN(n20158) );
  AOI22_X1 U23283 ( .A1(n20159), .A2(n20269), .B1(n20158), .B2(n20235), .ZN(
        n20160) );
  OAI211_X1 U23284 ( .C1(n20933), .C2(n20162), .A(n20161), .B(n20160), .ZN(
        P2_U2837) );
  NAND2_X1 U23285 ( .A1(n20163), .A2(n20165), .ZN(n20164) );
  MUX2_X1 U23286 ( .A(n20165), .B(n20164), .S(n15144), .Z(n20168) );
  INV_X1 U23287 ( .A(n20166), .ZN(n20167) );
  NAND2_X1 U23288 ( .A1(n20168), .A2(n20167), .ZN(n20179) );
  OAI21_X1 U23289 ( .B1(n20249), .B2(n20977), .A(n20169), .ZN(n20170) );
  AOI21_X1 U23290 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20255), .A(
        n20170), .ZN(n20171) );
  OAI21_X1 U23291 ( .B1(n20266), .B2(n20172), .A(n20171), .ZN(n20173) );
  AOI21_X1 U23292 ( .B1(n20174), .B2(n20246), .A(n20173), .ZN(n20178) );
  AOI22_X1 U23293 ( .A1(n20176), .A2(n20235), .B1(n20175), .B2(n20269), .ZN(
        n20177) );
  OAI211_X1 U23294 ( .C1(n20933), .C2(n20179), .A(n20178), .B(n20177), .ZN(
        P2_U2839) );
  NOR2_X1 U23295 ( .A1(n20180), .A2(n20182), .ZN(n20181) );
  MUX2_X1 U23296 ( .A(n20182), .B(n20181), .S(n15144), .Z(n20184) );
  NAND2_X1 U23297 ( .A1(n20245), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n20186) );
  AOI21_X1 U23298 ( .B1(n20264), .B2(P2_REIP_REG_14__SCAN_IN), .A(n20263), 
        .ZN(n20185) );
  OAI211_X1 U23299 ( .C1(n20258), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        n20188) );
  AOI21_X1 U23300 ( .B1(n20189), .B2(n20246), .A(n20188), .ZN(n20194) );
  OAI22_X1 U23301 ( .A1(n20191), .A2(n20251), .B1(n20190), .B2(n20267), .ZN(
        n20192) );
  INV_X1 U23302 ( .A(n20192), .ZN(n20193) );
  OAI211_X1 U23303 ( .C1(n20933), .C2(n20195), .A(n20194), .B(n20193), .ZN(
        P2_U2841) );
  NAND2_X1 U23304 ( .A1(n20196), .A2(n10462), .ZN(n20197) );
  MUX2_X1 U23305 ( .A(n10462), .B(n20197), .S(n15144), .Z(n20199) );
  NAND2_X1 U23306 ( .A1(n20199), .A2(n9870), .ZN(n20210) );
  INV_X1 U23307 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n20201) );
  OAI222_X1 U23308 ( .A1(n20258), .A2(n20202), .B1(n20201), .B2(n20266), .C1(
        n20200), .C2(n20260), .ZN(n20203) );
  AOI211_X1 U23309 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n20264), .A(n20263), 
        .B(n20203), .ZN(n20209) );
  INV_X1 U23310 ( .A(n20204), .ZN(n20207) );
  INV_X1 U23311 ( .A(n20205), .ZN(n20206) );
  AOI22_X1 U23312 ( .A1(n20207), .A2(n20269), .B1(n20206), .B2(n20235), .ZN(
        n20208) );
  OAI211_X1 U23313 ( .C1(n20933), .C2(n20210), .A(n20209), .B(n20208), .ZN(
        P2_U2843) );
  INV_X1 U23314 ( .A(n20211), .ZN(n20214) );
  OR2_X1 U23315 ( .A1(n20212), .A2(n20211), .ZN(n20213) );
  MUX2_X1 U23316 ( .A(n20214), .B(n20213), .S(n15144), .Z(n20216) );
  NAND2_X1 U23317 ( .A1(n20216), .A2(n20215), .ZN(n20224) );
  OAI22_X1 U23318 ( .A1(n20217), .A2(n20260), .B1(n20266), .B2(n10371), .ZN(
        n20218) );
  INV_X1 U23319 ( .A(n20218), .ZN(n20219) );
  OAI211_X1 U23320 ( .C1(n20968), .C2(n20249), .A(n20219), .B(n12586), .ZN(
        n20220) );
  AOI21_X1 U23321 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20255), .A(
        n20220), .ZN(n20223) );
  AOI22_X1 U23322 ( .A1(n10444), .A2(n20269), .B1(n20221), .B2(n20235), .ZN(
        n20222) );
  OAI211_X1 U23323 ( .C1(n20933), .C2(n20224), .A(n20223), .B(n20222), .ZN(
        P2_U2845) );
  NAND2_X1 U23324 ( .A1(n20243), .A2(n20226), .ZN(n20225) );
  MUX2_X1 U23325 ( .A(n20226), .B(n20225), .S(n15144), .Z(n20229) );
  INV_X1 U23326 ( .A(n20227), .ZN(n20228) );
  NAND2_X1 U23327 ( .A1(n20229), .A2(n20228), .ZN(n20240) );
  INV_X1 U23328 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20232) );
  OAI222_X1 U23329 ( .A1(n20258), .A2(n20232), .B1(n20231), .B2(n20266), .C1(
        n20230), .C2(n20260), .ZN(n20233) );
  AOI211_X1 U23330 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n20264), .A(n20263), .B(
        n20233), .ZN(n20239) );
  INV_X1 U23331 ( .A(n20234), .ZN(n20236) );
  AOI22_X1 U23332 ( .A1(n20237), .A2(n20269), .B1(n20236), .B2(n20235), .ZN(
        n20238) );
  OAI211_X1 U23333 ( .C1(n20933), .C2(n20240), .A(n20239), .B(n20238), .ZN(
        P2_U2847) );
  NAND2_X1 U23334 ( .A1(n20241), .A2(n9774), .ZN(n20242) );
  MUX2_X1 U23335 ( .A(n9774), .B(n20242), .S(n15144), .Z(n20244) );
  NAND2_X1 U23336 ( .A1(n20244), .A2(n20243), .ZN(n20257) );
  AOI22_X1 U23337 ( .A1(n20247), .A2(n20246), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n20245), .ZN(n20248) );
  OAI211_X1 U23338 ( .C1(n20963), .C2(n20249), .A(n20248), .B(n12586), .ZN(
        n20254) );
  OAI22_X1 U23339 ( .A1(n20252), .A2(n20251), .B1(n20267), .B2(n20250), .ZN(
        n20253) );
  AOI211_X1 U23340 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20255), .A(
        n20254), .B(n20253), .ZN(n20256) );
  OAI21_X1 U23341 ( .B1(n20257), .B2(n20933), .A(n20256), .ZN(P2_U2848) );
  OAI22_X1 U23342 ( .A1(n20261), .A2(n20260), .B1(n20259), .B2(n20258), .ZN(
        n20262) );
  AOI211_X1 U23343 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n20264), .A(n20263), .B(
        n20262), .ZN(n20281) );
  OAI22_X1 U23344 ( .A1(n20292), .A2(n20267), .B1(n20266), .B2(n20265), .ZN(
        n20268) );
  INV_X1 U23345 ( .A(n20268), .ZN(n20280) );
  AOI22_X1 U23346 ( .A1(n20289), .A2(n20270), .B1(n20269), .B2(n20357), .ZN(
        n20279) );
  NAND2_X1 U23347 ( .A1(n20271), .A2(n20273), .ZN(n20272) );
  MUX2_X1 U23348 ( .A(n20273), .B(n20272), .S(n15144), .Z(n20277) );
  INV_X1 U23349 ( .A(n20274), .ZN(n20275) );
  NAND3_X1 U23350 ( .A1(n20277), .A2(n20276), .A3(n20275), .ZN(n20278) );
  NAND4_X1 U23351 ( .A1(n20281), .A2(n20280), .A3(n20279), .A4(n20278), .ZN(
        P2_U2851) );
  AOI211_X1 U23352 ( .C1(n20285), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        n20286) );
  AOI21_X1 U23353 ( .B1(n10444), .B2(n20291), .A(n20286), .ZN(n20287) );
  OAI21_X1 U23354 ( .B1(n20291), .B2(n10371), .A(n20287), .ZN(P2_U2877) );
  AOI22_X1 U23355 ( .A1(n20289), .A2(n20288), .B1(n20291), .B2(n20357), .ZN(
        n20290) );
  OAI21_X1 U23356 ( .B1(n20291), .B2(n20265), .A(n20290), .ZN(P2_U2883) );
  INV_X1 U23357 ( .A(n20292), .ZN(n20354) );
  AOI22_X1 U23358 ( .A1(n20354), .A2(n20307), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n20306), .ZN(n20298) );
  XNOR2_X1 U23359 ( .A(n20294), .B(n20293), .ZN(n20296) );
  NAND2_X1 U23360 ( .A1(n20296), .A2(n20295), .ZN(n20297) );
  OAI211_X1 U23361 ( .C1(n20388), .C2(n20315), .A(n20298), .B(n20297), .ZN(
        P2_U2915) );
  AOI22_X1 U23362 ( .A1(n21029), .A2(n20307), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n20306), .ZN(n20304) );
  AOI21_X1 U23363 ( .B1(n20301), .B2(n20300), .A(n20299), .ZN(n20302) );
  OR2_X1 U23364 ( .A1(n20302), .A2(n20311), .ZN(n20303) );
  OAI211_X1 U23365 ( .C1(n20305), .C2(n20315), .A(n20304), .B(n20303), .ZN(
        P2_U2916) );
  AOI22_X1 U23366 ( .A1(n20307), .A2(n21047), .B1(n20306), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n20314) );
  AOI21_X1 U23367 ( .B1(n20310), .B2(n20309), .A(n20308), .ZN(n20312) );
  OR2_X1 U23368 ( .A1(n20312), .A2(n20311), .ZN(n20313) );
  OAI211_X1 U23369 ( .C1(n20380), .C2(n20315), .A(n20314), .B(n20313), .ZN(
        P2_U2918) );
  NOR2_X1 U23370 ( .A1(n21709), .A2(n20323), .ZN(P2_U2920) );
  AOI22_X1 U23371 ( .A1(n13718), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20316) );
  OAI21_X1 U23372 ( .B1(n13553), .B2(n20348), .A(n20316), .ZN(P2_U2936) );
  AOI22_X1 U23373 ( .A1(n13718), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20317) );
  OAI21_X1 U23374 ( .B1(n20318), .B2(n20348), .A(n20317), .ZN(P2_U2937) );
  AOI22_X1 U23375 ( .A1(n13718), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n20319) );
  OAI21_X1 U23376 ( .B1(n20320), .B2(n20348), .A(n20319), .ZN(P2_U2938) );
  AOI22_X1 U23377 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n20321), .B1(n13718), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n20322) );
  OAI21_X1 U23378 ( .B1(n21660), .B2(n20323), .A(n20322), .ZN(P2_U2939) );
  AOI22_X1 U23379 ( .A1(n13718), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20324) );
  OAI21_X1 U23380 ( .B1(n20325), .B2(n20348), .A(n20324), .ZN(P2_U2940) );
  AOI22_X1 U23381 ( .A1(n13718), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20326) );
  OAI21_X1 U23382 ( .B1(n20327), .B2(n20348), .A(n20326), .ZN(P2_U2941) );
  AOI22_X1 U23383 ( .A1(n13718), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20328) );
  OAI21_X1 U23384 ( .B1(n20329), .B2(n20348), .A(n20328), .ZN(P2_U2942) );
  AOI22_X1 U23385 ( .A1(n13718), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20330) );
  OAI21_X1 U23386 ( .B1(n20331), .B2(n20348), .A(n20330), .ZN(P2_U2943) );
  AOI22_X1 U23387 ( .A1(n13718), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20332) );
  OAI21_X1 U23388 ( .B1(n20333), .B2(n20348), .A(n20332), .ZN(P2_U2944) );
  AOI22_X1 U23389 ( .A1(n13718), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20334) );
  OAI21_X1 U23390 ( .B1(n20335), .B2(n20348), .A(n20334), .ZN(P2_U2945) );
  INV_X1 U23391 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20337) );
  AOI22_X1 U23392 ( .A1(n13718), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n20336) );
  OAI21_X1 U23393 ( .B1(n20337), .B2(n20348), .A(n20336), .ZN(P2_U2946) );
  INV_X1 U23394 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20339) );
  AOI22_X1 U23395 ( .A1(n13718), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n20338) );
  OAI21_X1 U23396 ( .B1(n20339), .B2(n20348), .A(n20338), .ZN(P2_U2947) );
  INV_X1 U23397 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20341) );
  AOI22_X1 U23398 ( .A1(n13718), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n20340) );
  OAI21_X1 U23399 ( .B1(n20341), .B2(n20348), .A(n20340), .ZN(P2_U2948) );
  AOI22_X1 U23400 ( .A1(n13718), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n20342) );
  OAI21_X1 U23401 ( .B1(n20343), .B2(n20348), .A(n20342), .ZN(P2_U2949) );
  INV_X1 U23402 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20346) );
  AOI22_X1 U23403 ( .A1(n13718), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n20345) );
  OAI21_X1 U23404 ( .B1(n20346), .B2(n20348), .A(n20345), .ZN(P2_U2950) );
  INV_X1 U23405 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n20349) );
  AOI22_X1 U23406 ( .A1(n13718), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20344), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20347) );
  OAI21_X1 U23407 ( .B1(n20349), .B2(n20348), .A(n20347), .ZN(P2_U2951) );
  AOI22_X1 U23408 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n20351), .B1(n20350), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n20353) );
  NAND2_X1 U23409 ( .A1(n20353), .A2(n20352), .ZN(P2_U2979) );
  AOI22_X1 U23410 ( .A1(n20357), .A2(n20356), .B1(n20355), .B2(n20354), .ZN(
        n20367) );
  OAI22_X1 U23411 ( .A1(n20361), .A2(n20360), .B1(n20359), .B2(n20358), .ZN(
        n20362) );
  AOI221_X1 U23412 ( .B1(n20365), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n20364), .C2(n20363), .A(n20362), .ZN(n20366) );
  OAI211_X1 U23413 ( .C1(n12488), .C2(n12586), .A(n20367), .B(n20366), .ZN(
        P2_U3042) );
  INV_X1 U23414 ( .A(n20925), .ZN(n20395) );
  NAND2_X1 U23415 ( .A1(n20473), .A2(n21050), .ZN(n20416) );
  AOI22_X1 U23416 ( .A1(n20876), .A2(n20395), .B1(n20866), .B2(n20394), .ZN(
        n20378) );
  AOI21_X1 U23417 ( .B1(n20925), .B2(n20442), .A(n20814), .ZN(n20370) );
  NOR2_X1 U23418 ( .A1(n20370), .A2(n21065), .ZN(n20373) );
  AOI21_X1 U23419 ( .B1(n20374), .B2(n20821), .A(n21028), .ZN(n20371) );
  AOI21_X1 U23420 ( .B1(n20373), .B2(n20871), .A(n20371), .ZN(n20372) );
  OAI21_X1 U23421 ( .B1(n20372), .B2(n20394), .A(n20874), .ZN(n20412) );
  INV_X1 U23422 ( .A(n20871), .ZN(n20917) );
  OAI21_X1 U23423 ( .B1(n20917), .B2(n20394), .A(n20373), .ZN(n20376) );
  OAI21_X1 U23424 ( .B1(n20374), .B2(n20394), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20375) );
  AOI22_X1 U23425 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20412), .B1(
        n20867), .B2(n20411), .ZN(n20377) );
  OAI211_X1 U23426 ( .C1(n20879), .C2(n20442), .A(n20378), .B(n20377), .ZN(
        P2_U3048) );
  AOI22_X1 U23427 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20405), .ZN(n20885) );
  AOI22_X1 U23428 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20405), .ZN(n20751) );
  INV_X1 U23429 ( .A(n20880), .ZN(n20683) );
  INV_X1 U23430 ( .A(n20394), .ZN(n20408) );
  OAI22_X1 U23431 ( .A1(n20925), .A2(n20751), .B1(n20683), .B2(n20408), .ZN(
        n20379) );
  INV_X1 U23432 ( .A(n20379), .ZN(n20382) );
  NOR2_X2 U23433 ( .A1(n20823), .A2(n20380), .ZN(n20881) );
  AOI22_X1 U23434 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20412), .B1(
        n20881), .B2(n20411), .ZN(n20381) );
  OAI211_X1 U23435 ( .C1(n20885), .C2(n20442), .A(n20382), .B(n20381), .ZN(
        P2_U3049) );
  AOI22_X1 U23436 ( .A1(n20888), .A2(n20395), .B1(n20886), .B2(n20394), .ZN(
        n20384) );
  AOI22_X1 U23437 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20412), .B1(
        n20887), .B2(n20411), .ZN(n20383) );
  OAI211_X1 U23438 ( .C1(n20891), .C2(n20442), .A(n20384), .B(n20383), .ZN(
        P2_U3050) );
  AOI22_X1 U23439 ( .A1(n20894), .A2(n20395), .B1(n20892), .B2(n20394), .ZN(
        n20386) );
  AOI22_X1 U23440 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20412), .B1(
        n20893), .B2(n20411), .ZN(n20385) );
  OAI211_X1 U23441 ( .C1(n20897), .C2(n20442), .A(n20386), .B(n20385), .ZN(
        P2_U3051) );
  AOI22_X1 U23442 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20405), .ZN(n20903) );
  AOI22_X1 U23443 ( .A1(n20900), .A2(n20395), .B1(n20898), .B2(n20394), .ZN(
        n20390) );
  NOR2_X2 U23444 ( .A1(n20823), .A2(n20388), .ZN(n20899) );
  AOI22_X1 U23445 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20412), .B1(
        n20899), .B2(n20411), .ZN(n20389) );
  OAI211_X1 U23446 ( .C1(n20903), .C2(n20442), .A(n20390), .B(n20389), .ZN(
        P2_U3052) );
  AOI22_X1 U23447 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20405), .ZN(n20909) );
  AOI22_X1 U23448 ( .A1(n20906), .A2(n20395), .B1(n20904), .B2(n20394), .ZN(
        n20399) );
  INV_X1 U23449 ( .A(n20396), .ZN(n20397) );
  NOR2_X2 U23450 ( .A1(n20823), .A2(n20397), .ZN(n20905) );
  AOI22_X1 U23451 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20412), .B1(
        n20905), .B2(n20411), .ZN(n20398) );
  OAI211_X1 U23452 ( .C1(n20909), .C2(n20442), .A(n20399), .B(n20398), .ZN(
        P2_U3053) );
  AOI22_X1 U23453 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20405), .ZN(n20915) );
  AOI22_X1 U23454 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20405), .ZN(n20766) );
  INV_X1 U23455 ( .A(n20910), .ZN(n20697) );
  OAI22_X1 U23456 ( .A1(n20925), .A2(n20766), .B1(n20697), .B2(n20408), .ZN(
        n20401) );
  INV_X1 U23457 ( .A(n20401), .ZN(n20404) );
  NOR2_X2 U23458 ( .A1(n20823), .A2(n20402), .ZN(n20911) );
  AOI22_X1 U23459 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20412), .B1(
        n20911), .B2(n20411), .ZN(n20403) );
  OAI211_X1 U23460 ( .C1(n20915), .C2(n20442), .A(n20404), .B(n20403), .ZN(
        P2_U3054) );
  AOI22_X1 U23461 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20405), .ZN(n20926) );
  AOI22_X1 U23462 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20406), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20405), .ZN(n20773) );
  INV_X1 U23463 ( .A(n20916), .ZN(n20664) );
  OAI22_X1 U23464 ( .A1(n20925), .A2(n20773), .B1(n20664), .B2(n20408), .ZN(
        n20409) );
  INV_X1 U23465 ( .A(n20409), .ZN(n20414) );
  NOR2_X2 U23466 ( .A1(n20823), .A2(n20410), .ZN(n20918) );
  AOI22_X1 U23467 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20412), .B1(
        n20918), .B2(n20411), .ZN(n20413) );
  OAI211_X1 U23468 ( .C1(n20926), .C2(n20442), .A(n20414), .B(n20413), .ZN(
        P2_U3055) );
  INV_X1 U23469 ( .A(n20876), .ZN(n20748) );
  INV_X1 U23470 ( .A(n20473), .ZN(n20476) );
  NOR2_X1 U23471 ( .A1(n20672), .A2(n20476), .ZN(n20437) );
  INV_X1 U23472 ( .A(n20419), .ZN(n20415) );
  AOI211_X2 U23473 ( .C1(n20416), .C2(n20864), .A(n20571), .B(n20415), .ZN(
        n20438) );
  AOI22_X1 U23474 ( .A1(n20438), .A2(n20867), .B1(n20866), .B2(n20437), .ZN(
        n20424) );
  NAND2_X1 U23475 ( .A1(n20422), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20601) );
  OAI21_X1 U23476 ( .B1(n20601), .B2(n20674), .A(n20416), .ZN(n20420) );
  INV_X1 U23477 ( .A(n20437), .ZN(n20417) );
  NAND2_X1 U23478 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20417), .ZN(n20418) );
  NAND4_X1 U23479 ( .A1(n20420), .A2(n20874), .A3(n20419), .A4(n20418), .ZN(
        n20439) );
  NOR2_X2 U23480 ( .A1(n20674), .A2(n20598), .ZN(n20443) );
  AOI22_X1 U23481 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20828), .ZN(n20423) );
  OAI211_X1 U23482 ( .C1(n20748), .C2(n20442), .A(n20424), .B(n20423), .ZN(
        P2_U3056) );
  AOI22_X1 U23483 ( .A1(n20438), .A2(n20881), .B1(n20880), .B2(n20437), .ZN(
        n20426) );
  AOI22_X1 U23484 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20832), .ZN(n20425) );
  OAI211_X1 U23485 ( .C1(n20751), .C2(n20442), .A(n20426), .B(n20425), .ZN(
        P2_U3057) );
  AOI22_X1 U23486 ( .A1(n20438), .A2(n20887), .B1(n20886), .B2(n20437), .ZN(
        n20428) );
  AOI22_X1 U23487 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20835), .ZN(n20427) );
  OAI211_X1 U23488 ( .C1(n20754), .C2(n20442), .A(n20428), .B(n20427), .ZN(
        P2_U3058) );
  AOI22_X1 U23489 ( .A1(n20438), .A2(n20893), .B1(n20892), .B2(n20437), .ZN(
        n20430) );
  AOI22_X1 U23490 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20839), .ZN(n20429) );
  OAI211_X1 U23491 ( .C1(n20757), .C2(n20442), .A(n20430), .B(n20429), .ZN(
        P2_U3059) );
  AOI22_X1 U23492 ( .A1(n20438), .A2(n20899), .B1(n20898), .B2(n20437), .ZN(
        n20432) );
  AOI22_X1 U23493 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20843), .ZN(n20431) );
  OAI211_X1 U23494 ( .C1(n20760), .C2(n20442), .A(n20432), .B(n20431), .ZN(
        P2_U3060) );
  AOI22_X1 U23495 ( .A1(n20438), .A2(n20905), .B1(n20904), .B2(n20437), .ZN(
        n20434) );
  INV_X1 U23496 ( .A(n20909), .ZN(n20847) );
  AOI22_X1 U23497 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20847), .ZN(n20433) );
  OAI211_X1 U23498 ( .C1(n20763), .C2(n20442), .A(n20434), .B(n20433), .ZN(
        P2_U3061) );
  AOI22_X1 U23499 ( .A1(n20438), .A2(n20911), .B1(n20910), .B2(n20437), .ZN(
        n20436) );
  INV_X1 U23500 ( .A(n20915), .ZN(n20851) );
  AOI22_X1 U23501 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20851), .ZN(n20435) );
  OAI211_X1 U23502 ( .C1(n20766), .C2(n20442), .A(n20436), .B(n20435), .ZN(
        P2_U3062) );
  AOI22_X1 U23503 ( .A1(n20438), .A2(n20918), .B1(n20916), .B2(n20437), .ZN(
        n20441) );
  INV_X1 U23504 ( .A(n20926), .ZN(n20856) );
  AOI22_X1 U23505 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20439), .B1(
        n20443), .B2(n20856), .ZN(n20440) );
  OAI211_X1 U23506 ( .C1(n20773), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P2_U3063) );
  NOR2_X1 U23507 ( .A1(n20476), .A2(n20820), .ZN(n20467) );
  OAI21_X1 U23508 ( .B1(n20446), .B2(n20467), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20445) );
  AND2_X1 U23509 ( .A1(n20473), .A2(n20706), .ZN(n20448) );
  INV_X1 U23510 ( .A(n20448), .ZN(n20444) );
  NAND2_X1 U23511 ( .A1(n20445), .A2(n20444), .ZN(n20468) );
  AOI22_X1 U23512 ( .A1(n20468), .A2(n20867), .B1(n20866), .B2(n20467), .ZN(
        n20454) );
  AOI21_X1 U23513 ( .B1(n20446), .B2(n20821), .A(n20467), .ZN(n20451) );
  INV_X1 U23514 ( .A(n20569), .ZN(n20447) );
  INV_X1 U23515 ( .A(n20741), .ZN(n21024) );
  NAND2_X1 U23516 ( .A1(n20505), .A2(n20472), .ZN(n20449) );
  AOI21_X1 U23517 ( .B1(n20449), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20448), 
        .ZN(n20450) );
  MUX2_X1 U23518 ( .A(n20451), .B(n20450), .S(n21028), .Z(n20452) );
  AOI22_X1 U23519 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20828), .ZN(n20453) );
  OAI211_X1 U23520 ( .C1(n20748), .C2(n20472), .A(n20454), .B(n20453), .ZN(
        P2_U3064) );
  AOI22_X1 U23521 ( .A1(n20468), .A2(n20881), .B1(n20467), .B2(n20880), .ZN(
        n20456) );
  AOI22_X1 U23522 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20832), .ZN(n20455) );
  OAI211_X1 U23523 ( .C1(n20751), .C2(n20472), .A(n20456), .B(n20455), .ZN(
        P2_U3065) );
  AOI22_X1 U23524 ( .A1(n20468), .A2(n20887), .B1(n20886), .B2(n20467), .ZN(
        n20458) );
  AOI22_X1 U23525 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20835), .ZN(n20457) );
  OAI211_X1 U23526 ( .C1(n20754), .C2(n20472), .A(n20458), .B(n20457), .ZN(
        P2_U3066) );
  AOI22_X1 U23527 ( .A1(n20468), .A2(n20893), .B1(n20892), .B2(n20467), .ZN(
        n20460) );
  AOI22_X1 U23528 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20839), .ZN(n20459) );
  OAI211_X1 U23529 ( .C1(n20757), .C2(n20472), .A(n20460), .B(n20459), .ZN(
        P2_U3067) );
  AOI22_X1 U23530 ( .A1(n20468), .A2(n20899), .B1(n20467), .B2(n20898), .ZN(
        n20462) );
  AOI22_X1 U23531 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20843), .ZN(n20461) );
  OAI211_X1 U23532 ( .C1(n20760), .C2(n20472), .A(n20462), .B(n20461), .ZN(
        P2_U3068) );
  AOI22_X1 U23533 ( .A1(n20468), .A2(n20905), .B1(n20467), .B2(n20904), .ZN(
        n20464) );
  AOI22_X1 U23534 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20847), .ZN(n20463) );
  OAI211_X1 U23535 ( .C1(n20763), .C2(n20472), .A(n20464), .B(n20463), .ZN(
        P2_U3069) );
  AOI22_X1 U23536 ( .A1(n20468), .A2(n20911), .B1(n20467), .B2(n20910), .ZN(
        n20466) );
  AOI22_X1 U23537 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20851), .ZN(n20465) );
  OAI211_X1 U23538 ( .C1(n20766), .C2(n20472), .A(n20466), .B(n20465), .ZN(
        P2_U3070) );
  AOI22_X1 U23539 ( .A1(n20468), .A2(n20918), .B1(n20467), .B2(n20916), .ZN(
        n20471) );
  AOI22_X1 U23540 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20469), .B1(
        n20498), .B2(n20856), .ZN(n20470) );
  OAI211_X1 U23541 ( .C1(n20773), .C2(n20472), .A(n20471), .B(n20470), .ZN(
        P2_U3071) );
  OAI21_X1 U23542 ( .B1(n20601), .B2(n20741), .A(n21028), .ZN(n20483) );
  NAND2_X1 U23543 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20473), .ZN(
        n20482) );
  INV_X1 U23544 ( .A(n20482), .ZN(n20474) );
  OR2_X1 U23545 ( .A1(n20483), .A2(n20474), .ZN(n20479) );
  OAI21_X1 U23546 ( .B1(n12298), .B2(n20864), .A(n20821), .ZN(n20477) );
  NOR2_X1 U23547 ( .A1(n20476), .A2(n20475), .ZN(n20497) );
  INV_X1 U23548 ( .A(n20497), .ZN(n20504) );
  AOI21_X1 U23549 ( .B1(n20477), .B2(n20504), .A(n20823), .ZN(n20478) );
  INV_X1 U23550 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n21567) );
  AOI22_X1 U23551 ( .A1(n20535), .A2(n20828), .B1(n20866), .B2(n20497), .ZN(
        n20485) );
  OAI21_X1 U23552 ( .B1(n12298), .B2(n20497), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20481) );
  AOI22_X1 U23553 ( .A1(n20867), .A2(n20507), .B1(n20498), .B2(n20876), .ZN(
        n20484) );
  OAI211_X1 U23554 ( .C1(n20492), .C2(n21567), .A(n20485), .B(n20484), .ZN(
        P2_U3072) );
  OAI22_X1 U23555 ( .A1(n20505), .A2(n20751), .B1(n20504), .B2(n20683), .ZN(
        n20486) );
  INV_X1 U23556 ( .A(n20486), .ZN(n20488) );
  AOI22_X1 U23557 ( .A1(n20881), .A2(n20507), .B1(n20535), .B2(n20832), .ZN(
        n20487) );
  OAI211_X1 U23558 ( .C1(n20492), .C2(n12212), .A(n20488), .B(n20487), .ZN(
        P2_U3073) );
  AOI22_X1 U23559 ( .A1(n20535), .A2(n20835), .B1(n20886), .B2(n20497), .ZN(
        n20490) );
  AOI22_X1 U23560 ( .A1(n20887), .A2(n20507), .B1(n20498), .B2(n20888), .ZN(
        n20489) );
  OAI211_X1 U23561 ( .C1(n20492), .C2(n20491), .A(n20490), .B(n20489), .ZN(
        P2_U3074) );
  AOI22_X1 U23562 ( .A1(n20535), .A2(n20839), .B1(n20892), .B2(n20497), .ZN(
        n20494) );
  AOI22_X1 U23563 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20508), .B1(
        n20893), .B2(n20507), .ZN(n20493) );
  OAI211_X1 U23564 ( .C1(n20757), .C2(n20505), .A(n20494), .B(n20493), .ZN(
        P2_U3075) );
  AOI22_X1 U23565 ( .A1(n20900), .A2(n20498), .B1(n20497), .B2(n20898), .ZN(
        n20496) );
  AOI22_X1 U23566 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20508), .B1(
        n20899), .B2(n20507), .ZN(n20495) );
  OAI211_X1 U23567 ( .C1(n20903), .C2(n20513), .A(n20496), .B(n20495), .ZN(
        P2_U3076) );
  AOI22_X1 U23568 ( .A1(n20906), .A2(n20498), .B1(n20497), .B2(n20904), .ZN(
        n20500) );
  AOI22_X1 U23569 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20508), .B1(
        n20905), .B2(n20507), .ZN(n20499) );
  OAI211_X1 U23570 ( .C1(n20909), .C2(n20513), .A(n20500), .B(n20499), .ZN(
        P2_U3077) );
  OAI22_X1 U23571 ( .A1(n20505), .A2(n20766), .B1(n20504), .B2(n20697), .ZN(
        n20501) );
  INV_X1 U23572 ( .A(n20501), .ZN(n20503) );
  AOI22_X1 U23573 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20508), .B1(
        n20911), .B2(n20507), .ZN(n20502) );
  OAI211_X1 U23574 ( .C1(n20915), .C2(n20513), .A(n20503), .B(n20502), .ZN(
        P2_U3078) );
  OAI22_X1 U23575 ( .A1(n20505), .A2(n20773), .B1(n20504), .B2(n20664), .ZN(
        n20506) );
  INV_X1 U23576 ( .A(n20506), .ZN(n20510) );
  AOI22_X1 U23577 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20508), .B1(
        n20918), .B2(n20507), .ZN(n20509) );
  OAI211_X1 U23578 ( .C1(n20926), .C2(n20513), .A(n20510), .B(n20509), .ZN(
        P2_U3079) );
  NAND2_X1 U23579 ( .A1(n21552), .A2(n21050), .ZN(n20546) );
  NOR3_X1 U23580 ( .A1(n12291), .A2(n20533), .A3(n20864), .ZN(n20514) );
  NOR2_X1 U23581 ( .A1(n20511), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20518) );
  AOI21_X1 U23582 ( .B1(n20821), .B2(n20518), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20512) );
  AOI22_X1 U23583 ( .A1(n20534), .A2(n20867), .B1(n20866), .B2(n20533), .ZN(
        n20520) );
  AOI21_X1 U23584 ( .B1(n20513), .B2(n20562), .A(n20814), .ZN(n20517) );
  INV_X1 U23585 ( .A(n20533), .ZN(n20515) );
  AOI211_X1 U23586 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20515), .A(n20823), 
        .B(n20514), .ZN(n20516) );
  AOI22_X1 U23587 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20876), .ZN(n20519) );
  OAI211_X1 U23588 ( .C1(n20879), .C2(n20562), .A(n20520), .B(n20519), .ZN(
        P2_U3080) );
  AOI22_X1 U23589 ( .A1(n20534), .A2(n20881), .B1(n20880), .B2(n20533), .ZN(
        n20522) );
  INV_X1 U23590 ( .A(n20751), .ZN(n20882) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20882), .ZN(n20521) );
  OAI211_X1 U23592 ( .C1(n20885), .C2(n20562), .A(n20522), .B(n20521), .ZN(
        P2_U3081) );
  AOI22_X1 U23593 ( .A1(n20534), .A2(n20887), .B1(n20886), .B2(n20533), .ZN(
        n20524) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20888), .ZN(n20523) );
  OAI211_X1 U23595 ( .C1(n20891), .C2(n20562), .A(n20524), .B(n20523), .ZN(
        P2_U3082) );
  AOI22_X1 U23596 ( .A1(n20534), .A2(n20893), .B1(n20892), .B2(n20533), .ZN(
        n20526) );
  AOI22_X1 U23597 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20894), .ZN(n20525) );
  OAI211_X1 U23598 ( .C1(n20897), .C2(n20562), .A(n20526), .B(n20525), .ZN(
        P2_U3083) );
  AOI22_X1 U23599 ( .A1(n20534), .A2(n20899), .B1(n20898), .B2(n20533), .ZN(
        n20528) );
  AOI22_X1 U23600 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20900), .ZN(n20527) );
  OAI211_X1 U23601 ( .C1(n20903), .C2(n20562), .A(n20528), .B(n20527), .ZN(
        P2_U3084) );
  AOI22_X1 U23602 ( .A1(n20534), .A2(n20905), .B1(n20904), .B2(n20533), .ZN(
        n20530) );
  AOI22_X1 U23603 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20906), .ZN(n20529) );
  OAI211_X1 U23604 ( .C1(n20909), .C2(n20562), .A(n20530), .B(n20529), .ZN(
        P2_U3085) );
  AOI22_X1 U23605 ( .A1(n20534), .A2(n20911), .B1(n20910), .B2(n20533), .ZN(
        n20532) );
  INV_X1 U23606 ( .A(n20766), .ZN(n20912) );
  AOI22_X1 U23607 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20912), .ZN(n20531) );
  OAI211_X1 U23608 ( .C1(n20915), .C2(n20562), .A(n20532), .B(n20531), .ZN(
        P2_U3086) );
  AOI22_X1 U23609 ( .A1(n20534), .A2(n20918), .B1(n20916), .B2(n20533), .ZN(
        n20538) );
  INV_X1 U23610 ( .A(n20773), .ZN(n20920) );
  AOI22_X1 U23611 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20536), .B1(
        n20535), .B2(n20920), .ZN(n20537) );
  OAI211_X1 U23612 ( .C1(n20926), .C2(n20562), .A(n20538), .B(n20537), .ZN(
        P2_U3087) );
  INV_X1 U23613 ( .A(n21552), .ZN(n20570) );
  NOR2_X1 U23614 ( .A1(n20672), .A2(n20570), .ZN(n20563) );
  AOI22_X1 U23615 ( .A1(n20588), .A2(n20828), .B1(n20866), .B2(n20563), .ZN(
        n20549) );
  AOI21_X1 U23616 ( .B1(n9905), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20543) );
  INV_X1 U23617 ( .A(n20601), .ZN(n20541) );
  INV_X1 U23618 ( .A(n20539), .ZN(n20540) );
  AOI21_X1 U23619 ( .B1(n20541), .B2(n20540), .A(n21065), .ZN(n20544) );
  NAND2_X1 U23620 ( .A1(n20544), .A2(n20546), .ZN(n20542) );
  OAI211_X1 U23621 ( .C1(n20563), .C2(n20543), .A(n20542), .B(n20874), .ZN(
        n20566) );
  INV_X1 U23622 ( .A(n20544), .ZN(n20547) );
  OAI21_X1 U23623 ( .B1(n12320), .B2(n20563), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20545) );
  AOI22_X1 U23624 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20566), .B1(
        n20867), .B2(n20565), .ZN(n20548) );
  OAI211_X1 U23625 ( .C1(n20748), .C2(n20562), .A(n20549), .B(n20548), .ZN(
        P2_U3088) );
  AOI22_X1 U23626 ( .A1(n20588), .A2(n20832), .B1(n20563), .B2(n20880), .ZN(
        n20551) );
  AOI22_X1 U23627 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20566), .B1(
        n20881), .B2(n20565), .ZN(n20550) );
  OAI211_X1 U23628 ( .C1(n20751), .C2(n20562), .A(n20551), .B(n20550), .ZN(
        P2_U3089) );
  AOI22_X1 U23629 ( .A1(n20588), .A2(n20835), .B1(n20886), .B2(n20563), .ZN(
        n20553) );
  AOI22_X1 U23630 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20566), .B1(
        n20887), .B2(n20565), .ZN(n20552) );
  OAI211_X1 U23631 ( .C1(n20754), .C2(n20562), .A(n20553), .B(n20552), .ZN(
        P2_U3090) );
  AOI22_X1 U23632 ( .A1(n20588), .A2(n20839), .B1(n20892), .B2(n20563), .ZN(
        n20555) );
  AOI22_X1 U23633 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20566), .B1(
        n20893), .B2(n20565), .ZN(n20554) );
  OAI211_X1 U23634 ( .C1(n20757), .C2(n20562), .A(n20555), .B(n20554), .ZN(
        P2_U3091) );
  AOI22_X1 U23635 ( .A1(n20588), .A2(n20843), .B1(n20563), .B2(n20898), .ZN(
        n20557) );
  AOI22_X1 U23636 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20566), .B1(
        n20899), .B2(n20565), .ZN(n20556) );
  OAI211_X1 U23637 ( .C1(n20760), .C2(n20562), .A(n20557), .B(n20556), .ZN(
        P2_U3092) );
  AOI22_X1 U23638 ( .A1(n20906), .A2(n20564), .B1(n20563), .B2(n20904), .ZN(
        n20559) );
  AOI22_X1 U23639 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20566), .B1(
        n20905), .B2(n20565), .ZN(n20558) );
  OAI211_X1 U23640 ( .C1(n20909), .C2(n20597), .A(n20559), .B(n20558), .ZN(
        P2_U3093) );
  AOI22_X1 U23641 ( .A1(n20588), .A2(n20851), .B1(n20563), .B2(n20910), .ZN(
        n20561) );
  AOI22_X1 U23642 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20566), .B1(
        n20911), .B2(n20565), .ZN(n20560) );
  OAI211_X1 U23643 ( .C1(n20766), .C2(n20562), .A(n20561), .B(n20560), .ZN(
        P2_U3094) );
  AOI22_X1 U23644 ( .A1(n20564), .A2(n20920), .B1(n20563), .B2(n20916), .ZN(
        n20568) );
  AOI22_X1 U23645 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20566), .B1(
        n20918), .B2(n20565), .ZN(n20567) );
  OAI211_X1 U23646 ( .C1(n20926), .C2(n20597), .A(n20568), .B(n20567), .ZN(
        P2_U3095) );
  INV_X1 U23647 ( .A(n20622), .ZN(n20591) );
  NAND2_X1 U23648 ( .A1(n20818), .A2(n21552), .ZN(n20573) );
  NOR3_X1 U23649 ( .A1(n12296), .A2(n20592), .A3(n20864), .ZN(n20572) );
  AOI211_X2 U23650 ( .C1(n20864), .C2(n20573), .A(n20571), .B(n20572), .ZN(
        n20593) );
  AOI22_X1 U23651 ( .A1(n20593), .A2(n20867), .B1(n20866), .B2(n20592), .ZN(
        n20577) );
  OAI21_X1 U23652 ( .B1(n20588), .B2(n20622), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20574) );
  AOI211_X1 U23653 ( .C1(n20574), .C2(n20573), .A(n20823), .B(n20572), .ZN(
        n20575) );
  OAI21_X1 U23654 ( .B1(n20592), .B2(n20821), .A(n20575), .ZN(n20594) );
  AOI22_X1 U23655 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20594), .B1(
        n20588), .B2(n20876), .ZN(n20576) );
  OAI211_X1 U23656 ( .C1(n20879), .C2(n20591), .A(n20577), .B(n20576), .ZN(
        P2_U3096) );
  AOI22_X1 U23657 ( .A1(n20593), .A2(n20881), .B1(n20592), .B2(n20880), .ZN(
        n20579) );
  AOI22_X1 U23658 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20832), .ZN(n20578) );
  OAI211_X1 U23659 ( .C1(n20751), .C2(n20597), .A(n20579), .B(n20578), .ZN(
        P2_U3097) );
  AOI22_X1 U23660 ( .A1(n20593), .A2(n20887), .B1(n20886), .B2(n20592), .ZN(
        n20581) );
  AOI22_X1 U23661 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20835), .ZN(n20580) );
  OAI211_X1 U23662 ( .C1(n20754), .C2(n20597), .A(n20581), .B(n20580), .ZN(
        P2_U3098) );
  AOI22_X1 U23663 ( .A1(n20593), .A2(n20893), .B1(n20892), .B2(n20592), .ZN(
        n20583) );
  AOI22_X1 U23664 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20839), .ZN(n20582) );
  OAI211_X1 U23665 ( .C1(n20757), .C2(n20597), .A(n20583), .B(n20582), .ZN(
        P2_U3099) );
  AOI22_X1 U23666 ( .A1(n20593), .A2(n20899), .B1(n20592), .B2(n20898), .ZN(
        n20585) );
  AOI22_X1 U23667 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20843), .ZN(n20584) );
  OAI211_X1 U23668 ( .C1(n20760), .C2(n20597), .A(n20585), .B(n20584), .ZN(
        P2_U3100) );
  AOI22_X1 U23669 ( .A1(n20593), .A2(n20905), .B1(n20592), .B2(n20904), .ZN(
        n20587) );
  AOI22_X1 U23670 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20847), .ZN(n20586) );
  OAI211_X1 U23671 ( .C1(n20763), .C2(n20597), .A(n20587), .B(n20586), .ZN(
        P2_U3101) );
  AOI22_X1 U23672 ( .A1(n20593), .A2(n20911), .B1(n20592), .B2(n20910), .ZN(
        n20590) );
  AOI22_X1 U23673 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20594), .B1(
        n20588), .B2(n20912), .ZN(n20589) );
  OAI211_X1 U23674 ( .C1(n20915), .C2(n20591), .A(n20590), .B(n20589), .ZN(
        P2_U3102) );
  AOI22_X1 U23675 ( .A1(n20593), .A2(n20918), .B1(n20592), .B2(n20916), .ZN(
        n20596) );
  AOI22_X1 U23676 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20594), .B1(
        n20622), .B2(n20856), .ZN(n20595) );
  OAI211_X1 U23677 ( .C1(n20773), .C2(n20597), .A(n20596), .B(n20595), .ZN(
        P2_U3103) );
  NAND2_X1 U23678 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21552), .ZN(
        n20602) );
  AND2_X1 U23679 ( .A1(n20737), .A2(n21552), .ZN(n20630) );
  OAI21_X1 U23680 ( .B1(n20599), .B2(n20630), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20600) );
  AOI22_X1 U23681 ( .A1(n20621), .A2(n20867), .B1(n20866), .B2(n20630), .ZN(
        n20608) );
  NOR2_X1 U23682 ( .A1(n20601), .A2(n20869), .ZN(n21027) );
  INV_X1 U23683 ( .A(n20602), .ZN(n20606) );
  INV_X1 U23684 ( .A(n20630), .ZN(n20603) );
  OAI211_X1 U23685 ( .C1(n20604), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n21065), 
        .B(n20603), .ZN(n20605) );
  OAI211_X1 U23686 ( .C1(n21027), .C2(n20606), .A(n20874), .B(n20605), .ZN(
        n20623) );
  AOI22_X1 U23687 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20876), .ZN(n20607) );
  OAI211_X1 U23688 ( .C1(n20879), .C2(n20670), .A(n20608), .B(n20607), .ZN(
        P2_U3104) );
  AOI22_X1 U23689 ( .A1(n20621), .A2(n20881), .B1(n20630), .B2(n20880), .ZN(
        n20610) );
  AOI22_X1 U23690 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20882), .ZN(n20609) );
  OAI211_X1 U23691 ( .C1(n20885), .C2(n20670), .A(n20610), .B(n20609), .ZN(
        P2_U3105) );
  AOI22_X1 U23692 ( .A1(n20621), .A2(n20887), .B1(n20886), .B2(n20630), .ZN(
        n20612) );
  AOI22_X1 U23693 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20888), .ZN(n20611) );
  OAI211_X1 U23694 ( .C1(n20891), .C2(n20670), .A(n20612), .B(n20611), .ZN(
        P2_U3106) );
  AOI22_X1 U23695 ( .A1(n20621), .A2(n20893), .B1(n20892), .B2(n20630), .ZN(
        n20614) );
  AOI22_X1 U23696 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20894), .ZN(n20613) );
  OAI211_X1 U23697 ( .C1(n20897), .C2(n20670), .A(n20614), .B(n20613), .ZN(
        P2_U3107) );
  AOI22_X1 U23698 ( .A1(n20621), .A2(n20899), .B1(n20630), .B2(n20898), .ZN(
        n20616) );
  AOI22_X1 U23699 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20900), .ZN(n20615) );
  OAI211_X1 U23700 ( .C1(n20903), .C2(n20670), .A(n20616), .B(n20615), .ZN(
        P2_U3108) );
  AOI22_X1 U23701 ( .A1(n20621), .A2(n20905), .B1(n20630), .B2(n20904), .ZN(
        n20618) );
  AOI22_X1 U23702 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20906), .ZN(n20617) );
  OAI211_X1 U23703 ( .C1(n20909), .C2(n20670), .A(n20618), .B(n20617), .ZN(
        P2_U3109) );
  AOI22_X1 U23704 ( .A1(n20621), .A2(n20911), .B1(n20630), .B2(n20910), .ZN(
        n20620) );
  AOI22_X1 U23705 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20912), .ZN(n20619) );
  OAI211_X1 U23706 ( .C1(n20915), .C2(n20670), .A(n20620), .B(n20619), .ZN(
        P2_U3110) );
  AOI22_X1 U23707 ( .A1(n20621), .A2(n20918), .B1(n20630), .B2(n20916), .ZN(
        n20625) );
  AOI22_X1 U23708 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20623), .B1(
        n20622), .B2(n20920), .ZN(n20624) );
  OAI211_X1 U23709 ( .C1(n20926), .C2(n20670), .A(n20625), .B(n20624), .ZN(
        P2_U3111) );
  INV_X1 U23710 ( .A(n20866), .ZN(n20626) );
  NAND2_X1 U23711 ( .A1(n21692), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20740) );
  NOR2_X1 U23712 ( .A1(n20740), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20677) );
  INV_X1 U23713 ( .A(n20677), .ZN(n20679) );
  NOR2_X1 U23714 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20679), .ZN(
        n20634) );
  INV_X1 U23715 ( .A(n20634), .ZN(n20663) );
  OAI22_X1 U23716 ( .A1(n20705), .A2(n20879), .B1(n20626), .B2(n20663), .ZN(
        n20627) );
  INV_X1 U23717 ( .A(n20627), .ZN(n20640) );
  AOI21_X1 U23718 ( .B1(n12218), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20633) );
  INV_X1 U23719 ( .A(n20705), .ZN(n20689) );
  INV_X1 U23720 ( .A(n20670), .ZN(n20628) );
  OAI21_X1 U23721 ( .B1(n20689), .B2(n20628), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20629) );
  NAND2_X1 U23722 ( .A1(n20629), .A2(n21028), .ZN(n20638) );
  INV_X1 U23723 ( .A(n20638), .ZN(n20631) );
  NOR2_X1 U23724 ( .A1(n20634), .A2(n20630), .ZN(n20636) );
  NAND2_X1 U23725 ( .A1(n20631), .A2(n20636), .ZN(n20632) );
  OAI211_X1 U23726 ( .C1(n20634), .C2(n20633), .A(n20632), .B(n20874), .ZN(
        n20667) );
  OAI21_X1 U23727 ( .B1(n20635), .B2(n20634), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20637) );
  AOI22_X1 U23728 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20667), .B1(
        n20867), .B2(n20666), .ZN(n20639) );
  OAI211_X1 U23729 ( .C1(n20748), .C2(n20670), .A(n20640), .B(n20639), .ZN(
        P2_U3112) );
  OAI22_X1 U23730 ( .A1(n20705), .A2(n20885), .B1(n20683), .B2(n20663), .ZN(
        n20641) );
  INV_X1 U23731 ( .A(n20641), .ZN(n20643) );
  AOI22_X1 U23732 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20667), .B1(
        n20881), .B2(n20666), .ZN(n20642) );
  OAI211_X1 U23733 ( .C1(n20751), .C2(n20670), .A(n20643), .B(n20642), .ZN(
        P2_U3113) );
  INV_X1 U23734 ( .A(n20886), .ZN(n20644) );
  OAI22_X1 U23735 ( .A1(n20705), .A2(n20891), .B1(n20644), .B2(n20663), .ZN(
        n20645) );
  INV_X1 U23736 ( .A(n20645), .ZN(n20647) );
  AOI22_X1 U23737 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20667), .B1(
        n20887), .B2(n20666), .ZN(n20646) );
  OAI211_X1 U23738 ( .C1(n20754), .C2(n20670), .A(n20647), .B(n20646), .ZN(
        P2_U3114) );
  INV_X1 U23739 ( .A(n20892), .ZN(n20648) );
  OAI22_X1 U23740 ( .A1(n20705), .A2(n20897), .B1(n20648), .B2(n20663), .ZN(
        n20649) );
  INV_X1 U23741 ( .A(n20649), .ZN(n20651) );
  AOI22_X1 U23742 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20667), .B1(
        n20893), .B2(n20666), .ZN(n20650) );
  OAI211_X1 U23743 ( .C1(n20757), .C2(n20670), .A(n20651), .B(n20650), .ZN(
        P2_U3115) );
  INV_X1 U23744 ( .A(n20898), .ZN(n20652) );
  OAI22_X1 U23745 ( .A1(n20705), .A2(n20903), .B1(n20652), .B2(n20663), .ZN(
        n20653) );
  INV_X1 U23746 ( .A(n20653), .ZN(n20655) );
  AOI22_X1 U23747 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20667), .B1(
        n20899), .B2(n20666), .ZN(n20654) );
  OAI211_X1 U23748 ( .C1(n20760), .C2(n20670), .A(n20655), .B(n20654), .ZN(
        P2_U3116) );
  INV_X1 U23749 ( .A(n20904), .ZN(n20656) );
  OAI22_X1 U23750 ( .A1(n20705), .A2(n20909), .B1(n20656), .B2(n20663), .ZN(
        n20657) );
  INV_X1 U23751 ( .A(n20657), .ZN(n20659) );
  AOI22_X1 U23752 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20667), .B1(
        n20905), .B2(n20666), .ZN(n20658) );
  OAI211_X1 U23753 ( .C1(n20763), .C2(n20670), .A(n20659), .B(n20658), .ZN(
        P2_U3117) );
  OAI22_X1 U23754 ( .A1(n20705), .A2(n20915), .B1(n20697), .B2(n20663), .ZN(
        n20660) );
  INV_X1 U23755 ( .A(n20660), .ZN(n20662) );
  AOI22_X1 U23756 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20667), .B1(
        n20911), .B2(n20666), .ZN(n20661) );
  OAI211_X1 U23757 ( .C1(n20766), .C2(n20670), .A(n20662), .B(n20661), .ZN(
        P2_U3118) );
  OAI22_X1 U23758 ( .A1(n20705), .A2(n20926), .B1(n20664), .B2(n20663), .ZN(
        n20665) );
  INV_X1 U23759 ( .A(n20665), .ZN(n20669) );
  AOI22_X1 U23760 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20667), .B1(
        n20918), .B2(n20666), .ZN(n20668) );
  OAI211_X1 U23761 ( .C1(n20773), .C2(n20670), .A(n20669), .B(n20668), .ZN(
        P2_U3119) );
  NOR2_X1 U23762 ( .A1(n20672), .A2(n20740), .ZN(n20710) );
  AOI22_X1 U23763 ( .A1(n20876), .A2(n20689), .B1(n20866), .B2(n20710), .ZN(
        n20682) );
  INV_X1 U23764 ( .A(n20673), .ZN(n20870) );
  OAI21_X1 U23765 ( .B1(n20870), .B2(n20674), .A(n21028), .ZN(n20680) );
  INV_X1 U23766 ( .A(n20710), .ZN(n20696) );
  OAI211_X1 U23767 ( .C1(n20675), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n21065), 
        .B(n20696), .ZN(n20676) );
  OAI211_X1 U23768 ( .C1(n20680), .C2(n20677), .A(n20874), .B(n20676), .ZN(
        n20702) );
  OAI21_X1 U23769 ( .B1(n12299), .B2(n20710), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20678) );
  AOI22_X1 U23770 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20702), .B1(
        n20867), .B2(n20701), .ZN(n20681) );
  OAI211_X1 U23771 ( .C1(n20879), .C2(n20734), .A(n20682), .B(n20681), .ZN(
        P2_U3120) );
  OAI22_X1 U23772 ( .A1(n20705), .A2(n20751), .B1(n20683), .B2(n20696), .ZN(
        n20684) );
  INV_X1 U23773 ( .A(n20684), .ZN(n20686) );
  AOI22_X1 U23774 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20702), .B1(
        n20881), .B2(n20701), .ZN(n20685) );
  OAI211_X1 U23775 ( .C1(n20885), .C2(n20734), .A(n20686), .B(n20685), .ZN(
        P2_U3121) );
  AOI22_X1 U23776 ( .A1(n20711), .A2(n20835), .B1(n20886), .B2(n20710), .ZN(
        n20688) );
  AOI22_X1 U23777 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20702), .B1(
        n20887), .B2(n20701), .ZN(n20687) );
  OAI211_X1 U23778 ( .C1(n20754), .C2(n20705), .A(n20688), .B(n20687), .ZN(
        P2_U3122) );
  AOI22_X1 U23779 ( .A1(n20894), .A2(n20689), .B1(n20892), .B2(n20710), .ZN(
        n20691) );
  AOI22_X1 U23780 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20702), .B1(
        n20893), .B2(n20701), .ZN(n20690) );
  OAI211_X1 U23781 ( .C1(n20897), .C2(n20734), .A(n20691), .B(n20690), .ZN(
        P2_U3123) );
  AOI22_X1 U23782 ( .A1(n20711), .A2(n20843), .B1(n20710), .B2(n20898), .ZN(
        n20693) );
  AOI22_X1 U23783 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20702), .B1(
        n20899), .B2(n20701), .ZN(n20692) );
  OAI211_X1 U23784 ( .C1(n20760), .C2(n20705), .A(n20693), .B(n20692), .ZN(
        P2_U3124) );
  AOI22_X1 U23785 ( .A1(n20711), .A2(n20847), .B1(n20904), .B2(n20710), .ZN(
        n20695) );
  AOI22_X1 U23786 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20702), .B1(
        n20905), .B2(n20701), .ZN(n20694) );
  OAI211_X1 U23787 ( .C1(n20763), .C2(n20705), .A(n20695), .B(n20694), .ZN(
        P2_U3125) );
  OAI22_X1 U23788 ( .A1(n20705), .A2(n20766), .B1(n20697), .B2(n20696), .ZN(
        n20698) );
  INV_X1 U23789 ( .A(n20698), .ZN(n20700) );
  AOI22_X1 U23790 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20702), .B1(
        n20911), .B2(n20701), .ZN(n20699) );
  OAI211_X1 U23791 ( .C1(n20915), .C2(n20734), .A(n20700), .B(n20699), .ZN(
        P2_U3126) );
  AOI22_X1 U23792 ( .A1(n20711), .A2(n20856), .B1(n20916), .B2(n20710), .ZN(
        n20704) );
  AOI22_X1 U23793 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20702), .B1(
        n20918), .B2(n20701), .ZN(n20703) );
  OAI211_X1 U23794 ( .C1(n20773), .C2(n20705), .A(n20704), .B(n20703), .ZN(
        P2_U3127) );
  INV_X1 U23795 ( .A(n20706), .ZN(n20708) );
  NOR2_X1 U23796 ( .A1(n20820), .A2(n20740), .ZN(n20729) );
  OAI21_X1 U23797 ( .B1(n20709), .B2(n20729), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20707) );
  AOI22_X1 U23798 ( .A1(n20730), .A2(n20867), .B1(n20729), .B2(n20866), .ZN(
        n20716) );
  INV_X1 U23799 ( .A(n20709), .ZN(n20713) );
  AOI221_X1 U23800 ( .B1(n20711), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20735), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20710), .ZN(n20712) );
  AOI211_X1 U23801 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20713), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20712), .ZN(n20714) );
  OAI21_X1 U23802 ( .B1(n20714), .B2(n20729), .A(n20874), .ZN(n20731) );
  AOI22_X1 U23803 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20828), .ZN(n20715) );
  OAI211_X1 U23804 ( .C1(n20748), .C2(n20734), .A(n20716), .B(n20715), .ZN(
        P2_U3128) );
  AOI22_X1 U23805 ( .A1(n20730), .A2(n20881), .B1(n20729), .B2(n20880), .ZN(
        n20718) );
  AOI22_X1 U23806 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20832), .ZN(n20717) );
  OAI211_X1 U23807 ( .C1(n20751), .C2(n20734), .A(n20718), .B(n20717), .ZN(
        P2_U3129) );
  AOI22_X1 U23808 ( .A1(n20730), .A2(n20887), .B1(n20729), .B2(n20886), .ZN(
        n20720) );
  AOI22_X1 U23809 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20835), .ZN(n20719) );
  OAI211_X1 U23810 ( .C1(n20754), .C2(n20734), .A(n20720), .B(n20719), .ZN(
        P2_U3130) );
  AOI22_X1 U23811 ( .A1(n20730), .A2(n20893), .B1(n20729), .B2(n20892), .ZN(
        n20722) );
  AOI22_X1 U23812 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20839), .ZN(n20721) );
  OAI211_X1 U23813 ( .C1(n20757), .C2(n20734), .A(n20722), .B(n20721), .ZN(
        P2_U3131) );
  AOI22_X1 U23814 ( .A1(n20730), .A2(n20899), .B1(n20729), .B2(n20898), .ZN(
        n20724) );
  AOI22_X1 U23815 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20843), .ZN(n20723) );
  OAI211_X1 U23816 ( .C1(n20760), .C2(n20734), .A(n20724), .B(n20723), .ZN(
        P2_U3132) );
  AOI22_X1 U23817 ( .A1(n20730), .A2(n20905), .B1(n20729), .B2(n20904), .ZN(
        n20726) );
  AOI22_X1 U23818 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20847), .ZN(n20725) );
  OAI211_X1 U23819 ( .C1(n20763), .C2(n20734), .A(n20726), .B(n20725), .ZN(
        P2_U3133) );
  AOI22_X1 U23820 ( .A1(n20730), .A2(n20911), .B1(n20729), .B2(n20910), .ZN(
        n20728) );
  AOI22_X1 U23821 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20851), .ZN(n20727) );
  OAI211_X1 U23822 ( .C1(n20766), .C2(n20734), .A(n20728), .B(n20727), .ZN(
        P2_U3134) );
  AOI22_X1 U23823 ( .A1(n20730), .A2(n20918), .B1(n20729), .B2(n20916), .ZN(
        n20733) );
  AOI22_X1 U23824 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20731), .B1(
        n20735), .B2(n20856), .ZN(n20732) );
  OAI211_X1 U23825 ( .C1(n20773), .C2(n20734), .A(n20733), .B(n20732), .ZN(
        P2_U3135) );
  OR2_X1 U23826 ( .A1(n21050), .A2(n20740), .ZN(n20739) );
  INV_X1 U23827 ( .A(n20740), .ZN(n20736) );
  NAND2_X1 U23828 ( .A1(n20737), .A2(n20736), .ZN(n20742) );
  OAI21_X1 U23829 ( .B1(n12290), .B2(n20767), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20738) );
  OAI21_X1 U23830 ( .B1(n20739), .B2(n21065), .A(n20738), .ZN(n20768) );
  AOI22_X1 U23831 ( .A1(n20768), .A2(n20867), .B1(n20866), .B2(n20767), .ZN(
        n20747) );
  OAI22_X1 U23832 ( .A1(n20870), .A2(n20741), .B1(n20740), .B2(n21050), .ZN(
        n20745) );
  OAI211_X1 U23833 ( .C1(n20743), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n21065), 
        .B(n20742), .ZN(n20744) );
  NAND3_X1 U23834 ( .A1(n20745), .A2(n20874), .A3(n20744), .ZN(n20769) );
  AOI22_X1 U23835 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20828), .ZN(n20746) );
  OAI211_X1 U23836 ( .C1(n20748), .C2(n20772), .A(n20747), .B(n20746), .ZN(
        P2_U3136) );
  AOI22_X1 U23837 ( .A1(n20768), .A2(n20881), .B1(n20880), .B2(n20767), .ZN(
        n20750) );
  AOI22_X1 U23838 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20832), .ZN(n20749) );
  OAI211_X1 U23839 ( .C1(n20751), .C2(n20772), .A(n20750), .B(n20749), .ZN(
        P2_U3137) );
  AOI22_X1 U23840 ( .A1(n20768), .A2(n20887), .B1(n20886), .B2(n20767), .ZN(
        n20753) );
  AOI22_X1 U23841 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20835), .ZN(n20752) );
  OAI211_X1 U23842 ( .C1(n20754), .C2(n20772), .A(n20753), .B(n20752), .ZN(
        P2_U3138) );
  AOI22_X1 U23843 ( .A1(n20768), .A2(n20893), .B1(n20892), .B2(n20767), .ZN(
        n20756) );
  AOI22_X1 U23844 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20839), .ZN(n20755) );
  OAI211_X1 U23845 ( .C1(n20757), .C2(n20772), .A(n20756), .B(n20755), .ZN(
        P2_U3139) );
  AOI22_X1 U23846 ( .A1(n20768), .A2(n20899), .B1(n20898), .B2(n20767), .ZN(
        n20759) );
  AOI22_X1 U23847 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20843), .ZN(n20758) );
  OAI211_X1 U23848 ( .C1(n20760), .C2(n20772), .A(n20759), .B(n20758), .ZN(
        P2_U3140) );
  AOI22_X1 U23849 ( .A1(n20768), .A2(n20905), .B1(n20904), .B2(n20767), .ZN(
        n20762) );
  AOI22_X1 U23850 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20847), .ZN(n20761) );
  OAI211_X1 U23851 ( .C1(n20763), .C2(n20772), .A(n20762), .B(n20761), .ZN(
        P2_U3141) );
  AOI22_X1 U23852 ( .A1(n20768), .A2(n20911), .B1(n20910), .B2(n20767), .ZN(
        n20765) );
  AOI22_X1 U23853 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20851), .ZN(n20764) );
  OAI211_X1 U23854 ( .C1(n20766), .C2(n20772), .A(n20765), .B(n20764), .ZN(
        P2_U3142) );
  AOI22_X1 U23855 ( .A1(n20768), .A2(n20918), .B1(n20916), .B2(n20767), .ZN(
        n20771) );
  AOI22_X1 U23856 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20769), .B1(
        n20787), .B2(n20856), .ZN(n20770) );
  OAI211_X1 U23857 ( .C1(n20773), .C2(n20772), .A(n20771), .B(n20770), .ZN(
        P2_U3143) );
  AOI22_X1 U23858 ( .A1(n20786), .A2(n20881), .B1(n20785), .B2(n20880), .ZN(
        n20775) );
  AOI22_X1 U23859 ( .A1(n20787), .A2(n20882), .B1(n20808), .B2(n20832), .ZN(
        n20774) );
  OAI211_X1 U23860 ( .C1(n20790), .C2(n12216), .A(n20775), .B(n20774), .ZN(
        P2_U3145) );
  INV_X1 U23861 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23862 ( .A1(n20786), .A2(n20899), .B1(n20785), .B2(n20898), .ZN(
        n20777) );
  AOI22_X1 U23863 ( .A1(n20787), .A2(n20900), .B1(n20808), .B2(n20843), .ZN(
        n20776) );
  OAI211_X1 U23864 ( .C1(n20790), .C2(n20778), .A(n20777), .B(n20776), .ZN(
        P2_U3148) );
  INV_X1 U23865 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U23866 ( .A1(n20786), .A2(n20905), .B1(n20785), .B2(n20904), .ZN(
        n20780) );
  AOI22_X1 U23867 ( .A1(n20787), .A2(n20906), .B1(n20808), .B2(n20847), .ZN(
        n20779) );
  OAI211_X1 U23868 ( .C1(n20790), .C2(n20781), .A(n20780), .B(n20779), .ZN(
        P2_U3149) );
  INV_X1 U23869 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20784) );
  AOI22_X1 U23870 ( .A1(n20786), .A2(n20911), .B1(n20785), .B2(n20910), .ZN(
        n20783) );
  AOI22_X1 U23871 ( .A1(n20787), .A2(n20912), .B1(n20808), .B2(n20851), .ZN(
        n20782) );
  OAI211_X1 U23872 ( .C1(n20790), .C2(n20784), .A(n20783), .B(n20782), .ZN(
        P2_U3150) );
  AOI22_X1 U23873 ( .A1(n20786), .A2(n20918), .B1(n20785), .B2(n20916), .ZN(
        n20789) );
  AOI22_X1 U23874 ( .A1(n20787), .A2(n20920), .B1(n20808), .B2(n20856), .ZN(
        n20788) );
  OAI211_X1 U23875 ( .C1(n20790), .C2(n12354), .A(n20789), .B(n20788), .ZN(
        P2_U3151) );
  AOI22_X1 U23876 ( .A1(n20807), .A2(n20881), .B1(n20806), .B2(n20880), .ZN(
        n20792) );
  AOI22_X1 U23877 ( .A1(n20808), .A2(n20882), .B1(n20857), .B2(n20832), .ZN(
        n20791) );
  OAI211_X1 U23878 ( .C1(n20812), .C2(n12217), .A(n20792), .B(n20791), .ZN(
        P2_U3153) );
  INV_X1 U23879 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U23880 ( .A1(n20807), .A2(n20887), .B1(n20886), .B2(n20806), .ZN(
        n20794) );
  AOI22_X1 U23881 ( .A1(n20808), .A2(n20888), .B1(n20857), .B2(n20835), .ZN(
        n20793) );
  OAI211_X1 U23882 ( .C1(n20812), .C2(n20795), .A(n20794), .B(n20793), .ZN(
        P2_U3154) );
  INV_X1 U23883 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U23884 ( .A1(n20807), .A2(n20893), .B1(n20892), .B2(n20806), .ZN(
        n20797) );
  AOI22_X1 U23885 ( .A1(n20808), .A2(n20894), .B1(n20857), .B2(n20839), .ZN(
        n20796) );
  OAI211_X1 U23886 ( .C1(n20812), .C2(n20798), .A(n20797), .B(n20796), .ZN(
        P2_U3155) );
  INV_X1 U23887 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20801) );
  AOI22_X1 U23888 ( .A1(n20807), .A2(n20899), .B1(n20806), .B2(n20898), .ZN(
        n20800) );
  AOI22_X1 U23889 ( .A1(n20808), .A2(n20900), .B1(n20857), .B2(n20843), .ZN(
        n20799) );
  OAI211_X1 U23890 ( .C1(n20812), .C2(n20801), .A(n20800), .B(n20799), .ZN(
        P2_U3156) );
  AOI22_X1 U23891 ( .A1(n20807), .A2(n20905), .B1(n20806), .B2(n20904), .ZN(
        n20803) );
  AOI22_X1 U23892 ( .A1(n20808), .A2(n20906), .B1(n20857), .B2(n20847), .ZN(
        n20802) );
  OAI211_X1 U23893 ( .C1(n20812), .C2(n21707), .A(n20803), .B(n20802), .ZN(
        P2_U3157) );
  INV_X1 U23894 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n21652) );
  AOI22_X1 U23895 ( .A1(n20807), .A2(n20911), .B1(n20806), .B2(n20910), .ZN(
        n20805) );
  AOI22_X1 U23896 ( .A1(n20808), .A2(n20912), .B1(n20857), .B2(n20851), .ZN(
        n20804) );
  OAI211_X1 U23897 ( .C1(n20812), .C2(n21652), .A(n20805), .B(n20804), .ZN(
        P2_U3158) );
  INV_X1 U23898 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U23899 ( .A1(n20807), .A2(n20918), .B1(n20806), .B2(n20916), .ZN(
        n20810) );
  AOI22_X1 U23900 ( .A1(n20808), .A2(n20920), .B1(n20857), .B2(n20856), .ZN(
        n20809) );
  OAI211_X1 U23901 ( .C1(n20812), .C2(n20811), .A(n20810), .B(n20809), .ZN(
        P2_U3159) );
  INV_X1 U23902 ( .A(n20921), .ZN(n20816) );
  INV_X1 U23903 ( .A(n20857), .ZN(n20815) );
  AOI21_X1 U23904 ( .B1(n20816), .B2(n20815), .A(n20814), .ZN(n20817) );
  NOR2_X1 U23905 ( .A1(n20817), .A2(n21065), .ZN(n20824) );
  NAND2_X1 U23906 ( .A1(n20818), .A2(n20863), .ZN(n20826) );
  NOR2_X1 U23907 ( .A1(n20820), .A2(n20819), .ZN(n20855) );
  INV_X1 U23908 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U23909 ( .A1(n20876), .A2(n20857), .B1(n20866), .B2(n20855), .ZN(
        n20830) );
  INV_X1 U23910 ( .A(n20824), .ZN(n20827) );
  AOI22_X1 U23911 ( .A1(n20867), .A2(n20858), .B1(n20921), .B2(n20828), .ZN(
        n20829) );
  OAI211_X1 U23912 ( .C1(n20861), .C2(n20831), .A(n20830), .B(n20829), .ZN(
        P2_U3160) );
  AOI22_X1 U23913 ( .A1(n20921), .A2(n20832), .B1(n20855), .B2(n20880), .ZN(
        n20834) );
  AOI22_X1 U23914 ( .A1(n20881), .A2(n20858), .B1(n20857), .B2(n20882), .ZN(
        n20833) );
  OAI211_X1 U23915 ( .C1(n20861), .C2(n12204), .A(n20834), .B(n20833), .ZN(
        P2_U3161) );
  AOI22_X1 U23916 ( .A1(n20921), .A2(n20835), .B1(n20886), .B2(n20855), .ZN(
        n20837) );
  AOI22_X1 U23917 ( .A1(n20887), .A2(n20858), .B1(n20857), .B2(n20888), .ZN(
        n20836) );
  OAI211_X1 U23918 ( .C1(n20861), .C2(n20838), .A(n20837), .B(n20836), .ZN(
        P2_U3162) );
  INV_X1 U23919 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20842) );
  AOI22_X1 U23920 ( .A1(n20894), .A2(n20857), .B1(n20892), .B2(n20855), .ZN(
        n20841) );
  AOI22_X1 U23921 ( .A1(n20893), .A2(n20858), .B1(n20921), .B2(n20839), .ZN(
        n20840) );
  OAI211_X1 U23922 ( .C1(n20861), .C2(n20842), .A(n20841), .B(n20840), .ZN(
        P2_U3163) );
  INV_X1 U23923 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U23924 ( .A1(n20900), .A2(n20857), .B1(n20855), .B2(n20898), .ZN(
        n20845) );
  AOI22_X1 U23925 ( .A1(n20899), .A2(n20858), .B1(n20921), .B2(n20843), .ZN(
        n20844) );
  OAI211_X1 U23926 ( .C1(n20861), .C2(n20846), .A(n20845), .B(n20844), .ZN(
        P2_U3164) );
  INV_X1 U23927 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20850) );
  AOI22_X1 U23928 ( .A1(n20906), .A2(n20857), .B1(n20855), .B2(n20904), .ZN(
        n20849) );
  AOI22_X1 U23929 ( .A1(n20905), .A2(n20858), .B1(n20921), .B2(n20847), .ZN(
        n20848) );
  OAI211_X1 U23930 ( .C1(n20861), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        P2_U3165) );
  AOI22_X1 U23931 ( .A1(n20921), .A2(n20851), .B1(n20855), .B2(n20910), .ZN(
        n20853) );
  AOI22_X1 U23932 ( .A1(n20911), .A2(n20858), .B1(n20857), .B2(n20912), .ZN(
        n20852) );
  OAI211_X1 U23933 ( .C1(n20861), .C2(n20854), .A(n20853), .B(n20852), .ZN(
        P2_U3166) );
  AOI22_X1 U23934 ( .A1(n20921), .A2(n20856), .B1(n20855), .B2(n20916), .ZN(
        n20860) );
  AOI22_X1 U23935 ( .A1(n20918), .A2(n20858), .B1(n20857), .B2(n20920), .ZN(
        n20859) );
  OAI211_X1 U23936 ( .C1(n20861), .C2(n21637), .A(n20860), .B(n20859), .ZN(
        P2_U3167) );
  NAND2_X1 U23937 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20863), .ZN(
        n20868) );
  OAI21_X1 U23938 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20868), .A(n20864), 
        .ZN(n20865) );
  AOI22_X1 U23939 ( .A1(n20919), .A2(n20867), .B1(n20917), .B2(n20866), .ZN(
        n20878) );
  OAI21_X1 U23940 ( .B1(n20870), .B2(n20869), .A(n20868), .ZN(n20875) );
  NAND2_X1 U23941 ( .A1(n20871), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20872) );
  NAND4_X1 U23942 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20922) );
  AOI22_X1 U23943 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20876), .ZN(n20877) );
  OAI211_X1 U23944 ( .C1(n20879), .C2(n20925), .A(n20878), .B(n20877), .ZN(
        P2_U3168) );
  AOI22_X1 U23945 ( .A1(n20919), .A2(n20881), .B1(n20917), .B2(n20880), .ZN(
        n20884) );
  AOI22_X1 U23946 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20882), .ZN(n20883) );
  OAI211_X1 U23947 ( .C1(n20885), .C2(n20925), .A(n20884), .B(n20883), .ZN(
        P2_U3169) );
  AOI22_X1 U23948 ( .A1(n20919), .A2(n20887), .B1(n20917), .B2(n20886), .ZN(
        n20890) );
  AOI22_X1 U23949 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20888), .ZN(n20889) );
  OAI211_X1 U23950 ( .C1(n20891), .C2(n20925), .A(n20890), .B(n20889), .ZN(
        P2_U3170) );
  AOI22_X1 U23951 ( .A1(n20919), .A2(n20893), .B1(n20917), .B2(n20892), .ZN(
        n20896) );
  AOI22_X1 U23952 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20894), .ZN(n20895) );
  OAI211_X1 U23953 ( .C1(n20897), .C2(n20925), .A(n20896), .B(n20895), .ZN(
        P2_U3171) );
  AOI22_X1 U23954 ( .A1(n20919), .A2(n20899), .B1(n20917), .B2(n20898), .ZN(
        n20902) );
  AOI22_X1 U23955 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20900), .ZN(n20901) );
  OAI211_X1 U23956 ( .C1(n20903), .C2(n20925), .A(n20902), .B(n20901), .ZN(
        P2_U3172) );
  AOI22_X1 U23957 ( .A1(n20919), .A2(n20905), .B1(n20917), .B2(n20904), .ZN(
        n20908) );
  AOI22_X1 U23958 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20906), .ZN(n20907) );
  OAI211_X1 U23959 ( .C1(n20909), .C2(n20925), .A(n20908), .B(n20907), .ZN(
        P2_U3173) );
  AOI22_X1 U23960 ( .A1(n20919), .A2(n20911), .B1(n20917), .B2(n20910), .ZN(
        n20914) );
  AOI22_X1 U23961 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20912), .ZN(n20913) );
  OAI211_X1 U23962 ( .C1(n20915), .C2(n20925), .A(n20914), .B(n20913), .ZN(
        P2_U3174) );
  AOI22_X1 U23963 ( .A1(n20919), .A2(n20918), .B1(n20917), .B2(n20916), .ZN(
        n20924) );
  AOI22_X1 U23964 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20922), .B1(
        n20921), .B2(n20920), .ZN(n20923) );
  OAI211_X1 U23965 ( .C1(n20926), .C2(n20925), .A(n20924), .B(n20923), .ZN(
        P2_U3175) );
  NOR3_X1 U23966 ( .A1(n21071), .A2(n21075), .A3(n21025), .ZN(n20928) );
  OAI21_X1 U23967 ( .B1(n20929), .B2(n20928), .A(n20927), .ZN(n20934) );
  OAI21_X1 U23968 ( .B1(n20931), .B2(n20930), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n20932) );
  NAND3_X1 U23969 ( .A1(n20934), .A2(n20933), .A3(n20932), .ZN(P2_U3177) );
  AND2_X1 U23970 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20935), .ZN(
        P2_U3179) );
  AND2_X1 U23971 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20935), .ZN(
        P2_U3180) );
  AND2_X1 U23972 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20935), .ZN(
        P2_U3181) );
  AND2_X1 U23973 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20935), .ZN(
        P2_U3182) );
  AND2_X1 U23974 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20935), .ZN(
        P2_U3183) );
  AND2_X1 U23975 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20935), .ZN(
        P2_U3184) );
  AND2_X1 U23976 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20935), .ZN(
        P2_U3185) );
  NOR2_X1 U23977 ( .A1(n21623), .A2(n21016), .ZN(P2_U3186) );
  AND2_X1 U23978 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20935), .ZN(
        P2_U3187) );
  AND2_X1 U23979 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20935), .ZN(
        P2_U3188) );
  AND2_X1 U23980 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20935), .ZN(
        P2_U3189) );
  AND2_X1 U23981 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20935), .ZN(
        P2_U3190) );
  AND2_X1 U23982 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20935), .ZN(
        P2_U3191) );
  NOR2_X1 U23983 ( .A1(n21497), .A2(n21016), .ZN(P2_U3192) );
  AND2_X1 U23984 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20935), .ZN(
        P2_U3193) );
  AND2_X1 U23985 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20935), .ZN(
        P2_U3194) );
  AND2_X1 U23986 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20935), .ZN(
        P2_U3195) );
  AND2_X1 U23987 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20935), .ZN(
        P2_U3196) );
  AND2_X1 U23988 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20935), .ZN(
        P2_U3197) );
  AND2_X1 U23989 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20935), .ZN(
        P2_U3198) );
  AND2_X1 U23990 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20935), .ZN(
        P2_U3199) );
  AND2_X1 U23991 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20935), .ZN(
        P2_U3200) );
  AND2_X1 U23992 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20935), .ZN(P2_U3201) );
  AND2_X1 U23993 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20935), .ZN(P2_U3202) );
  AND2_X1 U23994 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20935), .ZN(P2_U3203) );
  AND2_X1 U23995 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20935), .ZN(P2_U3204) );
  AND2_X1 U23996 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20935), .ZN(P2_U3205) );
  AND2_X1 U23997 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20935), .ZN(P2_U3206) );
  AND2_X1 U23998 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20935), .ZN(P2_U3207) );
  AND2_X1 U23999 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20935), .ZN(P2_U3208) );
  NOR2_X1 U24000 ( .A1(n20936), .A2(n21073), .ZN(n20948) );
  INV_X1 U24001 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21475) );
  OR3_X1 U24002 ( .A1(n20948), .A2(n21475), .A3(n20937), .ZN(n20939) );
  AOI211_X1 U24003 ( .C1(n21355), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n20949), .B(n20999), .ZN(n20938) );
  INV_X1 U24004 ( .A(NA), .ZN(n21353) );
  NOR2_X1 U24005 ( .A1(n21353), .A2(n20941), .ZN(n20954) );
  AOI211_X1 U24006 ( .C1(n20955), .C2(n20939), .A(n20938), .B(n20954), .ZN(
        n20940) );
  INV_X1 U24007 ( .A(n20940), .ZN(P2_U3209) );
  AOI21_X1 U24008 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21355), .A(n20955), 
        .ZN(n20946) );
  NOR2_X1 U24009 ( .A1(n21475), .A2(n20946), .ZN(n20942) );
  AOI21_X1 U24010 ( .B1(n20942), .B2(n20941), .A(n20948), .ZN(n20944) );
  INV_X1 U24011 ( .A(n21076), .ZN(n20943) );
  OAI211_X1 U24012 ( .C1(n21355), .C2(n20945), .A(n20944), .B(n20943), .ZN(
        P2_U3210) );
  AOI21_X1 U24013 ( .B1(n21071), .B2(n20947), .A(n20946), .ZN(n20953) );
  AOI22_X1 U24014 ( .A1(n21475), .A2(n20949), .B1(n21353), .B2(n20948), .ZN(
        n20950) );
  INV_X1 U24015 ( .A(n20950), .ZN(n20951) );
  OAI211_X1 U24016 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20951), .ZN(n20952) );
  OAI21_X1 U24017 ( .B1(n20954), .B2(n20953), .A(n20952), .ZN(P2_U3211) );
  NAND2_X2 U24018 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20999), .ZN(n21006) );
  NAND2_X2 U24019 ( .A1(n20999), .A2(n20955), .ZN(n21007) );
  OAI222_X1 U24020 ( .A1(n21006), .A2(n20957), .B1(n20956), .B2(n20999), .C1(
        n20959), .C2(n21007), .ZN(P2_U3212) );
  OAI222_X1 U24021 ( .A1(n21006), .A2(n20959), .B1(n20958), .B2(n20999), .C1(
        n12152), .C2(n21007), .ZN(P2_U3213) );
  OAI222_X1 U24022 ( .A1(n21006), .A2(n12152), .B1(n21453), .B2(n20999), .C1(
        n12488), .C2(n21007), .ZN(P2_U3214) );
  OAI222_X1 U24023 ( .A1(n21007), .A2(n12494), .B1(n21678), .B2(n20999), .C1(
        n12488), .C2(n21006), .ZN(P2_U3215) );
  OAI222_X1 U24024 ( .A1(n21007), .A2(n20961), .B1(n20960), .B2(n20999), .C1(
        n12494), .C2(n21006), .ZN(P2_U3216) );
  OAI222_X1 U24025 ( .A1(n21007), .A2(n20963), .B1(n20962), .B2(n20999), .C1(
        n20961), .C2(n21006), .ZN(P2_U3217) );
  OAI222_X1 U24026 ( .A1(n21007), .A2(n17077), .B1(n20964), .B2(n20999), .C1(
        n20963), .C2(n21006), .ZN(P2_U3218) );
  OAI222_X1 U24027 ( .A1(n21007), .A2(n20966), .B1(n20965), .B2(n20999), .C1(
        n17077), .C2(n21006), .ZN(P2_U3219) );
  OAI222_X1 U24028 ( .A1(n21007), .A2(n20968), .B1(n20967), .B2(n20999), .C1(
        n20966), .C2(n21006), .ZN(P2_U3220) );
  OAI222_X1 U24029 ( .A1(n21007), .A2(n12707), .B1(n20969), .B2(n20999), .C1(
        n20968), .C2(n21006), .ZN(P2_U3221) );
  OAI222_X1 U24030 ( .A1(n21007), .A2(n12476), .B1(n20970), .B2(n20999), .C1(
        n12707), .C2(n21006), .ZN(P2_U3222) );
  OAI222_X1 U24031 ( .A1(n21007), .A2(n21471), .B1(n20971), .B2(n20999), .C1(
        n12476), .C2(n21006), .ZN(P2_U3223) );
  OAI222_X1 U24032 ( .A1(n21007), .A2(n20973), .B1(n20972), .B2(n20999), .C1(
        n21471), .C2(n21006), .ZN(P2_U3224) );
  OAI222_X1 U24033 ( .A1(n21007), .A2(n20975), .B1(n20974), .B2(n20999), .C1(
        n20973), .C2(n21006), .ZN(P2_U3225) );
  OAI222_X1 U24034 ( .A1(n21007), .A2(n20977), .B1(n20976), .B2(n20999), .C1(
        n20975), .C2(n21006), .ZN(P2_U3226) );
  OAI222_X1 U24035 ( .A1(n21007), .A2(n20979), .B1(n20978), .B2(n20999), .C1(
        n20977), .C2(n21006), .ZN(P2_U3227) );
  OAI222_X1 U24036 ( .A1(n21007), .A2(n20981), .B1(n20980), .B2(n20999), .C1(
        n20979), .C2(n21006), .ZN(P2_U3228) );
  OAI222_X1 U24037 ( .A1(n21007), .A2(n20983), .B1(n20982), .B2(n20999), .C1(
        n20981), .C2(n21006), .ZN(P2_U3229) );
  OAI222_X1 U24038 ( .A1(n21007), .A2(n20985), .B1(n20984), .B2(n20999), .C1(
        n20983), .C2(n21006), .ZN(P2_U3230) );
  OAI222_X1 U24039 ( .A1(n21007), .A2(n20987), .B1(n20986), .B2(n20999), .C1(
        n20985), .C2(n21006), .ZN(P2_U3231) );
  OAI222_X1 U24040 ( .A1(n21007), .A2(n20989), .B1(n20988), .B2(n20999), .C1(
        n20987), .C2(n21006), .ZN(P2_U3232) );
  OAI222_X1 U24041 ( .A1(n21007), .A2(n20991), .B1(n20990), .B2(n20999), .C1(
        n20989), .C2(n21006), .ZN(P2_U3233) );
  OAI222_X1 U24042 ( .A1(n21007), .A2(n20993), .B1(n20992), .B2(n20999), .C1(
        n20991), .C2(n21006), .ZN(P2_U3234) );
  OAI222_X1 U24043 ( .A1(n21007), .A2(n20995), .B1(n20994), .B2(n20999), .C1(
        n20993), .C2(n21006), .ZN(P2_U3235) );
  OAI222_X1 U24044 ( .A1(n21007), .A2(n20997), .B1(n20996), .B2(n20999), .C1(
        n20995), .C2(n21006), .ZN(P2_U3236) );
  OAI222_X1 U24045 ( .A1(n21007), .A2(n21001), .B1(n20998), .B2(n20999), .C1(
        n20997), .C2(n21006), .ZN(P2_U3237) );
  INV_X1 U24046 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n21002) );
  OAI222_X1 U24047 ( .A1(n21006), .A2(n21001), .B1(n21000), .B2(n20999), .C1(
        n21002), .C2(n21007), .ZN(P2_U3238) );
  OAI222_X1 U24048 ( .A1(n21007), .A2(n21004), .B1(n21003), .B2(n20999), .C1(
        n21002), .C2(n21006), .ZN(P2_U3239) );
  OAI222_X1 U24049 ( .A1(n21007), .A2(n15174), .B1(n21005), .B2(n20999), .C1(
        n21004), .C2(n21006), .ZN(P2_U3240) );
  OAI222_X1 U24050 ( .A1(n21007), .A2(n12800), .B1(n21716), .B2(n20999), .C1(
        n15174), .C2(n21006), .ZN(P2_U3241) );
  INV_X1 U24051 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n21008) );
  AOI22_X1 U24052 ( .A1(n20999), .A2(n21009), .B1(n21008), .B2(n21085), .ZN(
        P2_U3585) );
  MUX2_X1 U24053 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20999), .Z(P2_U3586) );
  INV_X1 U24054 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U24055 ( .A1(n20999), .A2(n21632), .B1(n21010), .B2(n21085), .ZN(
        P2_U3587) );
  INV_X1 U24056 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n21011) );
  AOI22_X1 U24057 ( .A1(n20999), .A2(n21012), .B1(n21011), .B2(n21085), .ZN(
        P2_U3588) );
  OAI21_X1 U24058 ( .B1(n21016), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21014), 
        .ZN(n21013) );
  INV_X1 U24059 ( .A(n21013), .ZN(P2_U3591) );
  OAI21_X1 U24060 ( .B1(n21016), .B2(n21015), .A(n21014), .ZN(P2_U3592) );
  INV_X1 U24061 ( .A(n21017), .ZN(n21019) );
  OAI222_X1 U24062 ( .A1(n21036), .A2(n21021), .B1(n21020), .B2(n21019), .C1(
        n21025), .C2(n21018), .ZN(n21023) );
  MUX2_X1 U24063 ( .A(n21023), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n21022), .Z(P2_U3599) );
  NAND2_X1 U24064 ( .A1(n21024), .A2(n21045), .ZN(n21033) );
  NAND3_X1 U24065 ( .A1(n21043), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n21025), 
        .ZN(n21026) );
  NAND2_X1 U24066 ( .A1(n21026), .A2(n21040), .ZN(n21035) );
  NAND2_X1 U24067 ( .A1(n21033), .A2(n21035), .ZN(n21031) );
  AOI222_X1 U24068 ( .A1(n21031), .A2(n21030), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n21029), .C1(n21028), .C2(n21027), .ZN(n21032) );
  AOI22_X1 U24069 ( .A1(n21051), .A2(n21494), .B1(n21032), .B2(n21048), .ZN(
        P2_U3602) );
  INV_X1 U24070 ( .A(n21033), .ZN(n21038) );
  OAI22_X1 U24071 ( .A1(n21036), .A2(n21035), .B1(n21034), .B2(n20821), .ZN(
        n21037) );
  NOR2_X1 U24072 ( .A1(n21038), .A2(n21037), .ZN(n21039) );
  AOI22_X1 U24073 ( .A1(n21051), .A2(n21692), .B1(n21039), .B2(n21048), .ZN(
        P2_U3603) );
  INV_X1 U24074 ( .A(n21040), .ZN(n21042) );
  NOR2_X1 U24075 ( .A1(n21042), .A2(n21041), .ZN(n21044) );
  MUX2_X1 U24076 ( .A(n21045), .B(n21044), .S(n21043), .Z(n21046) );
  AOI21_X1 U24077 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n21047), .A(n21046), 
        .ZN(n21049) );
  AOI22_X1 U24078 ( .A1(n21051), .A2(n21050), .B1(n21049), .B2(n21048), .ZN(
        P2_U3604) );
  INV_X1 U24079 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n21052) );
  AOI22_X1 U24080 ( .A1(n20999), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n21052), 
        .B2(n21085), .ZN(P2_U3608) );
  INV_X1 U24081 ( .A(n21053), .ZN(n21062) );
  INV_X1 U24082 ( .A(n21054), .ZN(n21060) );
  INV_X1 U24083 ( .A(n21055), .ZN(n21058) );
  OAI21_X1 U24084 ( .B1(n21058), .B2(n21057), .A(n21056), .ZN(n21059) );
  OAI211_X1 U24085 ( .C1(n21062), .C2(n21061), .A(n21060), .B(n21059), .ZN(
        n21064) );
  MUX2_X1 U24086 ( .A(P2_MORE_REG_SCAN_IN), .B(n21064), .S(n21063), .Z(
        P2_U3609) );
  OAI21_X1 U24087 ( .B1(n21066), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n21065), 
        .ZN(n21067) );
  INV_X1 U24088 ( .A(n21067), .ZN(n21068) );
  OAI211_X1 U24089 ( .C1(n21071), .C2(n21070), .A(n21069), .B(n21068), .ZN(
        n21084) );
  AOI21_X1 U24090 ( .B1(n21073), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n21072), 
        .ZN(n21082) );
  AOI21_X1 U24091 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n21076), .A(n21074), 
        .ZN(n21080) );
  NOR3_X1 U24092 ( .A1(n21077), .A2(n21076), .A3(n21075), .ZN(n21079) );
  MUX2_X1 U24093 ( .A(n21080), .B(n21079), .S(n21078), .Z(n21081) );
  OAI21_X1 U24094 ( .B1(n21082), .B2(n21081), .A(n21084), .ZN(n21083) );
  OAI21_X1 U24095 ( .B1(n21084), .B2(n21475), .A(n21083), .ZN(P2_U3610) );
  INV_X1 U24096 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n21086) );
  AOI22_X1 U24097 ( .A1(n20999), .A2(n21087), .B1(n21086), .B2(n21085), .ZN(
        P2_U3611) );
  AOI21_X1 U24098 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21357), .A(n21345), 
        .ZN(n21348) );
  INV_X1 U24099 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21491) );
  NOR2_X4 U24100 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21341), .ZN(n21438) );
  AOI21_X1 U24101 ( .B1(n21348), .B2(n21491), .A(n21438), .ZN(P1_U2802) );
  INV_X1 U24102 ( .A(n21088), .ZN(n21090) );
  OAI21_X1 U24103 ( .B1(n21090), .B2(n21089), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n21091) );
  OAI21_X1 U24104 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21092), .A(n21091), 
        .ZN(P1_U2803) );
  NOR2_X1 U24105 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21349) );
  OAI21_X1 U24106 ( .B1(n21349), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21425), .ZN(
        n21093) );
  OAI21_X1 U24107 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21425), .A(n21093), 
        .ZN(P1_U2804) );
  OAI21_X1 U24108 ( .B1(BS16), .B2(n21349), .A(n21339), .ZN(n21413) );
  OAI21_X1 U24109 ( .B1(n21339), .B2(n21428), .A(n21413), .ZN(P1_U2805) );
  OAI21_X1 U24110 ( .B1(n21096), .B2(n21095), .A(n21094), .ZN(P1_U2806) );
  NOR2_X1 U24111 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21551) );
  AOI211_X1 U24112 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_3__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21097) );
  INV_X1 U24113 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n21338) );
  INV_X1 U24114 ( .A(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21645) );
  NAND4_X1 U24115 ( .A1(n21551), .A2(n21097), .A3(n21338), .A4(n21645), .ZN(
        n21105) );
  OR4_X1 U24116 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21104) );
  OR4_X1 U24117 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21103) );
  NOR4_X1 U24118 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n21101) );
  NOR4_X1 U24119 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21100) );
  NOR4_X1 U24120 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21099) );
  NOR4_X1 U24121 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21098) );
  NAND4_X1 U24122 ( .A1(n21101), .A2(n21100), .A3(n21099), .A4(n21098), .ZN(
        n21102) );
  NOR4_X2 U24123 ( .A1(n21105), .A2(n21104), .A3(n21103), .A4(n21102), .ZN(
        n21424) );
  INV_X1 U24124 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21411) );
  NOR3_X1 U24125 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n21107) );
  OAI21_X1 U24126 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n21107), .A(n21424), .ZN(
        n21106) );
  OAI21_X1 U24127 ( .B1(n21424), .B2(n21411), .A(n21106), .ZN(P1_U2807) );
  NAND2_X1 U24128 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21424), .ZN(n21420) );
  NOR2_X1 U24129 ( .A1(n21107), .A2(n21420), .ZN(n21109) );
  NOR2_X1 U24130 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(n21424), .ZN(n21108)
         );
  AOI211_X1 U24131 ( .C1(n21424), .C2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21109), 
        .B(n21108), .ZN(P1_U2808) );
  AOI22_X1 U24132 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n21182), .B1(n21176), .B2(
        n21110), .ZN(n21114) );
  NOR3_X1 U24133 ( .A1(n21173), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n21111), .ZN(
        n21112) );
  AOI211_X1 U24134 ( .C1(n21174), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n21163), .B(n21112), .ZN(n21113) );
  OAI211_X1 U24135 ( .C1(n21115), .C2(n21137), .A(n21114), .B(n21113), .ZN(
        n21116) );
  INV_X1 U24136 ( .A(n21116), .ZN(n21120) );
  AOI22_X1 U24137 ( .A1(n21118), .A2(n21185), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n21117), .ZN(n21119) );
  NAND2_X1 U24138 ( .A1(n21120), .A2(n21119), .ZN(P1_U2831) );
  OAI21_X1 U24139 ( .B1(n21149), .B2(n21121), .A(n21147), .ZN(n21125) );
  OAI22_X1 U24140 ( .A1(n21123), .A2(n21170), .B1(n21646), .B2(n21122), .ZN(
        n21124) );
  AOI211_X1 U24141 ( .C1(n21176), .C2(n21126), .A(n21125), .B(n21124), .ZN(
        n21133) );
  OR2_X1 U24142 ( .A1(n21127), .A2(n21129), .ZN(n21145) );
  OAI21_X1 U24143 ( .B1(n21129), .B2(n21128), .A(n21145), .ZN(n21140) );
  AOI22_X1 U24144 ( .A1(n21131), .A2(n21130), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n21140), .ZN(n21132) );
  OAI211_X1 U24145 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n21134), .A(n21133), .B(
        n21132), .ZN(P1_U2833) );
  AOI21_X1 U24146 ( .B1(n21174), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21163), .ZN(n21144) );
  AOI22_X1 U24147 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(n21182), .B1(n21176), .B2(
        n21135), .ZN(n21143) );
  OAI22_X1 U24148 ( .A1(n21138), .A2(n21137), .B1(n21136), .B2(n21170), .ZN(
        n21139) );
  AOI21_X1 U24149 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n21140), .A(n21139), .ZN(
        n21142) );
  NAND3_X1 U24150 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n21151), .A3(n21367), 
        .ZN(n21141) );
  NAND4_X1 U24151 ( .A1(n21144), .A2(n21143), .A3(n21142), .A4(n21141), .ZN(
        P1_U2834) );
  INV_X1 U24152 ( .A(n21145), .ZN(n21166) );
  AOI22_X1 U24153 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n21182), .B1(n21176), .B2(
        n21146), .ZN(n21148) );
  OAI211_X1 U24154 ( .C1(n21149), .C2(n21695), .A(n21148), .B(n21147), .ZN(
        n21150) );
  AOI221_X1 U24155 ( .B1(n21166), .B2(P1_REIP_REG_5__SCAN_IN), .C1(n21151), 
        .C2(n21584), .A(n21150), .ZN(n21155) );
  INV_X1 U24156 ( .A(n21152), .ZN(n21153) );
  NAND2_X1 U24157 ( .A1(n21187), .A2(n21153), .ZN(n21154) );
  OAI211_X1 U24158 ( .C1(n21170), .C2(n21156), .A(n21155), .B(n21154), .ZN(
        P1_U2835) );
  INV_X1 U24159 ( .A(n21178), .ZN(n21157) );
  AOI22_X1 U24160 ( .A1(n21158), .A2(n21157), .B1(n21182), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n21159) );
  OAI21_X1 U24161 ( .B1(n21161), .B2(n21160), .A(n21159), .ZN(n21162) );
  AOI211_X1 U24162 ( .C1(n21174), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21163), .B(n21162), .ZN(n21169) );
  OAI21_X1 U24163 ( .B1(n21173), .B2(n21164), .A(n21363), .ZN(n21165) );
  AOI22_X1 U24164 ( .A1(n21187), .A2(n21167), .B1(n21166), .B2(n21165), .ZN(
        n21168) );
  OAI211_X1 U24165 ( .C1(n21171), .C2(n21170), .A(n21169), .B(n21168), .ZN(
        P1_U2836) );
  NOR3_X1 U24166 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21173), .A3(n21172), .ZN(
        n21181) );
  AOI22_X1 U24167 ( .A1(n21176), .A2(n21175), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n21174), .ZN(n21177) );
  OAI21_X1 U24168 ( .B1(n21179), .B2(n21178), .A(n21177), .ZN(n21180) );
  AOI211_X1 U24169 ( .C1(n21182), .C2(P1_EBX_REG_3__SCAN_IN), .A(n21181), .B(
        n21180), .ZN(n21189) );
  INV_X1 U24170 ( .A(n21183), .ZN(n21184) );
  AOI22_X1 U24171 ( .A1(n21187), .A2(n21186), .B1(n21185), .B2(n21184), .ZN(
        n21188) );
  OAI211_X1 U24172 ( .C1(n21190), .C2(n13982), .A(n21189), .B(n21188), .ZN(
        P1_U2837) );
  INV_X1 U24173 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n21445) );
  INV_X1 U24174 ( .A(n21191), .ZN(n21193) );
  AOI22_X1 U24175 ( .A1(n13845), .A2(P1_DATAO_REG_20__SCAN_IN), .B1(n21193), 
        .B2(P1_EAX_REG_20__SCAN_IN), .ZN(n21192) );
  OAI21_X1 U24176 ( .B1(n21445), .B2(n21218), .A(n21192), .ZN(P1_U2916) );
  INV_X1 U24177 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n21684) );
  AOI22_X1 U24178 ( .A1(n21193), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n21435), .ZN(n21194) );
  OAI21_X1 U24179 ( .B1(n21684), .B2(n21221), .A(n21194), .ZN(P1_U2918) );
  AOI22_X1 U24180 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n21206), .B1(n13845), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n21195) );
  OAI21_X1 U24181 ( .B1(n21196), .B2(n21218), .A(n21195), .ZN(P1_U2921) );
  INV_X1 U24182 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21198) );
  AOI22_X1 U24183 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n21197) );
  OAI21_X1 U24184 ( .B1(n21198), .B2(n21220), .A(n21197), .ZN(P1_U2922) );
  INV_X1 U24185 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21200) );
  AOI22_X1 U24186 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n21199) );
  OAI21_X1 U24187 ( .B1(n21200), .B2(n21220), .A(n21199), .ZN(P1_U2923) );
  INV_X1 U24188 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21202) );
  AOI22_X1 U24189 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n21201) );
  OAI21_X1 U24190 ( .B1(n21202), .B2(n21220), .A(n21201), .ZN(P1_U2924) );
  AOI22_X1 U24191 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n21203) );
  OAI21_X1 U24192 ( .B1(n15631), .B2(n21220), .A(n21203), .ZN(P1_U2925) );
  INV_X1 U24193 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21205) );
  AOI22_X1 U24194 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n21204) );
  OAI21_X1 U24195 ( .B1(n21205), .B2(n21220), .A(n21204), .ZN(P1_U2926) );
  AOI22_X1 U24196 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n21206), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n21435), .ZN(n21207) );
  OAI21_X1 U24197 ( .B1(n21572), .B2(n21221), .A(n21207), .ZN(P1_U2927) );
  AOI22_X1 U24198 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n21208) );
  OAI21_X1 U24199 ( .B1(n15641), .B2(n21220), .A(n21208), .ZN(P1_U2928) );
  AOI22_X1 U24200 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n21209) );
  OAI21_X1 U24201 ( .B1(n11237), .B2(n21220), .A(n21209), .ZN(P1_U2929) );
  AOI22_X1 U24202 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n21210) );
  OAI21_X1 U24203 ( .B1(n11229), .B2(n21220), .A(n21210), .ZN(P1_U2930) );
  AOI22_X1 U24204 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n21211) );
  OAI21_X1 U24205 ( .B1(n11222), .B2(n21220), .A(n21211), .ZN(P1_U2931) );
  AOI22_X1 U24206 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n21212) );
  OAI21_X1 U24207 ( .B1(n21213), .B2(n21220), .A(n21212), .ZN(P1_U2932) );
  AOI22_X1 U24208 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n21214) );
  OAI21_X1 U24209 ( .B1(n11200), .B2(n21220), .A(n21214), .ZN(P1_U2933) );
  AOI22_X1 U24210 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21435), .B1(n13845), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n21215) );
  OAI21_X1 U24211 ( .B1(n11173), .B2(n21220), .A(n21215), .ZN(P1_U2934) );
  INV_X1 U24212 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n21636) );
  OAI222_X1 U24213 ( .A1(n21218), .A2(n21636), .B1(n21220), .B2(n21217), .C1(
        n21221), .C2(n21216), .ZN(P1_U2935) );
  INV_X1 U24214 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n21729) );
  INV_X1 U24215 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n21517) );
  OAI222_X1 U24216 ( .A1(n21221), .A2(n21729), .B1(n21220), .B2(n21219), .C1(
        n21218), .C2(n21517), .ZN(P1_U2936) );
  AOI22_X1 U24217 ( .A1(n21246), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n21245), .ZN(n21223) );
  NAND2_X1 U24218 ( .A1(n21231), .A2(n21222), .ZN(n21233) );
  NAND2_X1 U24219 ( .A1(n21223), .A2(n21233), .ZN(P1_U2945) );
  AOI22_X1 U24220 ( .A1(n21246), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n21225) );
  NAND2_X1 U24221 ( .A1(n21231), .A2(n21224), .ZN(n21239) );
  NAND2_X1 U24222 ( .A1(n21225), .A2(n21239), .ZN(P1_U2948) );
  AOI22_X1 U24223 ( .A1(n21246), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n21227) );
  NAND2_X1 U24224 ( .A1(n21231), .A2(n21226), .ZN(n21241) );
  NAND2_X1 U24225 ( .A1(n21227), .A2(n21241), .ZN(P1_U2949) );
  AOI22_X1 U24226 ( .A1(n21246), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n21229) );
  NAND2_X1 U24227 ( .A1(n21231), .A2(n21228), .ZN(n21243) );
  NAND2_X1 U24228 ( .A1(n21229), .A2(n21243), .ZN(P1_U2950) );
  AOI22_X1 U24229 ( .A1(n21246), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n21245), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n21232) );
  NAND2_X1 U24230 ( .A1(n21231), .A2(n21230), .ZN(n21247) );
  NAND2_X1 U24231 ( .A1(n21232), .A2(n21247), .ZN(P1_U2951) );
  AOI22_X1 U24232 ( .A1(n21246), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n21234) );
  NAND2_X1 U24233 ( .A1(n21234), .A2(n21233), .ZN(P1_U2960) );
  AOI22_X1 U24234 ( .A1(n21246), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n21245), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n21236) );
  NAND2_X1 U24235 ( .A1(n21236), .A2(n21235), .ZN(P1_U2961) );
  AOI22_X1 U24236 ( .A1(n21246), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n21245), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n21238) );
  NAND2_X1 U24237 ( .A1(n21238), .A2(n21237), .ZN(P1_U2962) );
  AOI22_X1 U24238 ( .A1(n21246), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n21245), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n21240) );
  NAND2_X1 U24239 ( .A1(n21240), .A2(n21239), .ZN(P1_U2963) );
  AOI22_X1 U24240 ( .A1(n21246), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n21245), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n21242) );
  NAND2_X1 U24241 ( .A1(n21242), .A2(n21241), .ZN(P1_U2964) );
  AOI22_X1 U24242 ( .A1(n21246), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n21245), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n21244) );
  NAND2_X1 U24243 ( .A1(n21244), .A2(n21243), .ZN(P1_U2965) );
  AOI22_X1 U24244 ( .A1(n21246), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n21245), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n21248) );
  NAND2_X1 U24245 ( .A1(n21248), .A2(n21247), .ZN(P1_U2966) );
  AOI22_X1 U24246 ( .A1(n21252), .A2(n21251), .B1(n21250), .B2(n21249), .ZN(
        n21257) );
  OAI22_X1 U24247 ( .A1(n21255), .A2(n21254), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21253), .ZN(n21256) );
  OAI211_X1 U24248 ( .C1(n13791), .C2(n17669), .A(n21257), .B(n21256), .ZN(
        P1_U3031) );
  AND2_X1 U24249 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21258), .ZN(
        P1_U3032) );
  INV_X1 U24250 ( .A(n21259), .ZN(n21264) );
  AOI22_X1 U24251 ( .A1(n21295), .A2(n21265), .B1(n21294), .B2(n21264), .ZN(
        n21261) );
  AOI22_X1 U24252 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n21266), .B2(n21296), .ZN(n21260) );
  OAI211_X1 U24253 ( .C1(n21299), .C2(n21270), .A(n21261), .B(n21260), .ZN(
        P1_U3107) );
  AOI22_X1 U24254 ( .A1(n21313), .A2(n21265), .B1(n21312), .B2(n21264), .ZN(
        n21263) );
  AOI22_X1 U24255 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n21266), .B2(n21314), .ZN(n21262) );
  OAI211_X1 U24256 ( .C1(n21317), .C2(n21270), .A(n21263), .B(n21262), .ZN(
        P1_U3110) );
  AOI22_X1 U24257 ( .A1(n21327), .A2(n21265), .B1(n21325), .B2(n21264), .ZN(
        n21269) );
  AOI22_X1 U24258 ( .A1(n21267), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n21266), .B2(n21328), .ZN(n21268) );
  OAI211_X1 U24259 ( .C1(n21334), .C2(n21270), .A(n21269), .B(n21268), .ZN(
        P1_U3112) );
  NOR2_X1 U24260 ( .A1(n21271), .A2(n21273), .ZN(n21326) );
  INV_X1 U24261 ( .A(n21272), .ZN(n21277) );
  INV_X1 U24262 ( .A(n21273), .ZN(n21282) );
  AOI22_X1 U24263 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21282), .B1(n21326), 
        .B2(n21274), .ZN(n21275) );
  AOI22_X1 U24264 ( .A1(n21279), .A2(n21326), .B1(n21278), .B2(n21324), .ZN(
        n21286) );
  AND2_X1 U24265 ( .A1(n21280), .A2(n14159), .ZN(n21283) );
  AOI22_X1 U24266 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n21329), .B2(n21284), .ZN(n21285) );
  OAI211_X1 U24267 ( .C1(n21287), .C2(n21333), .A(n21286), .B(n21285), .ZN(
        P1_U3137) );
  AOI22_X1 U24268 ( .A1(n21289), .A2(n21326), .B1(n21288), .B2(n21324), .ZN(
        n21292) );
  AOI22_X1 U24269 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n21329), .B2(n21290), .ZN(n21291) );
  OAI211_X1 U24270 ( .C1(n21293), .C2(n21333), .A(n21292), .B(n21291), .ZN(
        P1_U3138) );
  AOI22_X1 U24271 ( .A1(n21295), .A2(n21326), .B1(n21294), .B2(n21324), .ZN(
        n21298) );
  AOI22_X1 U24272 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n21329), .B2(n21296), .ZN(n21297) );
  OAI211_X1 U24273 ( .C1(n21299), .C2(n21333), .A(n21298), .B(n21297), .ZN(
        P1_U3139) );
  AOI22_X1 U24274 ( .A1(n21301), .A2(n21326), .B1(n21300), .B2(n21324), .ZN(
        n21304) );
  AOI22_X1 U24275 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n21329), .B2(n21302), .ZN(n21303) );
  OAI211_X1 U24276 ( .C1(n21305), .C2(n21333), .A(n21304), .B(n21303), .ZN(
        P1_U3140) );
  AOI22_X1 U24277 ( .A1(n21307), .A2(n21326), .B1(n21306), .B2(n21324), .ZN(
        n21310) );
  AOI22_X1 U24278 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n21329), .B2(n21308), .ZN(n21309) );
  OAI211_X1 U24279 ( .C1(n21311), .C2(n21333), .A(n21310), .B(n21309), .ZN(
        P1_U3141) );
  AOI22_X1 U24280 ( .A1(n21313), .A2(n21326), .B1(n21312), .B2(n21324), .ZN(
        n21316) );
  AOI22_X1 U24281 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n21329), .B2(n21314), .ZN(n21315) );
  OAI211_X1 U24282 ( .C1(n21317), .C2(n21333), .A(n21316), .B(n21315), .ZN(
        P1_U3142) );
  AOI22_X1 U24283 ( .A1(n21319), .A2(n21326), .B1(n21318), .B2(n21324), .ZN(
        n21322) );
  AOI22_X1 U24284 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n21329), .B2(n21320), .ZN(n21321) );
  OAI211_X1 U24285 ( .C1(n21323), .C2(n21333), .A(n21322), .B(n21321), .ZN(
        P1_U3143) );
  AOI22_X1 U24286 ( .A1(n21327), .A2(n21326), .B1(n21325), .B2(n21324), .ZN(
        n21332) );
  AOI22_X1 U24287 ( .A1(n21330), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n21329), .B2(n21328), .ZN(n21331) );
  OAI211_X1 U24288 ( .C1(n21334), .C2(n21333), .A(n21332), .B(n21331), .ZN(
        P1_U3144) );
  NOR2_X1 U24289 ( .A1(n21654), .A2(n21335), .ZN(n21337) );
  OAI21_X1 U24290 ( .B1(n21337), .B2(n14687), .A(n21336), .ZN(P1_U3163) );
  AND2_X1 U24291 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21416), .ZN(
        P1_U3164) );
  AND2_X1 U24292 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21416), .ZN(
        P1_U3165) );
  AND2_X1 U24293 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21416), .ZN(
        P1_U3166) );
  AND2_X1 U24294 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21416), .ZN(
        P1_U3167) );
  AND2_X1 U24295 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21416), .ZN(
        P1_U3168) );
  AND2_X1 U24296 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21416), .ZN(
        P1_U3169) );
  AND2_X1 U24297 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21416), .ZN(
        P1_U3170) );
  AND2_X1 U24298 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21416), .ZN(
        P1_U3171) );
  AND2_X1 U24299 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21416), .ZN(
        P1_U3172) );
  AND2_X1 U24300 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21416), .ZN(
        P1_U3173) );
  INV_X1 U24301 ( .A(P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21473) );
  NOR2_X1 U24302 ( .A1(n21339), .A2(n21473), .ZN(P1_U3174) );
  AND2_X1 U24303 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21416), .ZN(
        P1_U3175) );
  INV_X1 U24304 ( .A(P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21458) );
  NOR2_X1 U24305 ( .A1(n21339), .A2(n21458), .ZN(P1_U3176) );
  AND2_X1 U24306 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21416), .ZN(
        P1_U3177) );
  AND2_X1 U24307 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21416), .ZN(
        P1_U3178) );
  AND2_X1 U24308 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21416), .ZN(
        P1_U3179) );
  NOR2_X1 U24309 ( .A1(n21339), .A2(n21645), .ZN(P1_U3180) );
  AND2_X1 U24310 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21416), .ZN(
        P1_U3181) );
  AND2_X1 U24311 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21416), .ZN(
        P1_U3182) );
  AND2_X1 U24312 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21416), .ZN(
        P1_U3183) );
  AND2_X1 U24313 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21416), .ZN(
        P1_U3184) );
  AND2_X1 U24314 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21416), .ZN(
        P1_U3185) );
  AND2_X1 U24315 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21416), .ZN(P1_U3186) );
  AND2_X1 U24316 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21416), .ZN(P1_U3187) );
  AND2_X1 U24317 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21416), .ZN(P1_U3188) );
  AND2_X1 U24318 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21416), .ZN(P1_U3189) );
  AND2_X1 U24319 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21416), .ZN(P1_U3190) );
  AND2_X1 U24320 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21416), .ZN(P1_U3191) );
  AND2_X1 U24321 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21416), .ZN(P1_U3192) );
  NOR2_X1 U24322 ( .A1(n21339), .A2(n21338), .ZN(P1_U3193) );
  AOI21_X1 U24323 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21340), .A(n21345), 
        .ZN(n21350) );
  NAND2_X1 U24324 ( .A1(n21341), .A2(n21357), .ZN(n21343) );
  NAND2_X1 U24325 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(n21353), .ZN(
        n21351) );
  AOI22_X1 U24326 ( .A1(HOLD), .A2(n21343), .B1(n21342), .B2(n21351), .ZN(
        n21344) );
  OAI22_X1 U24327 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21350), .B1(n21438), 
        .B2(n21344), .ZN(P1_U3194) );
  NOR3_X1 U24328 ( .A1(NA), .A2(n21345), .A3(n21434), .ZN(n21347) );
  INV_X1 U24329 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21346) );
  OAI22_X1 U24330 ( .A1(n21348), .A2(n21347), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21346), .ZN(n21356) );
  AOI211_X1 U24331 ( .C1(n21357), .C2(n21351), .A(n21350), .B(n21349), .ZN(
        n21352) );
  OAI21_X1 U24332 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21353), .A(n21352), 
        .ZN(n21354) );
  OAI21_X1 U24333 ( .B1(n21356), .B2(n21355), .A(n21354), .ZN(P1_U3196) );
  NAND2_X2 U24334 ( .A1(n21438), .A2(n21357), .ZN(n21408) );
  INV_X1 U24335 ( .A(n21402), .ZN(n21406) );
  INV_X1 U24336 ( .A(n21406), .ZN(n21405) );
  OAI222_X1 U24337 ( .A1(n21408), .A2(n21361), .B1(n21359), .B2(n21438), .C1(
        n21358), .C2(n21405), .ZN(P1_U3197) );
  INV_X1 U24338 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21360) );
  OAI222_X1 U24339 ( .A1(n21402), .A2(n21361), .B1(n21360), .B2(n21438), .C1(
        n13982), .C2(n21408), .ZN(P1_U3198) );
  INV_X1 U24340 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21362) );
  OAI222_X1 U24341 ( .A1(n21405), .A2(n13982), .B1(n21362), .B2(n21438), .C1(
        n21363), .C2(n21408), .ZN(P1_U3199) );
  INV_X1 U24342 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21364) );
  OAI222_X1 U24343 ( .A1(n21408), .A2(n21584), .B1(n21364), .B2(n21438), .C1(
        n21363), .C2(n21405), .ZN(P1_U3200) );
  INV_X1 U24344 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21365) );
  OAI222_X1 U24345 ( .A1(n21408), .A2(n21367), .B1(n21365), .B2(n21438), .C1(
        n21584), .C2(n21405), .ZN(P1_U3201) );
  INV_X1 U24346 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21366) );
  OAI222_X1 U24347 ( .A1(n21402), .A2(n21367), .B1(n21366), .B2(n21438), .C1(
        n21369), .C2(n21408), .ZN(P1_U3202) );
  INV_X1 U24348 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21368) );
  OAI222_X1 U24349 ( .A1(n21402), .A2(n21369), .B1(n21368), .B2(n21438), .C1(
        n21564), .C2(n21408), .ZN(P1_U3203) );
  INV_X1 U24350 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21370) );
  OAI222_X1 U24351 ( .A1(n21402), .A2(n21564), .B1(n21370), .B2(n21438), .C1(
        n21372), .C2(n21408), .ZN(P1_U3204) );
  INV_X1 U24352 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21371) );
  INV_X1 U24353 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21374) );
  OAI222_X1 U24354 ( .A1(n21402), .A2(n21372), .B1(n21371), .B2(n21438), .C1(
        n21374), .C2(n21408), .ZN(P1_U3205) );
  INV_X1 U24355 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21373) );
  OAI222_X1 U24356 ( .A1(n21405), .A2(n21374), .B1(n21373), .B2(n21438), .C1(
        n21665), .C2(n21408), .ZN(P1_U3206) );
  INV_X1 U24357 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21375) );
  OAI222_X1 U24358 ( .A1(n21405), .A2(n21665), .B1(n21375), .B2(n21438), .C1(
        n21706), .C2(n21408), .ZN(P1_U3207) );
  INV_X1 U24359 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21376) );
  OAI222_X1 U24360 ( .A1(n21408), .A2(n21378), .B1(n21376), .B2(n21438), .C1(
        n21706), .C2(n21405), .ZN(P1_U3208) );
  INV_X1 U24361 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21377) );
  OAI222_X1 U24362 ( .A1(n21402), .A2(n21378), .B1(n21377), .B2(n21438), .C1(
        n21379), .C2(n21408), .ZN(P1_U3209) );
  INV_X1 U24363 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21380) );
  OAI222_X1 U24364 ( .A1(n21408), .A2(n21381), .B1(n21380), .B2(n21438), .C1(
        n21379), .C2(n21405), .ZN(P1_U3210) );
  INV_X1 U24365 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21468) );
  OAI222_X1 U24366 ( .A1(n21402), .A2(n21381), .B1(n21468), .B2(n21438), .C1(
        n21382), .C2(n21408), .ZN(P1_U3211) );
  INV_X1 U24367 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21527) );
  OAI222_X1 U24368 ( .A1(n21402), .A2(n21382), .B1(n21527), .B2(n21438), .C1(
        n21383), .C2(n21408), .ZN(P1_U3212) );
  INV_X1 U24369 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21384) );
  OAI222_X1 U24370 ( .A1(n21408), .A2(n21386), .B1(n21384), .B2(n21438), .C1(
        n21383), .C2(n21405), .ZN(P1_U3213) );
  AOI22_X1 U24371 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21425), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21403), .ZN(n21385) );
  OAI21_X1 U24372 ( .B1(n21386), .B2(n21405), .A(n21385), .ZN(P1_U3214) );
  INV_X1 U24373 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21389) );
  AOI22_X1 U24374 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21425), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21406), .ZN(n21387) );
  OAI21_X1 U24375 ( .B1(n21389), .B2(n21408), .A(n21387), .ZN(P1_U3215) );
  INV_X1 U24376 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21388) );
  OAI222_X1 U24377 ( .A1(n21402), .A2(n21389), .B1(n21388), .B2(n21438), .C1(
        n21391), .C2(n21408), .ZN(P1_U3216) );
  INV_X1 U24378 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21390) );
  OAI222_X1 U24379 ( .A1(n21402), .A2(n21391), .B1(n21390), .B2(n21438), .C1(
        n21393), .C2(n21408), .ZN(P1_U3217) );
  AOI22_X1 U24380 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21425), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21403), .ZN(n21392) );
  OAI21_X1 U24381 ( .B1(n21393), .B2(n21405), .A(n21392), .ZN(P1_U3218) );
  INV_X1 U24382 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21395) );
  AOI22_X1 U24383 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21425), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21406), .ZN(n21394) );
  OAI21_X1 U24384 ( .B1(n21395), .B2(n21408), .A(n21394), .ZN(P1_U3219) );
  INV_X1 U24385 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21586) );
  INV_X1 U24386 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21573) );
  OAI222_X1 U24387 ( .A1(n21405), .A2(n21395), .B1(n21586), .B2(n21438), .C1(
        n21573), .C2(n21408), .ZN(P1_U3220) );
  AOI22_X1 U24388 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21403), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21425), .ZN(n21396) );
  OAI21_X1 U24389 ( .B1(n21573), .B2(n21405), .A(n21396), .ZN(P1_U3221) );
  AOI22_X1 U24390 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n21406), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21425), .ZN(n21397) );
  OAI21_X1 U24391 ( .B1(n21399), .B2(n21408), .A(n21397), .ZN(P1_U3222) );
  INV_X1 U24392 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21398) );
  OAI222_X1 U24393 ( .A1(n21405), .A2(n21399), .B1(n21398), .B2(n21438), .C1(
        n21401), .C2(n21408), .ZN(P1_U3223) );
  INV_X1 U24394 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21400) );
  OAI222_X1 U24395 ( .A1(n21402), .A2(n21401), .B1(n21400), .B2(n21438), .C1(
        n21668), .C2(n21408), .ZN(P1_U3224) );
  AOI22_X1 U24396 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21403), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21425), .ZN(n21404) );
  OAI21_X1 U24397 ( .B1(n21668), .B2(n21405), .A(n21404), .ZN(P1_U3225) );
  AOI22_X1 U24398 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n21406), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21425), .ZN(n21407) );
  OAI21_X1 U24399 ( .B1(n21409), .B2(n21408), .A(n21407), .ZN(P1_U3226) );
  MUX2_X1 U24400 ( .A(P1_BE_N_REG_3__SCAN_IN), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n21438), .Z(P1_U3458) );
  MUX2_X1 U24401 ( .A(P1_BE_N_REG_2__SCAN_IN), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .S(n21438), .Z(P1_U3459) );
  INV_X1 U24402 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21410) );
  AOI22_X1 U24403 ( .A1(n21438), .A2(n21411), .B1(n21410), .B2(n21425), .ZN(
        P1_U3460) );
  INV_X1 U24404 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21422) );
  INV_X1 U24405 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21412) );
  AOI22_X1 U24406 ( .A1(n21438), .A2(n21422), .B1(n21412), .B2(n21425), .ZN(
        P1_U3461) );
  INV_X1 U24407 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21414) );
  INV_X1 U24408 ( .A(n21413), .ZN(n21415) );
  AOI21_X1 U24409 ( .B1(n21414), .B2(n21416), .A(n21415), .ZN(P1_U3464) );
  AOI21_X1 U24410 ( .B1(n21416), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21415), 
        .ZN(n21417) );
  INV_X1 U24411 ( .A(n21417), .ZN(P1_U3465) );
  AOI211_X1 U24412 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21418) );
  INV_X1 U24413 ( .A(n21424), .ZN(n21421) );
  AOI22_X1 U24414 ( .A1(n21424), .A2(n21418), .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n21421), .ZN(n21419) );
  OAI21_X1 U24415 ( .B1(n13791), .B2(n21420), .A(n21419), .ZN(P1_U3481) );
  NOR2_X1 U24416 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21423) );
  AOI22_X1 U24417 ( .A1(n21424), .A2(n21423), .B1(n21422), .B2(n21421), .ZN(
        P1_U3482) );
  AOI22_X1 U24418 ( .A1(n21438), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21426), 
        .B2(n21425), .ZN(P1_U3483) );
  AOI211_X1 U24419 ( .C1(n11047), .C2(n21428), .A(n14687), .B(n21427), .ZN(
        n21431) );
  NOR3_X1 U24420 ( .A1(n21431), .A2(n21430), .A3(n21429), .ZN(n21437) );
  AOI211_X1 U24421 ( .C1(n21435), .C2(n21434), .A(n21433), .B(n21432), .ZN(
        n21436) );
  MUX2_X1 U24422 ( .A(n21437), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21436), 
        .Z(P1_U3485) );
  MUX2_X1 U24423 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21438), .Z(P1_U3486) );
  INV_X1 U24424 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21440) );
  AOI22_X1 U24425 ( .A1(n21549), .A2(keyinput14), .B1(n21440), .B2(keyinput18), 
        .ZN(n21439) );
  OAI221_X1 U24426 ( .B1(n21549), .B2(keyinput14), .C1(n21440), .C2(keyinput18), .A(n21439), .ZN(n21450) );
  INV_X1 U24427 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21442) );
  AOI22_X1 U24428 ( .A1(n21443), .A2(keyinput109), .B1(keyinput37), .B2(n21442), .ZN(n21441) );
  OAI221_X1 U24429 ( .B1(n21443), .B2(keyinput109), .C1(n21442), .C2(
        keyinput37), .A(n21441), .ZN(n21449) );
  AOI22_X1 U24430 ( .A1(n21445), .A2(keyinput48), .B1(n21555), .B2(keyinput67), 
        .ZN(n21444) );
  OAI221_X1 U24431 ( .B1(n21445), .B2(keyinput48), .C1(n21555), .C2(keyinput67), .A(n21444), .ZN(n21448) );
  AOI22_X1 U24432 ( .A1(n18333), .A2(keyinput117), .B1(n21548), .B2(keyinput44), .ZN(n21446) );
  OAI221_X1 U24433 ( .B1(n18333), .B2(keyinput117), .C1(n21548), .C2(
        keyinput44), .A(n21446), .ZN(n21447) );
  NOR4_X1 U24434 ( .A1(n21450), .A2(n21449), .A3(n21448), .A4(n21447), .ZN(
        n21746) );
  NAND2_X1 U24435 ( .A1(n21452), .A2(keyinput32), .ZN(n21451) );
  OAI221_X1 U24436 ( .B1(n21453), .B2(keyinput85), .C1(n21452), .C2(keyinput32), .A(n21451), .ZN(n21465) );
  AOI22_X1 U24437 ( .A1(n21456), .A2(keyinput59), .B1(keyinput111), .B2(n21455), .ZN(n21454) );
  OAI221_X1 U24438 ( .B1(n21456), .B2(keyinput59), .C1(n21455), .C2(
        keyinput111), .A(n21454), .ZN(n21464) );
  INV_X1 U24439 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21550) );
  AOI22_X1 U24440 ( .A1(n21458), .A2(keyinput66), .B1(n21550), .B2(keyinput58), 
        .ZN(n21457) );
  OAI221_X1 U24441 ( .B1(n21458), .B2(keyinput66), .C1(n21550), .C2(keyinput58), .A(n21457), .ZN(n21463) );
  AOI22_X1 U24442 ( .A1(n21461), .A2(keyinput124), .B1(keyinput30), .B2(n21460), .ZN(n21459) );
  OAI221_X1 U24443 ( .B1(n21461), .B2(keyinput124), .C1(n21460), .C2(
        keyinput30), .A(n21459), .ZN(n21462) );
  NOR4_X1 U24444 ( .A1(n21465), .A2(n21464), .A3(n21463), .A4(n21462), .ZN(
        n21745) );
  AOI22_X1 U24445 ( .A1(n21468), .A2(keyinput51), .B1(n21467), .B2(keyinput63), 
        .ZN(n21466) );
  OAI221_X1 U24446 ( .B1(n21468), .B2(keyinput51), .C1(n21467), .C2(keyinput63), .A(n21466), .ZN(n21545) );
  AOI22_X1 U24447 ( .A1(n21471), .A2(keyinput15), .B1(keyinput11), .B2(n21470), 
        .ZN(n21469) );
  OAI221_X1 U24448 ( .B1(n21471), .B2(keyinput15), .C1(n21470), .C2(keyinput11), .A(n21469), .ZN(n21544) );
  OAI22_X1 U24449 ( .A1(n13611), .A2(keyinput36), .B1(n21473), .B2(keyinput1), 
        .ZN(n21472) );
  AOI221_X1 U24450 ( .B1(n13611), .B2(keyinput36), .C1(keyinput1), .C2(n21473), 
        .A(n21472), .ZN(n21487) );
  OAI22_X1 U24451 ( .A1(n21554), .A2(keyinput13), .B1(n21475), .B2(keyinput101), .ZN(n21474) );
  AOI221_X1 U24452 ( .B1(n21554), .B2(keyinput13), .C1(keyinput101), .C2(
        n21475), .A(n21474), .ZN(n21486) );
  AOI22_X1 U24453 ( .A1(n21565), .A2(keyinput82), .B1(n21567), .B2(keyinput19), 
        .ZN(n21476) );
  OAI221_X1 U24454 ( .B1(n21565), .B2(keyinput82), .C1(n21567), .C2(keyinput19), .A(n21476), .ZN(n21484) );
  AOI22_X1 U24455 ( .A1(n21566), .A2(keyinput16), .B1(n13190), .B2(keyinput25), 
        .ZN(n21477) );
  OAI221_X1 U24456 ( .B1(n21566), .B2(keyinput16), .C1(n13190), .C2(keyinput25), .A(n21477), .ZN(n21483) );
  XNOR2_X1 U24457 ( .A(n21563), .B(keyinput8), .ZN(n21482) );
  XOR2_X1 U24458 ( .A(n21564), .B(keyinput69), .Z(n21480) );
  XNOR2_X1 U24459 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B(keyinput65), .ZN(
        n21479) );
  XNOR2_X1 U24460 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B(keyinput74), .ZN(
        n21478) );
  NAND3_X1 U24461 ( .A1(n21480), .A2(n21479), .A3(n21478), .ZN(n21481) );
  NOR4_X1 U24462 ( .A1(n21484), .A2(n21483), .A3(n21482), .A4(n21481), .ZN(
        n21485) );
  NAND3_X1 U24463 ( .A1(n21487), .A2(n21486), .A3(n21485), .ZN(n21543) );
  INV_X1 U24464 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n21489) );
  AOI22_X1 U24465 ( .A1(n21489), .A2(keyinput72), .B1(n12850), .B2(keyinput23), 
        .ZN(n21488) );
  OAI221_X1 U24466 ( .B1(n21489), .B2(keyinput72), .C1(n12850), .C2(keyinput23), .A(n21488), .ZN(n21501) );
  INV_X1 U24467 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21574) );
  AOI22_X1 U24468 ( .A1(n21491), .A2(keyinput113), .B1(n21574), .B2(keyinput96), .ZN(n21490) );
  OAI221_X1 U24469 ( .B1(n21491), .B2(keyinput113), .C1(n21574), .C2(
        keyinput96), .A(n21490), .ZN(n21500) );
  INV_X1 U24470 ( .A(DATAI_27_), .ZN(n21493) );
  AOI22_X1 U24471 ( .A1(n21494), .A2(keyinput89), .B1(keyinput99), .B2(n21493), 
        .ZN(n21492) );
  OAI221_X1 U24472 ( .B1(n21494), .B2(keyinput89), .C1(n21493), .C2(keyinput99), .A(n21492), .ZN(n21499) );
  AOI22_X1 U24473 ( .A1(n21497), .A2(keyinput81), .B1(keyinput123), .B2(n21496), .ZN(n21495) );
  OAI221_X1 U24474 ( .B1(n21497), .B2(keyinput81), .C1(n21496), .C2(
        keyinput123), .A(n21495), .ZN(n21498) );
  NOR4_X1 U24475 ( .A1(n21501), .A2(n21500), .A3(n21499), .A4(n21498), .ZN(
        n21541) );
  AOI22_X1 U24476 ( .A1(n21573), .A2(keyinput83), .B1(keyinput2), .B2(n21572), 
        .ZN(n21502) );
  OAI221_X1 U24477 ( .B1(n21573), .B2(keyinput83), .C1(n21572), .C2(keyinput2), 
        .A(n21502), .ZN(n21513) );
  AOI22_X1 U24478 ( .A1(n21576), .A2(keyinput88), .B1(keyinput22), .B2(n21504), 
        .ZN(n21503) );
  OAI221_X1 U24479 ( .B1(n21576), .B2(keyinput88), .C1(n21504), .C2(keyinput22), .A(n21503), .ZN(n21512) );
  AOI22_X1 U24480 ( .A1(n21507), .A2(keyinput10), .B1(keyinput75), .B2(n21506), 
        .ZN(n21505) );
  OAI221_X1 U24481 ( .B1(n21507), .B2(keyinput10), .C1(n21506), .C2(keyinput75), .A(n21505), .ZN(n21511) );
  XNOR2_X1 U24482 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B(keyinput78), .ZN(
        n21509) );
  XNOR2_X1 U24483 ( .A(keyinput94), .B(P2_EBX_REG_1__SCAN_IN), .ZN(n21508) );
  NAND2_X1 U24484 ( .A1(n21509), .A2(n21508), .ZN(n21510) );
  NOR4_X1 U24485 ( .A1(n21513), .A2(n21512), .A3(n21511), .A4(n21510), .ZN(
        n21540) );
  INV_X1 U24486 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21585) );
  AOI22_X1 U24487 ( .A1(n21569), .A2(keyinput107), .B1(n21585), .B2(keyinput24), .ZN(n21514) );
  OAI221_X1 U24488 ( .B1(n21569), .B2(keyinput107), .C1(n21585), .C2(
        keyinput24), .A(n21514), .ZN(n21523) );
  AOI22_X1 U24489 ( .A1(n21568), .A2(keyinput4), .B1(n14687), .B2(keyinput28), 
        .ZN(n21515) );
  OAI221_X1 U24490 ( .B1(n21568), .B2(keyinput4), .C1(n14687), .C2(keyinput28), 
        .A(n21515), .ZN(n21522) );
  AOI22_X1 U24491 ( .A1(n21517), .A2(keyinput115), .B1(n21584), .B2(keyinput40), .ZN(n21516) );
  OAI221_X1 U24492 ( .B1(n21517), .B2(keyinput115), .C1(n21584), .C2(
        keyinput40), .A(n21516), .ZN(n21521) );
  AOI22_X1 U24493 ( .A1(n21519), .A2(keyinput46), .B1(n21586), .B2(keyinput34), 
        .ZN(n21518) );
  OAI221_X1 U24494 ( .B1(n21519), .B2(keyinput46), .C1(n21586), .C2(keyinput34), .A(n21518), .ZN(n21520) );
  NOR4_X1 U24495 ( .A1(n21523), .A2(n21522), .A3(n21521), .A4(n21520), .ZN(
        n21539) );
  INV_X1 U24496 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21525) );
  AOI22_X1 U24497 ( .A1(n21570), .A2(keyinput62), .B1(n21525), .B2(keyinput100), .ZN(n21524) );
  OAI221_X1 U24498 ( .B1(n21570), .B2(keyinput62), .C1(n21525), .C2(
        keyinput100), .A(n21524), .ZN(n21537) );
  AOI22_X1 U24499 ( .A1(n21528), .A2(keyinput112), .B1(n21527), .B2(keyinput98), .ZN(n21526) );
  OAI221_X1 U24500 ( .B1(n21528), .B2(keyinput112), .C1(n21527), .C2(
        keyinput98), .A(n21526), .ZN(n21536) );
  INV_X1 U24501 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21571) );
  AOI22_X1 U24502 ( .A1(n21571), .A2(keyinput121), .B1(keyinput47), .B2(n21530), .ZN(n21529) );
  OAI221_X1 U24503 ( .B1(n21571), .B2(keyinput121), .C1(n21530), .C2(
        keyinput47), .A(n21529), .ZN(n21535) );
  AOI22_X1 U24504 ( .A1(n21533), .A2(keyinput35), .B1(keyinput97), .B2(n21532), 
        .ZN(n21531) );
  OAI221_X1 U24505 ( .B1(n21533), .B2(keyinput35), .C1(n21532), .C2(keyinput97), .A(n21531), .ZN(n21534) );
  NOR4_X1 U24506 ( .A1(n21537), .A2(n21536), .A3(n21535), .A4(n21534), .ZN(
        n21538) );
  NAND4_X1 U24507 ( .A1(n21541), .A2(n21540), .A3(n21539), .A4(n21538), .ZN(
        n21542) );
  NOR4_X1 U24508 ( .A1(n21545), .A2(n21544), .A3(n21543), .A4(n21542), .ZN(
        n21744) );
  NAND4_X1 U24509 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_EBX_REG_11__SCAN_IN), .A3(P3_REIP_REG_5__SCAN_IN), .A4(
        P3_ADDRESS_REG_8__SCAN_IN), .ZN(n21546) );
  NOR4_X1 U24510 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(n21547), .A4(n21546), .ZN(n21562)
         );
  NOR4_X1 U24511 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__6__SCAN_IN), .A3(P1_UWORD_REG_4__SCAN_IN), .A4(
        n21548), .ZN(n21561) );
  NOR4_X1 U24512 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__0__SCAN_IN), .A3(n21550), .A4(n21549), .ZN(n21560)
         );
  NAND4_X1 U24513 ( .A1(n21553), .A2(n21552), .A3(n21551), .A4(n21731), .ZN(
        n21558) );
  NOR4_X1 U24514 ( .A1(BUF1_REG_9__SCAN_IN), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .A3(n21555), .A4(n21554), .ZN(n21556) );
  NAND3_X1 U24515 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(n21556), .ZN(n21557) );
  NOR4_X1 U24516 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(BUF2_REG_20__SCAN_IN), 
        .A3(n21558), .A4(n21557), .ZN(n21559) );
  NAND4_X1 U24517 ( .A1(n21562), .A2(n21561), .A3(n21560), .A4(n21559), .ZN(
        n21615) );
  NOR4_X1 U24518 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .A3(n21564), .A4(n21563), .ZN(n21613) );
  NOR4_X1 U24519 ( .A1(n21567), .A2(n13190), .A3(n21566), .A4(n21565), .ZN(
        n21612) );
  NAND4_X1 U24520 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P2_CODEFETCH_REG_SCAN_IN), .A3(n21569), .A4(n21568), .ZN(n21583) );
  NAND4_X1 U24521 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(
        P3_LWORD_REG_6__SCAN_IN), .A3(n21571), .A4(n21570), .ZN(n21582) );
  NOR4_X1 U24522 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21573), .A4(n21572), .ZN(n21580) );
  NOR4_X1 U24523 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_18__SCAN_IN), .A3(n12850), .A4(n21574), .ZN(n21579)
         );
  NOR4_X1 U24524 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(DATAI_27_), .A3(
        P3_ADDRESS_REG_2__SCAN_IN), .A4(P3_DATAO_REG_23__SCAN_IN), .ZN(n21578)
         );
  NOR4_X1 U24525 ( .A1(n21576), .A2(n21575), .A3(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .A4(P3_DATAO_REG_24__SCAN_IN), .ZN(
        n21577) );
  NAND4_X1 U24526 ( .A1(n21580), .A2(n21579), .A3(n21578), .A4(n21577), .ZN(
        n21581) );
  NOR3_X1 U24527 ( .A1(n21583), .A2(n21582), .A3(n21581), .ZN(n21611) );
  NAND4_X1 U24528 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(
        P3_EAX_REG_21__SCAN_IN), .A3(n21621), .A4(n21584), .ZN(n21609) );
  NAND4_X1 U24529 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P1_LWORD_REG_0__SCAN_IN), .A3(n21586), .A4(n21585), .ZN(n21608) );
  INV_X1 U24530 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n21649) );
  NAND4_X1 U24531 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(n21652), .A4(n21649), .ZN(n21590)
         );
  INV_X1 U24532 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21639) );
  NAND4_X1 U24533 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_7__6__SCAN_IN), .A3(P1_LWORD_REG_1__SCAN_IN), .A4(
        n21639), .ZN(n21589) );
  NAND4_X1 U24534 ( .A1(DATAI_31_), .A2(P1_REIP_REG_11__SCAN_IN), .A3(
        P2_DATAO_REG_12__SCAN_IN), .A4(n15610), .ZN(n21588) );
  NAND4_X1 U24535 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(BUF1_REG_5__SCAN_IN), 
        .A3(n21651), .A4(n16815), .ZN(n21587) );
  NOR4_X1 U24536 ( .A1(n21590), .A2(n21589), .A3(n21588), .A4(n21587), .ZN(
        n21593) );
  NOR4_X1 U24537 ( .A1(DATAI_8_), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .A3(
        n11410), .A4(n21637), .ZN(n21592) );
  NOR4_X1 U24538 ( .A1(n14111), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A3(
        P2_REIP_REG_8__SCAN_IN), .A4(P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21591) );
  NAND3_X1 U24539 ( .A1(n21593), .A2(n21592), .A3(n21591), .ZN(n21607) );
  NAND4_X1 U24540 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        BUF1_REG_17__SCAN_IN), .A3(P1_DATAO_REG_0__SCAN_IN), .A4(n21728), .ZN(
        n21594) );
  NOR3_X1 U24541 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21722), .A3(
        n21594), .ZN(n21605) );
  NOR4_X1 U24542 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAO_REG_31__SCAN_IN), .A4(
        n11013), .ZN(n21595) );
  NAND3_X1 U24543 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_12__0__SCAN_IN), .A3(n21595), .ZN(n21603) );
  NOR4_X1 U24544 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(
        P2_ADDRESS_REG_3__SCAN_IN), .A3(n15243), .A4(n21684), .ZN(n21601) );
  NAND4_X1 U24545 ( .A1(n21596), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21599) );
  NOR4_X1 U24546 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P1_REIP_REG_29__SCAN_IN), .A3(BUF1_REG_3__SCAN_IN), .A4(n21681), .ZN(
        n21597) );
  NAND3_X1 U24547 ( .A1(n21698), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        n21597), .ZN(n21598) );
  NOR4_X1 U24548 ( .A1(n21599), .A2(n21598), .A3(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(P2_EAX_REG_31__SCAN_IN), .ZN(
        n21600) );
  NAND2_X1 U24549 ( .A1(n21601), .A2(n21600), .ZN(n21602) );
  NOR4_X1 U24550 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P1_REIP_REG_12__SCAN_IN), .A3(n21603), .A4(n21602), .ZN(n21604) );
  NAND4_X1 U24551 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n21605), .A3(n21604), 
        .A4(n21715), .ZN(n21606) );
  NOR4_X1 U24552 ( .A1(n21609), .A2(n21608), .A3(n21607), .A4(n21606), .ZN(
        n21610) );
  NAND4_X1 U24553 ( .A1(n21613), .A2(n21612), .A3(n21611), .A4(n21610), .ZN(
        n21614) );
  OAI21_X1 U24554 ( .B1(n21615), .B2(n21614), .A(P2_ADDRESS_REG_2__SCAN_IN), 
        .ZN(n21742) );
  INV_X1 U24555 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21617) );
  AOI22_X1 U24556 ( .A1(n21617), .A2(keyinput87), .B1(keyinput90), .B2(n11410), 
        .ZN(n21616) );
  OAI221_X1 U24557 ( .B1(n21617), .B2(keyinput87), .C1(n11410), .C2(keyinput90), .A(n21616), .ZN(n21629) );
  AOI22_X1 U24558 ( .A1(n21619), .A2(keyinput33), .B1(n17077), .B2(keyinput6), 
        .ZN(n21618) );
  OAI221_X1 U24559 ( .B1(n21619), .B2(keyinput33), .C1(n17077), .C2(keyinput6), 
        .A(n21618), .ZN(n21628) );
  AOI22_X1 U24560 ( .A1(n21622), .A2(keyinput77), .B1(n21621), .B2(keyinput93), 
        .ZN(n21620) );
  OAI221_X1 U24561 ( .B1(n21622), .B2(keyinput77), .C1(n21621), .C2(keyinput93), .A(n21620), .ZN(n21627) );
  XOR2_X1 U24562 ( .A(n21623), .B(keyinput71), .Z(n21625) );
  XNOR2_X1 U24563 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput119), 
        .ZN(n21624) );
  NAND2_X1 U24564 ( .A1(n21625), .A2(n21624), .ZN(n21626) );
  NOR4_X1 U24565 ( .A1(n21629), .A2(n21628), .A3(n21627), .A4(n21626), .ZN(
        n21676) );
  AOI22_X1 U24566 ( .A1(n21632), .A2(keyinput20), .B1(n21631), .B2(keyinput21), 
        .ZN(n21630) );
  OAI221_X1 U24567 ( .B1(n21632), .B2(keyinput20), .C1(n21631), .C2(keyinput21), .A(n21630), .ZN(n21643) );
  AOI22_X1 U24568 ( .A1(n21634), .A2(keyinput122), .B1(n12394), .B2(keyinput91), .ZN(n21633) );
  OAI221_X1 U24569 ( .B1(n21634), .B2(keyinput122), .C1(n12394), .C2(
        keyinput91), .A(n21633), .ZN(n21642) );
  AOI22_X1 U24570 ( .A1(n21637), .A2(keyinput56), .B1(keyinput102), .B2(n21636), .ZN(n21635) );
  OAI221_X1 U24571 ( .B1(n21637), .B2(keyinput56), .C1(n21636), .C2(
        keyinput102), .A(n21635), .ZN(n21641) );
  AOI22_X1 U24572 ( .A1(n21639), .A2(keyinput61), .B1(keyinput0), .B2(n18387), 
        .ZN(n21638) );
  OAI221_X1 U24573 ( .B1(n21639), .B2(keyinput61), .C1(n18387), .C2(keyinput0), 
        .A(n21638), .ZN(n21640) );
  NOR4_X1 U24574 ( .A1(n21643), .A2(n21642), .A3(n21641), .A4(n21640), .ZN(
        n21675) );
  AOI22_X1 U24575 ( .A1(n21646), .A2(keyinput80), .B1(keyinput92), .B2(n21645), 
        .ZN(n21644) );
  OAI221_X1 U24576 ( .B1(n21646), .B2(keyinput80), .C1(n21645), .C2(keyinput92), .A(n21644), .ZN(n21658) );
  AOI22_X1 U24577 ( .A1(n21649), .A2(keyinput73), .B1(n21648), .B2(keyinput64), 
        .ZN(n21647) );
  OAI221_X1 U24578 ( .B1(n21649), .B2(keyinput73), .C1(n21648), .C2(keyinput64), .A(n21647), .ZN(n21657) );
  AOI22_X1 U24579 ( .A1(n21652), .A2(keyinput108), .B1(keyinput53), .B2(n21651), .ZN(n21650) );
  OAI221_X1 U24580 ( .B1(n21652), .B2(keyinput108), .C1(n21651), .C2(
        keyinput53), .A(n21650), .ZN(n21656) );
  AOI22_X1 U24581 ( .A1(n21654), .A2(keyinput9), .B1(keyinput42), .B2(n16815), 
        .ZN(n21653) );
  OAI221_X1 U24582 ( .B1(n21654), .B2(keyinput9), .C1(n16815), .C2(keyinput42), 
        .A(n21653), .ZN(n21655) );
  NOR4_X1 U24583 ( .A1(n21658), .A2(n21657), .A3(n21656), .A4(n21655), .ZN(
        n21674) );
  AOI22_X1 U24584 ( .A1(n21661), .A2(keyinput3), .B1(keyinput54), .B2(n21660), 
        .ZN(n21659) );
  OAI221_X1 U24585 ( .B1(n21661), .B2(keyinput3), .C1(n21660), .C2(keyinput54), 
        .A(n21659), .ZN(n21672) );
  INV_X1 U24586 ( .A(DATAI_31_), .ZN(n21663) );
  AOI22_X1 U24587 ( .A1(n15610), .A2(keyinput95), .B1(keyinput5), .B2(n21663), 
        .ZN(n21662) );
  OAI221_X1 U24588 ( .B1(n15610), .B2(keyinput95), .C1(n21663), .C2(keyinput5), 
        .A(n21662), .ZN(n21671) );
  AOI22_X1 U24589 ( .A1(n21665), .A2(keyinput31), .B1(keyinput114), .B2(n13579), .ZN(n21664) );
  OAI221_X1 U24590 ( .B1(n21665), .B2(keyinput31), .C1(n13579), .C2(
        keyinput114), .A(n21664), .ZN(n21670) );
  INV_X1 U24591 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21667) );
  AOI22_X1 U24592 ( .A1(n21668), .A2(keyinput49), .B1(n21667), .B2(keyinput116), .ZN(n21666) );
  OAI221_X1 U24593 ( .B1(n21668), .B2(keyinput49), .C1(n21667), .C2(
        keyinput116), .A(n21666), .ZN(n21669) );
  NOR4_X1 U24594 ( .A1(n21672), .A2(n21671), .A3(n21670), .A4(n21669), .ZN(
        n21673) );
  NAND4_X1 U24595 ( .A1(n21676), .A2(n21675), .A3(n21674), .A4(n21673), .ZN(
        n21741) );
  AOI22_X1 U24596 ( .A1(n15243), .A2(keyinput39), .B1(n21678), .B2(keyinput29), 
        .ZN(n21677) );
  OAI221_X1 U24597 ( .B1(n15243), .B2(keyinput39), .C1(n21678), .C2(keyinput29), .A(n21677), .ZN(n21690) );
  INV_X1 U24598 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21680) );
  AOI22_X1 U24599 ( .A1(n21681), .A2(keyinput76), .B1(n21680), .B2(keyinput127), .ZN(n21679) );
  OAI221_X1 U24600 ( .B1(n21681), .B2(keyinput76), .C1(n21680), .C2(
        keyinput127), .A(n21679), .ZN(n21689) );
  AOI22_X1 U24601 ( .A1(n21684), .A2(keyinput79), .B1(n21683), .B2(keyinput103), .ZN(n21682) );
  OAI221_X1 U24602 ( .B1(n21684), .B2(keyinput79), .C1(n21683), .C2(
        keyinput103), .A(n21682), .ZN(n21688) );
  XNOR2_X1 U24603 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B(keyinput106), 
        .ZN(n21686) );
  XNOR2_X1 U24604 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput57), .ZN(
        n21685) );
  NAND2_X1 U24605 ( .A1(n21686), .A2(n21685), .ZN(n21687) );
  NOR4_X1 U24606 ( .A1(n21690), .A2(n21689), .A3(n21688), .A4(n21687), .ZN(
        n21739) );
  AOI22_X1 U24607 ( .A1(n21692), .A2(keyinput70), .B1(keyinput12), .B2(n11013), 
        .ZN(n21691) );
  OAI221_X1 U24608 ( .B1(n21692), .B2(keyinput70), .C1(n11013), .C2(keyinput12), .A(n21691), .ZN(n21704) );
  AOI22_X1 U24609 ( .A1(n21695), .A2(keyinput68), .B1(keyinput120), .B2(n21694), .ZN(n21693) );
  OAI221_X1 U24610 ( .B1(n21695), .B2(keyinput68), .C1(n21694), .C2(
        keyinput120), .A(n21693), .ZN(n21703) );
  INV_X1 U24611 ( .A(P2_EAX_REG_31__SCAN_IN), .ZN(n21697) );
  AOI22_X1 U24612 ( .A1(n21698), .A2(keyinput45), .B1(n21697), .B2(keyinput125), .ZN(n21696) );
  OAI221_X1 U24613 ( .B1(n21698), .B2(keyinput45), .C1(n21697), .C2(
        keyinput125), .A(n21696), .ZN(n21702) );
  XNOR2_X1 U24614 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(keyinput41), 
        .ZN(n21700) );
  XNOR2_X1 U24615 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B(keyinput38), .ZN(
        n21699) );
  NAND2_X1 U24616 ( .A1(n21700), .A2(n21699), .ZN(n21701) );
  NOR4_X1 U24617 ( .A1(n21704), .A2(n21703), .A3(n21702), .A4(n21701), .ZN(
        n21738) );
  AOI22_X1 U24618 ( .A1(n21707), .A2(keyinput55), .B1(keyinput110), .B2(n21706), .ZN(n21705) );
  OAI221_X1 U24619 ( .B1(n21707), .B2(keyinput55), .C1(n21706), .C2(
        keyinput110), .A(n21705), .ZN(n21720) );
  AOI22_X1 U24620 ( .A1(n21710), .A2(keyinput26), .B1(keyinput60), .B2(n21709), 
        .ZN(n21708) );
  OAI221_X1 U24621 ( .B1(n21710), .B2(keyinput26), .C1(n21709), .C2(keyinput60), .A(n21708), .ZN(n21719) );
  INV_X1 U24622 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n21713) );
  INV_X1 U24623 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n21712) );
  AOI22_X1 U24624 ( .A1(n21713), .A2(keyinput126), .B1(keyinput118), .B2(
        n21712), .ZN(n21711) );
  OAI221_X1 U24625 ( .B1(n21713), .B2(keyinput126), .C1(n21712), .C2(
        keyinput118), .A(n21711), .ZN(n21718) );
  AOI22_X1 U24626 ( .A1(n21716), .A2(keyinput105), .B1(keyinput52), .B2(n21715), .ZN(n21714) );
  OAI221_X1 U24627 ( .B1(n21716), .B2(keyinput105), .C1(n21715), .C2(
        keyinput52), .A(n21714), .ZN(n21717) );
  NOR4_X1 U24628 ( .A1(n21720), .A2(n21719), .A3(n21718), .A4(n21717), .ZN(
        n21737) );
  AOI22_X1 U24629 ( .A1(n21723), .A2(keyinput43), .B1(n21722), .B2(keyinput27), 
        .ZN(n21721) );
  OAI221_X1 U24630 ( .B1(n21723), .B2(keyinput43), .C1(n21722), .C2(keyinput27), .A(n21721), .ZN(n21735) );
  INV_X1 U24631 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n21726) );
  AOI22_X1 U24632 ( .A1(n21726), .A2(keyinput50), .B1(keyinput17), .B2(n21725), 
        .ZN(n21724) );
  OAI221_X1 U24633 ( .B1(n21726), .B2(keyinput50), .C1(n21725), .C2(keyinput17), .A(n21724), .ZN(n21734) );
  AOI22_X1 U24634 ( .A1(n21729), .A2(keyinput86), .B1(n21728), .B2(keyinput104), .ZN(n21727) );
  OAI221_X1 U24635 ( .B1(n21729), .B2(keyinput86), .C1(n21728), .C2(
        keyinput104), .A(n21727), .ZN(n21733) );
  AOI22_X1 U24636 ( .A1(n16863), .A2(keyinput84), .B1(n21731), .B2(keyinput7), 
        .ZN(n21730) );
  OAI221_X1 U24637 ( .B1(n16863), .B2(keyinput84), .C1(n21731), .C2(keyinput7), 
        .A(n21730), .ZN(n21732) );
  NOR4_X1 U24638 ( .A1(n21735), .A2(n21734), .A3(n21733), .A4(n21732), .ZN(
        n21736) );
  NAND4_X1 U24639 ( .A1(n21739), .A2(n21738), .A3(n21737), .A4(n21736), .ZN(
        n21740) );
  AOI211_X1 U24640 ( .C1(keyinput85), .C2(n21742), .A(n21741), .B(n21740), 
        .ZN(n21743) );
  NAND4_X1 U24641 ( .A1(n21746), .A2(n21745), .A3(n21744), .A4(n21743), .ZN(
        n21760) );
  OAI22_X1 U24642 ( .A1(n21750), .A2(n21749), .B1(n21748), .B2(n21747), .ZN(
        n21751) );
  AOI21_X1 U24643 ( .B1(n21753), .B2(n21752), .A(n21751), .ZN(n21756) );
  NAND2_X1 U24644 ( .A1(n21754), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n21755) );
  OAI211_X1 U24645 ( .C1(n21758), .C2(n21757), .A(n21756), .B(n21755), .ZN(
        n21759) );
  XNOR2_X1 U24646 ( .A(n21760), .B(n21759), .ZN(P1_U3123) );
  OR2_X1 U12213 ( .A1(n20215), .A2(n17038), .ZN(n20196) );
  OR2_X1 U18779 ( .A1(n16578), .A2(n16990), .ZN(n20163) );
  AND2_X1 U18748 ( .A1(n16667), .A2(n16652), .ZN(n16637) );
  NOR2_X2 U11452 ( .A1(n9870), .A2(n9869), .ZN(n20180) );
  AOI21_X2 U12818 ( .B1(n16450), .B2(n15144), .A(n15153), .ZN(n16433) );
  NAND2_X2 U11277 ( .A1(n10709), .A2(n10708), .ZN(n15557) );
  BUF_X1 U11282 ( .A(n11769), .Z(n18497) );
  BUF_X1 U11335 ( .A(n10837), .Z(n11575) );
  NAND2_X1 U13311 ( .A1(n10425), .A2(n10702), .ZN(n10846) );
  CLKBUF_X1 U11159 ( .A(n10846), .Z(n11652) );
  CLKBUF_X1 U11186 ( .A(n11258), .Z(n11698) );
  INV_X2 U11197 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10289) );
  CLKBUF_X1 U11211 ( .A(n11740), .Z(n9729) );
  CLKBUF_X1 U11212 ( .A(n10777), .Z(n10868) );
  NOR2_X1 U11223 ( .A1(n20243), .A2(n20226), .ZN(n20227) );
  NAND2_X1 U11260 ( .A1(n13744), .A2(n12612), .ZN(n12624) );
  CLKBUF_X1 U11270 ( .A(n10883), .Z(n14697) );
  CLKBUF_X1 U11325 ( .A(n13782), .Z(n9720) );
  OR2_X1 U11346 ( .A1(n20149), .A2(n20130), .ZN(n20132) );
  OR2_X1 U11465 ( .A1(n20146), .A2(n20148), .ZN(n20149) );
  OR2_X1 U11888 ( .A1(n20241), .A2(n9774), .ZN(n20243) );
  CLKBUF_X1 U12203 ( .A(n18882), .Z(n18904) );
  INV_X1 U12621 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n21075) );
  AOI211_X1 U12753 ( .C1(n16690), .C2(n20269), .A(n16442), .B(n16441), .ZN(
        n16443) );
  OR3_X1 U12926 ( .A1(n10691), .A2(n10690), .A3(n10689), .ZN(P3_U2640) );
endmodule

