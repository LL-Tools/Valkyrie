

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6537, n6538, n6540,
         n6541, n6542, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6603, n6604, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15975;

  AOI211_X1 U7277 ( .C1(n15835), .C2(n14538), .A(n14537), .B(n14536), .ZN(
        n14622) );
  INV_X1 U7278 ( .A(n15224), .ZN(n15244) );
  NAND2_X1 U7279 ( .A1(n9492), .A2(n9491), .ZN(n13674) );
  INV_X1 U7280 ( .A(n13864), .ZN(n13799) );
  CLKBUF_X3 U7281 ( .A(n15975), .Z(n6552) );
  NAND4_X1 U7282 ( .A1(n9045), .A2(n9046), .A3(n6910), .A4(n6909), .ZN(n15866)
         );
  AND2_X1 U7283 ( .A1(n9025), .A2(n9024), .ZN(n9065) );
  MUX2_X1 U7284 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n6544), .Z(n11054) );
  INV_X2 U7285 ( .A(n6538), .ZN(n8277) );
  INV_X1 U7286 ( .A(n13727), .ZN(n13319) );
  INV_X1 U7287 ( .A(n15557), .ZN(n10156) );
  CLKBUF_X2 U7288 ( .A(n7827), .Z(n8442) );
  AND4_X1 U7289 ( .A1(n7831), .A2(n7830), .A3(n7829), .A4(n7828), .ZN(n15629)
         );
  CLKBUF_X2 U7290 ( .A(n7859), .Z(n8182) );
  BUF_X2 U7291 ( .A(n9815), .Z(n6550) );
  INV_X1 U7292 ( .A(n7309), .ZN(n10798) );
  BUF_X2 U7293 ( .A(n9722), .Z(n9914) );
  NAND2_X1 U7294 ( .A1(n7714), .A2(n7715), .ZN(n12696) );
  NAND2_X1 U7295 ( .A1(n6777), .A2(n6718), .ZN(n7763) );
  AND2_X1 U7296 ( .A1(n6876), .A2(n6874), .ZN(n6529) );
  NOR2_X1 U7297 ( .A1(n9726), .A2(n9725), .ZN(n9727) );
  CLKBUF_X2 U7298 ( .A(n8543), .Z(n6596) );
  INV_X1 U7299 ( .A(P2_U3088), .ZN(n6530) );
  INV_X1 U7300 ( .A(n6530), .ZN(n6531) );
  INV_X1 U7301 ( .A(n12625), .ZN(n12507) );
  OR2_X1 U7302 ( .A1(n7284), .A2(n6654), .ZN(n6881) );
  INV_X1 U7303 ( .A(n12850), .ZN(n12838) );
  BUF_X1 U7304 ( .A(n9722), .Z(n6595) );
  INV_X1 U7306 ( .A(n9066), .ZN(n9437) );
  AND2_X1 U7307 ( .A1(n9025), .A2(n13723), .ZN(n9052) );
  AND2_X1 U7308 ( .A1(n9590), .A2(n13383), .ZN(n13407) );
  NAND2_X1 U7309 ( .A1(n13534), .A2(n12877), .ZN(n13518) );
  NAND2_X1 U7310 ( .A1(n9035), .A2(n9034), .ZN(n13727) );
  INV_X2 U7312 ( .A(n14752), .ZN(n15276) );
  NOR2_X2 U7313 ( .A1(n7438), .A2(n12057), .ZN(n15201) );
  NAND2_X1 U7314 ( .A1(n13531), .A2(n12870), .ZN(n13564) );
  AND2_X1 U7315 ( .A1(n8516), .A2(n12319), .ZN(n8557) );
  AND2_X1 U7316 ( .A1(n8592), .A2(n8591), .ZN(n11520) );
  INV_X1 U7317 ( .A(n11370), .ZN(n15804) );
  NAND2_X1 U7318 ( .A1(n7839), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7779) );
  AND2_X1 U7319 ( .A1(n15141), .A2(n15315), .ZN(n15124) );
  NAND2_X1 U7320 ( .A1(n15527), .A2(n15529), .ZN(n11499) );
  NAND2_X1 U7321 ( .A1(n14995), .A2(n10142), .ZN(n15232) );
  INV_X1 U7322 ( .A(n12526), .ZN(n15659) );
  AND4_X1 U7323 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(n11803)
         );
  NAND2_X1 U7324 ( .A1(n12929), .A2(n12925), .ZN(n12914) );
  NAND2_X1 U7325 ( .A1(n12746), .A2(n12745), .ZN(n13664) );
  NAND2_X2 U7326 ( .A1(n8777), .A2(n8776), .ZN(n14557) );
  NAND2_X2 U7328 ( .A1(n8807), .A2(n8806), .ZN(n14543) );
  INV_X1 U7329 ( .A(n12592), .ZN(n15325) );
  NAND2_X1 U7330 ( .A1(n7972), .A2(n7971), .ZN(n15389) );
  CLKBUF_X3 U7331 ( .A(n7832), .Z(n10638) );
  INV_X1 U7332 ( .A(n15346), .ZN(n15211) );
  XNOR2_X1 U7333 ( .A(n8028), .B(n8027), .ZN(n10683) );
  INV_X2 U7334 ( .A(n6821), .ZN(n13285) );
  INV_X1 U7335 ( .A(n12755), .ZN(n12801) );
  INV_X1 U7336 ( .A(n12790), .ZN(n11659) );
  INV_X2 U7337 ( .A(n14499), .ZN(n14484) );
  INV_X1 U7338 ( .A(n8917), .ZN(n11772) );
  INV_X1 U7339 ( .A(n15131), .ZN(n15309) );
  INV_X1 U7340 ( .A(n15252), .ZN(n15223) );
  INV_X1 U7341 ( .A(n14688), .ZN(n15057) );
  INV_X2 U7342 ( .A(n15178), .ZN(n15584) );
  AND2_X1 U7344 ( .A1(n7401), .A2(n6576), .ZN(n6532) );
  AND3_X1 U7345 ( .A1(n8487), .A2(n8486), .A3(n8586), .ZN(n6533) );
  XOR2_X1 U7346 ( .A(n13614), .B(n12385), .Z(n6534) );
  XOR2_X1 U7347 ( .A(n14218), .B(n13865), .Z(n6535) );
  NAND2_X2 U7348 ( .A1(n12100), .A2(n10124), .ZN(n12099) );
  NAND2_X1 U7349 ( .A1(n7742), .A2(n6895), .ZN(n7747) );
  NAND2_X2 U7350 ( .A1(n8663), .A2(n8662), .ZN(n14598) );
  NOR2_X2 U7351 ( .A1(n8238), .A2(n14703), .ZN(n6889) );
  NAND2_X2 U7352 ( .A1(n6776), .A2(n6684), .ZN(n11423) );
  XNOR2_X2 U7353 ( .A(n7741), .B(n7738), .ZN(n12430) );
  BUF_X4 U7356 ( .A(n7794), .Z(n6538) );
  NAND2_X2 U7357 ( .A1(n10565), .A2(n12491), .ZN(n7794) );
  OR2_X2 U7358 ( .A1(n11454), .A2(n11455), .ZN(n11761) );
  NOR4_X2 U7359 ( .A1(n15120), .A2(n15156), .A3(n15138), .A4(n12666), .ZN(
        n12667) );
  INV_X4 U7360 ( .A(n9516), .ZN(n9490) );
  AOI21_X2 U7361 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10011) );
  OAI21_X2 U7362 ( .B1(n8082), .B2(n8081), .A(n8080), .ZN(n8085) );
  NAND2_X2 U7363 ( .A1(n8060), .A2(n8050), .ZN(n8082) );
  XNOR2_X2 U7364 ( .A(n14040), .B(n15804), .ZN(n11368) );
  INV_X1 U7365 ( .A(n15076), .ZN(n7418) );
  OR2_X2 U7366 ( .A1(n7763), .A2(n12434), .ZN(n6660) );
  NAND2_X2 U7367 ( .A1(n14331), .A2(n8963), .ZN(n14317) );
  NOR4_X2 U7368 ( .A1(n12663), .A2(n10124), .A3(n12662), .A4(n12661), .ZN(
        n12665) );
  INV_X1 U7370 ( .A(n6552), .ZN(n6540) );
  OAI21_X4 U7371 ( .B1(n12426), .B2(n6540), .A(n6636), .ZN(n14968) );
  NAND2_X2 U7372 ( .A1(n9938), .A2(n9937), .ZN(n12426) );
  AOI21_X2 U7373 ( .B1(n11499), .B2(n10162), .A(n7637), .ZN(n15511) );
  AND2_X2 U7374 ( .A1(n11659), .A2(n13316), .ZN(n12937) );
  OAI21_X2 U7375 ( .B1(n8773), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8775) );
  INV_X2 U7376 ( .A(n8266), .ZN(n6541) );
  OAI21_X2 U7377 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n10059), .A(n15965), .ZN(
        n15956) );
  NOR2_X2 U7378 ( .A1(n15154), .A2(n12597), .ZN(n15139) );
  XNOR2_X2 U7379 ( .A(n10067), .B(n10064), .ZN(n15444) );
  NOR2_X2 U7380 ( .A1(n13217), .A2(n13216), .ZN(n13219) );
  OAI21_X2 U7381 ( .B1(n13518), .B2(n7247), .A(n7244), .ZN(n13438) );
  AOI21_X2 U7382 ( .B1(n15171), .B2(n10179), .A(n10178), .ZN(n15153) );
  NAND2_X2 U7383 ( .A1(n12279), .A2(n10177), .ZN(n15171) );
  NAND2_X2 U7384 ( .A1(n15958), .A2(n10063), .ZN(n10067) );
  OAI211_X2 U7385 ( .C1(n7191), .C2(n9111), .A(n7189), .B(n9164), .ZN(n9173)
         );
  NAND2_X2 U7386 ( .A1(n9108), .A2(n9107), .ZN(n9111) );
  OAI21_X2 U7387 ( .B1(n8026), .B2(n8025), .A(n12288), .ZN(n14762) );
  NAND2_X2 U7388 ( .A1(n7564), .A2(n7561), .ZN(n12288) );
  OAI211_X2 U7389 ( .C1(n14384), .C2(n7284), .A(n6881), .B(n9987), .ZN(n14331)
         );
  NAND2_X2 U7390 ( .A1(n8958), .A2(n14373), .ZN(n14384) );
  BUF_X4 U7391 ( .A(n9052), .Z(n6542) );
  AOI21_X2 U7392 ( .B1(n8109), .B2(n7422), .A(n7420), .ZN(n7419) );
  NAND2_X2 U7393 ( .A1(n8085), .A2(n8084), .ZN(n8109) );
  OAI222_X1 U7394 ( .A1(n11978), .A2(n12426), .B1(n12703), .B2(P2_U3088), .C1(
        n12739), .C2(n12702), .ZN(P2_U3297) );
  AND2_X1 U7395 ( .A1(n12703), .A2(n7602), .ZN(n8536) );
  NAND3_X2 U7396 ( .A1(n8527), .A2(n8528), .A3(n8526), .ZN(n8529) );
  OR2_X1 U7397 ( .A1(n9939), .A2(n10615), .ZN(n8528) );
  NAND2_X2 U7398 ( .A1(n8514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8511) );
  OAI22_X2 U7400 ( .A1(n7316), .A2(n11288), .B1(n7314), .B2(n7312), .ZN(n11459) );
  XNOR2_X2 U7401 ( .A(n8910), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8917) );
  XNOR2_X2 U7402 ( .A(n13674), .B(n13343), .ZN(n13365) );
  NAND4_X4 U7403 ( .A1(n8541), .A2(n8540), .A3(n8538), .A4(n8539), .ZN(n9670)
         );
  NAND2_X1 U7404 ( .A1(n9035), .A2(n9034), .ZN(n6544) );
  NAND2_X1 U7405 ( .A1(n9035), .A2(n9034), .ZN(n6545) );
  BUF_X8 U7407 ( .A(n11225), .Z(n13864) );
  NOR2_X2 U7408 ( .A1(n11459), .A2(n11458), .ZN(n11460) );
  XNOR2_X2 U7409 ( .A(n8494), .B(n8493), .ZN(n12399) );
  NAND2_X2 U7410 ( .A1(n8549), .A2(n8548), .ZN(n14041) );
  XNOR2_X2 U7411 ( .A(n14823), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n6982) );
  INV_X4 U7412 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14823) );
  NAND2_X2 U7413 ( .A1(n15962), .A2(n10071), .ZN(n15447) );
  AND2_X1 U7414 ( .A1(n7603), .A2(n6735), .ZN(n14234) );
  NAND2_X1 U7415 ( .A1(n10141), .A2(n7432), .ZN(n14995) );
  OAI21_X1 U7416 ( .B1(n13926), .B2(n6565), .A(n6562), .ZN(n6567) );
  NAND2_X1 U7417 ( .A1(n7107), .A2(n6729), .ZN(n10141) );
  NAND2_X1 U7418 ( .A1(n6868), .A2(n15026), .ZN(n7107) );
  NAND2_X1 U7419 ( .A1(n6917), .A2(n6916), .ZN(n13369) );
  AND2_X1 U7420 ( .A1(n7272), .A2(n6548), .ZN(n13366) );
  AND2_X1 U7421 ( .A1(n6548), .A2(n12761), .ZN(n13372) );
  NAND2_X1 U7422 ( .A1(n14328), .A2(n14334), .ZN(n14330) );
  INV_X1 U7423 ( .A(n14241), .ZN(n6930) );
  AND2_X1 U7424 ( .A1(n8390), .A2(n8389), .ZN(n15003) );
  AND2_X1 U7425 ( .A1(n8372), .A2(n8371), .ZN(n15261) );
  NAND2_X1 U7426 ( .A1(n13972), .A2(n13747), .ZN(n13880) );
  AND2_X1 U7427 ( .A1(n8316), .A2(n8315), .ZN(n14752) );
  INV_X1 U7428 ( .A(n14334), .ZN(n9987) );
  NAND2_X1 U7429 ( .A1(n11933), .A2(n11930), .ZN(n13173) );
  NAND2_X1 U7430 ( .A1(n11763), .A2(n11762), .ZN(n11933) );
  AOI21_X1 U7431 ( .B1(n6710), .B2(n7076), .A(n6905), .ZN(n6906) );
  NAND2_X1 U7432 ( .A1(n11761), .A2(n11760), .ZN(n11763) );
  NAND2_X1 U7433 ( .A1(n8762), .A2(n8761), .ZN(n14562) );
  NAND2_X1 U7434 ( .A1(n11604), .A2(n6552), .ZN(n8213) );
  NAND2_X1 U7435 ( .A1(n12254), .A2(n6690), .ZN(n12305) );
  NAND2_X1 U7436 ( .A1(n7494), .A2(n7489), .ZN(n15452) );
  INV_X1 U7437 ( .A(n12098), .ZN(n6549) );
  INV_X2 U7438 ( .A(n15372), .ZN(n12062) );
  AND2_X1 U7439 ( .A1(n8066), .A2(n8065), .ZN(n15346) );
  CLKBUF_X1 U7440 ( .A(n7988), .Z(n7991) );
  INV_X2 U7441 ( .A(n15531), .ZN(n12338) );
  NOR2_X1 U7442 ( .A1(n8715), .A2(n14008), .ZN(n8693) );
  INV_X1 U7443 ( .A(n15793), .ZN(n15764) );
  INV_X4 U7444 ( .A(n6595), .ZN(n6546) );
  INV_X1 U7445 ( .A(n15667), .ZN(n11652) );
  INV_X1 U7446 ( .A(n15562), .ZN(n15486) );
  NAND2_X1 U7447 ( .A1(n11576), .A2(n8266), .ZN(n7931) );
  INV_X4 U7448 ( .A(n12385), .ZN(n11664) );
  NOR2_X2 U7449 ( .A1(n15866), .A2(n9554), .ZN(n11665) );
  NAND2_X2 U7450 ( .A1(n8635), .A2(n8660), .ZN(n15718) );
  NAND2_X1 U7451 ( .A1(n8620), .A2(n8632), .ZN(n14129) );
  BUF_X2 U7452 ( .A(n8536), .Z(n6598) );
  BUF_X2 U7453 ( .A(n8536), .Z(n6597) );
  BUF_X2 U7454 ( .A(n7825), .Z(n8396) );
  BUF_X4 U7455 ( .A(n9668), .Z(n6547) );
  NAND4_X1 U7456 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n13150)
         );
  NAND2_X1 U7457 ( .A1(n6946), .A2(n6944), .ZN(n11662) );
  INV_X4 U7458 ( .A(n8448), .ZN(n10208) );
  OR2_X1 U7459 ( .A1(n8619), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8632) );
  NAND3_X2 U7460 ( .A1(n10646), .A2(n12026), .A3(n11904), .ZN(n10565) );
  BUF_X1 U7461 ( .A(n8916), .Z(n10005) );
  INV_X2 U7462 ( .A(n9603), .ZN(n9359) );
  INV_X1 U7463 ( .A(n11605), .ZN(n6553) );
  INV_X1 U7464 ( .A(n12430), .ZN(n12645) );
  XNOR2_X1 U7465 ( .A(n8907), .B(n8906), .ZN(n11605) );
  OAI21_X1 U7466 ( .B1(n9631), .B2(P3_IR_REG_23__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9633) );
  XNOR2_X1 U7467 ( .A(n7674), .B(SI_5_), .ZN(n7878) );
  XNOR2_X1 U7468 ( .A(n9545), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12755) );
  AND2_X1 U7469 ( .A1(n8686), .A2(n6588), .ZN(n8873) );
  NAND4_X2 U7470 ( .A1(n9041), .A2(n9008), .A3(n7072), .A4(n7071), .ZN(n9095)
         );
  INV_X2 U7471 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7472 ( .A1(n6784), .A2(n9795), .ZN(n9802) );
  AND2_X1 U7473 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  OAI21_X1 U7474 ( .B1(n10529), .B2(n10528), .A(n10527), .ZN(n10530) );
  OR2_X1 U7475 ( .A1(n7277), .A2(n8995), .ZN(n8997) );
  OR2_X1 U7476 ( .A1(n7277), .A2(n9003), .ZN(n9005) );
  AND3_X1 U7477 ( .A1(n12487), .A2(n12488), .A3(n12486), .ZN(n12639) );
  XNOR2_X1 U7478 ( .A(n6566), .B(n6535), .ZN(n13872) );
  OAI21_X1 U7479 ( .B1(n15006), .B2(n7552), .A(n7549), .ZN(n10206) );
  AND2_X1 U7480 ( .A1(n12634), .A2(n12633), .ZN(n12635) );
  NAND2_X1 U7481 ( .A1(n6567), .A2(n6817), .ZN(n6566) );
  NAND2_X1 U7482 ( .A1(n6561), .A2(n7385), .ZN(n13861) );
  NAND2_X1 U7483 ( .A1(n14234), .A2(n14241), .ZN(n14233) );
  AOI21_X1 U7484 ( .B1(n8986), .B2(n8985), .A(n13870), .ZN(n14212) );
  NAND2_X1 U7485 ( .A1(n13926), .A2(n7386), .ZN(n6561) );
  AND2_X1 U7486 ( .A1(n14775), .A2(n6778), .ZN(n14745) );
  AND2_X1 U7487 ( .A1(n13331), .A2(n13333), .ZN(n12935) );
  OR2_X1 U7488 ( .A1(n13609), .A2(n13608), .ZN(n13678) );
  NAND2_X1 U7489 ( .A1(n12753), .A2(n12752), .ZN(n13331) );
  NAND2_X1 U7490 ( .A1(n7306), .A2(n6692), .ZN(n8986) );
  NAND3_X1 U7491 ( .A1(n13792), .A2(n13791), .A3(n13790), .ZN(n13926) );
  NAND2_X1 U7492 ( .A1(n13664), .A2(n12930), .ZN(n12927) );
  NOR2_X1 U7493 ( .A1(n13340), .A2(n7088), .ZN(n7087) );
  AOI21_X1 U7494 ( .B1(n10272), .B2(n15757), .A(n13810), .ZN(n14232) );
  NAND2_X1 U7495 ( .A1(n6558), .A2(n6678), .ZN(n7603) );
  NOR2_X1 U7496 ( .A1(n12467), .A2(n12466), .ZN(n12476) );
  OAI21_X1 U7497 ( .B1(n12459), .B2(n12453), .A(n12451), .ZN(n12467) );
  AND2_X1 U7498 ( .A1(n10245), .A2(n10244), .ZN(n10102) );
  OR2_X1 U7499 ( .A1(n9664), .A2(n13345), .ZN(n12929) );
  NAND2_X1 U7500 ( .A1(n14288), .A2(n8827), .ZN(n14274) );
  AOI21_X1 U7501 ( .B1(n7385), .B2(n6564), .A(n6563), .ZN(n6562) );
  AND2_X1 U7502 ( .A1(n12704), .A2(n10538), .ZN(n12721) );
  INV_X1 U7503 ( .A(n7385), .ZN(n6565) );
  AND2_X1 U7504 ( .A1(n13789), .A2(n13788), .ZN(n13825) );
  NAND2_X1 U7505 ( .A1(n12916), .A2(n12918), .ZN(n13338) );
  OR2_X1 U7506 ( .A1(n9525), .A2(n13358), .ZN(n12916) );
  NAND2_X1 U7507 ( .A1(n6801), .A2(n9896), .ZN(n12395) );
  NAND2_X1 U7508 ( .A1(n7551), .A2(n7550), .ZN(n7549) );
  OAI22_X1 U7509 ( .A1(n15220), .A2(n12625), .B1(n12447), .B2(n12446), .ZN(
        n12453) );
  NAND2_X1 U7510 ( .A1(n12641), .A2(n12640), .ZN(n15215) );
  OAI21_X1 U7511 ( .B1(n13874), .B2(n13873), .A(n6590), .ZN(n13789) );
  NAND2_X1 U7512 ( .A1(n14694), .A2(n8205), .ZN(n14754) );
  NAND2_X1 U7513 ( .A1(n7587), .A2(n7588), .ZN(n14694) );
  INV_X1 U7514 ( .A(n7386), .ZN(n6564) );
  NAND2_X1 U7515 ( .A1(n13945), .A2(n13781), .ZN(n13874) );
  OAI21_X1 U7516 ( .B1(n14315), .B2(n7623), .A(n7622), .ZN(n14290) );
  INV_X1 U7517 ( .A(n14968), .ZN(n15220) );
  INV_X1 U7518 ( .A(n12908), .ZN(n6548) );
  INV_X1 U7519 ( .A(n13860), .ZN(n6563) );
  INV_X1 U7520 ( .A(n10546), .ZN(n10552) );
  NAND2_X1 U7521 ( .A1(n13946), .A2(n13947), .ZN(n13945) );
  NAND2_X1 U7522 ( .A1(n14330), .A2(n8796), .ZN(n14315) );
  NOR2_X1 U7523 ( .A1(n6929), .A2(n6925), .ZN(n6924) );
  XNOR2_X1 U7524 ( .A(n9895), .B(n9894), .ZN(n14657) );
  CLKBUF_X1 U7525 ( .A(n13901), .Z(n6864) );
  INV_X1 U7526 ( .A(n15237), .ZN(n12448) );
  AND2_X1 U7527 ( .A1(n7531), .A2(n10201), .ZN(n7530) );
  XNOR2_X1 U7528 ( .A(n12722), .B(n11213), .ZN(n10546) );
  NAND2_X1 U7529 ( .A1(n13858), .A2(n13859), .ZN(n6817) );
  NAND2_X1 U7530 ( .A1(n7119), .A2(n7120), .ZN(n7117) );
  AND2_X1 U7531 ( .A1(n10144), .A2(n10143), .ZN(n15237) );
  NAND2_X1 U7532 ( .A1(n13813), .A2(n6884), .ZN(n13901) );
  NAND2_X1 U7533 ( .A1(n14350), .A2(n8786), .ZN(n14328) );
  OR2_X1 U7534 ( .A1(n9936), .A2(n9935), .ZN(n9938) );
  NAND2_X1 U7535 ( .A1(n9904), .A2(n9903), .ZN(n12722) );
  NAND2_X1 U7536 ( .A1(n13070), .A2(n13069), .ZN(n13068) );
  NAND2_X1 U7537 ( .A1(n7384), .A2(n7382), .ZN(n13813) );
  AND2_X1 U7538 ( .A1(n7498), .A2(n6986), .ZN(n6983) );
  AND2_X1 U7539 ( .A1(n8438), .A2(n8437), .ZN(n15224) );
  NAND2_X1 U7540 ( .A1(n6932), .A2(n6935), .ZN(n6931) );
  NAND2_X1 U7541 ( .A1(n8859), .A2(n8858), .ZN(n14218) );
  NAND2_X1 U7542 ( .A1(n7618), .A2(n7617), .ZN(n14350) );
  AND2_X1 U7543 ( .A1(n6584), .A2(n6583), .ZN(n7119) );
  AND2_X1 U7544 ( .A1(n9488), .A2(n7168), .ZN(n12320) );
  NOR2_X1 U7545 ( .A1(n7413), .A2(n7412), .ZN(n7123) );
  NAND2_X1 U7546 ( .A1(n8837), .A2(n8836), .ZN(n14519) );
  OR2_X1 U7547 ( .A1(n7120), .A2(n10134), .ZN(n6584) );
  AND2_X1 U7548 ( .A1(n15108), .A2(n10133), .ZN(n10134) );
  NAND2_X1 U7549 ( .A1(n9460), .A2(n9459), .ZN(n13399) );
  OR2_X1 U7550 ( .A1(n13784), .A2(n13783), .ZN(n6590) );
  NAND2_X1 U7551 ( .A1(n14399), .A2(n8734), .ZN(n8747) );
  INV_X1 U7552 ( .A(n7417), .ZN(n7412) );
  NAND2_X1 U7553 ( .A1(n13610), .A2(n12975), .ZN(n13383) );
  OR2_X1 U7554 ( .A1(n13610), .A2(n12975), .ZN(n9590) );
  OAI21_X1 U7555 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9901) );
  XNOR2_X1 U7556 ( .A(n14527), .B(n14020), .ZN(n14254) );
  NAND2_X1 U7557 ( .A1(n7418), .A2(n15089), .ZN(n7417) );
  NAND2_X2 U7558 ( .A1(n8496), .A2(n8495), .ZN(n14527) );
  AND2_X1 U7559 ( .A1(n8346), .A2(n8345), .ZN(n15267) );
  NAND2_X1 U7560 ( .A1(n13051), .A2(n13050), .ZN(n12356) );
  OAI21_X1 U7561 ( .B1(n14504), .B2(n7608), .A(n7606), .ZN(n14399) );
  NAND2_X1 U7562 ( .A1(n13166), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13193) );
  NOR2_X1 U7563 ( .A1(n13765), .A2(n7368), .ZN(n7367) );
  XNOR2_X1 U7564 ( .A(n14543), .B(n14287), .ZN(n14299) );
  NAND2_X1 U7565 ( .A1(n15458), .A2(n10082), .ZN(n15462) );
  AND2_X1 U7566 ( .A1(n6586), .A2(n6734), .ZN(n13974) );
  XNOR2_X1 U7567 ( .A(n15091), .B(n15098), .ZN(n15082) );
  NAND2_X2 U7568 ( .A1(n8829), .A2(n8828), .ZN(n14532) );
  NAND2_X1 U7569 ( .A1(n12125), .A2(n12124), .ZN(n12129) );
  NAND2_X1 U7570 ( .A1(n13933), .A2(n6585), .ZN(n6586) );
  NAND2_X1 U7571 ( .A1(n13933), .A2(n13739), .ZN(n13836) );
  NAND2_X1 U7572 ( .A1(n15434), .A2(n10638), .ZN(n15076) );
  NAND2_X2 U7573 ( .A1(n8798), .A2(n8797), .ZN(n14548) );
  NAND2_X2 U7574 ( .A1(n8237), .A2(n8236), .ZN(n15091) );
  OAI21_X1 U7575 ( .B1(n7350), .B2(n6907), .A(n6906), .ZN(n13471) );
  AOI21_X1 U7576 ( .B1(n14410), .B2(n7299), .A(n7303), .ZN(n7298) );
  NAND2_X1 U7577 ( .A1(n8341), .A2(n8340), .ZN(n8367) );
  XNOR2_X1 U7578 ( .A(n8284), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U7579 ( .A1(n8185), .A2(n8184), .ZN(n15131) );
  NAND2_X1 U7580 ( .A1(n7586), .A2(n7584), .ZN(n12125) );
  NAND2_X1 U7581 ( .A1(n11980), .A2(n11984), .ZN(n11982) );
  XNOR2_X1 U7582 ( .A(n8314), .B(n8313), .ZN(n11903) );
  XNOR2_X1 U7583 ( .A(n14557), .B(n14337), .ZN(n14351) );
  NAND2_X1 U7584 ( .A1(n6904), .A2(n8787), .ZN(n14553) );
  NAND2_X1 U7585 ( .A1(n13733), .A2(n13732), .ZN(n13934) );
  XNOR2_X1 U7586 ( .A(n8235), .B(n8234), .ZN(n11879) );
  XNOR2_X1 U7587 ( .A(n8311), .B(n8263), .ZN(n11546) );
  NAND2_X1 U7588 ( .A1(n8337), .A2(n8334), .ZN(n8314) );
  XNOR2_X1 U7589 ( .A(n8283), .B(n8282), .ZN(n8805) );
  XNOR2_X1 U7590 ( .A(n13628), .B(n13482), .ZN(n13470) );
  INV_X1 U7591 ( .A(n15332), .ZN(n15183) );
  NAND2_X1 U7592 ( .A1(n8262), .A2(n7165), .ZN(n8337) );
  AND2_X2 U7593 ( .A1(n8165), .A2(n8164), .ZN(n15315) );
  NAND2_X1 U7594 ( .A1(n8692), .A2(n8691), .ZN(n14573) );
  XNOR2_X1 U7595 ( .A(n8230), .B(n8254), .ZN(n11604) );
  NAND2_X2 U7596 ( .A1(n9379), .A2(n9378), .ZN(n13628) );
  AND2_X1 U7597 ( .A1(n6587), .A2(n13739), .ZN(n6585) );
  NAND2_X1 U7598 ( .A1(n8752), .A2(n8751), .ZN(n14568) );
  NAND2_X1 U7599 ( .A1(n11176), .A2(n9902), .ZN(n8692) );
  NAND2_X1 U7600 ( .A1(n6579), .A2(n11528), .ZN(n11857) );
  NAND2_X1 U7601 ( .A1(n6555), .A2(n8593), .ZN(n11549) );
  XNOR2_X1 U7602 ( .A(n8231), .B(n11484), .ZN(n8230) );
  NAND2_X1 U7603 ( .A1(n11512), .A2(n11513), .ZN(n6555) );
  NAND2_X1 U7604 ( .A1(n8950), .A2(n8949), .ZN(n14593) );
  OAI21_X1 U7605 ( .B1(n12336), .B2(n12333), .A(n12334), .ZN(n7892) );
  NAND2_X1 U7606 ( .A1(n11388), .A2(n11387), .ZN(n11389) );
  NAND2_X1 U7607 ( .A1(n8703), .A2(n8702), .ZN(n14578) );
  XNOR2_X1 U7608 ( .A(n8155), .B(n8156), .ZN(n11198) );
  OR2_X1 U7609 ( .A1(n14583), .A2(n14589), .ZN(n7520) );
  OAI21_X1 U7610 ( .B1(n11388), .B2(n6578), .A(n6532), .ZN(n6579) );
  XNOR2_X1 U7611 ( .A(n8137), .B(n7650), .ZN(n11176) );
  OR2_X1 U7612 ( .A1(n11463), .A2(n11464), .ZN(n7336) );
  NAND2_X1 U7613 ( .A1(n6922), .A2(n8211), .ZN(n8231) );
  NAND2_X1 U7614 ( .A1(n8116), .A2(n8115), .ZN(n12585) );
  NAND2_X1 U7615 ( .A1(n6556), .A2(n8577), .ZN(n11512) );
  NAND2_X1 U7616 ( .A1(n8713), .A2(n8712), .ZN(n14583) );
  NAND2_X1 U7617 ( .A1(n7869), .A2(n11423), .ZN(n12336) );
  NAND2_X1 U7618 ( .A1(n8011), .A2(n8010), .ZN(n15372) );
  NAND2_X1 U7619 ( .A1(n8725), .A2(n8724), .ZN(n14589) );
  NAND2_X1 U7620 ( .A1(n8036), .A2(n8035), .ZN(n15352) );
  NAND2_X1 U7621 ( .A1(n8649), .A2(n8648), .ZN(n13842) );
  OAI21_X1 U7622 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n10029), .A(n10028), .ZN(
        n10084) );
  NAND2_X1 U7623 ( .A1(n11275), .A2(n11274), .ZN(n11310) );
  NAND2_X1 U7624 ( .A1(n8638), .A2(n8637), .ZN(n14604) );
  OAI21_X1 U7625 ( .B1(n11269), .B2(n7056), .A(n7054), .ZN(n11473) );
  NAND2_X1 U7626 ( .A1(n6575), .A2(n7426), .ZN(n8060) );
  NAND2_X1 U7627 ( .A1(n6571), .A2(n7688), .ZN(n7988) );
  NAND2_X1 U7628 ( .A1(n8608), .A2(n8607), .ZN(n15834) );
  NOR2_X1 U7629 ( .A1(n15443), .A2(n10068), .ZN(n10070) );
  NAND2_X1 U7630 ( .A1(n8544), .A2(n6559), .ZN(n15761) );
  NAND2_X1 U7631 ( .A1(n7949), .A2(n7948), .ZN(n12548) );
  NOR2_X1 U7632 ( .A1(n15444), .A2(n15445), .ZN(n15443) );
  NAND2_X1 U7633 ( .A1(n11333), .A2(n9977), .ZN(n6559) );
  NAND2_X1 U7634 ( .A1(n7919), .A2(n7918), .ZN(n12530) );
  AND3_X1 U7636 ( .A1(n6677), .A2(n6943), .A3(n6942), .ZN(n11748) );
  NOR2_X1 U7637 ( .A1(n13862), .A2(n11335), .ZN(n11298) );
  CLKBUF_X1 U7638 ( .A(n13110), .Z(n13130) );
  NAND2_X1 U7640 ( .A1(n7182), .A2(n7183), .ZN(n9292) );
  NAND2_X1 U7641 ( .A1(n15622), .A2(n12492), .ZN(n15565) );
  NAND2_X1 U7642 ( .A1(n10025), .A2(n10026), .ZN(n10044) );
  NAND3_X1 U7643 ( .A1(n8565), .A2(n8566), .A3(n7404), .ZN(n11370) );
  AND2_X1 U7644 ( .A1(n8576), .A2(n8575), .ZN(n15811) );
  NAND2_X1 U7645 ( .A1(n15960), .A2(n15959), .ZN(n15958) );
  AND3_X2 U7646 ( .A1(n8554), .A2(n8553), .A3(n8552), .ZN(n15793) );
  NAND2_X2 U7647 ( .A1(n7203), .A2(n7204), .ZN(n9722) );
  NAND2_X1 U7648 ( .A1(n10992), .A2(n10991), .ZN(n11225) );
  NAND2_X1 U7649 ( .A1(n7912), .A2(n7677), .ZN(n7408) );
  AND2_X1 U7650 ( .A1(n7865), .A2(n7864), .ZN(n12519) );
  BUF_X4 U7651 ( .A(n12507), .Z(n12619) );
  XNOR2_X1 U7652 ( .A(n10060), .B(n10061), .ZN(n15960) );
  NAND2_X1 U7653 ( .A1(n7806), .A2(n6669), .ZN(n15562) );
  NOR2_X4 U7654 ( .A1(n11401), .A2(n11047), .ZN(n12802) );
  NAND2_X1 U7655 ( .A1(n6580), .A2(n7675), .ZN(n7912) );
  NAND2_X1 U7656 ( .A1(n8537), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U7657 ( .A1(n7407), .A2(n6581), .ZN(n6580) );
  NAND2_X1 U7658 ( .A1(n7764), .A2(n15207), .ZN(n11576) );
  AND4_X1 U7659 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n10153)
         );
  INV_X2 U7660 ( .A(n9940), .ZN(n8846) );
  NAND2_X1 U7661 ( .A1(n8557), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U7662 ( .A1(n8542), .A2(n10567), .ZN(n9940) );
  NAND2_X1 U7663 ( .A1(n6582), .A2(n7673), .ZN(n7407) );
  INV_X1 U7664 ( .A(n7826), .ZN(n8219) );
  NAND4_X1 U7665 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n11047)
         );
  XNOR2_X1 U7666 ( .A(n8775), .B(n8774), .ZN(n9668) );
  AND2_X1 U7668 ( .A1(n11772), .A2(n11880), .ZN(n6591) );
  NAND2_X1 U7669 ( .A1(n8516), .A2(n7602), .ZN(n8530) );
  NAND2_X1 U7670 ( .A1(n11147), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11146) );
  CLKBUF_X2 U7671 ( .A(n7873), .Z(n7976) );
  CLKBUF_X1 U7672 ( .A(n7812), .Z(n8064) );
  INV_X1 U7673 ( .A(n6538), .ZN(n6551) );
  INV_X1 U7674 ( .A(n12490), .ZN(n12492) );
  NAND2_X1 U7675 ( .A1(n7752), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8012) );
  INV_X1 U7676 ( .A(n6573), .ZN(n6572) );
  AND2_X1 U7677 ( .A1(n11128), .A2(n11091), .ZN(n11147) );
  NAND2_X1 U7678 ( .A1(n7359), .A2(n7357), .ZN(n9210) );
  CLKBUF_X3 U7679 ( .A(n9166), .Z(n12751) );
  INV_X1 U7680 ( .A(n15428), .ZN(n7749) );
  NAND2_X1 U7681 ( .A1(n7746), .A2(n7747), .ZN(n15428) );
  OAI21_X1 U7682 ( .B1(n7686), .B2(n6574), .A(n6728), .ZN(n6573) );
  NAND2_X1 U7683 ( .A1(n8916), .A2(n11605), .ZN(n10991) );
  INV_X1 U7684 ( .A(n7997), .ZN(n7752) );
  AND2_X1 U7685 ( .A1(n7731), .A2(n7730), .ZN(n10646) );
  MUX2_X1 U7686 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8513), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8515) );
  NAND2_X1 U7687 ( .A1(n6557), .A2(n8510), .ZN(n8514) );
  NAND2_X1 U7688 ( .A1(n9629), .A2(n9628), .ZN(n12323) );
  INV_X1 U7689 ( .A(n7878), .ZN(n6581) );
  NAND2_X1 U7690 ( .A1(n7663), .A2(n6569), .ZN(n7810) );
  AND2_X1 U7691 ( .A1(n8699), .A2(n8688), .ZN(n8749) );
  XNOR2_X1 U7692 ( .A(n7737), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11904) );
  OR2_X1 U7693 ( .A1(n7951), .A2(n7950), .ZN(n7974) );
  INV_X1 U7694 ( .A(n8512), .ZN(n6557) );
  NAND2_X1 U7695 ( .A1(n9030), .A2(n9032), .ZN(n12424) );
  NAND2_X1 U7696 ( .A1(n15420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7558) );
  XNOR2_X1 U7697 ( .A(n9129), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11283) );
  NAND2_X1 U7698 ( .A1(n8886), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8911) );
  MUX2_X1 U7699 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7762), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n12438) );
  NAND2_X1 U7700 ( .A1(n6660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7758) );
  XNOR2_X1 U7701 ( .A(n7740), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7760) );
  OAI21_X1 U7702 ( .B1(n8427), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7736) );
  NAND2_X1 U7703 ( .A1(n7711), .A2(n7557), .ZN(n15420) );
  NAND2_X2 U7704 ( .A1(n10581), .A2(n6531), .ZN(n11978) );
  XNOR2_X1 U7705 ( .A(n7678), .B(SI_6_), .ZN(n7913) );
  XNOR2_X1 U7706 ( .A(n9358), .B(n9357), .ZN(n13316) );
  NAND2_X1 U7707 ( .A1(n7791), .A2(n6570), .ZN(n7774) );
  XNOR2_X1 U7708 ( .A(n7683), .B(SI_8_), .ZN(n7942) );
  XNOR2_X1 U7709 ( .A(n9543), .B(P3_IR_REG_20__SCAN_IN), .ZN(n12790) );
  AND2_X1 U7710 ( .A1(n8873), .A2(n8687), .ZN(n8699) );
  NAND2_X1 U7711 ( .A1(n8491), .A2(n7626), .ZN(n8512) );
  OAI21_X1 U7712 ( .B1(n10050), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6653), .ZN(
        n10019) );
  MUX2_X1 U7713 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9033), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n9035) );
  MUX2_X1 U7714 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7713), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n7715) );
  INV_X1 U7715 ( .A(n8492), .ZN(n8491) );
  INV_X2 U7716 ( .A(n11545), .ZN(n6554) );
  INV_X2 U7717 ( .A(n7658), .ZN(n10581) );
  NAND2_X2 U7718 ( .A1(n10575), .A2(P1_U3086), .ZN(n15433) );
  AOI21_X1 U7719 ( .B1(n7375), .B2(n7374), .A(n7373), .ZN(n7372) );
  AND2_X1 U7720 ( .A1(n8686), .A2(n8685), .ZN(n7230) );
  OAI21_X1 U7721 ( .B1(n7676), .B2(n7665), .A(n7664), .ZN(n7667) );
  NAND2_X1 U7722 ( .A1(n7658), .A2(n7657), .ZN(n7791) );
  INV_X1 U7723 ( .A(n8160), .ZN(n6777) );
  NAND2_X1 U7724 ( .A1(n7676), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U7725 ( .A1(n7676), .A2(SI_0_), .ZN(n10572) );
  NAND4_X1 U7726 ( .A1(n7281), .A2(n7280), .A3(n6616), .A4(n7278), .ZN(n8492)
         );
  OR2_X1 U7727 ( .A1(n8563), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8585) );
  AND2_X1 U7728 ( .A1(n6560), .A2(n6533), .ZN(n7280) );
  AND2_X1 U7729 ( .A1(n7279), .A2(n8673), .ZN(n7278) );
  AND2_X1 U7730 ( .A1(n8872), .A2(n8478), .ZN(n7281) );
  NOR2_X1 U7731 ( .A1(n9615), .A2(n9017), .ZN(n9018) );
  NAND2_X1 U7732 ( .A1(n6898), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U7733 ( .A1(n7150), .A2(n10252), .ZN(n7149) );
  AND2_X1 U7734 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n6568) );
  AND3_X1 U7735 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n6560) );
  AND2_X1 U7736 ( .A1(n8685), .A2(n6589), .ZN(n6588) );
  AND2_X1 U7737 ( .A1(n7507), .A2(n7506), .ZN(n8673) );
  AND4_X1 U7738 ( .A1(n6589), .A2(n8685), .A3(n8906), .A4(n8488), .ZN(n6616)
         );
  INV_X1 U7739 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8140) );
  NOR2_X1 U7740 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n9011) );
  INV_X1 U7741 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14967) );
  INV_X1 U7742 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6903) );
  XNOR2_X1 U7743 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9047) );
  INV_X1 U7744 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8161) );
  INV_X4 U7745 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7746 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8482) );
  NOR2_X1 U7747 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n8483) );
  NOR2_X1 U7748 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8481) );
  NOR2_X1 U7749 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8479) );
  NOR2_X1 U7750 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8485) );
  INV_X1 U7751 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8096) );
  NOR2_X1 U7752 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8480) );
  INV_X1 U7753 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6835) );
  NOR2_X1 U7754 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8484) );
  INV_X1 U7755 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8906) );
  INV_X1 U7756 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8032) );
  INV_X2 U7757 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9041) );
  INV_X1 U7758 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U7759 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n9009) );
  CLKBUF_X1 U7760 ( .A(P1_IR_REG_5__SCAN_IN), .Z(n7880) );
  INV_X1 U7761 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7734) );
  INV_X1 U7762 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9112) );
  NOR2_X1 U7763 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7757) );
  OR2_X1 U7764 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n8887) );
  INV_X1 U7765 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7106) );
  XOR2_X1 U7766 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n10051) );
  INV_X2 U7767 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NAND2_X1 U7768 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7871) );
  NOR2_X1 U7769 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n7507) );
  NAND2_X1 U7770 ( .A1(n11318), .A2(n8928), .ZN(n6556) );
  INV_X1 U7771 ( .A(n14504), .ZN(n8671) );
  INV_X1 U7772 ( .A(n14274), .ZN(n6558) );
  XNOR2_X2 U7773 ( .A(n8535), .B(n8543), .ZN(n9977) );
  INV_X2 U7774 ( .A(n8529), .ZN(n8535) );
  NAND3_X1 U7775 ( .A1(n6560), .A2(n8673), .A3(n6533), .ZN(n8684) );
  AND3_X1 U7776 ( .A1(n8478), .A2(n6560), .A3(n8673), .ZN(n7283) );
  NAND2_X1 U7777 ( .A1(n7660), .A2(n7774), .ZN(n6569) );
  NAND2_X1 U7778 ( .A1(n7965), .A2(n7686), .ZN(n6571) );
  OAI21_X1 U7779 ( .B1(n7965), .B2(n6574), .A(n6572), .ZN(n6575) );
  INV_X1 U7780 ( .A(n7688), .ZN(n6574) );
  NAND2_X1 U7781 ( .A1(n11390), .A2(n6577), .ZN(n6576) );
  INV_X1 U7782 ( .A(n11387), .ZN(n6577) );
  INV_X1 U7783 ( .A(n11390), .ZN(n6578) );
  NAND2_X1 U7784 ( .A1(n11389), .A2(n11390), .ZN(n11435) );
  NAND2_X1 U7785 ( .A1(n7671), .A2(n7670), .ZN(n6582) );
  NOR2_X1 U7786 ( .A1(n7412), .A2(n15082), .ZN(n6583) );
  NAND2_X1 U7787 ( .A1(n13974), .A2(n13973), .ZN(n13972) );
  INV_X1 U7788 ( .A(n13837), .ZN(n6587) );
  INV_X1 U7789 ( .A(n7230), .ZN(n8720) );
  NAND2_X2 U7790 ( .A1(n6547), .A2(n10957), .ZN(n13862) );
  AND3_X2 U7791 ( .A1(n11772), .A2(n11880), .A3(n11605), .ZN(n10957) );
  NAND3_X1 U7792 ( .A1(n11214), .A2(n10994), .A3(n10995), .ZN(n6592) );
  NAND2_X1 U7793 ( .A1(n10994), .A2(n10995), .ZN(n11168) );
  NAND3_X1 U7794 ( .A1(n11219), .A2(n11218), .A3(n6592), .ZN(n6838) );
  XNOR2_X1 U7795 ( .A(n7758), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7767) );
  INV_X2 U7796 ( .A(n15539), .ZN(n7442) );
  NAND2_X1 U7797 ( .A1(n11857), .A2(n11856), .ZN(n11862) );
  NAND2_X1 U7798 ( .A1(n8536), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U7799 ( .A1(n7610), .A2(n7612), .ZN(n11581) );
  AND3_X4 U7800 ( .A1(n7815), .A2(n7814), .A3(n7813), .ZN(n12508) );
  NAND2_X2 U7801 ( .A1(n12904), .A2(n12905), .ZN(n13391) );
  INV_X1 U7803 ( .A(n12497), .ZN(n15622) );
  NOR4_X1 U7804 ( .A1(n12677), .A2(n15228), .A3(n12671), .A4(n12672), .ZN(
        n12673) );
  NAND2_X1 U7805 ( .A1(n7784), .A2(n7783), .ZN(n7800) );
  NOR2_X2 U7806 ( .A1(n15565), .A2(n11489), .ZN(n15554) );
  NAND2_X1 U7807 ( .A1(n8939), .A2(n8938), .ZN(n11583) );
  NOR2_X1 U7808 ( .A1(n8160), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n7732) );
  INV_X1 U7809 ( .A(n9668), .ZN(n7203) );
  AOI21_X2 U7810 ( .B1(n11460), .B2(n15887), .A(n11461), .ZN(n15885) );
  NOR2_X2 U7811 ( .A1(n11460), .A2(n15887), .ZN(n11461) );
  AOI211_X2 U7812 ( .C1(n15835), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        n14614) );
  OAI21_X2 U7813 ( .B1(n14251), .B2(n14461), .A(n14250), .ZN(n14525) );
  NAND2_X1 U7814 ( .A1(n10929), .A2(n10928), .ZN(n10927) );
  NAND2_X1 U7815 ( .A1(n9679), .A2(n6870), .ZN(n9687) );
  NOR2_X2 U7816 ( .A1(n7517), .A2(n14481), .ZN(n14392) );
  OR2_X2 U7817 ( .A1(n14480), .A2(n14593), .ZN(n14481) );
  NAND2_X2 U7818 ( .A1(n14317), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U7819 ( .A1(n8542), .A2(n10567), .ZN(n6594) );
  NAND2_X1 U7820 ( .A1(n8759), .A2(n8758), .ZN(n8773) );
  NAND2_X2 U7821 ( .A1(n12058), .A2(n12062), .ZN(n12057) );
  NAND2_X1 U7822 ( .A1(n10992), .A2(n10991), .ZN(n6599) );
  AND2_X2 U7823 ( .A1(n12144), .A2(n15378), .ZN(n12058) );
  INV_X2 U7824 ( .A(n9722), .ZN(n9787) );
  NOR2_X2 U7825 ( .A1(n14394), .A2(n14562), .ZN(n14368) );
  AND2_X1 U7826 ( .A1(n12703), .A2(n12319), .ZN(n8569) );
  OR2_X1 U7827 ( .A1(n11002), .A2(n7760), .ZN(n6601) );
  NOR2_X2 U7828 ( .A1(n7526), .A2(n7724), .ZN(n7708) );
  OAI21_X2 U7829 ( .B1(n14458), .B2(n8956), .A(n8955), .ZN(n14437) );
  OAI21_X2 U7830 ( .B1(n11583), .B2(n11582), .A(n8940), .ZN(n11983) );
  NOR2_X4 U7831 ( .A1(n15102), .A2(n10129), .ZN(n15103) );
  NAND2_X1 U7833 ( .A1(n11576), .A2(n8266), .ZN(n6603) );
  BUF_X4 U7834 ( .A(n7839), .Z(n6604) );
  INV_X1 U7835 ( .A(n7859), .ZN(n7839) );
  INV_X1 U7837 ( .A(n7309), .ZN(n6606) );
  NAND2_X1 U7838 ( .A1(n12923), .A2(n7652), .ZN(n7006) );
  OR2_X1 U7839 ( .A1(n13614), .A2(n13447), .ZN(n13381) );
  OR2_X1 U7840 ( .A1(n9410), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9445) );
  INV_X1 U7841 ( .A(n7352), .ZN(n7351) );
  OAI21_X1 U7842 ( .B1(n13564), .B2(n7353), .A(n9574), .ZN(n7352) );
  OR2_X1 U7843 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  INV_X1 U7844 ( .A(n12946), .ZN(n12800) );
  NAND2_X1 U7845 ( .A1(n9018), .A2(n7256), .ZN(n7255) );
  NOR2_X1 U7846 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7256) );
  NAND2_X1 U7847 ( .A1(n10623), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U7848 ( .A1(n8367), .A2(n8366), .ZN(n8369) );
  NAND2_X1 U7849 ( .A1(n12800), .A2(n12801), .ZN(n15928) );
  NAND2_X1 U7850 ( .A1(n9173), .A2(n7360), .ZN(n7359) );
  NOR2_X1 U7851 ( .A1(n9190), .A2(n7361), .ZN(n7360) );
  INV_X1 U7852 ( .A(n9172), .ZN(n7361) );
  AOI21_X1 U7853 ( .B1(n6928), .B2(n6931), .A(n6702), .ZN(n6927) );
  OAI21_X1 U7854 ( .B1(n9815), .B2(n8535), .A(n9669), .ZN(n9681) );
  OAI21_X1 U7855 ( .B1(n12523), .B2(n12522), .A(n12521), .ZN(n12525) );
  INV_X1 U7856 ( .A(n9724), .ZN(n6810) );
  AOI21_X1 U7857 ( .B1(n12828), .B2(n12827), .A(n12826), .ZN(n12837) );
  OAI21_X1 U7858 ( .B1(n12582), .B2(n7462), .A(n7461), .ZN(n12586) );
  NAND2_X1 U7859 ( .A1(n12583), .A2(n12584), .ZN(n7461) );
  OR2_X1 U7860 ( .A1(n7463), .A2(n12581), .ZN(n7462) );
  INV_X1 U7861 ( .A(n12595), .ZN(n7482) );
  INV_X1 U7862 ( .A(n12596), .ZN(n7481) );
  MUX2_X1 U7863 ( .A(n12853), .B(n12852), .S(n9602), .Z(n12855) );
  AND2_X1 U7864 ( .A1(n7017), .A2(n6748), .ZN(n7013) );
  INV_X1 U7865 ( .A(n12879), .ZN(n7017) );
  NAND2_X1 U7866 ( .A1(n12609), .A2(n6697), .ZN(n7464) );
  AOI21_X1 U7867 ( .B1(n7218), .B2(n7216), .A(n7215), .ZN(n7214) );
  INV_X1 U7868 ( .A(n9794), .ZN(n7215) );
  OR2_X1 U7869 ( .A1(n13674), .A2(n12910), .ZN(n12911) );
  OAI21_X1 U7870 ( .B1(n7181), .B2(n12909), .A(n13365), .ZN(n12912) );
  NOR2_X1 U7871 ( .A1(n7002), .A2(n6651), .ZN(n7001) );
  INV_X1 U7872 ( .A(n7006), .ZN(n7005) );
  NAND2_X1 U7873 ( .A1(n7398), .A2(n13027), .ZN(n12866) );
  INV_X1 U7874 ( .A(n13583), .ZN(n7398) );
  AND2_X1 U7875 ( .A1(n9842), .A2(n7224), .ZN(n7223) );
  NAND2_X1 U7876 ( .A1(n7225), .A2(n9811), .ZN(n7224) );
  AND2_X1 U7877 ( .A1(n9850), .A2(n9841), .ZN(n9842) );
  NOR2_X1 U7878 ( .A1(n12465), .A2(n12452), .ZN(n12466) );
  NAND2_X1 U7879 ( .A1(n6980), .A2(n13357), .ZN(n6979) );
  OR2_X1 U7880 ( .A1(n13118), .A2(n6975), .ZN(n6974) );
  INV_X1 U7881 ( .A(n12384), .ZN(n6980) );
  NOR2_X1 U7882 ( .A1(n9216), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9230) );
  NOR2_X2 U7883 ( .A1(n13331), .A2(n13333), .ZN(n7002) );
  INV_X1 U7884 ( .A(n13723), .ZN(n9024) );
  OR2_X1 U7885 ( .A1(n9481), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9495) );
  INV_X1 U7886 ( .A(n9298), .ZN(n9285) );
  NOR2_X1 U7887 ( .A1(n15866), .A2(n12407), .ZN(n11663) );
  AND2_X1 U7888 ( .A1(n9603), .A2(n10581), .ZN(n9166) );
  AND2_X1 U7889 ( .A1(n12300), .A2(n9621), .ZN(n9630) );
  NOR2_X1 U7890 ( .A1(n9387), .A2(n7178), .ZN(n7177) );
  INV_X1 U7891 ( .A(n9376), .ZN(n7178) );
  NAND2_X1 U7892 ( .A1(n10627), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9107) );
  INV_X1 U7893 ( .A(n13766), .ZN(n7365) );
  AND2_X1 U7894 ( .A1(n13815), .A2(n13814), .ZN(n6884) );
  XNOR2_X1 U7895 ( .A(n12395), .B(n14015), .ZN(n9994) );
  NOR2_X1 U7896 ( .A1(n14218), .A2(n14225), .ZN(n7525) );
  INV_X1 U7897 ( .A(n9990), .ZN(n7305) );
  INV_X1 U7898 ( .A(n14273), .ZN(n6925) );
  NAND2_X1 U7899 ( .A1(n6930), .A2(n6931), .ZN(n6929) );
  INV_X1 U7900 ( .A(n14289), .ZN(n7296) );
  NOR2_X1 U7901 ( .A1(n14299), .A2(n7295), .ZN(n7294) );
  INV_X1 U7902 ( .A(n8965), .ZN(n7295) );
  AND2_X1 U7903 ( .A1(n7229), .A2(n8906), .ZN(n7228) );
  AND2_X1 U7904 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  NOR2_X1 U7905 ( .A1(n8348), .A2(n8347), .ZN(n8394) );
  AOI21_X1 U7906 ( .B1(n7597), .B2(n7644), .A(n6709), .ZN(n7596) );
  AND2_X1 U7907 ( .A1(n7536), .A2(n7535), .ZN(n7534) );
  AND2_X1 U7908 ( .A1(n10199), .A2(n15024), .ZN(n7536) );
  NAND2_X1 U7909 ( .A1(n6640), .A2(n10198), .ZN(n7535) );
  INV_X1 U7910 ( .A(n10136), .ZN(n7120) );
  OR2_X1 U7911 ( .A1(n10129), .A2(n15129), .ZN(n10136) );
  NOR2_X1 U7912 ( .A1(n10132), .A2(n7649), .ZN(n10133) );
  INV_X1 U7913 ( .A(n10130), .ZN(n10132) );
  INV_X1 U7914 ( .A(n7135), .ZN(n7130) );
  NAND2_X1 U7915 ( .A1(n14752), .A2(n15057), .ZN(n6869) );
  NAND2_X1 U7916 ( .A1(n8337), .A2(n8336), .ZN(n8341) );
  AND2_X1 U7917 ( .A1(n8368), .A2(n8344), .ZN(n8366) );
  NAND2_X1 U7918 ( .A1(n8231), .A2(n8252), .ZN(n8281) );
  NAND2_X1 U7919 ( .A1(n7421), .A2(n8138), .ZN(n7420) );
  NAND2_X1 U7920 ( .A1(n7422), .A2(n7424), .ZN(n7421) );
  INV_X1 U7921 ( .A(n7423), .ZN(n7422) );
  NAND2_X1 U7922 ( .A1(n7695), .A2(n10663), .ZN(n8050) );
  AOI21_X1 U7923 ( .B1(n6958), .B2(n6956), .A(n6711), .ZN(n6955) );
  INV_X1 U7924 ( .A(n6647), .ZN(n6956) );
  INV_X1 U7925 ( .A(n12979), .ZN(n11676) );
  OAI21_X1 U7926 ( .B1(n6754), .B2(n6611), .A(n7453), .ZN(n7452) );
  NAND2_X1 U7927 ( .A1(n6611), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U7928 ( .A1(n6652), .A2(n7456), .ZN(n7454) );
  NAND2_X1 U7929 ( .A1(n9474), .A2(n12904), .ZN(n13371) );
  OAI21_X1 U7930 ( .B1(n13607), .B2(n13433), .A(n13394), .ZN(n6819) );
  AND2_X1 U7931 ( .A1(n9470), .A2(n9469), .ZN(n13410) );
  OR2_X1 U7932 ( .A1(n13459), .A2(n13474), .ZN(n13440) );
  NAND2_X1 U7933 ( .A1(n13453), .A2(n9584), .ZN(n13445) );
  AND2_X1 U7934 ( .A1(n13440), .A2(n13439), .ZN(n13456) );
  OR2_X1 U7935 ( .A1(n7073), .A2(n6908), .ZN(n6907) );
  INV_X1 U7936 ( .A(n12777), .ZN(n6905) );
  AOI21_X1 U7937 ( .B1(n6659), .B2(n7265), .A(n7259), .ZN(n7258) );
  INV_X1 U7938 ( .A(n12856), .ZN(n7259) );
  XNOR2_X1 U7939 ( .A(n12847), .B(n13087), .ZN(n12850) );
  XNOR2_X1 U7940 ( .A(n13147), .B(n15935), .ZN(n12829) );
  NAND2_X1 U7941 ( .A1(n10231), .A2(n9601), .ZN(n13562) );
  INV_X1 U7942 ( .A(n9516), .ZN(n9335) );
  NAND2_X2 U7943 ( .A1(n9603), .A2(n10567), .ZN(n9516) );
  OR2_X1 U7944 ( .A1(n9022), .A2(n9019), .ZN(n9020) );
  OAI21_X1 U7945 ( .B1(n9292), .B2(n9291), .A(n9279), .ZN(n9314) );
  NOR2_X1 U7946 ( .A1(n6759), .A2(n7358), .ZN(n7357) );
  INV_X1 U7947 ( .A(n9189), .ZN(n7358) );
  INV_X1 U7948 ( .A(n9161), .ZN(n7373) );
  AND2_X1 U7949 ( .A1(n9172), .A2(n9163), .ZN(n9164) );
  AND2_X1 U7950 ( .A1(n7379), .A2(n7380), .ZN(n7375) );
  INV_X1 U7951 ( .A(n9144), .ZN(n7379) );
  AND2_X1 U7952 ( .A1(n7392), .A2(n7390), .ZN(n7389) );
  INV_X1 U7953 ( .A(n13995), .ZN(n7390) );
  INV_X1 U7954 ( .A(n9945), .ZN(n8866) );
  NAND2_X1 U7955 ( .A1(n7034), .A2(n7037), .ZN(n14199) );
  NAND2_X1 U7956 ( .A1(n9942), .A2(n9941), .ZN(n12705) );
  OR2_X1 U7957 ( .A1(n12426), .A2(n9939), .ZN(n9942) );
  NAND2_X1 U7958 ( .A1(n6786), .A2(n6620), .ZN(n14270) );
  NOR2_X1 U7959 ( .A1(n14532), .A2(n14538), .ZN(n7508) );
  OR2_X1 U7960 ( .A1(n14543), .A2(n14287), .ZN(n7297) );
  NAND2_X1 U7961 ( .A1(n8967), .A2(n8826), .ZN(n14289) );
  OR2_X1 U7962 ( .A1(n14538), .A2(n14268), .ZN(n8826) );
  AND2_X1 U7963 ( .A1(n14351), .A2(n8772), .ZN(n7617) );
  INV_X1 U7964 ( .A(n9939), .ZN(n8594) );
  NAND2_X1 U7965 ( .A1(n8972), .A2(n8971), .ZN(n15757) );
  OR2_X1 U7966 ( .A1(n8982), .A2(n8981), .ZN(n14473) );
  XNOR2_X1 U7967 ( .A(n14532), .B(n14021), .ZN(n14273) );
  AND2_X1 U7968 ( .A1(n14467), .A2(n8657), .ZN(n12014) );
  NAND2_X1 U7969 ( .A1(n10589), .A2(n6552), .ZN(n7900) );
  OR2_X1 U7970 ( .A1(n8318), .A2(n8317), .ZN(n8348) );
  INV_X1 U7971 ( .A(n8394), .ZN(n8392) );
  INV_X1 U7972 ( .A(n8396), .ZN(n8464) );
  XNOR2_X1 U7973 ( .A(n12448), .B(n15241), .ZN(n15228) );
  NAND2_X1 U7974 ( .A1(n10203), .A2(n10202), .ZN(n15006) );
  XNOR2_X1 U7975 ( .A(n15255), .B(n15016), .ZN(n15007) );
  AOI21_X1 U7976 ( .B1(n15026), .B2(n7109), .A(n6708), .ZN(n7108) );
  INV_X1 U7977 ( .A(n10138), .ZN(n7109) );
  AND2_X1 U7978 ( .A1(n7415), .A2(n7414), .ZN(n7413) );
  XNOR2_X1 U7979 ( .A(n15076), .B(n15294), .ZN(n15069) );
  OR2_X1 U7980 ( .A1(n15091), .A2(n15098), .ZN(n7414) );
  INV_X1 U7981 ( .A(n15003), .ZN(n15255) );
  INV_X1 U7982 ( .A(n15665), .ZN(n15630) );
  OR2_X1 U7983 ( .A1(n12643), .A2(n10710), .ZN(n15628) );
  NAND2_X1 U7984 ( .A1(n7739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U7985 ( .A1(n6777), .A2(n6624), .ZN(n7739) );
  NAND2_X1 U7986 ( .A1(n7487), .A2(n6689), .ZN(n10060) );
  AOI21_X1 U7987 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n10825), .A(n10031), .ZN(
        n10086) );
  NOR2_X1 U7988 ( .A1(n10084), .A2(n10083), .ZN(n10031) );
  INV_X1 U7989 ( .A(n13428), .ZN(n12975) );
  INV_X1 U7990 ( .A(n13013), .ZN(n13482) );
  NAND2_X1 U7991 ( .A1(n7446), .A2(n6667), .ZN(n12991) );
  AND2_X1 U7992 ( .A1(n9417), .A2(n9416), .ZN(n13458) );
  NAND2_X1 U7993 ( .A1(n11705), .A2(n13553), .ZN(n15870) );
  XNOR2_X1 U7994 ( .A(n13372), .B(n13371), .ZN(n13605) );
  INV_X1 U7995 ( .A(n12705), .ZN(n14515) );
  INV_X1 U7996 ( .A(n15045), .ZN(n15273) );
  INV_X1 U7997 ( .A(n14818), .ZN(n15098) );
  INV_X1 U7998 ( .A(n10027), .ZN(n10077) );
  OR2_X1 U7999 ( .A1(n9695), .A2(n9697), .ZN(n7209) );
  NOR2_X1 U8000 ( .A1(n12625), .A2(n7639), .ZN(n12493) );
  OR2_X1 U8001 ( .A1(n12528), .A2(n7486), .ZN(n7485) );
  INV_X1 U8002 ( .A(n12527), .ZN(n7486) );
  NAND2_X1 U8003 ( .A1(n9742), .A2(n9741), .ZN(n9748) );
  OR3_X1 U8004 ( .A1(n12575), .A2(n12574), .A3(n12573), .ZN(n12576) );
  AND2_X1 U8005 ( .A1(n12577), .A2(n7470), .ZN(n7467) );
  NAND2_X1 U8006 ( .A1(n12586), .A2(n12587), .ZN(n12591) );
  AND2_X1 U8007 ( .A1(n12594), .A2(n7479), .ZN(n7478) );
  NAND2_X1 U8008 ( .A1(n7482), .A2(n7481), .ZN(n7479) );
  NOR2_X1 U8009 ( .A1(n7011), .A2(n7016), .ZN(n7010) );
  AOI21_X1 U8010 ( .B1(n7013), .B2(n7014), .A(n7012), .ZN(n7011) );
  AOI21_X1 U8011 ( .B1(n12605), .B2(n12604), .A(n15120), .ZN(n6886) );
  INV_X1 U8012 ( .A(n9784), .ZN(n7219) );
  NAND2_X1 U8013 ( .A1(n9779), .A2(n9778), .ZN(n9785) );
  AND2_X1 U8014 ( .A1(n9786), .A2(n7219), .ZN(n7218) );
  INV_X1 U8015 ( .A(n7763), .ZN(n7474) );
  NAND2_X1 U8016 ( .A1(n6799), .A2(n6798), .ZN(n12459) );
  NAND2_X1 U8017 ( .A1(n12444), .A2(n12642), .ZN(n6798) );
  NAND2_X1 U8018 ( .A1(n15220), .A2(n12625), .ZN(n6799) );
  NOR2_X1 U8019 ( .A1(n11463), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U8020 ( .A1(n11765), .A2(n7333), .ZN(n7332) );
  INV_X1 U8021 ( .A(n11464), .ZN(n7333) );
  NAND2_X1 U8022 ( .A1(n13388), .A2(n9592), .ZN(n7356) );
  INV_X1 U8023 ( .A(n9589), .ZN(n6919) );
  AND2_X1 U8024 ( .A1(n7356), .A2(n7354), .ZN(n6918) );
  NOR2_X1 U8025 ( .A1(n14376), .A2(n14351), .ZN(n6834) );
  INV_X1 U8026 ( .A(n14459), .ZN(n6829) );
  NAND2_X1 U8027 ( .A1(n6832), .A2(n14254), .ZN(n6831) );
  NOR2_X1 U8028 ( .A1(n6833), .A2(n14299), .ZN(n6832) );
  NAND2_X1 U8029 ( .A1(n14273), .A2(n9987), .ZN(n6833) );
  INV_X1 U8030 ( .A(n7608), .ZN(n7607) );
  OAI21_X1 U8031 ( .B1(n8670), .B2(n7609), .A(n14475), .ZN(n7608) );
  INV_X1 U8032 ( .A(n8672), .ZN(n7609) );
  NAND2_X1 U8033 ( .A1(n12646), .A2(n12445), .ZN(n12442) );
  NAND2_X1 U8034 ( .A1(n7475), .A2(n12645), .ZN(n12443) );
  INV_X1 U8035 ( .A(n12445), .ZN(n7475) );
  NOR2_X1 U8036 ( .A1(n12478), .A2(n12477), .ZN(n12479) );
  NAND2_X1 U8037 ( .A1(n8077), .A2(SI_14_), .ZN(n8078) );
  INV_X1 U8038 ( .A(n8076), .ZN(n8081) );
  OAI21_X1 U8039 ( .B1(n10575), .B2(n10623), .A(n6867), .ZN(n7681) );
  NAND2_X1 U8040 ( .A1(n10575), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6867) );
  AND2_X1 U8041 ( .A1(n7855), .A2(n7836), .ZN(n7668) );
  OAI21_X1 U8042 ( .B1(n7676), .B2(P2_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n7661) );
  INV_X1 U8043 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10016) );
  AND2_X1 U8044 ( .A1(n9634), .A2(n6945), .ZN(n6944) );
  INV_X1 U8045 ( .A(n11657), .ZN(n6945) );
  INV_X1 U8046 ( .A(n7458), .ZN(n7457) );
  OAI21_X1 U8047 ( .B1(n7460), .B2(n7459), .A(n12177), .ZN(n7458) );
  NAND2_X1 U8048 ( .A1(n11676), .A2(n11681), .ZN(n6950) );
  INV_X1 U8049 ( .A(n7000), .ZN(n6790) );
  NAND2_X1 U8050 ( .A1(n6719), .A2(n7275), .ZN(n6789) );
  INV_X1 U8051 ( .A(n11469), .ZN(n7056) );
  INV_X1 U8052 ( .A(n7329), .ZN(n7327) );
  NOR2_X1 U8053 ( .A1(n11938), .A2(n11921), .ZN(n7329) );
  OAI21_X1 U8054 ( .B1(n12920), .B2(n7276), .A(n12918), .ZN(n7273) );
  NAND2_X1 U8055 ( .A1(n9494), .A2(n9493), .ZN(n9518) );
  AND2_X1 U8056 ( .A1(n13385), .A2(n7093), .ZN(n12908) );
  NAND2_X1 U8057 ( .A1(n9462), .A2(n9461), .ZN(n9481) );
  INV_X1 U8058 ( .A(n9463), .ZN(n9462) );
  NAND2_X1 U8059 ( .A1(n13606), .A2(n13119), .ZN(n12904) );
  NOR2_X1 U8060 ( .A1(n9445), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7092) );
  AND2_X1 U8061 ( .A1(n13381), .A2(n9588), .ZN(n13420) );
  INV_X1 U8062 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7098) );
  AND2_X1 U8063 ( .A1(n9284), .A2(n7102), .ZN(n7101) );
  INV_X1 U8064 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7102) );
  NOR2_X1 U8065 ( .A1(n9307), .A2(n7240), .ZN(n7239) );
  INV_X1 U8066 ( .A(n12865), .ZN(n7240) );
  NAND2_X1 U8067 ( .A1(n13583), .A2(n13568), .ZN(n12865) );
  INV_X1 U8068 ( .A(n12860), .ZN(n7243) );
  OR2_X1 U8069 ( .A1(n13095), .A2(n13144), .ZN(n12856) );
  AND2_X1 U8070 ( .A1(n12838), .A2(n7268), .ZN(n7267) );
  NAND2_X1 U8071 ( .A1(n9187), .A2(n12845), .ZN(n7268) );
  INV_X1 U8072 ( .A(n12830), .ZN(n7234) );
  NOR2_X1 U8073 ( .A1(n7235), .A2(n11817), .ZN(n7232) );
  NAND2_X1 U8074 ( .A1(n9120), .A2(n12796), .ZN(n11812) );
  OAI211_X1 U8075 ( .C1(n9119), .C2(SI_2_), .A(n9044), .B(n9043), .ZN(n11670)
         );
  NAND2_X1 U8076 ( .A1(n12946), .A2(n12755), .ZN(n12926) );
  NAND2_X1 U8077 ( .A1(n7085), .A2(n7089), .ZN(n7084) );
  INV_X1 U8078 ( .A(n7087), .ZN(n7085) );
  INV_X1 U8079 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U8080 ( .A1(n6947), .A2(n6948), .ZN(n6946) );
  NOR2_X1 U8081 ( .A1(n12323), .A2(P3_D_REG_0__SCAN_IN), .ZN(n6947) );
  OAI21_X1 U8082 ( .B1(n9442), .B2(n9441), .A(n9426), .ZN(n9429) );
  NAND2_X1 U8083 ( .A1(n9541), .A2(n9536), .ZN(n9544) );
  INV_X1 U8084 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9536) );
  CLKBUF_X1 U8085 ( .A(n9174), .Z(n9175) );
  INV_X1 U8086 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9322) );
  INV_X1 U8087 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9240) );
  NOR2_X1 U8088 ( .A1(n9141), .A2(n7378), .ZN(n7377) );
  NAND2_X1 U8089 ( .A1(n7072), .A2(n7071), .ZN(n9040) );
  INV_X1 U8090 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9036) );
  AND2_X1 U8091 ( .A1(n9813), .A2(n7227), .ZN(n7226) );
  INV_X1 U8092 ( .A(n9811), .ZN(n7227) );
  AND2_X1 U8093 ( .A1(n9994), .A2(n9912), .ZN(n9933) );
  NAND2_X1 U8094 ( .A1(n7041), .A2(n7043), .ZN(n7040) );
  AND2_X1 U8095 ( .A1(n14410), .A2(n8957), .ZN(n7304) );
  OR2_X1 U8096 ( .A1(n8640), .A2(n8639), .ZN(n8651) );
  AND2_X1 U8097 ( .A1(n11733), .A2(n11552), .ZN(n7611) );
  INV_X1 U8098 ( .A(n8602), .ZN(n7613) );
  INV_X1 U8099 ( .A(n8986), .ZN(n10548) );
  OR2_X1 U8100 ( .A1(n14218), .A2(n14017), .ZN(n10524) );
  INV_X1 U8101 ( .A(n7569), .ZN(n7567) );
  INV_X1 U8102 ( .A(n8450), .ZN(n8404) );
  INV_X1 U8103 ( .A(n14669), .ZN(n7601) );
  NAND2_X1 U8104 ( .A1(n7600), .A2(n14763), .ZN(n7599) );
  OR2_X1 U8105 ( .A1(n7944), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7967) );
  AND2_X1 U8106 ( .A1(n8394), .A2(n8393), .ZN(n8439) );
  NAND2_X1 U8107 ( .A1(n6650), .A2(n7133), .ZN(n7128) );
  INV_X1 U8108 ( .A(n15172), .ZN(n7126) );
  NOR2_X1 U8109 ( .A1(n15352), .A2(n12098), .ZN(n7439) );
  INV_X1 U8110 ( .A(n12057), .ZN(n7440) );
  INV_X1 U8111 ( .A(n10163), .ZN(n7547) );
  NAND2_X1 U8112 ( .A1(n11507), .A2(n15659), .ZN(n7445) );
  NAND2_X1 U8113 ( .A1(n10211), .A2(n12519), .ZN(n15539) );
  AND2_X2 U8114 ( .A1(n7748), .A2(n15428), .ZN(n7827) );
  NAND2_X1 U8115 ( .A1(n6800), .A2(n7158), .ZN(n9887) );
  AOI21_X1 U8116 ( .B1(n7160), .B2(n7162), .A(n6764), .ZN(n7158) );
  XNOR2_X1 U8117 ( .A(n9883), .B(SI_28_), .ZN(n9886) );
  NOR2_X1 U8118 ( .A1(n8386), .A2(n7164), .ZN(n7163) );
  INV_X1 U8119 ( .A(n8368), .ZN(n7164) );
  INV_X1 U8120 ( .A(n7427), .ZN(n7426) );
  OAI21_X1 U8121 ( .B1(n7429), .B2(n7428), .A(n8027), .ZN(n7427) );
  AND2_X1 U8122 ( .A1(n7430), .A2(n7690), .ZN(n7429) );
  INV_X1 U8123 ( .A(n8006), .ZN(n7430) );
  INV_X1 U8124 ( .A(n7679), .ZN(n7156) );
  INV_X1 U8125 ( .A(n7913), .ZN(n7677) );
  INV_X1 U8126 ( .A(n10051), .ZN(n7495) );
  NOR2_X1 U8127 ( .A1(n13118), .A2(n6977), .ZN(n6976) );
  INV_X1 U8128 ( .A(n13035), .ZN(n6977) );
  AOI21_X1 U8129 ( .B1(n6969), .B2(n6973), .A(n6622), .ZN(n6967) );
  AOI21_X1 U8130 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6969) );
  INV_X1 U8131 ( .A(n6976), .ZN(n6971) );
  INV_X1 U8132 ( .A(n12959), .ZN(n6970) );
  AND2_X1 U8133 ( .A1(n11047), .A2(n15869), .ZN(n11668) );
  AND2_X1 U8134 ( .A1(n13059), .A2(n11678), .ZN(n7460) );
  NAND2_X1 U8135 ( .A1(n12203), .A2(n12202), .ZN(n12254) );
  NAND2_X1 U8136 ( .A1(n9363), .A2(n9362), .ZN(n9380) );
  INV_X1 U8137 ( .A(n12304), .ZN(n6960) );
  NAND2_X1 U8138 ( .A1(n9230), .A2(n6673), .ZN(n9298) );
  INV_X1 U8139 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7090) );
  XNOR2_X1 U8140 ( .A(n6787), .B(n13316), .ZN(n12789) );
  NOR2_X1 U8141 ( .A1(n7002), .A2(n12935), .ZN(n12788) );
  OAI21_X1 U8142 ( .B1(n12792), .B2(n12791), .A(n12790), .ZN(n12793) );
  OR2_X1 U8143 ( .A1(n12716), .A2(n9531), .ZN(n12033) );
  AND4_X1 U8144 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(n12180)
         );
  INV_X1 U8145 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n11151) );
  XNOR2_X1 U8146 ( .A(n11077), .B(n11076), .ZN(n11148) );
  OAI21_X1 U8147 ( .B1(n7340), .B2(n11097), .A(n7339), .ZN(n11285) );
  AOI21_X1 U8148 ( .B1(n11252), .B2(n7341), .A(n6771), .ZN(n7339) );
  INV_X1 U8149 ( .A(n11250), .ZN(n7068) );
  NOR2_X1 U8150 ( .A1(n9337), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8151 ( .A1(n13270), .A2(n6863), .ZN(n13295) );
  OR2_X1 U8152 ( .A1(n13272), .A2(n13271), .ZN(n6863) );
  XNOR2_X1 U8153 ( .A(n13295), .B(n13294), .ZN(n13299) );
  NAND2_X1 U8154 ( .A1(n9517), .A2(n10342), .ZN(n12716) );
  INV_X1 U8155 ( .A(n9518), .ZN(n9517) );
  INV_X1 U8156 ( .A(n13402), .ZN(n13421) );
  NAND2_X1 U8157 ( .A1(n13429), .A2(n9589), .ZN(n13386) );
  OR2_X1 U8158 ( .A1(n13386), .A2(n13407), .ZN(n13409) );
  NAND2_X1 U8159 ( .A1(n13445), .A2(n9585), .ZN(n9587) );
  AOI21_X1 U8160 ( .B1(n7246), .B2(n12883), .A(n7245), .ZN(n7244) );
  INV_X1 U8161 ( .A(n12889), .ZN(n7245) );
  INV_X1 U8162 ( .A(n13456), .ZN(n9583) );
  NAND2_X1 U8163 ( .A1(n13471), .A2(n13470), .ZN(n9582) );
  INV_X1 U8164 ( .A(n13140), .ZN(n13474) );
  AOI21_X1 U8165 ( .B1(n12882), .B2(n9372), .A(n7251), .ZN(n7250) );
  OR2_X1 U8166 ( .A1(n9349), .A2(n9348), .ZN(n9372) );
  INV_X1 U8167 ( .A(n12885), .ZN(n7251) );
  OAI21_X1 U8168 ( .B1(n6614), .B2(n7077), .A(n9580), .ZN(n7076) );
  NAND2_X1 U8169 ( .A1(n7078), .A2(n9576), .ZN(n7073) );
  OR2_X1 U8170 ( .A1(n13643), .A2(n13527), .ZN(n13489) );
  CLKBUF_X1 U8171 ( .A(n13518), .Z(n6836) );
  OR2_X1 U8172 ( .A1(n13651), .A2(n13565), .ZN(n13533) );
  AND2_X1 U8173 ( .A1(n12876), .A2(n12877), .ZN(n13535) );
  AND2_X1 U8174 ( .A1(n7349), .A2(n9575), .ZN(n7079) );
  NAND2_X1 U8175 ( .A1(n7351), .A2(n7353), .ZN(n7349) );
  NAND2_X1 U8176 ( .A1(n13561), .A2(n13564), .ZN(n13563) );
  AOI21_X1 U8177 ( .B1(n7267), .B2(n7264), .A(n7263), .ZN(n7262) );
  INV_X1 U8178 ( .A(n12843), .ZN(n7263) );
  INV_X1 U8179 ( .A(n12845), .ZN(n7264) );
  INV_X1 U8180 ( .A(n7267), .ZN(n7265) );
  OR2_X1 U8181 ( .A1(n12192), .A2(n12251), .ZN(n12845) );
  NAND2_X1 U8182 ( .A1(n9171), .A2(n12841), .ZN(n12039) );
  INV_X1 U8183 ( .A(n13145), .ZN(n12251) );
  NAND2_X1 U8184 ( .A1(n11812), .A2(n12765), .ZN(n11814) );
  INV_X1 U8185 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9100) );
  AND4_X1 U8186 ( .A1(n9126), .A2(n9125), .A3(n9124), .A4(n9123), .ZN(n12183)
         );
  NAND2_X1 U8187 ( .A1(n9558), .A2(n6688), .ZN(n7080) );
  INV_X1 U8188 ( .A(n13509), .ZN(n13567) );
  INV_X1 U8189 ( .A(n13399), .ZN(n13606) );
  INV_X1 U8190 ( .A(n13511), .ZN(n13566) );
  NOR2_X1 U8191 ( .A1(n9630), .A2(n12323), .ZN(n10752) );
  INV_X1 U8192 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7253) );
  INV_X1 U8193 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9623) );
  INV_X1 U8194 ( .A(n9625), .ZN(n9627) );
  OR2_X1 U8195 ( .A1(n9618), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n9622) );
  NOR2_X1 U8196 ( .A1(n9544), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9540) );
  AOI21_X1 U8197 ( .B1(n9373), .B2(n7177), .A(n6762), .ZN(n7175) );
  INV_X1 U8198 ( .A(n7177), .ZN(n7176) );
  NAND2_X1 U8199 ( .A1(n9356), .A2(n9355), .ZN(n9375) );
  INV_X1 U8200 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9338) );
  INV_X1 U8201 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9294) );
  AOI21_X1 U8202 ( .B1(n7184), .B2(n7187), .A(n6763), .ZN(n7183) );
  XNOR2_X1 U8203 ( .A(n9276), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9254) );
  INV_X1 U8204 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U8205 ( .A1(n9210), .A2(n9209), .ZN(n9223) );
  NAND2_X1 U8206 ( .A1(n7190), .A2(n7372), .ZN(n7189) );
  NAND2_X1 U8207 ( .A1(n9110), .A2(n7375), .ZN(n7190) );
  NAND2_X1 U8208 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7381), .ZN(n7380) );
  INV_X1 U8209 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7381) );
  NAND2_X1 U8210 ( .A1(n9128), .A2(n7377), .ZN(n7376) );
  NAND2_X1 U8211 ( .A1(n9161), .A2(n9143), .ZN(n9144) );
  XNOR2_X1 U8212 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n9140) );
  NAND2_X1 U8213 ( .A1(n9111), .A2(n9110), .ZN(n9128) );
  OR2_X1 U8214 ( .A1(n9093), .A2(n9092), .ZN(n9108) );
  INV_X1 U8215 ( .A(n9040), .ZN(n9039) );
  NAND2_X1 U8216 ( .A1(n9057), .A2(n9047), .ZN(n7406) );
  NAND2_X1 U8217 ( .A1(n10614), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7405) );
  AND2_X1 U8218 ( .A1(n9036), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9057) );
  INV_X1 U8219 ( .A(n11434), .ZN(n7402) );
  XNOR2_X1 U8220 ( .A(n8181), .B(n8180), .ZN(n11480) );
  NAND2_X1 U8221 ( .A1(n11862), .A2(n7403), .ZN(n13733) );
  AND2_X1 U8222 ( .A1(n11868), .A2(n11861), .ZN(n7403) );
  XNOR2_X1 U8223 ( .A(n6599), .B(n8529), .ZN(n11164) );
  NAND2_X1 U8224 ( .A1(n7367), .A2(n7370), .ZN(n7362) );
  AND2_X1 U8225 ( .A1(n7364), .A2(n7371), .ZN(n7363) );
  NAND2_X1 U8226 ( .A1(n13880), .A2(n13881), .ZN(n7384) );
  AND4_X1 U8227 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n13958)
         );
  AND4_X1 U8228 ( .A1(n8616), .A2(n8615), .A3(n8614), .A4(n8613), .ZN(n11873)
         );
  INV_X1 U8229 ( .A(n12703), .ZN(n8516) );
  NAND2_X1 U8230 ( .A1(n14151), .A2(n7053), .ZN(n7052) );
  OR2_X1 U8231 ( .A1(n14155), .A2(n11349), .ZN(n7053) );
  INV_X1 U8232 ( .A(n7040), .ZN(n7036) );
  NAND2_X1 U8233 ( .A1(n7043), .A2(n7038), .ZN(n7037) );
  NOR2_X1 U8234 ( .A1(n14167), .A2(n14189), .ZN(n7038) );
  OAI21_X1 U8235 ( .B1(n7044), .B2(n14167), .A(n14189), .ZN(n7035) );
  OR2_X1 U8236 ( .A1(n14169), .A2(n7039), .ZN(n7034) );
  OR2_X1 U8237 ( .A1(n7040), .A2(n14189), .ZN(n7039) );
  NAND2_X1 U8238 ( .A1(n14657), .A2(n9902), .ZN(n6801) );
  AND2_X1 U8239 ( .A1(n10524), .A2(n10521), .ZN(n9990) );
  INV_X1 U8240 ( .A(n14519), .ZN(n8844) );
  OR2_X1 U8241 ( .A1(n14254), .A2(n6736), .ZN(n7604) );
  AOI21_X1 U8242 ( .B1(n7291), .B2(n7290), .A(n7289), .ZN(n7288) );
  INV_X1 U8243 ( .A(n8967), .ZN(n7289) );
  INV_X1 U8244 ( .A(n7294), .ZN(n7290) );
  NAND2_X1 U8245 ( .A1(n8966), .A2(n7294), .ZN(n7293) );
  NAND2_X1 U8246 ( .A1(n7287), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8247 ( .A1(n8961), .A2(n14351), .ZN(n7287) );
  NAND2_X1 U8248 ( .A1(n8962), .A2(n7286), .ZN(n7285) );
  INV_X1 U8249 ( .A(n8960), .ZN(n7286) );
  AND2_X1 U8250 ( .A1(n8746), .A2(n7619), .ZN(n7616) );
  NOR2_X1 U8251 ( .A1(n8769), .A2(n14374), .ZN(n7619) );
  AND2_X1 U8252 ( .A1(n8795), .A2(n8794), .ZN(n14349) );
  XNOR2_X1 U8253 ( .A(n14573), .B(n14029), .ZN(n14410) );
  OR2_X1 U8254 ( .A1(n14427), .A2(n14430), .ZN(n14428) );
  NAND2_X1 U8255 ( .A1(n8501), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8664) );
  INV_X1 U8256 ( .A(n8651), .ZN(n8501) );
  INV_X1 U8257 ( .A(n10957), .ZN(n14482) );
  INV_X1 U8258 ( .A(n8928), .ZN(n11326) );
  INV_X1 U8259 ( .A(n14471), .ZN(n14496) );
  INV_X1 U8260 ( .A(n15757), .ZN(n14461) );
  NAND2_X1 U8261 ( .A1(n12722), .A2(n15835), .ZN(n12723) );
  NAND2_X1 U8262 ( .A1(n14212), .A2(n8993), .ZN(n7277) );
  AND2_X1 U8263 ( .A1(n14215), .A2(n8992), .ZN(n8993) );
  NAND2_X1 U8264 ( .A1(n14218), .A2(n15835), .ZN(n8992) );
  NAND2_X1 U8265 ( .A1(n8848), .A2(n8847), .ZN(n14225) );
  NAND2_X1 U8266 ( .A1(n12301), .A2(n9902), .ZN(n8848) );
  OR2_X1 U8267 ( .A1(n14538), .A2(n14022), .ZN(n8827) );
  OR2_X1 U8268 ( .A1(n14274), .A2(n14273), .ZN(n7605) );
  NOR2_X1 U8269 ( .A1(n7628), .A2(n7621), .ZN(n7625) );
  NAND2_X1 U8270 ( .A1(n11604), .A2(n9902), .ZN(n6904) );
  NAND2_X1 U8271 ( .A1(n11982), .A2(n7620), .ZN(n12005) );
  AND2_X1 U8272 ( .A1(n8658), .A2(n8646), .ZN(n7620) );
  AND2_X1 U8273 ( .A1(n10563), .A2(n10799), .ZN(n10948) );
  NAND2_X1 U8274 ( .A1(n8489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7345) );
  INV_X1 U8275 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8908) );
  AND2_X1 U8276 ( .A1(n14695), .A2(n14693), .ZN(n8201) );
  AOI21_X1 U8277 ( .B1(n14754), .B2(n14753), .A(n8229), .ZN(n14677) );
  AOI21_X1 U8278 ( .B1(n6617), .B2(n7577), .A(n7572), .ZN(n7571) );
  INV_X1 U8279 ( .A(n14743), .ZN(n7572) );
  AOI21_X1 U8280 ( .B1(n11596), .B2(n7964), .A(n7585), .ZN(n7584) );
  NAND2_X1 U8281 ( .A1(n8038), .A2(n8037), .ZN(n8067) );
  NAND2_X1 U8282 ( .A1(n7570), .A2(n6757), .ZN(n7569) );
  INV_X1 U8283 ( .A(n12065), .ZN(n7570) );
  NAND2_X1 U8284 ( .A1(n7592), .A2(n7593), .ZN(n7591) );
  INV_X1 U8285 ( .A(n14732), .ZN(n7592) );
  NAND2_X1 U8286 ( .A1(n7591), .A2(n7590), .ZN(n14784) );
  NAND2_X1 U8287 ( .A1(n8102), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8168) );
  INV_X1 U8288 ( .A(n6890), .ZN(n8187) );
  INV_X1 U8289 ( .A(n12643), .ZN(n10637) );
  NOR2_X1 U8290 ( .A1(n14983), .A2(n7554), .ZN(n7553) );
  INV_X1 U8291 ( .A(n10204), .ZN(n7554) );
  NAND2_X1 U8292 ( .A1(n7534), .A2(n7532), .ZN(n7531) );
  INV_X1 U8293 ( .A(n7534), .ZN(n7533) );
  NAND2_X1 U8294 ( .A1(n15073), .A2(n7441), .ZN(n15042) );
  NOR2_X1 U8295 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  INV_X1 U8296 ( .A(n15082), .ZN(n7409) );
  OR2_X1 U8297 ( .A1(n14778), .A2(n8464), .ZN(n8294) );
  NAND2_X1 U8298 ( .A1(n15100), .A2(n10136), .ZN(n7410) );
  NAND2_X1 U8299 ( .A1(n10135), .A2(n10134), .ZN(n15100) );
  AND2_X1 U8300 ( .A1(n7127), .A2(n7136), .ZN(n7132) );
  NOR2_X1 U8301 ( .A1(n7636), .A2(n6642), .ZN(n7135) );
  AOI21_X1 U8302 ( .B1(n7540), .B2(n10167), .A(n6705), .ZN(n7539) );
  INV_X1 U8303 ( .A(n10166), .ZN(n7540) );
  NOR2_X2 U8304 ( .A1(n11912), .A2(n15389), .ZN(n12144) );
  NAND2_X1 U8305 ( .A1(n10618), .A2(n6552), .ZN(n7949) );
  NAND2_X1 U8306 ( .A1(n10113), .A2(n10112), .ZN(n11610) );
  INV_X1 U8307 ( .A(n15530), .ZN(n7116) );
  INV_X1 U8308 ( .A(n15574), .ZN(n15540) );
  NAND2_X1 U8309 ( .A1(n12511), .A2(n10157), .ZN(n7544) );
  AND2_X2 U8310 ( .A1(n7748), .A2(n7749), .ZN(n7825) );
  NAND2_X1 U8311 ( .A1(n10212), .A2(n14976), .ZN(n15235) );
  INV_X1 U8312 ( .A(n6856), .ZN(n6855) );
  OAI21_X1 U8313 ( .B1(n15682), .B2(n15237), .A(n15236), .ZN(n6856) );
  AND2_X1 U8314 ( .A1(n15228), .A2(n15225), .ZN(n7435) );
  INV_X1 U8315 ( .A(n15651), .ZN(n15568) );
  XNOR2_X1 U8316 ( .A(n9887), .B(n9886), .ZN(n14664) );
  XNOR2_X1 U8317 ( .A(n8387), .B(n8370), .ZN(n12157) );
  NAND2_X1 U8318 ( .A1(n8369), .A2(n8368), .ZN(n8387) );
  NAND2_X1 U8319 ( .A1(n8281), .A2(n8259), .ZN(n8262) );
  AND2_X1 U8320 ( .A1(n8280), .A2(n8258), .ZN(n8259) );
  NAND2_X1 U8321 ( .A1(n8281), .A2(n8280), .ZN(n8283) );
  INV_X1 U8322 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U8323 ( .A1(n10053), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U8324 ( .B1(n6982), .B2(n10054), .A(n7137), .ZN(n7496) );
  NAND2_X1 U8325 ( .A1(n14823), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8326 ( .A1(n10069), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10025) );
  INV_X1 U8327 ( .A(n6815), .ZN(n10024) );
  NAND2_X1 U8328 ( .A1(n10039), .A2(n10040), .ZN(n10028) );
  NAND2_X1 U8329 ( .A1(n6997), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6996) );
  OAI21_X1 U8330 ( .B1(n10086), .B2(n10085), .A(n7145), .ZN(n7144) );
  NAND2_X1 U8331 ( .A1(n10032), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n7145) );
  XNOR2_X1 U8332 ( .A(n10099), .B(n10098), .ZN(n10095) );
  OR2_X1 U8333 ( .A1(n15457), .A2(n7501), .ZN(n7499) );
  INV_X1 U8334 ( .A(n7503), .ZN(n7501) );
  XNOR2_X1 U8335 ( .A(n6534), .B(n13447), .ZN(n6812) );
  INV_X1 U8336 ( .A(n12980), .ZN(n6949) );
  NAND2_X1 U8337 ( .A1(n9391), .A2(n9390), .ZN(n13459) );
  NAND2_X1 U8338 ( .A1(n12981), .A2(n7460), .ZN(n13057) );
  NAND2_X1 U8339 ( .A1(n13043), .A2(n12352), .ZN(n13051) );
  NOR2_X1 U8340 ( .A1(n6621), .A2(n15867), .ZN(n7449) );
  NAND2_X1 U8341 ( .A1(n7452), .A2(n7455), .ZN(n7451) );
  NAND2_X1 U8342 ( .A1(n6611), .A2(n7456), .ZN(n7455) );
  AOI21_X1 U8343 ( .B1(n13076), .B2(n13458), .A(n12416), .ZN(n12417) );
  NAND2_X1 U8344 ( .A1(n12991), .A2(n12361), .ZN(n13070) );
  NAND2_X1 U8345 ( .A1(n9326), .A2(n9325), .ZN(n13492) );
  NOR2_X1 U8346 ( .A1(n11701), .A2(n11700), .ZN(n13110) );
  NAND2_X1 U8347 ( .A1(n12320), .A2(n9490), .ZN(n7167) );
  NAND2_X1 U8348 ( .A1(n11699), .A2(n11700), .ZN(n15874) );
  AOI21_X1 U8349 ( .B1(n12757), .B2(n12929), .A(n7274), .ZN(n12758) );
  NAND2_X1 U8350 ( .A1(n6701), .A2(n7275), .ZN(n7274) );
  NAND2_X1 U8351 ( .A1(n9440), .A2(n9439), .ZN(n13428) );
  NAND2_X1 U8352 ( .A1(n9386), .A2(n9385), .ZN(n13013) );
  NAND4_X1 U8353 ( .A1(n9208), .A2(n9207), .A3(n9206), .A4(n9205), .ZN(n13087)
         );
  NAND4_X1 U8354 ( .A1(n9139), .A2(n9138), .A3(n9137), .A4(n9136), .ZN(n13147)
         );
  NAND2_X1 U8355 ( .A1(n9066), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n6909) );
  OR2_X1 U8356 ( .A1(n11090), .A2(n11152), .ZN(n11091) );
  NAND2_X1 U8357 ( .A1(n7321), .A2(n6612), .ZN(n7319) );
  AND2_X1 U8358 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  AND2_X1 U8359 ( .A1(n7320), .A2(n13307), .ZN(n7318) );
  INV_X1 U8360 ( .A(n13326), .ZN(n7197) );
  NAND2_X1 U8361 ( .A1(n13327), .A2(n15895), .ZN(n7201) );
  AND2_X1 U8362 ( .A1(n6722), .A2(n6879), .ZN(n13604) );
  AOI21_X1 U8363 ( .B1(n13374), .B2(n13562), .A(n13373), .ZN(n6879) );
  NAND2_X1 U8364 ( .A1(n9444), .A2(n9443), .ZN(n13614) );
  INV_X1 U8365 ( .A(n13580), .ZN(n13574) );
  INV_X1 U8366 ( .A(n13588), .ZN(n13551) );
  OR2_X1 U8367 ( .A1(n11702), .A2(n11414), .ZN(n13553) );
  OR2_X1 U8368 ( .A1(n6938), .A2(n6939), .ZN(n6774) );
  INV_X1 U8369 ( .A(n13348), .ZN(n6938) );
  NAND2_X1 U8370 ( .A1(n6893), .A2(n13347), .ZN(n6939) );
  NAND2_X1 U8371 ( .A1(n9202), .A2(n9201), .ZN(n12847) );
  OR2_X1 U8372 ( .A1(n15941), .A2(n15928), .ZN(n13711) );
  OR2_X1 U8373 ( .A1(n7389), .A2(n7387), .ZN(n7385) );
  NOR2_X1 U8374 ( .A1(n7388), .A2(n7387), .ZN(n7386) );
  XNOR2_X1 U8375 ( .A(n13858), .B(n13857), .ZN(n13860) );
  AND2_X1 U8376 ( .A1(n8815), .A2(n8814), .ZN(n14287) );
  NAND2_X1 U8377 ( .A1(n11879), .A2(n9902), .ZN(n8798) );
  NAND2_X1 U8378 ( .A1(n11903), .A2(n9902), .ZN(n8829) );
  AND2_X1 U8379 ( .A1(n8785), .A2(n8784), .ZN(n14337) );
  INV_X1 U8380 ( .A(n14014), .ZN(n14000) );
  NAND2_X1 U8381 ( .A1(n8856), .A2(n8855), .ZN(n14018) );
  NAND2_X1 U8382 ( .A1(n8522), .A2(n8521), .ZN(n14020) );
  OR2_X1 U8383 ( .A1(n14257), .A2(n8975), .ZN(n8522) );
  NAND2_X1 U8384 ( .A1(n14047), .A2(n14048), .ZN(n14060) );
  NOR2_X1 U8385 ( .A1(n11963), .A2(n11962), .ZN(n14169) );
  OAI21_X1 U8386 ( .B1(n14210), .B2(n14197), .A(n7026), .ZN(n7025) );
  INV_X1 U8387 ( .A(n14208), .ZN(n7026) );
  NAND2_X1 U8388 ( .A1(n7030), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U8389 ( .A1(n14209), .A2(n15744), .ZN(n7029) );
  NAND2_X1 U8390 ( .A1(n14210), .A2(n15734), .ZN(n7030) );
  NAND2_X1 U8391 ( .A1(n12710), .A2(n12709), .ZN(n14518) );
  AND2_X1 U8392 ( .A1(n12707), .A2(n10957), .ZN(n12710) );
  OR2_X1 U8393 ( .A1(n12706), .A2(n14515), .ZN(n12707) );
  INV_X1 U8394 ( .A(n15759), .ZN(n14486) );
  NOR2_X1 U8395 ( .A1(n14520), .A2(n14521), .ZN(n6882) );
  INV_X1 U8396 ( .A(n14522), .ZN(n6883) );
  NAND2_X1 U8397 ( .A1(n12301), .A2(n6552), .ZN(n8390) );
  AND2_X1 U8398 ( .A1(n14684), .A2(n14685), .ZN(n6778) );
  AND2_X1 U8399 ( .A1(n8348), .A2(n8319), .ZN(n15044) );
  INV_X1 U8400 ( .A(n14808), .ZN(n14779) );
  OR2_X1 U8401 ( .A1(n15029), .A2(n8464), .ZN(n8355) );
  AND2_X1 U8402 ( .A1(n8432), .A2(n8431), .ZN(n15491) );
  OR2_X1 U8403 ( .A1(n11647), .A2(n15682), .ZN(n14809) );
  INV_X1 U8404 ( .A(n15495), .ZN(n14813) );
  INV_X1 U8405 ( .A(n15274), .ZN(n15015) );
  NAND2_X1 U8406 ( .A1(n8273), .A2(n8272), .ZN(n15045) );
  OR2_X1 U8407 ( .A1(n15058), .A2(n8464), .ZN(n8273) );
  OAI21_X1 U8408 ( .B1(n15085), .B2(n8464), .A(n8244), .ZN(n14818) );
  NAND2_X1 U8409 ( .A1(n8222), .A2(n8221), .ZN(n15306) );
  OR2_X1 U8410 ( .A1(n15104), .A2(n8464), .ZN(n8222) );
  INV_X1 U8411 ( .A(n14766), .ZN(n15354) );
  OAI21_X1 U8412 ( .B1(n14967), .B2(n15509), .A(n14966), .ZN(n6843) );
  AOI21_X1 U8413 ( .B1(n15006), .B2(n15007), .A(n15005), .ZN(n15258) );
  NAND2_X1 U8414 ( .A1(n15040), .A2(n15039), .ZN(n6897) );
  NAND2_X1 U8415 ( .A1(n11879), .A2(n6552), .ZN(n8237) );
  OR2_X1 U8416 ( .A1(n10219), .A2(n10213), .ZN(n15185) );
  INV_X1 U8417 ( .A(n15185), .ZN(n15582) );
  OR2_X1 U8418 ( .A1(n15584), .A2(n15563), .ZN(n15552) );
  NAND2_X1 U8419 ( .A1(n6848), .A2(n15655), .ZN(n6847) );
  INV_X1 U8420 ( .A(n15293), .ZN(n6848) );
  NAND2_X1 U8421 ( .A1(n6981), .A2(n6825), .ZN(n7487) );
  INV_X1 U8422 ( .A(n15956), .ZN(n6981) );
  AND2_X1 U8423 ( .A1(n7490), .A2(n15453), .ZN(n7489) );
  NAND2_X1 U8424 ( .A1(n6995), .A2(n6648), .ZN(n6994) );
  INV_X1 U8425 ( .A(n15462), .ZN(n6995) );
  NAND2_X1 U8426 ( .A1(n15480), .A2(n7505), .ZN(n7503) );
  XNOR2_X1 U8427 ( .A(n10095), .B(n10341), .ZN(n15457) );
  OR2_X1 U8428 ( .A1(n15480), .A2(n7505), .ZN(n7504) );
  INV_X1 U8429 ( .A(n7499), .ZN(n7500) );
  INV_X1 U8430 ( .A(n9681), .ZN(n6871) );
  NAND2_X1 U8431 ( .A1(n9695), .A2(n9697), .ZN(n7210) );
  OR2_X1 U8432 ( .A1(n15566), .A2(n12625), .ZN(n12496) );
  NAND2_X1 U8433 ( .A1(n9711), .A2(n6875), .ZN(n6874) );
  INV_X1 U8434 ( .A(n9712), .ZN(n6875) );
  OR2_X1 U8435 ( .A1(n12527), .A2(n12529), .ZN(n7484) );
  NAND2_X1 U8436 ( .A1(n9731), .A2(n6629), .ZN(n7211) );
  AND2_X1 U8437 ( .A1(n12564), .A2(n6749), .ZN(n7469) );
  NOR2_X1 U8438 ( .A1(n12583), .A2(n12584), .ZN(n7463) );
  INV_X1 U8439 ( .A(n9757), .ZN(n7207) );
  INV_X1 U8440 ( .A(n13549), .ZN(n7014) );
  INV_X1 U8441 ( .A(n12878), .ZN(n7012) );
  AOI21_X1 U8442 ( .B1(n7478), .B2(n7480), .A(n12599), .ZN(n7477) );
  NOR2_X1 U8443 ( .A1(n7482), .A2(n7481), .ZN(n7480) );
  INV_X1 U8444 ( .A(n7009), .ZN(n7008) );
  OAI21_X1 U8445 ( .B1(n6609), .B2(n6712), .A(n6625), .ZN(n7009) );
  NAND2_X1 U8446 ( .A1(n12610), .A2(n7466), .ZN(n7465) );
  MUX2_X1 U8447 ( .A(n14988), .B(n12448), .S(n12642), .Z(n12454) );
  NAND2_X1 U8448 ( .A1(n13372), .A2(n12906), .ZN(n7018) );
  NAND2_X1 U8449 ( .A1(n12898), .A2(n6623), .ZN(n7019) );
  NOR2_X1 U8450 ( .A1(n14475), .A2(n6828), .ZN(n6827) );
  NAND2_X1 U8451 ( .A1(n12014), .A2(n6758), .ZN(n6828) );
  OAI21_X1 U8452 ( .B1(n9785), .B2(n7218), .A(n6820), .ZN(n9795) );
  NOR2_X1 U8453 ( .A1(n7217), .A2(n9794), .ZN(n6820) );
  OR2_X1 U8454 ( .A1(n9869), .A2(n9825), .ZN(n9875) );
  NOR2_X1 U8455 ( .A1(n9845), .A2(n9837), .ZN(n9850) );
  NAND2_X1 U8456 ( .A1(n12440), .A2(n7472), .ZN(n12445) );
  NAND2_X1 U8457 ( .A1(n12438), .A2(n7473), .ZN(n7472) );
  NOR2_X1 U8458 ( .A1(n7474), .A2(n12441), .ZN(n7473) );
  INV_X1 U8459 ( .A(n7634), .ZN(n6975) );
  INV_X1 U8460 ( .A(n12934), .ZN(n7004) );
  OAI21_X1 U8461 ( .B1(n7002), .B2(n12933), .A(n7003), .ZN(n7000) );
  INV_X1 U8462 ( .A(n12935), .ZN(n7003) );
  NAND2_X1 U8463 ( .A1(n13535), .A2(n6894), .ZN(n9308) );
  INV_X1 U8464 ( .A(n13533), .ZN(n6894) );
  NAND2_X1 U8465 ( .A1(n9080), .A2(n12985), .ZN(n12812) );
  NAND2_X1 U8466 ( .A1(n9525), .A2(n13138), .ZN(n7089) );
  INV_X1 U8467 ( .A(n8174), .ZN(n8179) );
  INV_X1 U8468 ( .A(n10006), .ZN(n7204) );
  NAND2_X1 U8469 ( .A1(n8710), .A2(n14403), .ZN(n8735) );
  OR2_X1 U8470 ( .A1(n14573), .A2(n14029), .ZN(n8710) );
  INV_X1 U8471 ( .A(n14753), .ZN(n7575) );
  AND2_X1 U8472 ( .A1(n8306), .A2(n14742), .ZN(n8307) );
  OR2_X1 U8473 ( .A1(n10190), .A2(n15069), .ZN(n10192) );
  INV_X1 U8474 ( .A(n7161), .ZN(n7160) );
  OAI21_X1 U8475 ( .B1(n7163), .B2(n7162), .A(n8433), .ZN(n7161) );
  INV_X1 U8476 ( .A(n8385), .ZN(n7162) );
  INV_X1 U8477 ( .A(n8206), .ZN(n8210) );
  INV_X1 U8478 ( .A(n8156), .ZN(n6921) );
  OAI21_X1 U8479 ( .B1(n7648), .B2(n7424), .A(n7650), .ZN(n7423) );
  INV_X1 U8480 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n7699) );
  OAI21_X1 U8481 ( .B1(n7680), .B2(n6639), .A(n7682), .ZN(n7153) );
  NOR2_X1 U8482 ( .A1(n7156), .A2(n6639), .ZN(n7155) );
  AND2_X1 U8483 ( .A1(n10016), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10017) );
  AND2_X1 U8484 ( .A1(n9362), .A2(n7100), .ZN(n7099) );
  INV_X1 U8485 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7100) );
  INV_X1 U8486 ( .A(n9364), .ZN(n9363) );
  INV_X1 U8487 ( .A(n12965), .ZN(n6954) );
  NOR2_X1 U8488 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_REG3_REG_12__SCAN_IN), 
        .ZN(n7091) );
  NAND2_X1 U8489 ( .A1(n9039), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11087) );
  OR2_X1 U8490 ( .A1(n11096), .A2(n11248), .ZN(n11097) );
  AOI21_X1 U8491 ( .B1(n11250), .B2(n7067), .A(n7066), .ZN(n7064) );
  INV_X1 U8492 ( .A(n11262), .ZN(n7066) );
  NOR2_X1 U8493 ( .A1(n6633), .A2(n11928), .ZN(n7335) );
  NAND2_X1 U8494 ( .A1(n13220), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7344) );
  AOI21_X1 U8495 ( .B1(n13295), .B2(n6638), .A(n6772), .ZN(n7059) );
  INV_X1 U8496 ( .A(n13312), .ZN(n7060) );
  INV_X1 U8497 ( .A(n9590), .ZN(n12899) );
  NAND2_X1 U8498 ( .A1(n6721), .A2(n7356), .ZN(n6916) );
  NOR2_X1 U8499 ( .A1(n13420), .A2(n7355), .ZN(n7354) );
  INV_X1 U8500 ( .A(n9586), .ZN(n7355) );
  INV_X1 U8501 ( .A(n12778), .ZN(n6908) );
  INV_X1 U8502 ( .A(n9573), .ZN(n7353) );
  OR2_X1 U8503 ( .A1(n13707), .A2(n13545), .ZN(n13531) );
  NAND2_X1 U8504 ( .A1(n7400), .A2(n12242), .ZN(n7399) );
  INV_X1 U8505 ( .A(n12774), .ZN(n7400) );
  INV_X1 U8506 ( .A(n12854), .ZN(n7260) );
  OAI21_X1 U8507 ( .B1(n11804), .B2(n9561), .A(n9560), .ZN(n9563) );
  INV_X1 U8508 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7104) );
  INV_X1 U8509 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9132) );
  INV_X1 U8510 ( .A(n9134), .ZN(n9133) );
  INV_X1 U8511 ( .A(n12762), .ZN(n12815) );
  INV_X1 U8512 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n9081) );
  AND2_X1 U8513 ( .A1(n12812), .A2(n12813), .ZN(n11790) );
  AND3_X1 U8514 ( .A1(n9051), .A2(n9050), .A3(n9049), .ZN(n9554) );
  OR2_X1 U8515 ( .A1(n9602), .A2(n9657), .ZN(n11409) );
  INV_X1 U8516 ( .A(n9599), .ZN(n7088) );
  OR2_X1 U8517 ( .A1(n11702), .A2(n11048), .ZN(n11698) );
  INV_X1 U8518 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9016) );
  AND3_X1 U8519 ( .A1(n7083), .A2(n9174), .A3(n6737), .ZN(n9541) );
  AND2_X1 U8520 ( .A1(n7185), .A2(n9277), .ZN(n7184) );
  NAND2_X1 U8521 ( .A1(n7186), .A2(n9275), .ZN(n7185) );
  INV_X1 U8522 ( .A(n9241), .ZN(n7186) );
  INV_X1 U8523 ( .A(n9275), .ZN(n7187) );
  NAND2_X1 U8524 ( .A1(n9239), .A2(n9238), .ZN(n9242) );
  INV_X1 U8525 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9198) );
  INV_X1 U8526 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9148) );
  INV_X1 U8527 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7655) );
  INV_X1 U8528 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7656) );
  NOR2_X1 U8529 ( .A1(n13773), .A2(n13850), .ZN(n7371) );
  INV_X1 U8530 ( .A(n13848), .ZN(n7368) );
  XNOR2_X1 U8531 ( .A(n14568), .B(n13864), .ZN(n13767) );
  NOR2_X1 U8532 ( .A1(n13890), .A2(n7395), .ZN(n7394) );
  INV_X1 U8533 ( .A(n13925), .ZN(n7395) );
  NOR2_X1 U8534 ( .A1(n6831), .A2(n14318), .ZN(n6830) );
  NOR2_X1 U8535 ( .A1(n14241), .A2(n6933), .ZN(n6928) );
  NOR2_X1 U8536 ( .A1(n8969), .A2(n6934), .ZN(n6933) );
  INV_X1 U8537 ( .A(n8968), .ZN(n6934) );
  NOR2_X1 U8538 ( .A1(n7301), .A2(n7300), .ZN(n7299) );
  INV_X1 U8539 ( .A(n8957), .ZN(n7300) );
  INV_X1 U8540 ( .A(n14382), .ZN(n7303) );
  NOR2_X1 U8541 ( .A1(n13842), .A2(n7511), .ZN(n7510) );
  INV_X1 U8542 ( .A(n7512), .ZN(n7511) );
  NAND2_X1 U8543 ( .A1(n8500), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8640) );
  INV_X1 U8544 ( .A(n8624), .ZN(n8500) );
  NOR2_X1 U8545 ( .A1(n14604), .A2(n11876), .ZN(n7512) );
  NAND2_X1 U8546 ( .A1(n8499), .A2(n8498), .ZN(n8624) );
  AND2_X1 U8547 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8498) );
  INV_X1 U8548 ( .A(n8611), .ZN(n8499) );
  NAND2_X1 U8549 ( .A1(n8931), .A2(n7307), .ZN(n11551) );
  NOR2_X1 U8550 ( .A1(n8932), .A2(n7308), .ZN(n7307) );
  INV_X1 U8551 ( .A(n8930), .ZN(n7308) );
  NOR2_X1 U8552 ( .A1(n13807), .A2(n8857), .ZN(n10519) );
  AOI21_X1 U8553 ( .B1(n7607), .B2(n7609), .A(n6691), .ZN(n7606) );
  INV_X1 U8554 ( .A(n11320), .ZN(n8987) );
  NAND2_X1 U8555 ( .A1(n6547), .A2(n8919), .ZN(n10992) );
  INV_X1 U8556 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7282) );
  INV_X1 U8557 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8487) );
  INV_X1 U8558 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8486) );
  INV_X1 U8559 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8586) );
  AND2_X1 U8560 ( .A1(n8406), .A2(n8405), .ZN(n8407) );
  XNOR2_X1 U8561 ( .A(n8247), .B(n10208), .ZN(n14678) );
  AND2_X1 U8562 ( .A1(n8358), .A2(n8357), .ZN(n8360) );
  OR2_X1 U8563 ( .A1(n15267), .A2(n6537), .ZN(n8358) );
  AND2_X1 U8564 ( .A1(n8328), .A2(n8327), .ZN(n8330) );
  OR2_X1 U8565 ( .A1(n14752), .A2(n6537), .ZN(n8328) );
  INV_X1 U8566 ( .A(n14678), .ZN(n14682) );
  INV_X1 U8567 ( .A(n8299), .ZN(n14681) );
  OR2_X1 U8568 ( .A1(n15076), .A2(n6537), .ZN(n8297) );
  NOR2_X1 U8569 ( .A1(n8168), .A2(n8167), .ZN(n6890) );
  XOR2_X1 U8570 ( .A(n14971), .B(n15215), .Z(n12677) );
  AND2_X1 U8571 ( .A1(n12470), .A2(n12471), .ZN(n12488) );
  NOR2_X1 U8572 ( .A1(n12462), .A2(n12461), .ZN(n12471) );
  NOR2_X1 U8573 ( .A1(n12474), .A2(n12468), .ZN(n12469) );
  AND2_X1 U8574 ( .A1(n12481), .A2(n12480), .ZN(n6824) );
  NAND2_X1 U8575 ( .A1(n7530), .A2(n7533), .ZN(n7528) );
  INV_X1 U8576 ( .A(n6640), .ZN(n7532) );
  NOR2_X1 U8577 ( .A1(n15276), .A2(n15062), .ZN(n7441) );
  INV_X1 U8578 ( .A(n15055), .ZN(n7122) );
  AND2_X1 U8579 ( .A1(n15096), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U8580 ( .A1(n15309), .A2(n15145), .ZN(n6900) );
  NOR2_X1 U8581 ( .A1(n10172), .A2(n7556), .ZN(n7555) );
  INV_X1 U8582 ( .A(n10168), .ZN(n7556) );
  NAND2_X1 U8583 ( .A1(n12099), .A2(n10168), .ZN(n12213) );
  OR2_X1 U8584 ( .A1(n10124), .A2(n12088), .ZN(n12090) );
  NOR2_X1 U8585 ( .A1(n7541), .A2(n12657), .ZN(n7538) );
  INV_X1 U8586 ( .A(n10167), .ZN(n7541) );
  AND2_X1 U8587 ( .A1(n10157), .A2(n10154), .ZN(n7542) );
  XNOR2_X1 U8588 ( .A(n15562), .B(n12508), .ZN(n11485) );
  INV_X1 U8589 ( .A(n12491), .ZN(n10209) );
  NOR2_X1 U8590 ( .A1(n8310), .A2(n7166), .ZN(n7165) );
  INV_X1 U8591 ( .A(n8261), .ZN(n7166) );
  AOI22_X1 U8592 ( .A1(n8257), .A2(n8256), .B1(n8255), .B2(SI_21_), .ZN(n8280)
         );
  INV_X1 U8593 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7702) );
  XNOR2_X1 U8594 ( .A(n8051), .B(n10815), .ZN(n8076) );
  AND2_X1 U8595 ( .A1(n8050), .A2(n7697), .ZN(n8027) );
  NAND2_X1 U8596 ( .A1(n7694), .A2(n7693), .ZN(n8006) );
  XNOR2_X1 U8597 ( .A(n7689), .B(n10630), .ZN(n7989) );
  INV_X1 U8598 ( .A(n7966), .ZN(n7686) );
  XNOR2_X1 U8599 ( .A(n7687), .B(SI_9_), .ZN(n7966) );
  OAI21_X1 U8600 ( .B1(n10567), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n7662), .ZN(
        n7663) );
  INV_X1 U8601 ( .A(n7661), .ZN(n7662) );
  OR2_X1 U8602 ( .A1(n10023), .A2(n6816), .ZN(n6815) );
  AND2_X1 U8603 ( .A1(n10840), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8604 ( .A1(n7141), .A2(n7140), .ZN(n10042) );
  NAND2_X1 U8605 ( .A1(n10044), .A2(n11281), .ZN(n7140) );
  OAI21_X1 U8606 ( .B1(n10044), .B2(n11281), .A(P1_ADDR_REG_8__SCAN_IN), .ZN(
        n7141) );
  AND2_X1 U8607 ( .A1(n7147), .A2(n7146), .ZN(n10039) );
  NAND2_X1 U8608 ( .A1(n10853), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U8609 ( .A1(n10027), .A2(n7148), .ZN(n7147) );
  INV_X1 U8610 ( .A(n10076), .ZN(n7148) );
  OAI22_X1 U8611 ( .A1(n7144), .A2(n7143), .B1(P3_ADDR_REG_14__SCAN_IN), .B2(
        n10975), .ZN(n10091) );
  INV_X1 U8612 ( .A(n10088), .ZN(n7143) );
  XNOR2_X1 U8613 ( .A(n10097), .B(n7142), .ZN(n10099) );
  INV_X1 U8614 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U8615 ( .A1(n12356), .A2(n6679), .ZN(n7446) );
  INV_X1 U8616 ( .A(n12355), .ZN(n7447) );
  NAND2_X1 U8617 ( .A1(n12305), .A2(n12304), .ZN(n13021) );
  INV_X1 U8618 ( .A(n6754), .ZN(n7456) );
  NAND2_X1 U8619 ( .A1(n9363), .A2(n7099), .ZN(n9392) );
  NAND2_X1 U8620 ( .A1(n9230), .A2(n7091), .ZN(n9269) );
  NAND2_X1 U8621 ( .A1(n9230), .A2(n9229), .ZN(n9247) );
  OR2_X1 U8622 ( .A1(n9203), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9216) );
  OAI21_X1 U8623 ( .B1(n12980), .B2(n6950), .A(n7457), .ZN(n6951) );
  AND2_X1 U8624 ( .A1(n12033), .A2(n9608), .ZN(n12930) );
  AND4_X1 U8625 ( .A1(n9160), .A2(n9159), .A3(n9158), .A4(n9157), .ZN(n12193)
         );
  NAND2_X1 U8626 ( .A1(n6542), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9068) );
  NAND2_X1 U8627 ( .A1(n6542), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8628 ( .A1(n7058), .A2(n7057), .ZN(n11116) );
  OR2_X1 U8629 ( .A1(n11088), .A2(n9023), .ZN(n7058) );
  NAND2_X1 U8630 ( .A1(n11088), .A2(n9023), .ZN(n7057) );
  NAND2_X1 U8631 ( .A1(n6768), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U8632 ( .A1(n7315), .A2(n7316), .ZN(n7314) );
  NOR2_X1 U8633 ( .A1(n7055), .A2(n6681), .ZN(n7054) );
  NOR2_X1 U8634 ( .A1(n11268), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8635 ( .A1(n11450), .A2(n11449), .ZN(n15884) );
  AOI21_X1 U8636 ( .B1(n11757), .B2(n11928), .A(n11920), .ZN(n11758) );
  AND3_X1 U8637 ( .A1(n7336), .A2(n6633), .A3(n7337), .ZN(n11757) );
  NAND3_X1 U8638 ( .A1(n7324), .A2(n7325), .A3(n7326), .ZN(n13166) );
  OR2_X1 U8639 ( .A1(n13185), .A2(n7327), .ZN(n7326) );
  OR2_X1 U8640 ( .A1(n13165), .A2(n6766), .ZN(n7325) );
  AND2_X1 U8641 ( .A1(n7328), .A2(n13185), .ZN(n13190) );
  NAND2_X1 U8642 ( .A1(n13173), .A2(n13172), .ZN(n13204) );
  NAND2_X1 U8643 ( .A1(n13204), .A2(n6793), .ZN(n13225) );
  NOR2_X1 U8644 ( .A1(n6795), .A2(n6794), .ZN(n6793) );
  INV_X1 U8645 ( .A(n13203), .ZN(n6794) );
  INV_X1 U8646 ( .A(n13202), .ZN(n6795) );
  NAND2_X1 U8647 ( .A1(n13218), .A2(n13226), .ZN(n13258) );
  OR2_X1 U8648 ( .A1(n7344), .A2(n7343), .ZN(n13260) );
  INV_X1 U8649 ( .A(n13258), .ZN(n7343) );
  NAND2_X1 U8650 ( .A1(n13266), .A2(n6873), .ZN(n13267) );
  OR2_X1 U8651 ( .A1(n13272), .A2(n13539), .ZN(n6873) );
  NAND2_X1 U8652 ( .A1(n6612), .A2(n7323), .ZN(n13292) );
  INV_X1 U8653 ( .A(n13290), .ZN(n7322) );
  XNOR2_X1 U8654 ( .A(n7063), .B(n7062), .ZN(n13327) );
  INV_X1 U8655 ( .A(n13321), .ZN(n7062) );
  OAI21_X1 U8656 ( .B1(n13299), .B2(n7061), .A(n7059), .ZN(n7063) );
  NAND2_X1 U8657 ( .A1(n13312), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7061) );
  OAI21_X1 U8658 ( .B1(n13371), .B2(n7270), .A(n7269), .ZN(n12757) );
  INV_X1 U8659 ( .A(n7271), .ZN(n7270) );
  AND2_X1 U8660 ( .A1(n6618), .A2(n12916), .ZN(n7271) );
  NAND2_X1 U8661 ( .A1(n9597), .A2(n9596), .ZN(n13354) );
  INV_X1 U8662 ( .A(n7092), .ZN(n9447) );
  NAND2_X1 U8663 ( .A1(n7092), .A2(n9433), .ZN(n9463) );
  AND2_X1 U8664 ( .A1(n13407), .A2(n13381), .ZN(n13382) );
  NAND2_X1 U8665 ( .A1(n9587), .A2(n7354), .ZN(n13429) );
  OR2_X1 U8666 ( .A1(n13492), .A2(n13512), .ZN(n13477) );
  INV_X1 U8667 ( .A(n12881), .ZN(n13496) );
  NAND2_X1 U8668 ( .A1(n9285), .A2(n6761), .ZN(n9344) );
  OR2_X1 U8669 ( .A1(n9344), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9364) );
  AND2_X1 U8670 ( .A1(n13489), .A2(n9577), .ZN(n13517) );
  NAND2_X1 U8671 ( .A1(n7074), .A2(n9576), .ZN(n13508) );
  NAND2_X1 U8672 ( .A1(n7350), .A2(n6614), .ZN(n7074) );
  OR2_X1 U8673 ( .A1(n7238), .A2(n7239), .ZN(n7236) );
  INV_X1 U8674 ( .A(n9311), .ZN(n7238) );
  AND2_X1 U8675 ( .A1(n12861), .A2(n12860), .ZN(n12774) );
  NAND2_X1 U8676 ( .A1(n9133), .A2(n7103), .ZN(n9203) );
  AND2_X1 U8677 ( .A1(n6657), .A2(n9180), .ZN(n7103) );
  INV_X1 U8678 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U8679 ( .A1(n12829), .A2(n7234), .ZN(n7233) );
  NAND2_X1 U8680 ( .A1(n9133), .A2(n6657), .ZN(n9181) );
  NAND2_X1 U8681 ( .A1(n9133), .A2(n9132), .ZN(n9155) );
  OR2_X1 U8682 ( .A1(n9121), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9134) );
  INV_X1 U8683 ( .A(n12763), .ZN(n12821) );
  NAND2_X1 U8684 ( .A1(n9082), .A2(n9081), .ZN(n9101) );
  NAND2_X1 U8685 ( .A1(n12402), .A2(n9555), .ZN(n11777) );
  INV_X1 U8686 ( .A(n9554), .ZN(n12407) );
  NAND2_X1 U8687 ( .A1(n11692), .A2(n13713), .ZN(n11702) );
  NAND2_X1 U8688 ( .A1(n12798), .A2(n12403), .ZN(n12402) );
  AOI21_X1 U8689 ( .B1(n13422), .B2(n13430), .A(n13421), .ZN(n13616) );
  NAND2_X1 U8690 ( .A1(n9361), .A2(n9360), .ZN(n12990) );
  NAND2_X1 U8691 ( .A1(n9323), .A2(n7082), .ZN(n9034) );
  AND2_X1 U8692 ( .A1(n9018), .A2(n7254), .ZN(n7082) );
  INV_X1 U8693 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7254) );
  AOI21_X1 U8694 ( .B1(n6634), .B2(n7176), .A(n7172), .ZN(n7171) );
  INV_X1 U8695 ( .A(n9401), .ZN(n7172) );
  NAND2_X1 U8696 ( .A1(n6892), .A2(n6891), .ZN(n9259) );
  INV_X1 U8697 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n6891) );
  OR2_X1 U8698 ( .A1(n9195), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9197) );
  INV_X1 U8699 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9150) );
  OR2_X1 U8700 ( .A1(n9115), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9147) );
  OAI21_X1 U8701 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9093) );
  NAND2_X1 U8702 ( .A1(n10585), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9088) );
  AND2_X1 U8703 ( .A1(n10577), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U8704 ( .A1(n9107), .A2(n9091), .ZN(n9092) );
  INV_X1 U8705 ( .A(n7394), .ZN(n7388) );
  INV_X1 U8706 ( .A(n13804), .ZN(n7387) );
  NAND2_X1 U8707 ( .A1(n13862), .A2(n6596), .ZN(n11165) );
  OR2_X1 U8708 ( .A1(n8753), .A2(n14170), .ZN(n8779) );
  NOR2_X1 U8709 ( .A1(n13955), .A2(n7383), .ZN(n7382) );
  INV_X1 U8710 ( .A(n13882), .ZN(n7383) );
  NAND2_X1 U8711 ( .A1(n6782), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8726) );
  INV_X1 U8712 ( .A(n8678), .ZN(n6782) );
  NAND2_X1 U8713 ( .A1(n8505), .A2(n8504), .ZN(n8818) );
  INV_X1 U8714 ( .A(n8809), .ZN(n8505) );
  NAND2_X1 U8715 ( .A1(n8497), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8611) );
  INV_X1 U8716 ( .A(n8579), .ZN(n8497) );
  AND2_X1 U8717 ( .A1(n8917), .A2(n10005), .ZN(n10954) );
  INV_X1 U8718 ( .A(n7393), .ZN(n7392) );
  OAI22_X1 U8719 ( .A1(n13890), .A2(n7397), .B1(n13797), .B2(n13798), .ZN(
        n7393) );
  NAND2_X1 U8720 ( .A1(n13926), .A2(n7394), .ZN(n7391) );
  AND2_X1 U8721 ( .A1(n6547), .A2(n10002), .ZN(n6866) );
  AND2_X1 U8722 ( .A1(n9933), .A2(n7630), .ZN(n9927) );
  NOR2_X1 U8723 ( .A1(n7651), .A2(n9965), .ZN(n9966) );
  AND3_X1 U8724 ( .A1(n9933), .A2(n9932), .A3(n9931), .ZN(n7651) );
  NAND2_X1 U8725 ( .A1(n8918), .A2(n11772), .ZN(n10006) );
  INV_X1 U8726 ( .A(n10991), .ZN(n8918) );
  AND2_X1 U8727 ( .A1(n8870), .A2(n8869), .ZN(n10551) );
  NOR2_X1 U8728 ( .A1(n7050), .A2(n7049), .ZN(n7048) );
  INV_X1 U8729 ( .A(n10883), .ZN(n7049) );
  INV_X1 U8730 ( .A(n15717), .ZN(n7050) );
  OR2_X1 U8731 ( .A1(n10889), .A2(n10888), .ZN(n15733) );
  AOI22_X1 U8732 ( .A1(n11565), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11568), 
        .B2(n7052), .ZN(n11958) );
  AND2_X1 U8733 ( .A1(n14236), .A2(n7521), .ZN(n12708) );
  NOR2_X1 U8734 ( .A1(n7523), .A2(n12705), .ZN(n7521) );
  AOI21_X1 U8735 ( .B1(n8973), .B2(n9990), .A(n14461), .ZN(n8985) );
  NAND2_X1 U8736 ( .A1(n7306), .A2(n7646), .ZN(n8973) );
  INV_X1 U8737 ( .A(n14254), .ZN(n6932) );
  AND2_X1 U8738 ( .A1(n14235), .A2(n8844), .ZN(n14236) );
  NOR2_X1 U8739 ( .A1(n14270), .A2(n14527), .ZN(n14235) );
  AND2_X1 U8740 ( .A1(n8860), .A2(n8839), .ZN(n14238) );
  OR2_X1 U8741 ( .A1(n14316), .A2(n6662), .ZN(n7623) );
  OR2_X1 U8742 ( .A1(n7625), .A2(n6662), .ZN(n7622) );
  NOR3_X1 U8743 ( .A1(n6610), .A2(n14543), .A3(n14548), .ZN(n14305) );
  NOR2_X1 U8744 ( .A1(n6610), .A2(n14548), .ZN(n14304) );
  NAND2_X1 U8745 ( .A1(n14365), .A2(n8960), .ZN(n14346) );
  NAND2_X1 U8746 ( .A1(n7516), .A2(n7519), .ZN(n14420) );
  OR2_X1 U8747 ( .A1(n8726), .A2(n14154), .ZN(n8728) );
  OR2_X1 U8748 ( .A1(n8728), .A2(n13820), .ZN(n8715) );
  NOR2_X1 U8749 ( .A1(n14481), .A2(n14589), .ZN(n14452) );
  NAND2_X1 U8750 ( .A1(n6783), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8678) );
  INV_X1 U8751 ( .A(n8664), .ZN(n6783) );
  AND2_X1 U8752 ( .A1(n8989), .A2(n7510), .ZN(n14506) );
  NAND2_X1 U8753 ( .A1(n8989), .A2(n8988), .ZN(n11989) );
  AOI21_X1 U8754 ( .B1(n7613), .B2(n11733), .A(n6703), .ZN(n7612) );
  INV_X1 U8755 ( .A(n11738), .ZN(n8989) );
  NOR2_X1 U8756 ( .A1(n11321), .A2(n7515), .ZN(n11737) );
  NAND2_X1 U8757 ( .A1(n11520), .A2(n11561), .ZN(n7515) );
  NAND2_X1 U8758 ( .A1(n7514), .A2(n11520), .ZN(n11558) );
  NAND2_X1 U8759 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8579) );
  NAND2_X1 U8760 ( .A1(n6606), .A2(n14058), .ZN(n7404) );
  NOR2_X1 U8761 ( .A1(n15763), .A2(n15764), .ZN(n11369) );
  NAND2_X1 U8762 ( .A1(n8535), .A2(n11335), .ZN(n15763) );
  INV_X1 U8763 ( .A(n14473), .ZN(n14494) );
  INV_X1 U8764 ( .A(n6596), .ZN(n11158) );
  CLKBUF_X1 U8765 ( .A(n10992), .Z(n8920) );
  AND2_X1 U8766 ( .A1(n8493), .A2(n8489), .ZN(n7626) );
  INV_X1 U8767 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8493) );
  INV_X1 U8768 ( .A(n8886), .ZN(n8875) );
  OR2_X1 U8769 ( .A1(n8879), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8881) );
  AND2_X1 U8770 ( .A1(n8872), .A2(n6589), .ZN(n7229) );
  INV_X1 U8771 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8758) );
  INV_X1 U8772 ( .A(n8757), .ZN(n8759) );
  OR2_X1 U8773 ( .A1(n8617), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8619) );
  OR2_X1 U8774 ( .A1(n8589), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8603) );
  AND2_X1 U8775 ( .A1(n7911), .A2(n7910), .ZN(n11842) );
  NAND2_X1 U8776 ( .A1(n7751), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7923) );
  INV_X1 U8777 ( .A(n7921), .ZN(n7751) );
  NAND2_X1 U8778 ( .A1(n6889), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8288) );
  AND2_X1 U8779 ( .A1(n8408), .A2(n8407), .ZN(n8456) );
  INV_X1 U8780 ( .A(n6889), .ZN(n8286) );
  NOR2_X1 U8781 ( .A1(n6619), .A2(n6706), .ZN(n7565) );
  AND2_X1 U8782 ( .A1(n12229), .A2(n7570), .ZN(n7568) );
  NAND2_X1 U8783 ( .A1(n10586), .A2(n15975), .ZN(n7885) );
  NAND2_X1 U8784 ( .A1(n7750), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7921) );
  INV_X1 U8785 ( .A(n7871), .ZN(n7750) );
  AOI21_X1 U8786 ( .B1(n7596), .B2(n7598), .A(n6716), .ZN(n7595) );
  OR2_X1 U8787 ( .A1(n8133), .A2(n14723), .ZN(n8135) );
  AND2_X1 U8788 ( .A1(n8144), .A2(n8143), .ZN(n12592) );
  NAND2_X1 U8789 ( .A1(n8267), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8318) );
  INV_X1 U8790 ( .A(n8288), .ZN(n8267) );
  NOR2_X1 U8791 ( .A1(n6684), .A2(n7582), .ZN(n7581) );
  INV_X1 U8792 ( .A(n7847), .ZN(n7582) );
  INV_X1 U8793 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7973) );
  OR2_X1 U8794 ( .A1(n8214), .A2(n14755), .ZN(n8238) );
  NAND2_X1 U8795 ( .A1(n6890), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8214) );
  OAI21_X1 U8796 ( .B1(n14762), .B2(n7598), .A(n7596), .ZN(n14720) );
  AND2_X1 U8797 ( .A1(n8470), .A2(n8469), .ZN(n15241) );
  AND4_X1 U8798 ( .A1(n8072), .A2(n8071), .A3(n8070), .A4(n8069), .ZN(n14766)
         );
  INV_X1 U8799 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10013) );
  AND2_X1 U8800 ( .A1(n14878), .A2(n10694), .ZN(n14893) );
  INV_X1 U8801 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10840) );
  OR2_X1 U8802 ( .A1(n10837), .A2(n10836), .ZN(n14911) );
  OR2_X1 U8803 ( .A1(n10849), .A2(n10850), .ZN(n10708) );
  OR2_X1 U8804 ( .A1(n10822), .A2(n10823), .ZN(n10979) );
  OR2_X1 U8805 ( .A1(n11629), .A2(n11628), .ZN(n11632) );
  OR2_X1 U8806 ( .A1(n11637), .A2(n11638), .ZN(n12110) );
  INV_X1 U8807 ( .A(n7553), .ZN(n7551) );
  INV_X1 U8808 ( .A(n10205), .ZN(n7550) );
  AND2_X1 U8809 ( .A1(n15244), .A2(n15223), .ZN(n10205) );
  AND2_X1 U8810 ( .A1(n8395), .A2(n8440), .ZN(n14999) );
  NOR2_X1 U8811 ( .A1(n7434), .A2(n7433), .ZN(n7432) );
  INV_X1 U8812 ( .A(n10140), .ZN(n7433) );
  OAI21_X1 U8813 ( .B1(n15053), .B2(n10198), .A(n6640), .ZN(n15040) );
  OR2_X1 U8814 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  NAND2_X1 U8815 ( .A1(n15073), .A2(n15285), .ZN(n15041) );
  CLKBUF_X1 U8816 ( .A(n15115), .Z(n15136) );
  NOR2_X2 U8817 ( .A1(n7638), .A2(n15325), .ZN(n15141) );
  NAND2_X1 U8818 ( .A1(n7125), .A2(n6649), .ZN(n7124) );
  NAND2_X1 U8819 ( .A1(n7439), .A2(n15346), .ZN(n7438) );
  NAND2_X1 U8820 ( .A1(n7440), .A2(n7439), .ZN(n15198) );
  NAND2_X1 U8821 ( .A1(n7440), .A2(n6549), .ZN(n12218) );
  INV_X1 U8822 ( .A(n8038), .ZN(n8040) );
  XNOR2_X1 U8823 ( .A(n12562), .B(n14820), .ZN(n12660) );
  AOI21_X1 U8824 ( .B1(n7548), .B2(n7546), .A(n6666), .ZN(n10165) );
  NOR2_X1 U8825 ( .A1(n6671), .A2(n7547), .ZN(n7546) );
  NAND2_X1 U8826 ( .A1(n10165), .A2(n10164), .ZN(n11906) );
  NOR2_X1 U8827 ( .A1(n7445), .A2(n12548), .ZN(n7443) );
  NAND2_X1 U8828 ( .A1(n6888), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7951) );
  INV_X1 U8829 ( .A(n7923), .ZN(n6888) );
  NAND2_X1 U8830 ( .A1(n15511), .A2(n15512), .ZN(n7548) );
  INV_X1 U8831 ( .A(n7112), .ZN(n7111) );
  OAI21_X1 U8832 ( .B1(n6655), .B2(n7113), .A(n10110), .ZN(n7112) );
  NAND2_X1 U8833 ( .A1(n7442), .A2(n7444), .ZN(n15522) );
  NOR2_X1 U8834 ( .A1(n7445), .A2(n12538), .ZN(n7444) );
  NOR2_X1 U8835 ( .A1(n6850), .A2(n7445), .ZN(n15523) );
  INV_X1 U8836 ( .A(n15162), .ZN(n15192) );
  CLKBUF_X1 U8837 ( .A(n15539), .Z(n6850) );
  OAI22_X1 U8838 ( .A1(n11487), .A2(n11485), .B1(n12508), .B2(n15562), .ZN(
        n15547) );
  NAND2_X1 U8839 ( .A1(n10155), .A2(n10154), .ZN(n15545) );
  INV_X1 U8840 ( .A(n12511), .ZN(n15546) );
  INV_X1 U8841 ( .A(n15566), .ZN(n12495) );
  OR2_X1 U8842 ( .A1(n14986), .A2(n8464), .ZN(n8447) );
  AND2_X1 U8843 ( .A1(n8378), .A2(n8377), .ZN(n15251) );
  NAND2_X1 U8844 ( .A1(n10139), .A2(n10138), .ZN(n15027) );
  AND3_X1 U8845 ( .A1(n8172), .A2(n8171), .A3(n8170), .ZN(n15322) );
  AND2_X1 U8846 ( .A1(n11007), .A2(n10147), .ZN(n15395) );
  NAND2_X1 U8847 ( .A1(n9938), .A2(n9892), .ZN(n9895) );
  NOR2_X1 U8848 ( .A1(n7743), .A2(n15419), .ZN(n6895) );
  XNOR2_X1 U8849 ( .A(n9901), .B(n9900), .ZN(n12318) );
  NAND2_X1 U8850 ( .A1(n7159), .A2(n8385), .ZN(n8434) );
  NAND2_X1 U8851 ( .A1(n8369), .A2(n7163), .ZN(n7159) );
  NAND2_X1 U8852 ( .A1(n8233), .A2(n8232), .ZN(n8235) );
  XNOR2_X1 U8853 ( .A(n8159), .B(n8158), .ZN(n11402) );
  AND2_X1 U8854 ( .A1(n8062), .A2(n8034), .ZN(n10981) );
  OR2_X1 U8855 ( .A1(n8008), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7721) );
  XNOR2_X1 U8856 ( .A(n8007), .B(n8006), .ZN(n10657) );
  NAND2_X1 U8857 ( .A1(n7431), .A2(n7690), .ZN(n8007) );
  OAI21_X1 U8858 ( .B1(n7408), .B2(n7894), .A(n7157), .ZN(n7943) );
  AOI21_X1 U8859 ( .B1(n7680), .B2(n7156), .A(n6639), .ZN(n7157) );
  OR2_X1 U8860 ( .A1(n7914), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U8861 ( .A1(n7408), .A2(n7679), .ZN(n7893) );
  XNOR2_X1 U8862 ( .A(n6982), .B(n10055), .ZN(n10057) );
  NAND2_X1 U8863 ( .A1(n6653), .A2(n10015), .ZN(n10050) );
  INV_X1 U8864 ( .A(n10060), .ZN(n10062) );
  XNOR2_X1 U8865 ( .A(n6815), .B(n11309), .ZN(n10069) );
  OAI22_X1 U8866 ( .A1(n10042), .A2(n10041), .B1(n15899), .B2(
        P1_ADDR_REG_9__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U8867 ( .A1(n7488), .A2(n7492), .ZN(n6988) );
  OR2_X1 U8868 ( .A1(n15450), .A2(n7491), .ZN(n7488) );
  NAND2_X1 U8869 ( .A1(n7493), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U8870 ( .A1(n15452), .A2(n6988), .ZN(n10081) );
  AOI21_X1 U8871 ( .B1(n13349), .B2(n9524), .A(n9523), .ZN(n13358) );
  NAND2_X1 U8872 ( .A1(n6968), .A2(n6972), .ZN(n12958) );
  OAI21_X1 U8873 ( .B1(n12305), .B2(n6957), .A(n6955), .ZN(n12966) );
  AND4_X1 U8874 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(n13085)
         );
  NAND2_X1 U8875 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  AND2_X1 U8876 ( .A1(n7446), .A2(n6656), .ZN(n12993) );
  OAI21_X1 U8877 ( .B1(n6967), .B2(n6978), .A(n6963), .ZN(n6962) );
  NAND2_X1 U8878 ( .A1(n6967), .A2(n6964), .ZN(n6963) );
  NAND2_X1 U8879 ( .A1(n6965), .A2(n12387), .ZN(n6964) );
  INV_X1 U8880 ( .A(n6969), .ZN(n6965) );
  NAND2_X1 U8881 ( .A1(n6967), .A2(n12387), .ZN(n6966) );
  NAND2_X1 U8882 ( .A1(n11748), .A2(n11669), .ZN(n11747) );
  NAND2_X1 U8883 ( .A1(n13068), .A2(n12364), .ZN(n13011) );
  NAND2_X1 U8884 ( .A1(n13125), .A2(n12349), .ZN(n13042) );
  AND2_X1 U8885 ( .A1(n12981), .A2(n11678), .ZN(n13058) );
  NAND2_X1 U8886 ( .A1(n6959), .A2(n12309), .ZN(n12345) );
  NAND2_X1 U8887 ( .A1(n12305), .A2(n6647), .ZN(n6959) );
  NAND2_X1 U8888 ( .A1(n9409), .A2(n9408), .ZN(n13080) );
  INV_X1 U8889 ( .A(n13143), .ZN(n13090) );
  NAND2_X1 U8890 ( .A1(n11716), .A2(n11717), .ZN(n11715) );
  NAND2_X1 U8891 ( .A1(n12356), .A2(n12355), .ZN(n13098) );
  NAND2_X1 U8892 ( .A1(n12789), .A2(n12801), .ZN(n12795) );
  AND2_X1 U8893 ( .A1(n12033), .A2(n12032), .ZN(n13333) );
  AND2_X1 U8894 ( .A1(n12033), .A2(n9535), .ZN(n13345) );
  NAND2_X1 U8895 ( .A1(n9502), .A2(n9501), .ZN(n13343) );
  NAND2_X1 U8896 ( .A1(n13375), .A2(n9524), .ZN(n7094) );
  INV_X1 U8897 ( .A(n13410), .ZN(n13119) );
  NAND2_X1 U8898 ( .A1(n9399), .A2(n9398), .ZN(n13140) );
  NAND2_X1 U8899 ( .A1(n9370), .A2(n9369), .ZN(n13499) );
  INV_X1 U8900 ( .A(P3_U3897), .ZN(n13142) );
  OR2_X1 U8901 ( .A1(n11181), .A2(n12410), .ZN(n11183) );
  NAND2_X1 U8902 ( .A1(n11064), .A2(n11063), .ZN(n11125) );
  NAND2_X1 U8903 ( .A1(n11093), .A2(n11127), .ZN(n11131) );
  NAND2_X1 U8904 ( .A1(n7195), .A2(n11246), .ZN(n11271) );
  NAND2_X1 U8905 ( .A1(n7065), .A2(n11250), .ZN(n11263) );
  NAND2_X1 U8906 ( .A1(n11247), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7065) );
  OAI21_X1 U8907 ( .B1(n15884), .B2(n15880), .A(n15881), .ZN(n11454) );
  XNOR2_X1 U8908 ( .A(n11918), .B(n11928), .ZN(n7070) );
  INV_X1 U8909 ( .A(n6892), .ZN(n9243) );
  NOR2_X1 U8910 ( .A1(n11765), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7069) );
  OAI22_X1 U8911 ( .A1(n13242), .A2(n13241), .B1(n13247), .B2(n13240), .ZN(
        n13244) );
  NAND2_X1 U8912 ( .A1(n7319), .A2(n7320), .ZN(n13308) );
  OAI22_X1 U8913 ( .A1(n13299), .A2(n13298), .B1(n13296), .B2(n13297), .ZN(
        n13313) );
  INV_X1 U8914 ( .A(n13295), .ZN(n13296) );
  NAND2_X1 U8915 ( .A1(n12297), .A2(n9490), .ZN(n9460) );
  NAND2_X1 U8916 ( .A1(n13393), .A2(n6818), .ZN(n13609) );
  INV_X1 U8917 ( .A(n6819), .ZN(n6818) );
  AND2_X1 U8918 ( .A1(n13574), .A2(n11776), .ZN(n13418) );
  NAND2_X1 U8919 ( .A1(n9582), .A2(n9581), .ZN(n13455) );
  NAND2_X1 U8920 ( .A1(n7249), .A2(n7246), .ZN(n13465) );
  NAND2_X1 U8921 ( .A1(n6836), .A2(n12882), .ZN(n7249) );
  OAI22_X1 U8922 ( .A1(n7350), .A2(n7073), .B1(n7075), .B2(n9579), .ZN(n13479)
         );
  INV_X1 U8923 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U8924 ( .A1(n9341), .A2(n9340), .ZN(n13643) );
  NAND2_X1 U8925 ( .A1(n9283), .A2(n9282), .ZN(n13541) );
  NAND2_X1 U8926 ( .A1(n7350), .A2(n7079), .ZN(n13526) );
  NAND2_X1 U8927 ( .A1(n9297), .A2(n9296), .ZN(n13651) );
  NAND2_X1 U8928 ( .A1(n13563), .A2(n9573), .ZN(n13544) );
  NAND2_X1 U8929 ( .A1(n9215), .A2(n9214), .ZN(n13095) );
  NAND2_X1 U8930 ( .A1(n7261), .A2(n7262), .ZN(n12080) );
  OR2_X1 U8931 ( .A1(n12039), .A2(n7265), .ZN(n7261) );
  NAND2_X1 U8932 ( .A1(n7266), .A2(n12845), .ZN(n11995) );
  OR2_X1 U8933 ( .A1(n12039), .A2(n9187), .ZN(n7266) );
  NAND2_X1 U8934 ( .A1(n11814), .A2(n12830), .ZN(n11948) );
  INV_X1 U8935 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U8936 ( .A1(n13574), .A2(n12082), .ZN(n13588) );
  INV_X1 U8937 ( .A(n13553), .ZN(n13579) );
  INV_X1 U8938 ( .A(n13582), .ZN(n13557) );
  INV_X1 U8939 ( .A(n13601), .ZN(n13660) );
  INV_X1 U8940 ( .A(n13331), .ZN(n13663) );
  NAND2_X1 U8941 ( .A1(n13604), .A2(n6877), .ZN(n13677) );
  INV_X1 U8942 ( .A(n6878), .ZN(n6877) );
  OAI21_X1 U8943 ( .B1(n13605), .B2(n15930), .A(n13603), .ZN(n6878) );
  INV_X1 U8944 ( .A(n13080), .ZN(n13687) );
  NAND2_X1 U8945 ( .A1(n9246), .A2(n9245), .ZN(n13583) );
  AND2_X1 U8946 ( .A1(n9179), .A2(n9178), .ZN(n12192) );
  INV_X1 U8947 ( .A(n13711), .ZN(n13675) );
  AND2_X1 U8948 ( .A1(n11069), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13713) );
  INV_X1 U8949 ( .A(n9025), .ZN(n12742) );
  NAND2_X1 U8950 ( .A1(n6837), .A2(n6857), .ZN(n13723) );
  NOR2_X1 U8951 ( .A1(n9627), .A2(n9626), .ZN(n9628) );
  OR2_X1 U8952 ( .A1(n9624), .A2(n9623), .ZN(n9629) );
  NOR2_X1 U8953 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n9626) );
  NAND2_X1 U8954 ( .A1(n7170), .A2(n7169), .ZN(n7168) );
  INV_X1 U8955 ( .A(n9478), .ZN(n7169) );
  INV_X1 U8956 ( .A(n9479), .ZN(n7170) );
  NAND2_X1 U8957 ( .A1(n9619), .A2(n9622), .ZN(n12300) );
  AND2_X1 U8958 ( .A1(n9476), .A2(n9458), .ZN(n12297) );
  OR2_X1 U8959 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U8960 ( .A1(n9430), .A2(n7194), .ZN(n9453) );
  AND2_X1 U8961 ( .A1(n7020), .A2(n9631), .ZN(n12946) );
  NAND2_X1 U8962 ( .A1(n7174), .A2(n7175), .ZN(n9402) );
  OR2_X1 U8963 ( .A1(n9375), .A2(n7176), .ZN(n7174) );
  NAND2_X1 U8964 ( .A1(n7179), .A2(n9376), .ZN(n9388) );
  NAND2_X1 U8965 ( .A1(n9375), .A2(n9374), .ZN(n7179) );
  INV_X1 U8966 ( .A(SI_11_), .ZN(n10651) );
  INV_X1 U8967 ( .A(SI_10_), .ZN(n10630) );
  NAND2_X1 U8968 ( .A1(n7359), .A2(n9189), .ZN(n9192) );
  NAND2_X1 U8969 ( .A1(n7188), .A2(n7372), .ZN(n9165) );
  NAND2_X1 U8970 ( .A1(n9111), .A2(n7192), .ZN(n7188) );
  INV_X1 U8971 ( .A(n7190), .ZN(n7192) );
  NAND2_X1 U8972 ( .A1(n7376), .A2(n7375), .ZN(n9162) );
  NAND2_X1 U8973 ( .A1(n7376), .A2(n7380), .ZN(n9145) );
  NAND2_X1 U8974 ( .A1(n9127), .A2(n9128), .ZN(n9142) );
  NAND2_X1 U8975 ( .A1(n9039), .A2(n9041), .ZN(n9076) );
  NAND2_X1 U8976 ( .A1(n7406), .A2(n7405), .ZN(n9071) );
  NOR2_X1 U8977 ( .A1(n11525), .A2(n7402), .ZN(n7401) );
  AND4_X1 U8978 ( .A1(n8645), .A2(n8644), .A3(n8643), .A4(n8642), .ZN(n13839)
         );
  NAND2_X1 U8979 ( .A1(n11862), .A2(n11861), .ZN(n11871) );
  NAND2_X1 U8980 ( .A1(n10993), .A2(n7647), .ZN(n10994) );
  AOI21_X1 U8981 ( .B1(n13926), .B2(n13925), .A(n7396), .ZN(n13891) );
  INV_X1 U8982 ( .A(n13765), .ZN(n7366) );
  NAND2_X1 U8983 ( .A1(n6864), .A2(n13766), .ZN(n7369) );
  AND2_X1 U8984 ( .A1(n8825), .A2(n8824), .ZN(n14268) );
  INV_X1 U8985 ( .A(n11234), .ZN(n11231) );
  INV_X1 U8986 ( .A(n13862), .ZN(n13800) );
  NAND2_X1 U8987 ( .A1(n7384), .A2(n13882), .ZN(n13956) );
  CLKBUF_X1 U8988 ( .A(n13824), .Z(n13965) );
  AND4_X1 U8989 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), .ZN(n13977)
         );
  NAND2_X1 U8990 ( .A1(n11435), .A2(n11434), .ZN(n11524) );
  NAND2_X1 U8991 ( .A1(n7391), .A2(n7392), .ZN(n13996) );
  NAND2_X1 U8992 ( .A1(n12157), .A2(n9902), .ZN(n8837) );
  AND2_X1 U8993 ( .A1(n10953), .A2(n14406), .ZN(n14014) );
  INV_X1 U8994 ( .A(n14002), .ZN(n14004) );
  AOI21_X1 U8995 ( .B1(n10009), .B2(n11605), .A(n10004), .ZN(n10010) );
  AND2_X1 U8996 ( .A1(n8980), .A2(n8979), .ZN(n11213) );
  INV_X1 U8997 ( .A(n10551), .ZN(n14017) );
  INV_X1 U8998 ( .A(n13958), .ZN(n14495) );
  AND3_X1 U8999 ( .A1(n8547), .A2(n8546), .A3(n8545), .ZN(n8548) );
  NAND2_X1 U9000 ( .A1(n14060), .A2(n14059), .ZN(n10870) );
  NAND2_X1 U9001 ( .A1(n10881), .A2(n10880), .ZN(n14134) );
  NAND2_X1 U9002 ( .A1(n7048), .A2(n14134), .ZN(n15716) );
  OAI22_X1 U9003 ( .A1(n7048), .A2(n7047), .B1(n7046), .B2(n7045), .ZN(n14147)
         );
  INV_X1 U9004 ( .A(n10885), .ZN(n7047) );
  NAND2_X1 U9005 ( .A1(n10880), .A2(n10885), .ZN(n7045) );
  INV_X1 U9006 ( .A(n10881), .ZN(n7046) );
  OR2_X1 U9007 ( .A1(n14138), .A2(n14139), .ZN(n14140) );
  NAND2_X1 U9008 ( .A1(n14153), .A2(n14152), .ZN(n14151) );
  OR2_X1 U9009 ( .A1(n14159), .A2(n14158), .ZN(n14160) );
  XNOR2_X1 U9010 ( .A(n7052), .B(n7051), .ZN(n11565) );
  OAI21_X1 U9011 ( .B1(n14169), .B2(n6637), .A(n14167), .ZN(n14181) );
  AOI21_X1 U9012 ( .B1(n14169), .B2(n7033), .A(n7032), .ZN(n7031) );
  INV_X1 U9013 ( .A(n7035), .ZN(n7033) );
  OAI21_X1 U9014 ( .B1(n7035), .B2(n7036), .A(n7037), .ZN(n7032) );
  INV_X1 U9015 ( .A(n14211), .ZN(n7022) );
  NAND2_X1 U9016 ( .A1(n14664), .A2(n9902), .ZN(n8859) );
  NAND2_X1 U9017 ( .A1(n7615), .A2(n10271), .ZN(n14223) );
  NAND2_X1 U9018 ( .A1(n6936), .A2(n8968), .ZN(n14249) );
  NAND2_X1 U9019 ( .A1(n7603), .A2(n7604), .ZN(n14253) );
  INV_X1 U9020 ( .A(n14270), .ZN(n8990) );
  NAND2_X1 U9021 ( .A1(n7293), .A2(n7297), .ZN(n14284) );
  NAND2_X1 U9022 ( .A1(n8966), .A2(n8965), .ZN(n14300) );
  AOI21_X1 U9023 ( .B1(n14384), .B2(n6654), .A(n7284), .ZN(n14333) );
  AND2_X1 U9024 ( .A1(n7618), .A2(n8772), .ZN(n14352) );
  AND2_X1 U9025 ( .A1(n14428), .A2(n8957), .ZN(n14411) );
  NAND2_X1 U9026 ( .A1(n14502), .A2(n8672), .ZN(n14476) );
  NAND2_X1 U9027 ( .A1(n8931), .A2(n8930), .ZN(n11515) );
  NAND2_X1 U9028 ( .A1(n15781), .A2(n10945), .ZN(n14406) );
  OR2_X1 U9029 ( .A1(n8542), .A2(n10867), .ZN(n8526) );
  NOR2_X1 U9030 ( .A1(n14484), .A2(n10541), .ZN(n15759) );
  NAND2_X1 U9031 ( .A1(n14518), .A2(n14517), .ZN(n14609) );
  OAI21_X1 U9032 ( .B1(n14515), .B2(n15843), .A(n14514), .ZN(n14516) );
  NAND2_X1 U9033 ( .A1(n12724), .A2(n12723), .ZN(n12725) );
  NAND2_X1 U9034 ( .A1(n7625), .A2(n7624), .ZN(n14297) );
  INV_X1 U9035 ( .A(n14314), .ZN(n7624) );
  NAND2_X1 U9036 ( .A1(n11982), .A2(n8646), .ZN(n12007) );
  AND2_X1 U9037 ( .A1(n10948), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15781) );
  INV_X1 U9038 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11177) );
  INV_X1 U9039 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11037) );
  INV_X1 U9040 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10939) );
  INV_X1 U9041 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10751) );
  INV_X1 U9042 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10659) );
  XNOR2_X1 U9043 ( .A(n8661), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11352) );
  INV_X1 U9044 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10591) );
  INV_X1 U9045 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10588) );
  INV_X1 U9046 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10596) );
  INV_X1 U9047 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10585) );
  INV_X1 U9048 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10593) );
  XNOR2_X1 U9049 ( .A(n8550), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14049) );
  INV_X1 U9050 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10614) );
  AND4_X1 U9051 ( .A1(n8045), .A2(n8044), .A3(n8043), .A4(n8042), .ZN(n14673)
         );
  NAND2_X1 U9052 ( .A1(n12129), .A2(n12126), .ZN(n12067) );
  AND2_X1 U9053 ( .A1(n8201), .A2(n7589), .ZN(n7588) );
  NAND2_X1 U9054 ( .A1(n7590), .A2(n8152), .ZN(n7589) );
  AND2_X1 U9055 ( .A1(n8457), .A2(n15491), .ZN(n6803) );
  INV_X1 U9056 ( .A(n15362), .ZN(n12565) );
  NOR2_X1 U9057 ( .A1(n7563), .A2(n7562), .ZN(n7561) );
  INV_X1 U9058 ( .A(n12289), .ZN(n7562) );
  INV_X1 U9059 ( .A(n7565), .ZN(n7563) );
  AND2_X1 U9060 ( .A1(n7564), .A2(n7565), .ZN(n12290) );
  AND3_X1 U9061 ( .A1(n8107), .A2(n8106), .A3(n8105), .ZN(n15321) );
  NOR2_X1 U9062 ( .A1(n14762), .A2(n14763), .ZN(n14761) );
  NAND3_X1 U9063 ( .A1(n14774), .A2(n14776), .A3(n14773), .ZN(n14775) );
  AND4_X1 U9064 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(n15384)
         );
  NAND2_X1 U9065 ( .A1(n7566), .A2(n7569), .ZN(n12230) );
  AND2_X1 U9066 ( .A1(n7591), .A2(n6663), .ZN(n14785) );
  XNOR2_X1 U9067 ( .A(n8392), .B(P1_REG3_REG_26__SCAN_IN), .ZN(n15017) );
  AND2_X1 U9068 ( .A1(n8459), .A2(n8458), .ZN(n12698) );
  INV_X1 U9069 ( .A(n12701), .ZN(n6781) );
  INV_X1 U9070 ( .A(n15242), .ZN(n15016) );
  INV_X1 U9071 ( .A(n14673), .ZN(n15363) );
  INV_X1 U9072 ( .A(n15629), .ZN(n15647) );
  NAND2_X1 U9073 ( .A1(n10690), .A2(n10689), .ZN(n14876) );
  AND2_X1 U9074 ( .A1(n14913), .A2(n10699), .ZN(n10787) );
  AND2_X1 U9075 ( .A1(n7970), .A2(n7992), .ZN(n14924) );
  INV_X1 U9076 ( .A(n14962), .ZN(n15504) );
  NAND2_X1 U9077 ( .A1(n15004), .A2(n10204), .ZN(n14982) );
  AND2_X1 U9078 ( .A1(n15004), .A2(n7553), .ZN(n14981) );
  NAND2_X1 U9079 ( .A1(n7529), .A2(n7530), .ZN(n15012) );
  OR2_X1 U9080 ( .A1(n15053), .A2(n7533), .ZN(n7529) );
  NAND2_X1 U9081 ( .A1(n7107), .A2(n7108), .ZN(n15011) );
  NAND2_X1 U9082 ( .A1(n7411), .A2(n7417), .ZN(n15056) );
  NAND2_X1 U9083 ( .A1(n7416), .A2(n7413), .ZN(n7411) );
  XNOR2_X1 U9084 ( .A(n6849), .B(n7415), .ZN(n15070) );
  NAND2_X1 U9085 ( .A1(n7416), .A2(n7414), .ZN(n6849) );
  AOI21_X1 U9086 ( .B1(n7437), .B2(n15091), .A(n15574), .ZN(n15084) );
  INV_X1 U9087 ( .A(n15103), .ZN(n7437) );
  INV_X1 U9088 ( .A(n7410), .ZN(n15080) );
  NAND2_X1 U9089 ( .A1(n10187), .A2(n10186), .ZN(n15109) );
  NAND2_X1 U9090 ( .A1(n11480), .A2(n6552), .ZN(n8185) );
  NOR2_X1 U9091 ( .A1(n7135), .A2(n12274), .ZN(n7134) );
  AOI21_X1 U9092 ( .B1(n10128), .B2(n7636), .A(n6642), .ZN(n12275) );
  INV_X1 U9093 ( .A(n15552), .ZN(n15212) );
  CLKBUF_X1 U9094 ( .A(n12048), .Z(n12049) );
  NAND2_X1 U9095 ( .A1(n10653), .A2(n6552), .ZN(n7995) );
  NAND2_X1 U9096 ( .A1(n10149), .A2(n10645), .ZN(n15549) );
  NAND2_X1 U9097 ( .A1(n7115), .A2(n10109), .ZN(n11501) );
  NAND2_X1 U9098 ( .A1(n7116), .A2(n6655), .ZN(n7115) );
  NAND2_X1 U9099 ( .A1(n10594), .A2(n15975), .ZN(n7865) );
  NAND2_X1 U9100 ( .A1(n10219), .A2(n15549), .ZN(n15178) );
  CLKBUF_X1 U9101 ( .A(n12495), .Z(n6804) );
  INV_X1 U9102 ( .A(n15714), .ZN(n15711) );
  NAND2_X1 U9103 ( .A1(n15216), .A2(n6853), .ZN(n15396) );
  INV_X1 U9104 ( .A(n6854), .ZN(n6853) );
  OAI21_X1 U9105 ( .B1(n15217), .B2(n15682), .A(n15218), .ZN(n6854) );
  NAND2_X1 U9106 ( .A1(n15219), .A2(n6807), .ZN(n15397) );
  INV_X1 U9107 ( .A(n6808), .ZN(n6807) );
  OAI21_X1 U9108 ( .B1(n15220), .B2(n15682), .A(n15218), .ZN(n6808) );
  AOI21_X1 U9109 ( .B1(n15281), .B2(n15568), .A(n15280), .ZN(n15282) );
  AND2_X1 U9110 ( .A1(n7710), .A2(n7743), .ZN(n7557) );
  INV_X1 U9111 ( .A(n7714), .ZN(n7711) );
  NAND2_X1 U9112 ( .A1(n8262), .A2(n8261), .ZN(n8311) );
  NAND2_X1 U9113 ( .A1(n8805), .A2(n10567), .ZN(n8284) );
  INV_X1 U9114 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11178) );
  INV_X1 U9115 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11038) );
  INV_X1 U9116 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10661) );
  INV_X1 U9117 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10619) );
  INV_X1 U9118 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10625) );
  INV_X1 U9119 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10627) );
  INV_X1 U9120 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10577) );
  OAI21_X1 U9121 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7811) );
  XNOR2_X1 U9122 ( .A(n10057), .B(n10056), .ZN(n15970) );
  INV_X1 U9123 ( .A(n7496), .ZN(n10052) );
  XNOR2_X1 U9124 ( .A(n10044), .B(n10043), .ZN(n15448) );
  NAND2_X1 U9125 ( .A1(n6990), .A2(n6991), .ZN(n15470) );
  AOI21_X1 U9126 ( .B1(n6993), .B2(n6992), .A(n6717), .ZN(n6991) );
  INV_X1 U9127 ( .A(n6648), .ZN(n6992) );
  INV_X1 U9128 ( .A(n7144), .ZN(n10089) );
  XNOR2_X1 U9129 ( .A(n12417), .B(n6812), .ZN(n12978) );
  NAND2_X1 U9130 ( .A1(n13057), .A2(n11681), .ZN(n12178) );
  NAND2_X1 U9131 ( .A1(n7451), .A2(n13128), .ZN(n7450) );
  NAND2_X1 U9132 ( .A1(n11269), .A2(n11268), .ZN(n11470) );
  AND2_X1 U9133 ( .A1(n7319), .A2(n7318), .ZN(n13310) );
  NAND2_X1 U9134 ( .A1(n10238), .A2(n15954), .ZN(n9667) );
  OAI21_X1 U9135 ( .B1(n13669), .B2(n15951), .A(n6940), .ZN(P3_U3487) );
  INV_X1 U9136 ( .A(n6941), .ZN(n6940) );
  INV_X1 U9137 ( .A(n6774), .ZN(n13669) );
  OAI22_X1 U9138 ( .A1(n13671), .A2(n13660), .B1(n15954), .B2(n13596), .ZN(
        n6941) );
  OAI21_X1 U9139 ( .B1(n10240), .B2(n13711), .A(n10239), .ZN(n10241) );
  OAI21_X1 U9140 ( .B1(n6774), .B2(n15941), .A(n6773), .ZN(n13670) );
  NAND2_X1 U9141 ( .A1(n15941), .A2(n13668), .ZN(n6773) );
  NOR2_X1 U9142 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  NAND2_X1 U9143 ( .A1(n7028), .A2(n6547), .ZN(n7027) );
  NAND2_X1 U9144 ( .A1(n7025), .A2(n14214), .ZN(n7024) );
  NAND2_X1 U9145 ( .A1(n6860), .A2(n6859), .ZN(P2_U3525) );
  NAND2_X1 U9146 ( .A1(n14613), .A2(n14590), .ZN(n6859) );
  INV_X1 U9147 ( .A(n14523), .ZN(n6860) );
  NAND2_X1 U9148 ( .A1(n6862), .A2(n6861), .ZN(P2_U3493) );
  NAND2_X1 U9149 ( .A1(n14613), .A2(n9001), .ZN(n6861) );
  INV_X1 U9150 ( .A(n14612), .ZN(n6862) );
  OAI21_X1 U9151 ( .B1(n15003), .B2(n14809), .A(n10265), .ZN(n10266) );
  OAI21_X1 U9152 ( .B1(n14747), .B2(n14746), .A(n15491), .ZN(n14751) );
  INV_X1 U9153 ( .A(n6843), .ZN(n6842) );
  NAND2_X1 U9154 ( .A1(n14965), .A2(n10213), .ZN(n6844) );
  NAND2_X1 U9155 ( .A1(n14964), .A2(n15207), .ZN(n6841) );
  AOI21_X1 U9156 ( .B1(n10226), .B2(n15582), .A(n10225), .ZN(n10227) );
  INV_X1 U9157 ( .A(n6839), .ZN(n15009) );
  OAI21_X1 U9158 ( .B1(n15258), .B2(n15214), .A(n6840), .ZN(n6839) );
  AOI21_X1 U9159 ( .B1(n15253), .B2(n15582), .A(n15008), .ZN(n6840) );
  NAND2_X1 U9160 ( .A1(n6852), .A2(n6851), .ZN(P1_U3527) );
  NAND2_X1 U9161 ( .A1(n15698), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U9162 ( .A1(n15396), .A2(n15700), .ZN(n6852) );
  NAND2_X1 U9163 ( .A1(n6806), .A2(n6805), .ZN(P1_U3526) );
  NAND2_X1 U9164 ( .A1(n15698), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U9165 ( .A1(n15397), .A2(n15700), .ZN(n6806) );
  NAND2_X1 U9166 ( .A1(n6846), .A2(n6845), .ZN(P1_U3518) );
  NAND2_X1 U9167 ( .A1(n15698), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6845) );
  INV_X1 U9168 ( .A(n7487), .ZN(n15955) );
  AND2_X1 U9169 ( .A1(n7494), .A2(n7490), .ZN(n15454) );
  NOR2_X1 U9170 ( .A1(n15462), .A2(n15463), .ZN(n15461) );
  NAND2_X1 U9171 ( .A1(n15467), .A2(n15466), .ZN(n15465) );
  AND2_X1 U9172 ( .A1(n6994), .A2(n6665), .ZN(n15467) );
  NAND2_X1 U9173 ( .A1(n15479), .A2(n15480), .ZN(n15478) );
  NAND2_X1 U9174 ( .A1(n7502), .A2(n7503), .ZN(n15456) );
  NAND2_X1 U9175 ( .A1(n15479), .A2(n7504), .ZN(n7502) );
  XNOR2_X1 U9176 ( .A(n10253), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n10254) );
  NAND2_X2 U9177 ( .A1(n8213), .A2(n8212), .ZN(n10129) );
  INV_X1 U9178 ( .A(n6610), .ZN(n6786) );
  OR2_X1 U9179 ( .A1(n12888), .A2(n7010), .ZN(n6609) );
  OR2_X1 U9180 ( .A1(n14338), .A2(n14553), .ZN(n6610) );
  XNOR2_X1 U9181 ( .A(n13428), .B(n12418), .ZN(n6611) );
  AND2_X1 U9182 ( .A1(n13291), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6612) );
  AND2_X1 U9183 ( .A1(n11661), .A2(n11660), .ZN(n6613) );
  INV_X1 U9184 ( .A(n13470), .ZN(n7248) );
  INV_X1 U9185 ( .A(n10244), .ZN(n6986) );
  INV_X1 U9186 ( .A(n12829), .ZN(n7235) );
  INV_X1 U9187 ( .A(n7598), .ZN(n7597) );
  NAND2_X1 U9188 ( .A1(n7601), .A2(n7599), .ZN(n7598) );
  AND2_X1 U9189 ( .A1(n7079), .A2(n6686), .ZN(n6614) );
  OR2_X1 U9190 ( .A1(n10341), .A2(n10095), .ZN(n6615) );
  INV_X1 U9191 ( .A(n7986), .ZN(n7585) );
  AND2_X1 U9192 ( .A1(n7574), .A2(n8309), .ZN(n6617) );
  AND2_X1 U9193 ( .A1(n13365), .A2(n6548), .ZN(n6618) );
  AND2_X1 U9194 ( .A1(n8194), .A2(n8193), .ZN(n15314) );
  AND2_X1 U9195 ( .A1(n12229), .A2(n7567), .ZN(n6619) );
  INV_X1 U9196 ( .A(n7002), .ZN(n7275) );
  AND2_X1 U9197 ( .A1(n7605), .A2(n6736), .ZN(n14252) );
  AND3_X1 U9198 ( .A1(n7509), .A2(n14310), .A3(n7508), .ZN(n6620) );
  INV_X1 U9199 ( .A(n15811), .ZN(n11324) );
  AND2_X1 U9200 ( .A1(n7452), .A2(n6675), .ZN(n6621) );
  AND2_X1 U9201 ( .A1(n12386), .A2(n13370), .ZN(n6622) );
  AND2_X1 U9202 ( .A1(n13407), .A2(n6695), .ZN(n6623) );
  INV_X1 U9203 ( .A(n7644), .ZN(n7600) );
  AND2_X1 U9204 ( .A1(n6718), .A2(n7738), .ZN(n6624) );
  AND2_X1 U9205 ( .A1(n7248), .A2(n12887), .ZN(n6625) );
  AND3_X1 U9206 ( .A1(n11520), .A2(n11741), .A3(n11561), .ZN(n6626) );
  INV_X1 U9207 ( .A(n15466), .ZN(n6997) );
  AND2_X1 U9208 ( .A1(n6958), .A2(n12965), .ZN(n6627) );
  AND2_X1 U9209 ( .A1(n15267), .A2(n7441), .ZN(n6628) );
  AND2_X1 U9210 ( .A1(n9729), .A2(n9728), .ZN(n6629) );
  NOR2_X1 U9211 ( .A1(n15372), .A2(n15362), .ZN(n6630) );
  AND2_X1 U9212 ( .A1(n7509), .A2(n14293), .ZN(n6631) );
  AND2_X1 U9213 ( .A1(n12350), .A2(n12349), .ZN(n6632) );
  NAND2_X1 U9214 ( .A1(n6756), .A2(n7283), .ZN(n8877) );
  NAND2_X1 U9215 ( .A1(n11756), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6633) );
  AND2_X1 U9216 ( .A1(n7175), .A2(n9400), .ZN(n6634) );
  AND2_X1 U9217 ( .A1(n7336), .A2(n7337), .ZN(n6635) );
  NAND2_X1 U9218 ( .A1(n11306), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11287) );
  NAND2_X1 U9219 ( .A1(n6604), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U9220 ( .A1(n14165), .A2(n11961), .ZN(n6637) );
  NOR2_X1 U9221 ( .A1(n13297), .A2(n7060), .ZN(n6638) );
  INV_X1 U9222 ( .A(n9345), .ZN(n9396) );
  CLKBUF_X3 U9223 ( .A(n8594), .Z(n9902) );
  INV_X1 U9224 ( .A(n6542), .ZN(n9467) );
  INV_X1 U9225 ( .A(n8216), .ZN(n8121) );
  AND2_X1 U9226 ( .A1(n7681), .A2(SI_7_), .ZN(n6639) );
  OR2_X1 U9227 ( .A1(n15285), .A2(n15273), .ZN(n6640) );
  AND2_X1 U9228 ( .A1(n9598), .A2(n9596), .ZN(n6641) );
  AND2_X1 U9229 ( .A1(n15346), .A2(n15354), .ZN(n6642) );
  INV_X1 U9230 ( .A(n13027), .ZN(n13568) );
  AND4_X1 U9231 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(n13027)
         );
  NAND2_X1 U9232 ( .A1(n7241), .A2(n12865), .ZN(n13529) );
  NAND2_X1 U9233 ( .A1(n8747), .A2(n8746), .ZN(n14372) );
  XNOR2_X1 U9234 ( .A(n13583), .B(n13027), .ZN(n9569) );
  NAND2_X1 U9235 ( .A1(n14428), .A2(n7304), .ZN(n14381) );
  OR2_X1 U9236 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n11073), .ZN(n6643) );
  INV_X1 U9237 ( .A(n13801), .ZN(n14019) );
  NAND2_X1 U9238 ( .A1(n7034), .A2(n7031), .ZN(n6644) );
  XNOR2_X1 U9239 ( .A(n14519), .B(n13801), .ZN(n14241) );
  OR2_X1 U9240 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6645) );
  INV_X1 U9241 ( .A(n9579), .ZN(n7078) );
  AND2_X1 U9242 ( .A1(n13533), .A2(n12873), .ZN(n13549) );
  AND2_X1 U9243 ( .A1(n15073), .A2(n6628), .ZN(n6646) );
  XNOR2_X1 U9244 ( .A(n14553), .B(n14349), .ZN(n14334) );
  NOR2_X1 U9245 ( .A1(n12310), .A2(n6960), .ZN(n6647) );
  NAND2_X1 U9246 ( .A1(n15463), .A2(n7497), .ZN(n6648) );
  AND2_X1 U9247 ( .A1(n7129), .A2(n7128), .ZN(n6649) );
  OR2_X1 U9248 ( .A1(n15332), .A2(n14819), .ZN(n6650) );
  OR2_X1 U9249 ( .A1(n12928), .A2(n12926), .ZN(n6651) );
  INV_X1 U9250 ( .A(n6607), .ZN(n8988) );
  NAND2_X1 U9251 ( .A1(n8622), .A2(n8621), .ZN(n11876) );
  INV_X1 U9252 ( .A(n10080), .ZN(n6989) );
  NOR2_X1 U9253 ( .A1(n6534), .A2(n13139), .ZN(n6652) );
  NAND2_X1 U9254 ( .A1(n7410), .A2(n7409), .ZN(n7416) );
  OR2_X1 U9255 ( .A1(n10014), .A2(n11151), .ZN(n6653) );
  NOR2_X1 U9256 ( .A1(n6937), .A2(n7255), .ZN(n9022) );
  AND2_X1 U9257 ( .A1(n8962), .A2(n8959), .ZN(n6654) );
  OR2_X1 U9258 ( .A1(n15659), .A2(n15666), .ZN(n6655) );
  NAND2_X1 U9259 ( .A1(n12357), .A2(n13512), .ZN(n6656) );
  INV_X1 U9260 ( .A(n15069), .ZN(n7415) );
  INV_X1 U9261 ( .A(n11561), .ZN(n15827) );
  AND2_X1 U9262 ( .A1(n8597), .A2(n8596), .ZN(n11561) );
  AND2_X1 U9263 ( .A1(n9132), .A2(n7104), .ZN(n6657) );
  NAND2_X1 U9264 ( .A1(n14384), .A2(n8959), .ZN(n14365) );
  NOR2_X1 U9265 ( .A1(n14761), .A2(n7644), .ZN(n6658) );
  NAND2_X1 U9266 ( .A1(n9530), .A2(n9529), .ZN(n9664) );
  AND2_X1 U9267 ( .A1(n7262), .A2(n7260), .ZN(n6659) );
  AND2_X1 U9268 ( .A1(n6615), .A2(n7504), .ZN(n6661) );
  INV_X1 U9269 ( .A(n11266), .ZN(n11307) );
  NAND2_X1 U9270 ( .A1(n8515), .A2(n8514), .ZN(n12319) );
  INV_X1 U9271 ( .A(n12319), .ZN(n7602) );
  NOR2_X1 U9272 ( .A1(n14315), .A2(n14316), .ZN(n14314) );
  AND3_X1 U9273 ( .A1(n8485), .A2(n8483), .A3(n8484), .ZN(n8872) );
  AND2_X1 U9274 ( .A1(n14543), .A2(n14023), .ZN(n6662) );
  INV_X1 U9275 ( .A(n12558), .ZN(n7471) );
  NAND2_X1 U9276 ( .A1(n8154), .A2(n8153), .ZN(n6663) );
  AND3_X1 U9277 ( .A1(n9029), .A2(n9026), .A3(n9028), .ZN(n6664) );
  OR2_X1 U9278 ( .A1(n15463), .A2(n7497), .ZN(n6665) );
  AND2_X1 U9279 ( .A1(n12548), .A2(n15514), .ZN(n6666) );
  INV_X1 U9280 ( .A(n10271), .ZN(n8970) );
  XNOR2_X1 U9281 ( .A(n14225), .B(n14018), .ZN(n10271) );
  AND2_X1 U9282 ( .A1(n12992), .A2(n6656), .ZN(n6667) );
  INV_X1 U9283 ( .A(n12463), .ZN(n12465) );
  OR2_X1 U9284 ( .A1(n12338), .A2(n12530), .ZN(n6668) );
  INV_X1 U9285 ( .A(n12722), .ZN(n7524) );
  AND3_X1 U9286 ( .A1(n7805), .A2(n7807), .A3(n7808), .ZN(n6669) );
  NOR2_X1 U9287 ( .A1(n10520), .A2(n10519), .ZN(n6670) );
  NOR2_X1 U9288 ( .A1(n12548), .A2(n15514), .ZN(n6671) );
  AND2_X1 U9289 ( .A1(n7369), .A2(n7366), .ZN(n6672) );
  INV_X1 U9290 ( .A(n15089), .ZN(n15294) );
  AND2_X1 U9291 ( .A1(n8294), .A2(n8293), .ZN(n15089) );
  AND2_X1 U9292 ( .A1(n7091), .A2(n7090), .ZN(n6673) );
  NOR2_X1 U9293 ( .A1(n7002), .A2(n12934), .ZN(n6674) );
  OR2_X1 U9294 ( .A1(n6611), .A2(n6652), .ZN(n6675) );
  AND2_X1 U9295 ( .A1(n7249), .A2(n7250), .ZN(n6676) );
  OR2_X1 U9296 ( .A1(n12385), .A2(n11666), .ZN(n6677) );
  INV_X1 U9297 ( .A(n12519), .ZN(n12520) );
  NOR2_X1 U9298 ( .A1(n14254), .A2(n14273), .ZN(n6678) );
  NOR2_X1 U9299 ( .A1(n12358), .A2(n7447), .ZN(n6679) );
  AND2_X1 U9300 ( .A1(n10141), .A2(n10140), .ZN(n6680) );
  INV_X1 U9301 ( .A(n7136), .ZN(n7133) );
  NAND2_X1 U9302 ( .A1(n15339), .A2(n15344), .ZN(n7136) );
  NOR2_X1 U9303 ( .A1(n11471), .A2(n12036), .ZN(n6681) );
  INV_X1 U9304 ( .A(n13849), .ZN(n7370) );
  AND2_X1 U9305 ( .A1(n6943), .A2(n6942), .ZN(n6682) );
  INV_X1 U9306 ( .A(n11681), .ZN(n7459) );
  AND2_X1 U9307 ( .A1(n7001), .A2(n7005), .ZN(n6683) );
  NAND2_X1 U9308 ( .A1(n7867), .A2(n7866), .ZN(n6684) );
  INV_X1 U9309 ( .A(n6973), .ZN(n6972) );
  NAND2_X1 U9310 ( .A1(n6974), .A2(n6979), .ZN(n6973) );
  INV_X1 U9311 ( .A(n9576), .ZN(n7077) );
  AND3_X1 U9312 ( .A1(n14373), .A2(n7301), .A3(n14410), .ZN(n6685) );
  NAND2_X1 U9313 ( .A1(n13541), .A2(n13546), .ZN(n6686) );
  AND2_X1 U9314 ( .A1(n8945), .A2(n14469), .ZN(n6687) );
  NAND2_X1 U9315 ( .A1(n11829), .A2(n9559), .ZN(n6688) );
  NAND2_X1 U9316 ( .A1(n10049), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n6689) );
  XNOR2_X1 U9317 ( .A(n7681), .B(SI_7_), .ZN(n7894) );
  AND2_X1 U9318 ( .A1(n12257), .A2(n12253), .ZN(n6690) );
  AND2_X1 U9319 ( .A1(n14593), .A2(n14495), .ZN(n6691) );
  NAND2_X2 U9320 ( .A1(n8817), .A2(n8816), .ZN(n14538) );
  AND2_X1 U9321 ( .A1(n7305), .A2(n7646), .ZN(n6692) );
  AND2_X1 U9322 ( .A1(n15235), .A2(n6855), .ZN(n6693) );
  INV_X1 U9323 ( .A(n7577), .ZN(n7576) );
  NAND2_X1 U9324 ( .A1(n7629), .A2(n7578), .ZN(n7577) );
  AND2_X1 U9325 ( .A1(n7727), .A2(n7106), .ZN(n6694) );
  AND2_X1 U9326 ( .A1(n12897), .A2(n13420), .ZN(n6695) );
  AND2_X1 U9327 ( .A1(n8970), .A2(n8845), .ZN(n6696) );
  OR2_X1 U9328 ( .A1(n7466), .A2(n12610), .ZN(n6697) );
  INV_X1 U9329 ( .A(n7694), .ZN(n7428) );
  NAND2_X1 U9330 ( .A1(n7691), .A2(n10651), .ZN(n7694) );
  AND2_X1 U9331 ( .A1(n14734), .A2(n14733), .ZN(n8152) );
  INV_X1 U9332 ( .A(n6896), .ZN(n15279) );
  NAND2_X1 U9333 ( .A1(n14527), .A2(n14020), .ZN(n6698) );
  INV_X1 U9334 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9357) );
  INV_X1 U9335 ( .A(n14225), .ZN(n13807) );
  XNOR2_X1 U9336 ( .A(n15020), .B(n15028), .ZN(n15013) );
  INV_X1 U9337 ( .A(n15261), .ZN(n15020) );
  AND2_X1 U9338 ( .A1(n7391), .A2(n7389), .ZN(n6699) );
  AND2_X1 U9339 ( .A1(n7293), .A2(n7291), .ZN(n6700) );
  AND3_X1 U9340 ( .A1(n12927), .A2(n12925), .A3(n12756), .ZN(n6701) );
  NOR2_X1 U9341 ( .A1(n8844), .A2(n14019), .ZN(n6702) );
  NOR2_X1 U9342 ( .A1(n14036), .A2(n15834), .ZN(n6703) );
  INV_X1 U9343 ( .A(n8969), .ZN(n6935) );
  AND2_X1 U9344 ( .A1(n9587), .A2(n9586), .ZN(n6704) );
  INV_X1 U9345 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7901) );
  INV_X1 U9346 ( .A(n7397), .ZN(n7396) );
  AND2_X1 U9347 ( .A1(n15378), .A2(n15384), .ZN(n6705) );
  AND2_X1 U9348 ( .A1(n8021), .A2(n8022), .ZN(n6706) );
  NAND2_X1 U9349 ( .A1(n12347), .A2(n13545), .ZN(n6707) );
  INV_X1 U9350 ( .A(n7523), .ZN(n7522) );
  NAND2_X1 U9351 ( .A1(n7525), .A2(n7524), .ZN(n7523) );
  INV_X1 U9352 ( .A(n15007), .ZN(n7434) );
  AND2_X1 U9353 ( .A1(n15034), .A2(n15274), .ZN(n6708) );
  NOR2_X1 U9354 ( .A1(n8075), .A2(n8074), .ZN(n6709) );
  NOR2_X1 U9355 ( .A1(n9579), .A2(n6908), .ZN(n6710) );
  AND2_X1 U9356 ( .A1(n12344), .A2(n13568), .ZN(n6711) );
  INV_X1 U9357 ( .A(n7016), .ZN(n7015) );
  NAND2_X1 U9358 ( .A1(n13496), .A2(n13517), .ZN(n7016) );
  AND2_X1 U9359 ( .A1(n7015), .A2(n7013), .ZN(n6712) );
  NAND2_X1 U9360 ( .A1(n10009), .A2(n10008), .ZN(n6713) );
  INV_X1 U9361 ( .A(n9711), .ZN(n7205) );
  INV_X1 U9362 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10623) );
  INV_X1 U9363 ( .A(n7247), .ZN(n7246) );
  NAND2_X1 U9364 ( .A1(n7250), .A2(n7248), .ZN(n7247) );
  NOR2_X1 U9365 ( .A1(n9253), .A2(n7243), .ZN(n7242) );
  INV_X1 U9366 ( .A(n7292), .ZN(n7291) );
  NAND2_X1 U9367 ( .A1(n7296), .A2(n7297), .ZN(n7292) );
  OR3_X1 U9368 ( .A1(n9845), .A2(n9844), .A3(n9843), .ZN(n6714) );
  AND2_X1 U9369 ( .A1(n7510), .A2(n14505), .ZN(n6715) );
  NAND2_X1 U9370 ( .A1(n8131), .A2(n8130), .ZN(n6716) );
  AND2_X1 U9371 ( .A1(n15466), .A2(n10087), .ZN(n6717) );
  AND2_X1 U9372 ( .A1(n7734), .A2(n8161), .ZN(n6718) );
  INV_X1 U9373 ( .A(n12761), .ZN(n12907) );
  AND2_X1 U9374 ( .A1(n7006), .A2(n7004), .ZN(n6719) );
  INV_X1 U9375 ( .A(n8229), .ZN(n7578) );
  AND2_X1 U9376 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  INV_X1 U9377 ( .A(n15267), .ZN(n15034) );
  AND2_X1 U9378 ( .A1(n6661), .A2(n10244), .ZN(n6720) );
  INV_X1 U9379 ( .A(n6958), .ZN(n6957) );
  AND2_X1 U9380 ( .A1(n6733), .A2(n12309), .ZN(n6958) );
  OR2_X1 U9381 ( .A1(n9593), .A2(n6919), .ZN(n6721) );
  INV_X1 U9382 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10629) );
  OR2_X1 U9383 ( .A1(n13605), .A2(n13433), .ZN(n6722) );
  AND2_X1 U9384 ( .A1(n6969), .A2(n6978), .ZN(n6723) );
  OR2_X1 U9385 ( .A1(n9731), .A2(n6629), .ZN(n6724) );
  OR2_X1 U9386 ( .A1(n9757), .A2(n9759), .ZN(n6725) );
  AND2_X1 U9387 ( .A1(n10188), .A2(n10186), .ZN(n6726) );
  AND3_X1 U9388 ( .A1(n12901), .A2(n12902), .A3(n12903), .ZN(n6727) );
  XNOR2_X1 U9389 ( .A(n9020), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9025) );
  AND2_X1 U9390 ( .A1(n9371), .A2(n12886), .ZN(n12882) );
  AND2_X1 U9391 ( .A1(n7989), .A2(n7694), .ZN(n6728) );
  AND2_X1 U9392 ( .A1(n15013), .A2(n7108), .ZN(n6729) );
  AND2_X1 U9393 ( .A1(n9311), .A2(n7242), .ZN(n6730) );
  NAND2_X1 U9394 ( .A1(n15372), .A2(n15362), .ZN(n6731) );
  AND2_X1 U9395 ( .A1(n7528), .A2(n15010), .ZN(n6732) );
  NAND2_X1 U9396 ( .A1(n12343), .A2(n13027), .ZN(n6733) );
  NAND2_X1 U9397 ( .A1(n13741), .A2(n13740), .ZN(n6734) );
  AND2_X1 U9398 ( .A1(n7604), .A2(n6698), .ZN(n6735) );
  NAND2_X1 U9399 ( .A1(n14532), .A2(n14021), .ZN(n6736) );
  AND2_X1 U9400 ( .A1(n9322), .A2(n9357), .ZN(n6737) );
  AND2_X1 U9401 ( .A1(n6641), .A2(n7089), .ZN(n6738) );
  AND2_X1 U9402 ( .A1(n9583), .A2(n9581), .ZN(n6739) );
  AND2_X1 U9403 ( .A1(n12365), .A2(n12364), .ZN(n6740) );
  AND2_X1 U9404 ( .A1(n6628), .A2(n15261), .ZN(n6741) );
  AND2_X1 U9405 ( .A1(n7500), .A2(n7502), .ZN(n6742) );
  AND2_X1 U9406 ( .A1(n10013), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n6743) );
  OR2_X1 U9407 ( .A1(n7207), .A2(n9758), .ZN(n6744) );
  AND2_X1 U9408 ( .A1(n7465), .A2(n12615), .ZN(n6745) );
  AND2_X1 U9409 ( .A1(n7233), .A2(n12832), .ZN(n6746) );
  AND2_X1 U9410 ( .A1(n12557), .A2(n7471), .ZN(n6747) );
  OAI21_X1 U9411 ( .B1(n6955), .B2(n6954), .A(n6707), .ZN(n6953) );
  OR2_X1 U9412 ( .A1(n12871), .A2(n7014), .ZN(n6748) );
  OR2_X1 U9413 ( .A1(n12557), .A2(n7471), .ZN(n6749) );
  INV_X1 U9414 ( .A(n12669), .ZN(n15026) );
  AND2_X1 U9415 ( .A1(n14786), .A2(n6663), .ZN(n7590) );
  INV_X1 U9416 ( .A(n12915), .ZN(n7276) );
  AND2_X1 U9417 ( .A1(n13674), .A2(n13370), .ZN(n12915) );
  OR2_X1 U9418 ( .A1(n10020), .A2(n11100), .ZN(n10021) );
  INV_X1 U9419 ( .A(n7114), .ZN(n7113) );
  AND2_X1 U9420 ( .A1(n6668), .A2(n10109), .ZN(n7114) );
  AND2_X1 U9421 ( .A1(n6996), .A2(n6665), .ZN(n6993) );
  INV_X1 U9422 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U9423 ( .A1(n7205), .A2(n9712), .ZN(n6750) );
  INV_X1 U9424 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U9425 ( .A1(n13356), .A2(n7087), .ZN(n6751) );
  AND2_X1 U9426 ( .A1(n12786), .A2(n12927), .ZN(n6752) );
  INV_X1 U9427 ( .A(n14430), .ZN(n7301) );
  NAND2_X1 U9428 ( .A1(n6715), .A2(n8989), .ZN(n14480) );
  NOR2_X1 U9429 ( .A1(n6850), .A2(n12526), .ZN(n6753) );
  INV_X1 U9430 ( .A(n12937), .ZN(n11661) );
  NAND2_X1 U9431 ( .A1(n8671), .A2(n8670), .ZN(n14502) );
  INV_X1 U9432 ( .A(n15091), .ZN(n7436) );
  AND2_X1 U9434 ( .A1(n6534), .A2(n13139), .ZN(n6754) );
  NAND2_X1 U9435 ( .A1(n7081), .A2(n7080), .ZN(n11804) );
  NAND2_X1 U9436 ( .A1(n9452), .A2(n9451), .ZN(n13139) );
  INV_X1 U9437 ( .A(n13139), .ZN(n13447) );
  INV_X1 U9438 ( .A(n14573), .ZN(n7518) );
  NOR2_X1 U9439 ( .A1(n6608), .A2(n7760), .ZN(n6755) );
  NAND2_X1 U9440 ( .A1(n11906), .A2(n10166), .ZN(n12143) );
  NAND2_X1 U9441 ( .A1(n7548), .A2(n10163), .ZN(n11609) );
  NAND2_X1 U9442 ( .A1(n7614), .A2(n8602), .ZN(n11726) );
  NAND2_X1 U9443 ( .A1(n7094), .A2(n9486), .ZN(n13385) );
  INV_X1 U9444 ( .A(n13385), .ZN(n13357) );
  AND4_X1 U9445 ( .A1(n6616), .A2(n8479), .A3(n6533), .A4(n8872), .ZN(n6756)
         );
  NOR2_X1 U9446 ( .A1(n14481), .A2(n7520), .ZN(n14419) );
  INV_X1 U9447 ( .A(n14548), .ZN(n7509) );
  NAND2_X1 U9448 ( .A1(n7167), .A2(n9480), .ZN(n9594) );
  INV_X1 U9449 ( .A(n9594), .ZN(n7093) );
  NOR2_X1 U9450 ( .A1(n8005), .A2(n8004), .ZN(n6757) );
  AND2_X1 U9451 ( .A1(n9981), .A2(n9982), .ZN(n6758) );
  INV_X1 U9452 ( .A(n14481), .ZN(n7516) );
  NAND2_X1 U9453 ( .A1(n8989), .A2(n7512), .ZN(n7513) );
  NAND2_X1 U9454 ( .A1(n9209), .A2(n9193), .ZN(n6759) );
  OR2_X1 U9455 ( .A1(n11928), .A2(n11919), .ZN(n6760) );
  INV_X1 U9456 ( .A(n7217), .ZN(n7216) );
  NOR2_X1 U9457 ( .A1(n9786), .A2(n7219), .ZN(n7217) );
  AND2_X1 U9458 ( .A1(n7101), .A2(n10474), .ZN(n6761) );
  AND2_X1 U9459 ( .A1(n11606), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6762) );
  AND2_X1 U9460 ( .A1(n10939), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n6763) );
  AND2_X1 U9461 ( .A1(n8436), .A2(SI_27_), .ZN(n6764) );
  AND2_X1 U9462 ( .A1(n7338), .A2(n11765), .ZN(n6765) );
  OR2_X1 U9463 ( .A1(n13199), .A2(n7329), .ZN(n6766) );
  INV_X1 U9464 ( .A(n8089), .ZN(n7424) );
  INV_X1 U9465 ( .A(n9813), .ZN(n7225) );
  AND2_X1 U9466 ( .A1(n7099), .A2(n7098), .ZN(n6767) );
  NAND2_X1 U9467 ( .A1(n7230), .A2(n7228), .ZN(n8886) );
  INV_X1 U9468 ( .A(n15867), .ZN(n13128) );
  NAND2_X1 U9469 ( .A1(n9268), .A2(n9267), .ZN(n13707) );
  AND2_X2 U9470 ( .A1(n11413), .A2(n9662), .ZN(n15954) );
  AND2_X1 U9471 ( .A1(n10807), .A2(n10802), .ZN(n15734) );
  NOR2_X1 U9472 ( .A1(n14182), .A2(n14183), .ZN(n7044) );
  NAND2_X1 U9473 ( .A1(n7759), .A2(n12430), .ZN(n11002) );
  AND2_X1 U9474 ( .A1(n11252), .A2(n11097), .ZN(n6768) );
  AND2_X1 U9475 ( .A1(n13287), .A2(n13294), .ZN(n6769) );
  NAND2_X1 U9476 ( .A1(n6949), .A2(n11676), .ZN(n12981) );
  INV_X1 U9477 ( .A(n7314), .ZN(n11306) );
  AND2_X1 U9478 ( .A1(n15137), .A2(n15674), .ZN(n15694) );
  AND2_X1 U9479 ( .A1(n11166), .A2(n11165), .ZN(n11215) );
  NAND2_X1 U9480 ( .A1(n7311), .A2(n11266), .ZN(n7316) );
  INV_X1 U9481 ( .A(n7044), .ZN(n7043) );
  AND2_X1 U9482 ( .A1(n14134), .A2(n10883), .ZN(n6770) );
  INV_X1 U9483 ( .A(n11568), .ZN(n7051) );
  INV_X1 U9484 ( .A(n14189), .ZN(n7042) );
  NAND2_X1 U9485 ( .A1(n12438), .A2(n7763), .ZN(n15207) );
  XOR2_X1 U9486 ( .A(n11283), .B(P3_REG2_REG_6__SCAN_IN), .Z(n6771) );
  INV_X1 U9487 ( .A(n6547), .ZN(n14214) );
  INV_X1 U9488 ( .A(n9022), .ZN(n6857) );
  INV_X1 U9489 ( .A(n6637), .ZN(n7041) );
  AND2_X1 U9490 ( .A1(n13311), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6772) );
  INV_X1 U9491 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7559) );
  INV_X1 U9492 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n10252) );
  INV_X1 U9493 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7067) );
  INV_X1 U9494 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U9495 ( .A1(n13267), .A2(n13294), .ZN(n13291) );
  AOI21_X1 U9496 ( .B1(n14982), .B2(n14983), .A(n14981), .ZN(n15248) );
  INV_X2 U9497 ( .A(n12653), .ZN(n11885) );
  NAND2_X1 U9498 ( .A1(n6814), .A2(n7434), .ZN(n15004) );
  NAND2_X1 U9499 ( .A1(n15066), .A2(n10191), .ZN(n10197) );
  NAND2_X1 U9500 ( .A1(n10184), .A2(n7653), .ZN(n10187) );
  INV_X1 U9501 ( .A(n15426), .ZN(n7748) );
  INV_X1 U9502 ( .A(n15006), .ZN(n6814) );
  NAND2_X1 U9503 ( .A1(n7537), .A2(n7539), .ZN(n12048) );
  AOI21_X2 U9504 ( .B1(n13360), .B2(n13562), .A(n13359), .ZN(n13599) );
  NAND3_X1 U9505 ( .A1(n6751), .A2(n13342), .A3(n13562), .ZN(n13348) );
  NAND2_X1 U9506 ( .A1(n13356), .A2(n9599), .ZN(n13341) );
  NAND2_X1 U9507 ( .A1(n10165), .A2(n7538), .ZN(n7537) );
  NAND2_X1 U9508 ( .A1(n10176), .A2(n10175), .ZN(n12279) );
  OAI21_X1 U9509 ( .B1(n12048), .B2(n6630), .A(n6731), .ZN(n6813) );
  NOR2_X1 U9510 ( .A1(n13278), .A2(n13279), .ZN(n13286) );
  AOI21_X1 U9511 ( .B1(n13248), .B2(n13247), .A(n13246), .ZN(n13277) );
  NAND2_X1 U9512 ( .A1(n9510), .A2(n9511), .ZN(n9527) );
  NAND2_X1 U9513 ( .A1(n9457), .A2(n9456), .ZN(n9476) );
  NAND2_X1 U9514 ( .A1(n9354), .A2(n9353), .ZN(n9356) );
  OAI22_X1 U9515 ( .A1(n12748), .A2(n12747), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n15425), .ZN(n12750) );
  NAND2_X1 U9516 ( .A1(n9225), .A2(n9224), .ZN(n9239) );
  INV_X1 U9517 ( .A(n7377), .ZN(n7374) );
  NAND2_X1 U9518 ( .A1(n10923), .A2(n6552), .ZN(n8036) );
  NAND2_X1 U9519 ( .A1(n15038), .A2(n6897), .ZN(n6896) );
  NOR2_X1 U9520 ( .A1(n13228), .A2(n13227), .ZN(n13246) );
  NOR2_X1 U9521 ( .A1(n13322), .A2(n7200), .ZN(n7199) );
  NOR2_X1 U9522 ( .A1(n13286), .A2(n6769), .ZN(n13324) );
  OAI21_X1 U9523 ( .B1(n13277), .B2(n13276), .A(n13275), .ZN(n13278) );
  NAND2_X1 U9524 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  NAND2_X1 U9525 ( .A1(n12476), .A2(n12469), .ZN(n12470) );
  NAND2_X1 U9526 ( .A1(n9721), .A2(n9720), .ZN(n9726) );
  NAND2_X1 U9527 ( .A1(n9957), .A2(n6775), .ZN(n9964) );
  OAI22_X1 U9528 ( .A1(n9968), .A2(n9969), .B1(n9956), .B2(n9955), .ZN(n6775)
         );
  NAND2_X1 U9529 ( .A1(n7583), .A2(n7847), .ZN(n6776) );
  NAND3_X1 U9530 ( .A1(n12126), .A2(n7568), .A3(n12129), .ZN(n7564) );
  NAND2_X1 U9531 ( .A1(n7941), .A2(n7940), .ZN(n11595) );
  NOR2_X1 U9532 ( .A1(n15485), .A2(n7580), .ZN(n7579) );
  AOI21_X4 U9533 ( .B1(n6608), .B2(n15207), .A(n12491), .ZN(n8448) );
  NAND3_X1 U9534 ( .A1(n7180), .A2(n6779), .A3(n12947), .ZN(P3_U3296) );
  NAND3_X1 U9535 ( .A1(n6880), .A2(n12760), .A3(n12941), .ZN(n6779) );
  NAND2_X1 U9536 ( .A1(n15054), .A2(n10137), .ZN(n15037) );
  NAND2_X1 U9537 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  AOI21_X1 U9538 ( .B1(n7019), .B2(n6727), .A(n7018), .ZN(n7181) );
  NAND4_X1 U9539 ( .A1(n6999), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n7095)
         );
  NAND2_X1 U9540 ( .A1(n14657), .A2(n6552), .ZN(n12641) );
  NAND2_X1 U9541 ( .A1(n8369), .A2(n7160), .ZN(n6800) );
  NAND2_X1 U9542 ( .A1(n6780), .A2(n12700), .ZN(P1_U3242) );
  OAI21_X1 U9543 ( .B1(n12695), .B2(n12694), .A(n6781), .ZN(n6780) );
  OR2_X2 U9544 ( .A1(n8838), .A2(n10380), .ZN(n8860) );
  NAND2_X1 U9545 ( .A1(n8693), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U9546 ( .A1(n14290), .A2(n14289), .ZN(n14288) );
  NAND2_X1 U9547 ( .A1(n8503), .A2(n8502), .ZN(n8788) );
  NAND2_X1 U9548 ( .A1(n9793), .A2(n9792), .ZN(n6784) );
  NAND2_X1 U9549 ( .A1(n6785), .A2(n7211), .ZN(n9737) );
  NAND3_X1 U9550 ( .A1(n6809), .A2(n7212), .A3(n6724), .ZN(n6785) );
  NAND3_X1 U9551 ( .A1(n8093), .A2(n8094), .A3(n7726), .ZN(n8160) );
  INV_X1 U9552 ( .A(n10010), .ZN(n6797) );
  INV_X1 U9553 ( .A(n7822), .ZN(n7580) );
  AOI21_X1 U9554 ( .B1(n10537), .B2(n12722), .A(n14482), .ZN(n10538) );
  NAND2_X1 U9555 ( .A1(n14368), .A2(n14361), .ZN(n14338) );
  NAND2_X1 U9556 ( .A1(n7519), .A2(n7518), .ZN(n7517) );
  INV_X1 U9557 ( .A(n12721), .ZN(n12724) );
  NAND2_X1 U9558 ( .A1(n7342), .A2(n13257), .ZN(n13266) );
  NOR2_X1 U9559 ( .A1(n6911), .A2(n10557), .ZN(n12731) );
  NOR2_X1 U9560 ( .A1(n12725), .A2(n10556), .ZN(n6912) );
  NAND2_X1 U9561 ( .A1(n15885), .A2(n7338), .ZN(n7337) );
  NAND2_X1 U9562 ( .A1(n12788), .A2(n6788), .ZN(n6787) );
  AND2_X1 U9563 ( .A1(n12787), .A2(n6752), .ZN(n6788) );
  NAND2_X1 U9564 ( .A1(n12795), .A2(n12794), .ZN(n12940) );
  NAND2_X1 U9565 ( .A1(n9476), .A2(n9475), .ZN(n9479) );
  NAND2_X1 U9566 ( .A1(n6792), .A2(n6674), .ZN(n6791) );
  NAND2_X1 U9567 ( .A1(n9316), .A2(n9315), .ZN(n9333) );
  NAND2_X1 U9568 ( .A1(n9507), .A2(n9506), .ZN(n9510) );
  NAND2_X1 U9569 ( .A1(n9424), .A2(n9423), .ZN(n9442) );
  NAND2_X1 U9570 ( .A1(n9429), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9430) );
  INV_X1 U9571 ( .A(n12924), .ZN(n6792) );
  NAND2_X1 U9572 ( .A1(n6796), .A2(n11060), .ZN(n11144) );
  NAND2_X1 U9573 ( .A1(n11108), .A2(n11109), .ZN(n6796) );
  AOI21_X1 U9574 ( .B1(n7198), .B2(n13154), .A(n6885), .ZN(n13328) );
  NAND3_X1 U9575 ( .A1(n10011), .A2(n6713), .A3(n6797), .ZN(P2_U3328) );
  NAND3_X1 U9576 ( .A1(n7633), .A2(n9882), .A3(n6714), .ZN(n7222) );
  AND2_X4 U9577 ( .A1(n7995), .A2(n7994), .ZN(n15378) );
  NAND2_X1 U9578 ( .A1(n8477), .A2(n6802), .ZN(P1_U3220) );
  NAND2_X1 U9579 ( .A1(n8453), .A2(n6803), .ZN(n6802) );
  NAND2_X1 U9580 ( .A1(n7576), .A2(n7575), .ZN(n7574) );
  OR2_X1 U9581 ( .A1(n9853), .A2(n9833), .ZN(n9845) );
  INV_X1 U9582 ( .A(n15420), .ZN(n7745) );
  NAND2_X1 U9583 ( .A1(n7573), .A2(n7571), .ZN(n14708) );
  NAND2_X1 U9584 ( .A1(n7367), .A2(n7365), .ZN(n7364) );
  XNOR2_X1 U9585 ( .A(n7781), .B(n8448), .ZN(n7801) );
  NAND2_X2 U9586 ( .A1(n15103), .A2(n7436), .ZN(n15083) );
  NAND2_X1 U9587 ( .A1(n6811), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U9588 ( .A1(n9726), .A2(n9725), .ZN(n6811) );
  NAND2_X1 U9589 ( .A1(n15201), .A2(n15339), .ZN(n15174) );
  NAND2_X1 U9590 ( .A1(n13009), .A2(n12368), .ZN(n12415) );
  AOI21_X1 U9591 ( .B1(n6952), .B2(n6627), .A(n6953), .ZN(n13126) );
  NAND2_X1 U9592 ( .A1(n10187), .A2(n6726), .ZN(n15111) );
  NAND2_X1 U9593 ( .A1(n7527), .A2(n6732), .ZN(n10203) );
  NAND2_X1 U9594 ( .A1(n11486), .A2(n11485), .ZN(n10155) );
  INV_X1 U9595 ( .A(n6813), .ZN(n12100) );
  NAND2_X1 U9596 ( .A1(n11184), .A2(n6643), .ZN(n11115) );
  AOI22_X1 U9597 ( .A1(n11755), .A2(n11754), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11756), .ZN(n11918) );
  OAI21_X1 U9598 ( .B1(n13215), .B2(n13214), .A(n13223), .ZN(n13239) );
  AOI22_X1 U9599 ( .A1(n13163), .A2(n13162), .B1(P3_REG1_REG_12__SCAN_IN), 
        .B2(n13167), .ZN(n13183) );
  NAND2_X1 U9600 ( .A1(n10035), .A2(n10036), .ZN(n10097) );
  NOR2_X1 U9601 ( .A1(n10246), .A2(n6987), .ZN(n10255) );
  NAND2_X1 U9602 ( .A1(n8747), .A2(n7616), .ZN(n7618) );
  INV_X1 U9603 ( .A(n7138), .ZN(n10066) );
  OAI21_X1 U9604 ( .B1(n7498), .B2(n6986), .A(P2_ADDR_REG_18__SCAN_IN), .ZN(
        n6985) );
  NOR2_X1 U9605 ( .A1(n10034), .A2(n10033), .ZN(n10037) );
  NAND2_X1 U9606 ( .A1(n9242), .A2(n9241), .ZN(n9276) );
  INV_X1 U9607 ( .A(n9127), .ZN(n7378) );
  NAND2_X1 U9608 ( .A1(n12494), .A2(n12493), .ZN(n12499) );
  NAND3_X1 U9609 ( .A1(n6823), .A2(n6822), .A3(n7478), .ZN(n7476) );
  NAND2_X1 U9610 ( .A1(n12589), .A2(n12588), .ZN(n6822) );
  NAND2_X1 U9611 ( .A1(n12591), .A2(n12590), .ZN(n6823) );
  NAND2_X1 U9612 ( .A1(n12634), .A2(n6824), .ZN(n12487) );
  NOR2_X2 U9613 ( .A1(n12482), .A2(n12479), .ZN(n12634) );
  NAND2_X1 U9614 ( .A1(n12731), .A2(n15864), .ZN(n6914) );
  NAND2_X1 U9615 ( .A1(n6914), .A2(n6913), .ZN(n12732) );
  NAND2_X1 U9616 ( .A1(n7096), .A2(n12941), .ZN(n7180) );
  NAND2_X1 U9617 ( .A1(n12738), .A2(n12737), .ZN(n12748) );
  NAND2_X1 U9618 ( .A1(n10081), .A2(n6989), .ZN(n10078) );
  NAND2_X1 U9619 ( .A1(n9428), .A2(n9427), .ZN(n7194) );
  NAND2_X2 U9620 ( .A1(n15475), .A2(n15473), .ZN(n15479) );
  NAND2_X1 U9621 ( .A1(n15460), .A2(n15459), .ZN(n15458) );
  INV_X1 U9622 ( .A(n10019), .ZN(n10048) );
  INV_X1 U9623 ( .A(n6826), .ZN(n10094) );
  INV_X1 U9624 ( .A(n15957), .ZN(n6825) );
  XNOR2_X1 U9625 ( .A(n10049), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15957) );
  OAI21_X1 U9626 ( .B1(n10090), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15469), .ZN(
        n6826) );
  NOR2_X2 U9627 ( .A1(n10246), .A2(n10102), .ZN(n10104) );
  NAND2_X1 U9628 ( .A1(n10079), .A2(n10078), .ZN(n15460) );
  NOR2_X1 U9629 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  NOR2_X1 U9630 ( .A1(n15967), .A2(n15966), .ZN(n10059) );
  NAND4_X1 U9631 ( .A1(n6829), .A2(n9983), .A3(n6827), .A4(n14503), .ZN(n9984)
         );
  NAND3_X1 U9632 ( .A1(n9988), .A2(n6830), .A3(n6930), .ZN(n9989) );
  XNOR2_X2 U9633 ( .A(n7991), .B(n7990), .ZN(n10653) );
  NAND3_X1 U9634 ( .A1(n9985), .A2(n6685), .A3(n6834), .ZN(n9986) );
  XNOR2_X1 U9635 ( .A(n11671), .B(n12809), .ZN(n9556) );
  NAND2_X1 U9636 ( .A1(n12239), .A2(n12774), .ZN(n12238) );
  NAND2_X1 U9637 ( .A1(n15037), .A2(n6869), .ZN(n10139) );
  NAND2_X1 U9638 ( .A1(n9323), .A2(n9018), .ZN(n9625) );
  AND2_X2 U9639 ( .A1(n7749), .A2(n15426), .ZN(n7826) );
  XNOR2_X2 U9640 ( .A(n7558), .B(n6835), .ZN(n15426) );
  NAND2_X1 U9641 ( .A1(n15139), .A2(n6899), .ZN(n10135) );
  NAND2_X1 U9642 ( .A1(n9552), .A2(n12802), .ZN(n11667) );
  NAND2_X1 U9643 ( .A1(n15530), .A2(n7114), .ZN(n7110) );
  NAND2_X1 U9644 ( .A1(n7111), .A2(n7110), .ZN(n15513) );
  NAND2_X1 U9645 ( .A1(n12653), .A2(n11884), .ZN(n10108) );
  NAND2_X1 U9646 ( .A1(n13594), .A2(n15905), .ZN(n6893) );
  MUX2_X1 U9647 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9021), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n6837) );
  AOI21_X2 U9648 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n10009) );
  OAI21_X1 U9649 ( .B1(n13826), .B2(n13827), .A(n13825), .ZN(n13791) );
  INV_X1 U9650 ( .A(n10165), .ZN(n11908) );
  NAND2_X1 U9651 ( .A1(n6838), .A2(n11224), .ZN(n11235) );
  OR2_X2 U9652 ( .A1(n7714), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7742) );
  OAI21_X1 U9653 ( .B1(n12622), .B2(n12621), .A(n12620), .ZN(n12624) );
  NAND3_X1 U9654 ( .A1(n6844), .A2(n6842), .A3(n6841), .ZN(P1_U3262) );
  INV_X1 U9655 ( .A(n7419), .ZN(n8155) );
  NOR2_X1 U9656 ( .A1(n15155), .A2(n15156), .ZN(n15154) );
  NAND2_X1 U9657 ( .A1(n11198), .A2(n6552), .ZN(n8144) );
  NAND3_X1 U9658 ( .A1(n7118), .A2(n7117), .A3(n7121), .ZN(n15054) );
  NAND2_X1 U9659 ( .A1(n9802), .A2(n9803), .ZN(n9801) );
  NAND2_X1 U9660 ( .A1(n6876), .A2(n6874), .ZN(n9717) );
  INV_X1 U9661 ( .A(n12603), .ZN(n6887) );
  NAND2_X1 U9662 ( .A1(n15405), .A2(n15700), .ZN(n6846) );
  NAND2_X1 U9663 ( .A1(n15292), .A2(n6847), .ZN(n15405) );
  INV_X1 U9664 ( .A(n10128), .ZN(n6902) );
  NAND2_X1 U9665 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  INV_X1 U9666 ( .A(n10139), .ZN(n6868) );
  NAND3_X1 U9667 ( .A1(n7406), .A2(n9072), .A3(n7405), .ZN(n9074) );
  NAND2_X1 U9668 ( .A1(n9488), .A2(n9487), .ZN(n9505) );
  NAND2_X1 U9669 ( .A1(n7193), .A2(n7194), .ZN(n9457) );
  NAND2_X1 U9670 ( .A1(n7231), .A2(n6746), .ZN(n11894) );
  NAND2_X1 U9671 ( .A1(n7173), .A2(n7171), .ZN(n9406) );
  INV_X1 U9672 ( .A(n12927), .ZN(n12928) );
  NAND2_X1 U9673 ( .A1(n7097), .A2(n12938), .ZN(n7096) );
  AND2_X2 U9674 ( .A1(n9027), .A2(n6664), .ZN(n11671) );
  NAND2_X1 U9675 ( .A1(n14233), .A2(n8845), .ZN(n7615) );
  AOI21_X1 U9676 ( .B1(n15248), .B2(n15655), .A(n15247), .ZN(n15249) );
  NAND2_X1 U9677 ( .A1(n14245), .A2(n14244), .ZN(n14522) );
  NAND2_X1 U9678 ( .A1(n6858), .A2(n8089), .ZN(n8137) );
  NAND2_X1 U9679 ( .A1(n8109), .A2(n7648), .ZN(n6858) );
  NAND2_X1 U9680 ( .A1(n6883), .A2(n6882), .ZN(n14611) );
  NAND2_X1 U9681 ( .A1(n9717), .A2(n9718), .ZN(n9716) );
  NAND2_X1 U9682 ( .A1(n6936), .A2(n6933), .ZN(n6926) );
  INV_X2 U9683 ( .A(n10153), .ZN(n15566) );
  NAND2_X1 U9684 ( .A1(n7201), .A2(n7197), .ZN(n6885) );
  NAND2_X1 U9685 ( .A1(n10683), .A2(n6552), .ZN(n7723) );
  AOI21_X1 U9686 ( .B1(n6887), .B2(n6886), .A(n12608), .ZN(n12609) );
  INV_X1 U9687 ( .A(n12454), .ZN(n12450) );
  OR2_X1 U9688 ( .A1(n6594), .A2(n10614), .ZN(n8527) );
  NAND2_X1 U9689 ( .A1(n7676), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U9690 ( .A1(n10632), .A2(n6552), .ZN(n7972) );
  NAND2_X1 U9691 ( .A1(n7823), .A2(n7579), .ZN(n7583) );
  INV_X1 U9692 ( .A(n7153), .ZN(n7152) );
  NAND2_X1 U9693 ( .A1(n6865), .A2(n9998), .ZN(n9999) );
  NAND2_X1 U9694 ( .A1(n9995), .A2(n6866), .ZN(n6865) );
  INV_X1 U9695 ( .A(n7894), .ZN(n7680) );
  NAND2_X1 U9696 ( .A1(n10580), .A2(n15975), .ZN(n7919) );
  NAND4_X1 U9697 ( .A1(n7708), .A2(n8094), .A3(n7727), .A4(n7707), .ZN(n7731)
         );
  NAND3_X1 U9698 ( .A1(n7543), .A2(n11885), .A3(n7544), .ZN(n10159) );
  OAI21_X1 U9699 ( .B1(n7419), .B2(n8176), .A(n6920), .ZN(n6922) );
  OR2_X1 U9700 ( .A1(n9875), .A2(n9829), .ZN(n9853) );
  AOI21_X1 U9701 ( .B1(n7223), .B2(n7226), .A(n7222), .ZN(n7221) );
  INV_X1 U9702 ( .A(n7311), .ZN(n11286) );
  NAND2_X1 U9703 ( .A1(n11285), .A2(n11284), .ZN(n7311) );
  NAND2_X1 U9704 ( .A1(n9687), .A2(n9688), .ZN(n9686) );
  NAND2_X1 U9705 ( .A1(n6872), .A2(n6871), .ZN(n6870) );
  INV_X1 U9706 ( .A(n9680), .ZN(n6872) );
  NAND3_X1 U9707 ( .A1(n9708), .A2(n9707), .A3(n6750), .ZN(n6876) );
  AND2_X2 U9708 ( .A1(n7083), .A2(n9174), .ZN(n9323) );
  NAND2_X1 U9709 ( .A1(n11812), .A2(n7232), .ZN(n7231) );
  NAND3_X1 U9710 ( .A1(n12938), .A2(n7097), .A3(n12940), .ZN(n6880) );
  INV_X1 U9711 ( .A(n7095), .ZN(n12939) );
  NAND2_X1 U9712 ( .A1(n6926), .A2(n6931), .ZN(n14242) );
  NAND2_X1 U9713 ( .A1(n8178), .A2(n8177), .ZN(n8209) );
  NAND2_X1 U9714 ( .A1(n11232), .A2(n11231), .ZN(n11388) );
  NAND2_X1 U9715 ( .A1(n11180), .A2(n13155), .ZN(n11057) );
  NAND2_X1 U9716 ( .A1(n12680), .A2(n12679), .ZN(n12693) );
  NAND2_X1 U9717 ( .A1(n12638), .A2(n12639), .ZN(n12680) );
  NOR2_X1 U9718 ( .A1(n7745), .A2(n7744), .ZN(n7746) );
  NAND2_X2 U9719 ( .A1(n10197), .A2(n10196), .ZN(n15053) );
  NAND2_X1 U9720 ( .A1(n7431), .A2(n7429), .ZN(n7425) );
  NAND2_X1 U9721 ( .A1(n7425), .A2(n7694), .ZN(n8028) );
  NAND4_X2 U9722 ( .A1(n7877), .A2(n7876), .A3(n7875), .A4(n7874), .ZN(n15666)
         );
  XNOR2_X2 U9723 ( .A(n15276), .B(n15057), .ZN(n15039) );
  NOR2_X2 U9724 ( .A1(n8012), .A2(n10744), .ZN(n8038) );
  AOI21_X1 U9725 ( .B1(n7272), .B2(n6618), .A(n12915), .ZN(n13339) );
  INV_X1 U9726 ( .A(n12651), .ZN(n15529) );
  NAND3_X1 U9727 ( .A1(n14967), .A2(n6903), .A3(n7655), .ZN(n6898) );
  NAND2_X1 U9728 ( .A1(n7124), .A2(n6901), .ZN(n15155) );
  NAND3_X1 U9729 ( .A1(n7132), .A2(n7126), .A3(n6902), .ZN(n6901) );
  NAND2_X1 U9730 ( .A1(n11176), .A2(n6552), .ZN(n8101) );
  NAND2_X1 U9731 ( .A1(n11036), .A2(n6552), .ZN(n8116) );
  NOR2_X1 U9732 ( .A1(n15753), .A2(n6903), .ZN(n7023) );
  AND2_X2 U9733 ( .A1(n12742), .A2(n13723), .ZN(n9066) );
  NAND2_X1 U9734 ( .A1(n10558), .A2(n10555), .ZN(n6915) );
  NAND2_X1 U9735 ( .A1(n10558), .A2(n6912), .ZN(n6911) );
  OR2_X1 U9736 ( .A1(n10557), .A2(n6915), .ZN(n12726) );
  OR2_X1 U9737 ( .A1(n15864), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U9738 ( .A1(n9587), .A2(n6918), .ZN(n6917) );
  NAND2_X1 U9739 ( .A1(n7419), .A2(n8156), .ZN(n8178) );
  AOI21_X1 U9740 ( .B1(n6921), .B2(n8177), .A(n8208), .ZN(n6920) );
  NAND2_X1 U9741 ( .A1(n14265), .A2(n14273), .ZN(n6936) );
  NAND2_X1 U9742 ( .A1(n6923), .A2(n6927), .ZN(n10270) );
  NAND2_X1 U9743 ( .A1(n14265), .A2(n6924), .ZN(n6923) );
  NAND2_X1 U9744 ( .A1(n9552), .A2(n9553), .ZN(n12798) );
  NAND3_X1 U9745 ( .A1(n7083), .A2(n9174), .A3(n7253), .ZN(n6937) );
  NAND2_X1 U9746 ( .A1(n13348), .A2(n13347), .ZN(n13595) );
  NAND2_X1 U9747 ( .A1(n11665), .A2(n12385), .ZN(n6942) );
  NAND2_X1 U9748 ( .A1(n11664), .A2(n11663), .ZN(n6943) );
  NAND2_X1 U9749 ( .A1(n6946), .A2(n9634), .ZN(n11658) );
  INV_X1 U9750 ( .A(n9630), .ZN(n6948) );
  NAND2_X1 U9751 ( .A1(n6951), .A2(n12182), .ZN(n13104) );
  NAND4_X1 U9752 ( .A1(n7083), .A2(n9175), .A3(n9322), .A4(n9616), .ZN(n9618)
         );
  NAND3_X1 U9753 ( .A1(n7083), .A2(n9175), .A3(n9322), .ZN(n9614) );
  INV_X1 U9754 ( .A(n12305), .ZN(n6952) );
  NAND2_X1 U9755 ( .A1(n13034), .A2(n6723), .ZN(n6961) );
  OAI211_X1 U9756 ( .C1(n13034), .C2(n6966), .A(n6962), .B(n6961), .ZN(n12392)
         );
  NAND2_X1 U9757 ( .A1(n13034), .A2(n6976), .ZN(n6968) );
  AOI21_X1 U9758 ( .B1(n13034), .B2(n13035), .A(n7634), .ZN(n13117) );
  INV_X1 U9759 ( .A(n12387), .ZN(n6978) );
  NAND2_X1 U9760 ( .A1(n15479), .A2(n6661), .ZN(n6984) );
  NAND2_X1 U9761 ( .A1(n6984), .A2(n7498), .ZN(n10245) );
  AND2_X2 U9762 ( .A1(n6984), .A2(n6983), .ZN(n10246) );
  AOI21_X1 U9763 ( .B1(n15479), .B2(n6720), .A(n6985), .ZN(n6987) );
  NAND3_X1 U9764 ( .A1(n15452), .A2(n6988), .A3(n10080), .ZN(n10079) );
  NAND2_X1 U9765 ( .A1(n15462), .A2(n6993), .ZN(n6990) );
  NAND2_X1 U9766 ( .A1(n6998), .A2(n15438), .ZN(n15967) );
  OAI21_X1 U9767 ( .B1(n15439), .B2(n15440), .A(n15441), .ZN(n6998) );
  NOR2_X2 U9768 ( .A1(n15969), .A2(n10058), .ZN(n15439) );
  NAND2_X1 U9769 ( .A1(n12924), .A2(n6683), .ZN(n6999) );
  NAND2_X1 U9770 ( .A1(n7007), .A2(n7008), .ZN(n12892) );
  OR2_X1 U9771 ( .A1(n12872), .A2(n6609), .ZN(n7007) );
  INV_X4 U9772 ( .A(n12926), .ZN(n9602) );
  MUX2_X1 U9773 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9538), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7020) );
  NAND3_X1 U9774 ( .A1(n7027), .A2(n7024), .A3(n7021), .ZN(P2_U3233) );
  MUX2_X1 U9775 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10864), .S(n14049), .Z(
        n14048) );
  XNOR2_X1 U9776 ( .A(n11473), .B(n15887), .ZN(n15879) );
  NAND2_X1 U9777 ( .A1(n11114), .A2(n11075), .ZN(n11077) );
  NAND2_X1 U9778 ( .A1(n11115), .A2(n11116), .ZN(n11114) );
  OAI21_X1 U9779 ( .B1(n7068), .B2(n11247), .A(n7064), .ZN(n11265) );
  XNOR2_X1 U9780 ( .A(n11249), .B(n11244), .ZN(n11247) );
  AOI21_X1 U9781 ( .B1(n11918), .B2(n6760), .A(n7069), .ZN(n13163) );
  XNOR2_X1 U9782 ( .A(n7070), .B(P3_REG1_REG_11__SCAN_IN), .ZN(n11770) );
  NAND3_X1 U9783 ( .A1(n9558), .A2(n11792), .A3(n11793), .ZN(n7081) );
  NOR2_X2 U9784 ( .A1(n9336), .A2(n9013), .ZN(n7083) );
  NOR2_X2 U9785 ( .A1(n9010), .A2(n9095), .ZN(n9174) );
  NAND2_X1 U9786 ( .A1(n9597), .A2(n6641), .ZN(n13356) );
  NAND2_X1 U9787 ( .A1(n7086), .A2(n7084), .ZN(n9600) );
  NAND2_X1 U9788 ( .A1(n9597), .A2(n6738), .ZN(n7086) );
  NAND2_X1 U9789 ( .A1(n7095), .A2(n12936), .ZN(n7097) );
  NAND2_X1 U9790 ( .A1(n9363), .A2(n6767), .ZN(n9410) );
  NAND2_X1 U9791 ( .A1(n9285), .A2(n7101), .ZN(n9342) );
  NAND2_X1 U9792 ( .A1(n9285), .A2(n9284), .ZN(n9300) );
  NAND3_X1 U9793 ( .A1(n9082), .A2(n9081), .A3(n9100), .ZN(n9121) );
  XNOR2_X2 U9794 ( .A(n15487), .B(n12519), .ZN(n12653) );
  AND3_X2 U9795 ( .A1(n7708), .A2(n8094), .A3(n7707), .ZN(n7105) );
  NAND2_X2 U9796 ( .A1(n7105), .A2(n6694), .ZN(n7714) );
  NAND2_X1 U9797 ( .A1(n7714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U9798 ( .A1(n15513), .A2(n10111), .ZN(n10113) );
  NAND2_X1 U9799 ( .A1(n10135), .A2(n7119), .ZN(n7118) );
  NAND2_X1 U9800 ( .A1(n15172), .A2(n6650), .ZN(n7125) );
  NAND3_X1 U9801 ( .A1(n7130), .A2(n6642), .A3(n12664), .ZN(n7127) );
  NAND3_X1 U9802 ( .A1(n7130), .A2(n6650), .A3(n12664), .ZN(n7129) );
  NAND2_X1 U9803 ( .A1(n7131), .A2(n7132), .ZN(n15173) );
  NAND2_X1 U9804 ( .A1(n10128), .A2(n7134), .ZN(n7131) );
  AOI21_X1 U9805 ( .B1(n7496), .B2(n7495), .A(n6743), .ZN(n10014) );
  OAI21_X1 U9806 ( .B1(n10046), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10021), .ZN(
        n7138) );
  NAND2_X1 U9807 ( .A1(n10021), .A2(n7139), .ZN(n10046) );
  NAND2_X1 U9808 ( .A1(n10020), .A2(n11100), .ZN(n7139) );
  INV_X2 U9809 ( .A(n7676), .ZN(n7658) );
  NAND2_X4 U9810 ( .A1(n7151), .A2(n7149), .ZN(n7676) );
  NAND3_X1 U9811 ( .A1(n7656), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U9812 ( .A1(n7408), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U9813 ( .A1(n7154), .A2(n7152), .ZN(n7685) );
  NAND2_X1 U9814 ( .A1(n9375), .A2(n6634), .ZN(n7173) );
  NAND2_X1 U9815 ( .A1(n9242), .A2(n7184), .ZN(n7182) );
  INV_X1 U9816 ( .A(n7372), .ZN(n7191) );
  NAND2_X1 U9817 ( .A1(n9430), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U9818 ( .A1(n11242), .A2(n11241), .ZN(n7195) );
  NAND2_X1 U9819 ( .A1(n7196), .A2(n11067), .ZN(n11242) );
  NAND2_X1 U9820 ( .A1(n11125), .A2(n11126), .ZN(n7196) );
  XNOR2_X1 U9821 ( .A(n7199), .B(n13325), .ZN(n7198) );
  AND2_X1 U9822 ( .A1(n13324), .A2(n13323), .ZN(n7200) );
  AND2_X1 U9823 ( .A1(n7202), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n13155) );
  MUX2_X1 U9824 ( .A(n11399), .B(n11415), .S(n13319), .Z(n7202) );
  NAND2_X1 U9825 ( .A1(n10958), .A2(n9787), .ZN(n9674) );
  NAND2_X1 U9826 ( .A1(n7206), .A2(n6744), .ZN(n9764) );
  NAND3_X1 U9827 ( .A1(n9753), .A2(n9752), .A3(n6725), .ZN(n7206) );
  NAND2_X1 U9828 ( .A1(n7208), .A2(n7210), .ZN(n9703) );
  NAND3_X1 U9829 ( .A1(n9692), .A2(n9691), .A3(n7209), .ZN(n7208) );
  INV_X1 U9830 ( .A(n9727), .ZN(n7212) );
  NAND2_X1 U9831 ( .A1(n9785), .A2(n7216), .ZN(n7213) );
  NAND2_X1 U9832 ( .A1(n7213), .A2(n7214), .ZN(n9793) );
  NAND2_X1 U9833 ( .A1(n7220), .A2(n7221), .ZN(n9928) );
  NAND2_X1 U9834 ( .A1(n9812), .A2(n7223), .ZN(n7220) );
  NAND2_X1 U9835 ( .A1(n7230), .A2(n7229), .ZN(n8905) );
  NAND2_X1 U9836 ( .A1(n12238), .A2(n6730), .ZN(n7237) );
  NAND2_X1 U9837 ( .A1(n12238), .A2(n7242), .ZN(n7241) );
  NAND2_X1 U9838 ( .A1(n7237), .A2(n7236), .ZN(n13534) );
  NAND2_X1 U9839 ( .A1(n12238), .A2(n12860), .ZN(n12324) );
  INV_X1 U9840 ( .A(n7255), .ZN(n7252) );
  NAND2_X1 U9841 ( .A1(n7252), .A2(n9323), .ZN(n9030) );
  NAND2_X1 U9842 ( .A1(n7257), .A2(n7258), .ZN(n12239) );
  NAND2_X1 U9843 ( .A1(n12039), .A2(n6659), .ZN(n7257) );
  NAND2_X1 U9844 ( .A1(n13371), .A2(n12761), .ZN(n7272) );
  AOI21_X1 U9845 ( .B1(n7271), .B2(n12907), .A(n7273), .ZN(n7269) );
  AND2_X1 U9846 ( .A1(n8479), .A2(n7282), .ZN(n7279) );
  OAI21_X2 U9847 ( .B1(n8966), .B2(n7292), .A(n7288), .ZN(n14265) );
  NAND2_X1 U9848 ( .A1(n7302), .A2(n7298), .ZN(n8958) );
  NAND2_X1 U9849 ( .A1(n14427), .A2(n7304), .ZN(n7302) );
  NAND2_X1 U9850 ( .A1(n10270), .A2(n10271), .ZN(n7306) );
  NAND2_X1 U9851 ( .A1(n6606), .A2(n14049), .ZN(n8553) );
  OAI21_X2 U9852 ( .B1(n7309), .B2(n7506), .A(n7310), .ZN(n11301) );
  NAND2_X1 U9853 ( .A1(n7309), .A2(n14668), .ZN(n7310) );
  OAI22_X1 U9854 ( .A1(n15718), .A2(n7309), .B1(n9940), .B2(n10633), .ZN(n8636) );
  OR2_X1 U9855 ( .A1(n11288), .A2(n7313), .ZN(n7312) );
  INV_X1 U9856 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U9857 ( .A1(n11286), .A2(n11307), .ZN(n7315) );
  INV_X1 U9858 ( .A(n13291), .ZN(n7317) );
  NAND2_X1 U9859 ( .A1(n7317), .A2(n7322), .ZN(n7320) );
  NAND2_X1 U9860 ( .A1(n7323), .A2(n13291), .ZN(n13269) );
  OR2_X1 U9861 ( .A1(n13267), .A2(n13294), .ZN(n7323) );
  NAND2_X1 U9862 ( .A1(n13165), .A2(n13199), .ZN(n7324) );
  OR2_X1 U9863 ( .A1(n13165), .A2(n7329), .ZN(n7328) );
  NAND2_X1 U9864 ( .A1(n7334), .A2(n7330), .ZN(n11920) );
  NOR2_X1 U9865 ( .A1(n7331), .A2(n7335), .ZN(n7330) );
  NAND2_X1 U9866 ( .A1(n15885), .A2(n6765), .ZN(n7334) );
  NAND2_X1 U9867 ( .A1(n15885), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11462) );
  NOR2_X1 U9868 ( .A1(n11464), .A2(n12076), .ZN(n7338) );
  INV_X1 U9869 ( .A(n11252), .ZN(n7340) );
  NAND2_X1 U9870 ( .A1(n13258), .A2(n7344), .ZN(n7342) );
  AND2_X1 U9871 ( .A1(n13258), .A2(n13220), .ZN(n13221) );
  NAND2_X1 U9872 ( .A1(n7346), .A2(n7345), .ZN(n8490) );
  NAND2_X1 U9873 ( .A1(n7347), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U9874 ( .A1(n7348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U9875 ( .A1(n8491), .A2(n8493), .ZN(n7348) );
  NAND2_X1 U9876 ( .A1(n13561), .A2(n7351), .ZN(n7350) );
  NAND2_X1 U9877 ( .A1(n13391), .A2(n13387), .ZN(n13388) );
  NAND2_X1 U9878 ( .A1(n9173), .A2(n9172), .ZN(n9191) );
  OAI22_X2 U9879 ( .A1(n13901), .A2(n7362), .B1(n7363), .B2(n13849), .ZN(
        n13946) );
  NAND2_X1 U9880 ( .A1(n9582), .A2(n6739), .ZN(n13453) );
  NAND2_X1 U9881 ( .A1(n13794), .A2(n13795), .ZN(n7397) );
  NOR2_X1 U9882 ( .A1(n7399), .A2(n9569), .ZN(n7643) );
  XNOR2_X1 U9883 ( .A(n7407), .B(n7878), .ZN(n10586) );
  NAND2_X1 U9884 ( .A1(n7988), .A2(n7989), .ZN(n7431) );
  NAND2_X1 U9885 ( .A1(n15232), .A2(n7435), .ZN(n15230) );
  AND2_X2 U9886 ( .A1(n15073), .A2(n6741), .ZN(n14997) );
  NAND3_X2 U9887 ( .A1(n7442), .A2(n15683), .A3(n7443), .ZN(n11912) );
  NAND2_X1 U9888 ( .A1(n13125), .A2(n6632), .ZN(n13043) );
  NAND2_X1 U9889 ( .A1(n13068), .A2(n6740), .ZN(n13009) );
  NAND2_X1 U9890 ( .A1(n12417), .A2(n7449), .ZN(n7448) );
  OAI211_X1 U9891 ( .C1(n12417), .C2(n7450), .A(n7448), .B(n12422), .ZN(
        P3_U3169) );
  NAND2_X1 U9892 ( .A1(n7464), .A2(n7465), .ZN(n12614) );
  NAND2_X1 U9893 ( .A1(n7464), .A2(n6745), .ZN(n12613) );
  INV_X1 U9894 ( .A(n12611), .ZN(n7466) );
  NAND2_X1 U9895 ( .A1(n12564), .A2(n6747), .ZN(n7470) );
  NAND3_X1 U9896 ( .A1(n7468), .A2(n12576), .A3(n7467), .ZN(n12579) );
  NAND3_X1 U9897 ( .A1(n12556), .A2(n12555), .A3(n7469), .ZN(n7468) );
  NAND2_X1 U9898 ( .A1(n7476), .A2(n7477), .ZN(n12602) );
  NAND2_X1 U9899 ( .A1(n7483), .A2(n7485), .ZN(n12533) );
  NAND3_X1 U9900 ( .A1(n12525), .A2(n12524), .A3(n7484), .ZN(n7483) );
  OR2_X2 U9901 ( .A1(n15450), .A2(n15730), .ZN(n7494) );
  INV_X1 U9902 ( .A(n10075), .ZN(n7490) );
  AOI21_X1 U9903 ( .B1(n10075), .B2(n7493), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7492) );
  INV_X1 U9904 ( .A(n15453), .ZN(n7493) );
  INV_X1 U9905 ( .A(n7494), .ZN(n15451) );
  INV_X1 U9906 ( .A(n10054), .ZN(n10055) );
  INV_X1 U9907 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U9908 ( .A1(n7499), .A2(n6615), .ZN(n7498) );
  INV_X1 U9909 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7505) );
  INV_X1 U9910 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7506) );
  NAND3_X1 U9911 ( .A1(n6631), .A2(n6786), .A3(n14310), .ZN(n14281) );
  INV_X1 U9912 ( .A(n7513), .ZN(n11988) );
  INV_X1 U9913 ( .A(n11321), .ZN(n7514) );
  NAND2_X1 U9914 ( .A1(n7514), .A2(n6626), .ZN(n11738) );
  NOR2_X2 U9915 ( .A1(n7520), .A2(n14578), .ZN(n7519) );
  NAND2_X1 U9916 ( .A1(n14236), .A2(n7522), .ZN(n12704) );
  NAND2_X1 U9917 ( .A1(n14236), .A2(n7525), .ZN(n10537) );
  NAND2_X1 U9918 ( .A1(n14236), .A2(n13807), .ZN(n10275) );
  NOR2_X1 U9919 ( .A1(n7526), .A2(n7725), .ZN(n8093) );
  NAND4_X1 U9920 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n8032), .ZN(n7526)
         );
  NAND2_X1 U9921 ( .A1(n15053), .A2(n7530), .ZN(n7527) );
  NAND2_X1 U9922 ( .A1(n10155), .A2(n7542), .ZN(n7543) );
  NAND2_X1 U9923 ( .A1(n7545), .A2(n10157), .ZN(n11886) );
  NAND2_X1 U9924 ( .A1(n15545), .A2(n15546), .ZN(n7545) );
  INV_X1 U9925 ( .A(n15487), .ZN(n15532) );
  AND2_X2 U9926 ( .A1(n15111), .A2(n10189), .ZN(n15066) );
  OR2_X1 U9927 ( .A1(n10205), .A2(n15007), .ZN(n7552) );
  NAND2_X1 U9928 ( .A1(n12099), .A2(n7555), .ZN(n10176) );
  NOR2_X2 U9929 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7560) );
  AND2_X2 U9930 ( .A1(n7560), .A2(n7559), .ZN(n7833) );
  NAND3_X1 U9931 ( .A1(n12129), .A2(n12126), .A3(n7570), .ZN(n7566) );
  NAND2_X1 U9932 ( .A1(n14754), .A2(n6617), .ZN(n7573) );
  NAND2_X1 U9933 ( .A1(n7581), .A2(n7583), .ZN(n11422) );
  NAND2_X1 U9934 ( .A1(n7823), .A2(n7822), .ZN(n15484) );
  OAI21_X1 U9935 ( .B1(n11595), .B2(n11596), .A(n7964), .ZN(n7985) );
  NAND2_X1 U9936 ( .A1(n11595), .A2(n7964), .ZN(n7586) );
  NAND2_X1 U9937 ( .A1(n14732), .A2(n7590), .ZN(n7587) );
  INV_X1 U9938 ( .A(n8152), .ZN(n7593) );
  NAND2_X1 U9939 ( .A1(n14762), .A2(n7596), .ZN(n7594) );
  NAND2_X1 U9940 ( .A1(n7594), .A2(n7595), .ZN(n8136) );
  INV_X2 U9941 ( .A(n8530), .ZN(n8849) );
  NAND3_X1 U9942 ( .A1(n8516), .A2(n7602), .A3(P2_REG3_REG_2__SCAN_IN), .ZN(
        n8547) );
  INV_X1 U9943 ( .A(n7605), .ZN(n14276) );
  NAND2_X1 U9944 ( .A1(n11549), .A2(n11552), .ZN(n7614) );
  NAND2_X1 U9945 ( .A1(n11549), .A2(n7611), .ZN(n7610) );
  NAND2_X2 U9946 ( .A1(n14233), .A2(n6696), .ZN(n14222) );
  NAND3_X1 U9947 ( .A1(n14222), .A2(n14223), .A3(n15797), .ZN(n10277) );
  INV_X1 U9948 ( .A(n14299), .ZN(n7621) );
  NOR2_X1 U9949 ( .A1(n14314), .A2(n7628), .ZN(n14298) );
  NAND2_X1 U9950 ( .A1(n8512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8513) );
  INV_X1 U9951 ( .A(n15235), .ZN(n10226) );
  INV_X1 U9952 ( .A(n10009), .ZN(n10001) );
  AOI21_X1 U9953 ( .B1(n9612), .B2(n13562), .A(n9611), .ZN(n12714) );
  NAND2_X1 U9954 ( .A1(n12091), .A2(n10126), .ZN(n10128) );
  NAND2_X1 U9955 ( .A1(n12185), .A2(n12184), .ZN(n13106) );
  NAND2_X1 U9956 ( .A1(n14998), .A2(n15224), .ZN(n14984) );
  AND2_X2 U9957 ( .A1(n14997), .A2(n15003), .ZN(n14998) );
  NAND2_X1 U9958 ( .A1(n15566), .A2(n7782), .ZN(n7784) );
  AND2_X1 U9959 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  NAND2_X1 U9960 ( .A1(n12415), .A2(n12371), .ZN(n12381) );
  XNOR2_X1 U9961 ( .A(n8911), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8916) );
  INV_X1 U9962 ( .A(n11235), .ZN(n11232) );
  INV_X1 U9963 ( .A(n12914), .ZN(n12923) );
  NAND2_X1 U9964 ( .A1(n8987), .A2(n15811), .ZN(n11321) );
  CLKBUF_X1 U9965 ( .A(n8463), .Z(n15430) );
  OR2_X1 U9966 ( .A1(n15564), .A2(n6538), .ZN(n7797) );
  OR2_X1 U9967 ( .A1(n6603), .A2(n15564), .ZN(n7793) );
  XNOR2_X1 U9968 ( .A(n7801), .B(n7800), .ZN(n11041) );
  AND4_X2 U9969 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n15564)
         );
  CLKBUF_X1 U9970 ( .A(n15527), .Z(n15528) );
  INV_X1 U9971 ( .A(n7985), .ZN(n7987) );
  XNOR2_X1 U9972 ( .A(n12415), .B(n12413), .ZN(n13076) );
  OAI21_X1 U9973 ( .B1(n12495), .B2(n6538), .A(n7780), .ZN(n7781) );
  INV_X1 U9974 ( .A(n14392), .ZN(n14405) );
  NAND2_X1 U9975 ( .A1(n14392), .A2(n13924), .ZN(n14394) );
  NAND2_X1 U9976 ( .A1(n11369), .A2(n15804), .ZN(n11320) );
  AND2_X1 U9977 ( .A1(n12014), .A2(n8941), .ZN(n7627) );
  NOR2_X1 U9978 ( .A1(n14548), .A2(n14024), .ZN(n7628) );
  AND3_X1 U9979 ( .A1(n8298), .A2(n14683), .A3(n14685), .ZN(n7629) );
  AND2_X1 U9980 ( .A1(n9926), .A2(n9925), .ZN(n7630) );
  AND3_X1 U9981 ( .A1(n14232), .A2(n14228), .A3(n10276), .ZN(n7631) );
  OR2_X1 U9982 ( .A1(n15239), .A2(n15214), .ZN(n7632) );
  INV_X1 U9983 ( .A(n14649), .ZN(n9001) );
  INV_X1 U9984 ( .A(n15864), .ZN(n8995) );
  NAND2_X1 U9985 ( .A1(n8749), .A2(n8748), .ZN(n8757) );
  AND4_X1 U9986 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9924), .ZN(n7633)
         );
  AND2_X1 U9987 ( .A1(n12383), .A2(n13410), .ZN(n7634) );
  AND2_X1 U9988 ( .A1(n8135), .A2(n8134), .ZN(n7635) );
  AND2_X1 U9989 ( .A1(n12580), .A2(n10127), .ZN(n7636) );
  NOR2_X1 U9990 ( .A1(n10161), .A2(n12655), .ZN(n7637) );
  OR2_X2 U9991 ( .A1(n15174), .A2(n15183), .ZN(n7638) );
  AND2_X1 U9992 ( .A1(n12492), .A2(n10209), .ZN(n7639) );
  AND2_X1 U9993 ( .A1(n9664), .A2(n13601), .ZN(n7640) );
  AND2_X1 U9994 ( .A1(n8455), .A2(n7654), .ZN(n7641) );
  NOR2_X1 U9995 ( .A1(n12244), .A2(n12774), .ZN(n7642) );
  AND2_X1 U9996 ( .A1(n8048), .A2(n8047), .ZN(n7644) );
  AND2_X1 U9997 ( .A1(n12578), .A2(n12642), .ZN(n7645) );
  OR2_X1 U9998 ( .A1(n13807), .A2(n14018), .ZN(n7646) );
  INV_X1 U9999 ( .A(n14457), .ZN(n14507) );
  NOR2_X1 U10000 ( .A1(n11338), .A2(n11298), .ZN(n7647) );
  INV_X1 U10001 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10045) );
  AND2_X1 U10002 ( .A1(n8089), .A2(n8088), .ZN(n7648) );
  NAND2_X1 U10003 ( .A1(n15563), .A2(n8429), .ZN(n15388) );
  INV_X1 U10004 ( .A(n15388), .ZN(n15682) );
  INV_X1 U10005 ( .A(n7976), .ZN(n8216) );
  AND2_X1 U10006 ( .A1(n10131), .A2(n15314), .ZN(n7649) );
  INV_X2 U10007 ( .A(n7676), .ZN(n10567) );
  AND2_X1 U10008 ( .A1(n8138), .A2(n8092), .ZN(n7650) );
  INV_X1 U10009 ( .A(n9065), .ZN(n9531) );
  AND2_X1 U10010 ( .A1(n12922), .A2(n12921), .ZN(n7652) );
  XNOR2_X1 U10011 ( .A(n8871), .B(n9990), .ZN(n14221) );
  AND2_X1 U10012 ( .A1(n15116), .A2(n10183), .ZN(n7653) );
  AND2_X1 U10013 ( .A1(n8454), .A2(n15491), .ZN(n7654) );
  NAND2_X1 U10014 ( .A1(n9690), .A2(n9689), .ZN(n9691) );
  AND2_X1 U10015 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  NAND2_X1 U10016 ( .A1(n6529), .A2(n9719), .ZN(n9720) );
  AND2_X1 U10017 ( .A1(n12572), .A2(n12563), .ZN(n12564) );
  INV_X1 U10018 ( .A(n12455), .ZN(n12449) );
  NAND2_X1 U10019 ( .A1(n12920), .A2(n12926), .ZN(n12921) );
  OR2_X1 U10020 ( .A1(n14604), .A2(n13839), .ZN(n8941) );
  NAND2_X1 U10021 ( .A1(n12614), .A2(n12616), .ZN(n12617) );
  NOR2_X1 U10022 ( .A1(n11471), .A2(n11944), .ZN(n11458) );
  INV_X1 U10023 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10024 ( .A1(n11659), .A2(n12755), .ZN(n11660) );
  OR2_X1 U10025 ( .A1(n9516), .A2(n9038), .ZN(n9044) );
  INV_X1 U10026 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9008) );
  INV_X1 U10027 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8639) );
  OAI21_X1 U10028 ( .B1(n9671), .B2(n11772), .A(n10006), .ZN(n8919) );
  INV_X1 U10029 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U10030 ( .A1(n15211), .A2(n14766), .ZN(n10127) );
  INV_X1 U10031 ( .A(n7942), .ZN(n7682) );
  NAND2_X1 U10032 ( .A1(n12413), .A2(n13427), .ZN(n12370) );
  OAI21_X1 U10033 ( .B1(n13827), .B2(n14022), .A(n13964), .ZN(n13786) );
  INV_X1 U10034 ( .A(n8830), .ZN(n8507) );
  OR2_X1 U10035 ( .A1(n6596), .A2(n8535), .ZN(n8922) );
  INV_X1 U10036 ( .A(n10555), .ZN(n10556) );
  INV_X1 U10037 ( .A(n14503), .ZN(n8670) );
  NAND2_X1 U10038 ( .A1(n7832), .A2(n10575), .ZN(n7859) );
  INV_X1 U10039 ( .A(n8439), .ZN(n8440) );
  OR2_X1 U10040 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  INV_X1 U10041 ( .A(n15329), .ZN(n15181) );
  INV_X1 U10042 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7950) );
  INV_X1 U10043 ( .A(n12508), .ZN(n11489) );
  INV_X1 U10044 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7710) );
  AND2_X1 U10045 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  AND2_X1 U10046 ( .A1(n8079), .A2(n8078), .ZN(n8080) );
  INV_X1 U10047 ( .A(n13012), .ZN(n12365) );
  INV_X1 U10048 ( .A(n13041), .ZN(n12350) );
  INV_X1 U10049 ( .A(n12793), .ZN(n12794) );
  INV_X1 U10050 ( .A(n13365), .ZN(n9598) );
  INV_X1 U10051 ( .A(n13381), .ZN(n13404) );
  OR2_X1 U10052 ( .A1(n11804), .A2(n12821), .ZN(n11819) );
  INV_X1 U10053 ( .A(n11670), .ZN(n12809) );
  AND2_X1 U10054 ( .A1(n11217), .A2(n11216), .ZN(n11219) );
  NAND2_X1 U10055 ( .A1(n8507), .A2(n8506), .ZN(n8838) );
  INV_X1 U10056 ( .A(n15797), .ZN(n10269) );
  INV_X1 U10057 ( .A(n10638), .ZN(n7812) );
  INV_X1 U10058 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10744) );
  INV_X1 U10059 ( .A(n12657), .ZN(n10164) );
  NAND2_X1 U10060 ( .A1(n10108), .A2(n10107), .ZN(n15530) );
  INV_X1 U10061 ( .A(n15108), .ZN(n10188) );
  NAND2_X1 U10062 ( .A1(n8086), .A2(n10813), .ZN(n8089) );
  NOR2_X1 U10063 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7698) );
  NOR2_X1 U10064 ( .A1(n10092), .A2(n10091), .ZN(n10033) );
  NOR2_X1 U10065 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  OR2_X1 U10066 ( .A1(n11698), .A2(n11697), .ZN(n11701) );
  INV_X1 U10067 ( .A(n13141), .ZN(n13512) );
  NAND2_X1 U10068 ( .A1(n15941), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10239) );
  INV_X1 U10069 ( .A(n13562), .ZN(n13507) );
  AND2_X1 U10070 ( .A1(n9551), .A2(n9656), .ZN(n13433) );
  NAND2_X1 U10071 ( .A1(n9527), .A2(n9526), .ZN(n12736) );
  NAND2_X1 U10072 ( .A1(n10625), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9127) );
  AND2_X1 U10073 ( .A1(n8676), .A2(n8675), .ZN(n8949) );
  OR2_X1 U10074 ( .A1(n8788), .A2(n13949), .ZN(n8809) );
  AND2_X1 U10075 ( .A1(n10957), .A2(n14214), .ZN(n10945) );
  INV_X1 U10076 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10890) );
  INV_X1 U10077 ( .A(n15850), .ZN(n9003) );
  NAND2_X1 U10078 ( .A1(n8909), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8910) );
  AND2_X1 U10079 ( .A1(n8365), .A2(n8363), .ZN(n14710) );
  AND2_X1 U10080 ( .A1(n14709), .A2(n8333), .ZN(n14743) );
  NAND2_X1 U10081 ( .A1(n8202), .A2(n8204), .ZN(n8205) );
  OR2_X1 U10082 ( .A1(n8462), .A2(n8461), .ZN(n8471) );
  INV_X1 U10083 ( .A(n14806), .ZN(n14798) );
  OR2_X1 U10084 ( .A1(n11016), .A2(n11017), .ZN(n11018) );
  NAND2_X1 U10085 ( .A1(n7873), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7770) );
  OR2_X1 U10086 ( .A1(n12224), .A2(n12223), .ZN(n12226) );
  NOR2_X1 U10087 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7744) );
  XNOR2_X1 U10088 ( .A(n8157), .B(n11009), .ZN(n8156) );
  XNOR2_X1 U10089 ( .A(n7667), .B(SI_2_), .ZN(n7809) );
  XNOR2_X1 U10090 ( .A(n12385), .B(n12829), .ZN(n12949) );
  INV_X1 U10091 ( .A(n13317), .ZN(n15886) );
  INV_X1 U10092 ( .A(n13329), .ZN(n15888) );
  AND2_X1 U10093 ( .A1(n11072), .A2(n13285), .ZN(n15895) );
  AND3_X1 U10094 ( .A1(n9154), .A2(n9153), .A3(n9152), .ZN(n15935) );
  NAND2_X1 U10095 ( .A1(n11419), .A2(n13553), .ZN(n13585) );
  AND2_X1 U10096 ( .A1(n9653), .A2(n9652), .ZN(n11413) );
  AND2_X1 U10097 ( .A1(n15954), .A2(n15936), .ZN(n13601) );
  AND2_X1 U10098 ( .A1(n13433), .A2(n15930), .ZN(n13630) );
  INV_X1 U10099 ( .A(n13630), .ZN(n15905) );
  INV_X1 U10100 ( .A(n11406), .ZN(n11410) );
  INV_X1 U10101 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9176) );
  AND2_X1 U10102 ( .A1(n9127), .A2(n9109), .ZN(n9110) );
  AND2_X1 U10103 ( .A1(n10963), .A2(n10962), .ZN(n13992) );
  INV_X1 U10104 ( .A(n14207), .ZN(n15744) );
  INV_X1 U10105 ( .A(n9977), .ZN(n11334) );
  NAND2_X1 U10106 ( .A1(n8995), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10278) );
  INV_X1 U10107 ( .A(n15835), .ZN(n15843) );
  AND2_X1 U10108 ( .A1(n15782), .A2(n8912), .ZN(n9000) );
  AND2_X1 U10109 ( .A1(n8891), .A2(n8914), .ZN(n15771) );
  INV_X1 U10110 ( .A(n8442), .ZN(n12429) );
  INV_X1 U10111 ( .A(n14960), .ZN(n15505) );
  INV_X1 U10112 ( .A(n15207), .ZN(n10213) );
  INV_X1 U10113 ( .A(n15013), .ZN(n15010) );
  AND2_X1 U10114 ( .A1(n10637), .A2(n10710), .ZN(n15665) );
  INV_X1 U10115 ( .A(n11485), .ZN(n12652) );
  INV_X1 U10116 ( .A(n15214), .ZN(n15581) );
  AND2_X1 U10117 ( .A1(n10151), .A2(n10150), .ZN(n15651) );
  INV_X1 U10118 ( .A(n15628), .ZN(n15668) );
  AND2_X1 U10119 ( .A1(n10647), .A2(n10565), .ZN(n10645) );
  INV_X1 U10120 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10056) );
  INV_X1 U10121 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10064) );
  AND2_X1 U10122 ( .A1(n11099), .A2(n11098), .ZN(n15865) );
  NAND2_X1 U10123 ( .A1(n11686), .A2(n11685), .ZN(n15867) );
  INV_X1 U10124 ( .A(n13458), .ZN(n13427) );
  INV_X1 U10125 ( .A(n13085), .ZN(n13144) );
  INV_X1 U10126 ( .A(n15865), .ZN(n15898) );
  INV_X1 U10127 ( .A(n15895), .ZN(n13237) );
  OR2_X1 U10128 ( .A1(n11419), .A2(n11418), .ZN(n13582) );
  INV_X2 U10129 ( .A(n13585), .ZN(n13580) );
  INV_X1 U10130 ( .A(n13418), .ZN(n13436) );
  NOR2_X1 U10131 ( .A1(n9665), .A2(n7640), .ZN(n9666) );
  INV_X1 U10132 ( .A(n15954), .ZN(n15951) );
  AND2_X1 U10133 ( .A1(n10237), .A2(n10236), .ZN(n15941) );
  INV_X1 U10134 ( .A(SI_13_), .ZN(n10815) );
  OR2_X1 U10135 ( .A1(n10960), .A2(n10956), .ZN(n14002) );
  AND2_X1 U10136 ( .A1(n14488), .A2(n10536), .ZN(n14465) );
  AND2_X2 U10137 ( .A1(n9000), .A2(n10943), .ZN(n15864) );
  NOR2_X1 U10138 ( .A1(n10531), .A2(n10530), .ZN(n12733) );
  INV_X1 U10139 ( .A(n15777), .ZN(n15778) );
  INV_X1 U10140 ( .A(n15062), .ZN(n15285) );
  INV_X1 U10141 ( .A(n15251), .ZN(n15028) );
  INV_X1 U10142 ( .A(n15322), .ZN(n15305) );
  OR2_X1 U10143 ( .A1(n15584), .A2(n15651), .ZN(n15095) );
  OR2_X1 U10144 ( .A1(n15584), .A2(n10210), .ZN(n15214) );
  INV_X1 U10145 ( .A(n15700), .ZN(n15698) );
  INV_X1 U10146 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11481) );
  INV_X1 U10147 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10937) );
  OAI211_X1 U10148 ( .C1(n10228), .C2(n15095), .A(n7632), .B(n10227), .ZN(
        P1_U3356) );
  XNOR2_X1 U10149 ( .A(n10104), .B(n10103), .ZN(SUB_1596_U62) );
  MUX2_X1 U10150 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10581), .Z(n7674) );
  AND2_X1 U10151 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7657) );
  INV_X1 U10152 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10578) );
  AOI21_X1 U10153 ( .B1(n7676), .B2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n7659) );
  OAI21_X1 U10154 ( .B1(n7676), .B2(n10578), .A(n7659), .ZN(n7660) );
  INV_X1 U10155 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7665) );
  INV_X1 U10156 ( .A(n7809), .ZN(n7666) );
  NAND2_X1 U10157 ( .A1(n7810), .A2(n7666), .ZN(n7837) );
  MUX2_X1 U10158 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7676), .Z(n7838) );
  NAND2_X1 U10159 ( .A1(n7838), .A2(SI_3_), .ZN(n7855) );
  NAND2_X1 U10160 ( .A1(n7667), .A2(SI_2_), .ZN(n7836) );
  NAND2_X1 U10161 ( .A1(n7837), .A2(n7668), .ZN(n7671) );
  MUX2_X1 U10162 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7676), .Z(n7672) );
  XNOR2_X1 U10163 ( .A(n7672), .B(SI_4_), .ZN(n7857) );
  NOR2_X1 U10164 ( .A1(n7838), .A2(SI_3_), .ZN(n7669) );
  NOR2_X1 U10165 ( .A1(n7857), .A2(n7669), .ZN(n7670) );
  NAND2_X1 U10166 ( .A1(n7672), .A2(SI_4_), .ZN(n7673) );
  NAND2_X1 U10167 ( .A1(n7674), .A2(SI_5_), .ZN(n7675) );
  BUF_X4 U10168 ( .A(n7676), .Z(n10575) );
  MUX2_X1 U10169 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10575), .Z(n7678) );
  NAND2_X1 U10170 ( .A1(n7678), .A2(SI_6_), .ZN(n7679) );
  MUX2_X1 U10171 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10575), .Z(n7683) );
  NAND2_X1 U10172 ( .A1(n7683), .A2(SI_8_), .ZN(n7684) );
  NAND2_X1 U10173 ( .A1(n7685), .A2(n7684), .ZN(n7965) );
  MUX2_X1 U10174 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10575), .Z(n7687) );
  NAND2_X1 U10175 ( .A1(n7687), .A2(SI_9_), .ZN(n7688) );
  MUX2_X1 U10176 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10575), .Z(n7689) );
  NAND2_X1 U10177 ( .A1(n7689), .A2(SI_10_), .ZN(n7690) );
  MUX2_X1 U10178 ( .A(n10661), .B(n10659), .S(n10581), .Z(n7691) );
  INV_X1 U10179 ( .A(n7691), .ZN(n7692) );
  NAND2_X1 U10180 ( .A1(n7692), .A2(SI_11_), .ZN(n7693) );
  MUX2_X1 U10181 ( .A(n9240), .B(n10751), .S(n10575), .Z(n7695) );
  INV_X1 U10182 ( .A(SI_12_), .ZN(n10663) );
  INV_X1 U10183 ( .A(n7695), .ZN(n7696) );
  NAND2_X1 U10184 ( .A1(n7696), .A2(SI_12_), .ZN(n7697) );
  AND2_X4 U10185 ( .A1(n7833), .A2(n7698), .ZN(n8094) );
  NOR2_X1 U10186 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n7701) );
  NOR2_X2 U10187 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7700) );
  NAND3_X1 U10188 ( .A1(n8096), .A2(n7702), .A3(n8140), .ZN(n7724) );
  INV_X2 U10189 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7945) );
  INV_X2 U10192 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7915) );
  NAND4_X1 U10193 ( .A1(n7968), .A2(n8029), .A3(n7945), .A4(n7915), .ZN(n7725)
         );
  NAND3_X1 U10194 ( .A1(n7734), .A2(n8161), .A3(n7703), .ZN(n7704) );
  NOR2_X1 U10195 ( .A1(n7725), .A2(n7704), .ZN(n7707) );
  NOR2_X1 U10196 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n7706) );
  NOR2_X1 U10197 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n7705) );
  AND3_X2 U10198 ( .A1(n7757), .A2(n7706), .A3(n7705), .ZN(n7727) );
  MUX2_X2 U10199 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7709), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n7712) );
  NAND2_X1 U10200 ( .A1(n7712), .A2(n7742), .ZN(n8463) );
  NAND2_X1 U10201 ( .A1(n7731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7713) );
  NAND2_X2 U10202 ( .A1(n8463), .A2(n12696), .ZN(n7832) );
  INV_X1 U10204 ( .A(n7880), .ZN(n7717) );
  NAND2_X1 U10205 ( .A1(n8094), .A2(n7717), .ZN(n7914) );
  INV_X1 U10206 ( .A(n7895), .ZN(n7718) );
  INV_X1 U10207 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10208 ( .A1(n7718), .A2(n7896), .ZN(n7944) );
  INV_X1 U10209 ( .A(n7967), .ZN(n7720) );
  NOR2_X1 U10210 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7719) );
  NAND2_X1 U10211 ( .A1(n7720), .A2(n7719), .ZN(n8008) );
  NAND2_X1 U10212 ( .A1(n7721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8030) );
  XNOR2_X1 U10213 ( .A(n8030), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U10214 ( .A1(n10977), .A2(n8064), .B1(n6604), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7722) );
  NAND2_X2 U10215 ( .A1(n7723), .A2(n7722), .ZN(n12098) );
  INV_X1 U10216 ( .A(n7724), .ZN(n7726) );
  INV_X1 U10217 ( .A(n7727), .ZN(n7728) );
  OAI21_X1 U10218 ( .B1(n7763), .B2(n7728), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7729) );
  MUX2_X1 U10219 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7729), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n7730) );
  INV_X1 U10220 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n12431) );
  INV_X1 U10221 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7733) );
  AND4_X1 U10222 ( .A1(n7757), .A2(n7734), .A3(n12431), .A4(n7733), .ZN(n7735)
         );
  NAND2_X1 U10223 ( .A1(n7732), .A2(n7735), .ZN(n8427) );
  XNOR2_X2 U10224 ( .A(n7736), .B(P1_IR_REG_25__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U10225 ( .A1(n8427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7737) );
  INV_X1 U10226 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10227 ( .A1(n7763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7741) );
  AND2_X2 U10228 ( .A1(n7760), .A2(n12430), .ZN(n12491) );
  INV_X1 U10229 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7743) );
  INV_X4 U10230 ( .A(n8219), .ZN(n10216) );
  NAND2_X1 U10231 ( .A1(n10216), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7756) );
  OR2_X2 U10232 ( .A1(n7974), .A2(n7973), .ZN(n7997) );
  XNOR2_X1 U10233 ( .A(n8040), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U10234 ( .A1(n8396), .A2(n12294), .ZN(n7755) );
  AND2_X2 U10235 ( .A1(n15426), .A2(n15428), .ZN(n7873) );
  NAND2_X1 U10236 ( .A1(n8145), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7754) );
  NAND2_X1 U10237 ( .A1(n8442), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7753) );
  NAND4_X1 U10238 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n15353) );
  INV_X1 U10239 ( .A(n15353), .ZN(n12217) );
  INV_X1 U10240 ( .A(n7757), .ZN(n12434) );
  INV_X1 U10241 ( .A(n7767), .ZN(n7759) );
  OR2_X4 U10242 ( .A1(n11002), .A2(n7760), .ZN(n15574) );
  INV_X1 U10243 ( .A(n15574), .ZN(n7764) );
  INV_X1 U10244 ( .A(n7732), .ZN(n7761) );
  NAND2_X1 U10245 ( .A1(n7761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7762) );
  AND2_X4 U10246 ( .A1(n10209), .A2(n10565), .ZN(n8266) );
  OAI22_X1 U10247 ( .A1(n6549), .A2(n6538), .B1(n12217), .B2(n8450), .ZN(n8024) );
  INV_X1 U10248 ( .A(n8024), .ZN(n8026) );
  NAND2_X1 U10249 ( .A1(n12098), .A2(n8266), .ZN(n7766) );
  NAND2_X1 U10250 ( .A1(n15353), .A2(n8277), .ZN(n7765) );
  NAND2_X1 U10251 ( .A1(n7766), .A2(n7765), .ZN(n7768) );
  XNOR2_X1 U10252 ( .A(n7768), .B(n10208), .ZN(n8023) );
  INV_X1 U10253 ( .A(n8023), .ZN(n8025) );
  NAND2_X1 U10254 ( .A1(n7827), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10255 ( .A1(n7825), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U10256 ( .A1(n7826), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10257 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7773) );
  XNOR2_X1 U10258 ( .A(n7773), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14825) );
  NAND2_X1 U10259 ( .A1(n7812), .A2(n14825), .ZN(n7778) );
  XNOR2_X1 U10260 ( .A(n7774), .B(SI_1_), .ZN(n7776) );
  MUX2_X1 U10261 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n10581), .Z(n7775) );
  XNOR2_X1 U10262 ( .A(n7776), .B(n7775), .ZN(n8523) );
  NAND2_X1 U10263 ( .A1(n15975), .A2(n8523), .ZN(n7777) );
  NAND3_X2 U10264 ( .A1(n7778), .A2(n7779), .A3(n7777), .ZN(n12497) );
  NAND2_X1 U10265 ( .A1(n12497), .A2(n8266), .ZN(n7780) );
  INV_X1 U10266 ( .A(n7931), .ZN(n7782) );
  NAND2_X1 U10267 ( .A1(n12497), .A2(n6551), .ZN(n7783) );
  NAND2_X1 U10268 ( .A1(n7873), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10269 ( .A1(n7826), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10270 ( .A1(n7825), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10271 ( .A1(n7827), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7785) );
  INV_X1 U10272 ( .A(SI_0_), .ZN(n7789) );
  INV_X1 U10273 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9058) );
  OAI21_X1 U10274 ( .B1(n10575), .B2(n7789), .A(n9058), .ZN(n7790) );
  AND2_X1 U10275 ( .A1(n7791), .A2(n7790), .ZN(n15435) );
  MUX2_X1 U10276 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15435), .S(n7832), .Z(n12490)
         );
  INV_X1 U10277 ( .A(n10565), .ZN(n7795) );
  AOI22_X1 U10278 ( .A1(n6551), .A2(n12490), .B1(n7795), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7792) );
  AND2_X1 U10279 ( .A1(n7793), .A2(n7792), .ZN(n10929) );
  AOI22_X1 U10280 ( .A1(n8266), .A2(n12490), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n7795), .ZN(n7796) );
  NAND2_X1 U10281 ( .A1(n7797), .A2(n7796), .ZN(n10928) );
  INV_X1 U10282 ( .A(n10928), .ZN(n7798) );
  NAND2_X1 U10283 ( .A1(n7798), .A2(n10208), .ZN(n7799) );
  NAND2_X1 U10284 ( .A1(n10927), .A2(n7799), .ZN(n11040) );
  NAND2_X1 U10285 ( .A1(n11041), .A2(n11040), .ZN(n7804) );
  INV_X1 U10286 ( .A(n7800), .ZN(n7802) );
  NAND2_X1 U10287 ( .A1(n7802), .A2(n7801), .ZN(n7803) );
  NAND2_X1 U10288 ( .A1(n7804), .A2(n7803), .ZN(n11029) );
  NAND2_X1 U10289 ( .A1(n7825), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10290 ( .A1(n7826), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10291 ( .A1(n7976), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U10292 ( .A1(n7827), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7805) );
  XNOR2_X1 U10293 ( .A(n7809), .B(n7810), .ZN(n10592) );
  NAND2_X1 U10294 ( .A1(n15975), .A2(n10592), .ZN(n7815) );
  NAND2_X1 U10295 ( .A1(n6604), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7814) );
  XNOR2_X1 U10296 ( .A(n7811), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U10297 ( .A1(n7812), .A2(n14844), .ZN(n7813) );
  OAI22_X1 U10298 ( .A1(n15486), .A2(n6537), .B1(n12508), .B2(n6541), .ZN(
        n7816) );
  XNOR2_X1 U10299 ( .A(n7816), .B(n8448), .ZN(n7821) );
  OR2_X1 U10300 ( .A1(n7931), .A2(n15486), .ZN(n7818) );
  NAND2_X1 U10301 ( .A1(n11489), .A2(n8277), .ZN(n7817) );
  NAND2_X1 U10302 ( .A1(n7818), .A2(n7817), .ZN(n7819) );
  XNOR2_X1 U10303 ( .A(n7821), .B(n7819), .ZN(n11030) );
  NAND2_X1 U10304 ( .A1(n11029), .A2(n11030), .ZN(n7823) );
  INV_X1 U10305 ( .A(n7819), .ZN(n7820) );
  NAND2_X1 U10306 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  INV_X1 U10307 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10308 ( .A1(n7825), .A2(n7824), .ZN(n7831) );
  NAND2_X1 U10309 ( .A1(n7826), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10310 ( .A1(n7873), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10311 ( .A1(n7827), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7828) );
  INV_X1 U10312 ( .A(n7833), .ZN(n7860) );
  NAND2_X1 U10313 ( .A1(n7860), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7835) );
  INV_X1 U10314 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U10315 ( .A(n7835), .B(n7834), .ZN(n14859) );
  NAND2_X1 U10316 ( .A1(n7837), .A2(n7836), .ZN(n7854) );
  XNOR2_X1 U10317 ( .A(n7838), .B(SI_3_), .ZN(n7852) );
  XNOR2_X1 U10318 ( .A(n7854), .B(n7852), .ZN(n10576) );
  NAND2_X1 U10319 ( .A1(n10576), .A2(n15975), .ZN(n7841) );
  NAND2_X1 U10320 ( .A1(n6604), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7840) );
  OAI211_X1 U10321 ( .C1(n10638), .C2(n14859), .A(n7841), .B(n7840), .ZN(
        n15557) );
  OAI22_X1 U10322 ( .A1(n15629), .A2(n6537), .B1(n10156), .B2(n6541), .ZN(
        n7842) );
  XNOR2_X1 U10323 ( .A(n7842), .B(n10208), .ZN(n7846) );
  OR2_X1 U10324 ( .A1(n7931), .A2(n15629), .ZN(n7844) );
  NAND2_X1 U10325 ( .A1(n8277), .A2(n15557), .ZN(n7843) );
  NAND2_X1 U10326 ( .A1(n7844), .A2(n7843), .ZN(n7845) );
  XNOR2_X1 U10327 ( .A(n7846), .B(n7845), .ZN(n15485) );
  NAND2_X1 U10328 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  OAI21_X1 U10329 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n7871), .ZN(n11430) );
  INV_X1 U10330 ( .A(n11430), .ZN(n11888) );
  NAND2_X1 U10331 ( .A1(n8396), .A2(n11888), .ZN(n7851) );
  NAND2_X1 U10332 ( .A1(n10216), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10333 ( .A1(n7976), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10334 ( .A1(n7827), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7848) );
  AND4_X2 U10335 ( .A1(n7851), .A2(n7850), .A3(n7849), .A4(n7848), .ZN(n15487)
         );
  OR2_X1 U10336 ( .A1(n8450), .A2(n15487), .ZN(n7867) );
  INV_X1 U10337 ( .A(n7852), .ZN(n7853) );
  NAND2_X1 U10338 ( .A1(n7854), .A2(n7853), .ZN(n7856) );
  NAND2_X1 U10339 ( .A1(n7856), .A2(n7855), .ZN(n7858) );
  XNOR2_X1 U10340 ( .A(n7858), .B(n7857), .ZN(n10594) );
  OAI21_X1 U10341 ( .B1(n7860), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7862) );
  INV_X1 U10342 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U10343 ( .A(n7862), .B(n7861), .ZN(n14873) );
  OAI22_X1 U10344 ( .A1(n8182), .A2(n10627), .B1(n10638), .B2(n14873), .ZN(
        n7863) );
  INV_X1 U10345 ( .A(n7863), .ZN(n7864) );
  NAND2_X1 U10346 ( .A1(n12520), .A2(n8277), .ZN(n7866) );
  OAI22_X1 U10347 ( .A1(n15487), .A2(n6537), .B1(n12519), .B2(n6541), .ZN(
        n7868) );
  XNOR2_X1 U10348 ( .A(n7868), .B(n10208), .ZN(n11424) );
  NAND2_X1 U10349 ( .A1(n11422), .A2(n11424), .ZN(n7869) );
  NAND2_X1 U10350 ( .A1(n10216), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7877) );
  INV_X1 U10351 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U10352 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  AND2_X1 U10353 ( .A1(n7921), .A2(n7872), .ZN(n15536) );
  NAND2_X1 U10354 ( .A1(n8396), .A2(n15536), .ZN(n7876) );
  NAND2_X1 U10355 ( .A1(n7873), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10356 ( .A1(n8442), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7874) );
  INV_X1 U10357 ( .A(n15666), .ZN(n11506) );
  OR2_X1 U10358 ( .A1(n11506), .A2(n8450), .ZN(n7887) );
  INV_X1 U10359 ( .A(n8094), .ZN(n7879) );
  NAND2_X1 U10360 ( .A1(n7879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7881) );
  MUX2_X1 U10361 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7881), .S(n7880), .Z(n7882)
         );
  NAND2_X1 U10362 ( .A1(n7882), .A2(n7914), .ZN(n14886) );
  OAI22_X1 U10363 ( .A1(n8182), .A2(n10625), .B1(n10638), .B2(n14886), .ZN(
        n7883) );
  INV_X1 U10364 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U10365 ( .A1(n7885), .A2(n7884), .ZN(n12526) );
  NAND2_X1 U10366 ( .A1(n12526), .A2(n8277), .ZN(n7886) );
  NAND2_X1 U10367 ( .A1(n7887), .A2(n7886), .ZN(n12333) );
  NAND2_X1 U10368 ( .A1(n15666), .A2(n8277), .ZN(n7889) );
  NAND2_X1 U10369 ( .A1(n8266), .A2(n12526), .ZN(n7888) );
  NAND2_X1 U10370 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  XNOR2_X1 U10371 ( .A(n7890), .B(n10208), .ZN(n12334) );
  NAND2_X1 U10372 ( .A1(n12336), .A2(n12333), .ZN(n7891) );
  NAND2_X1 U10373 ( .A1(n7892), .A2(n7891), .ZN(n11644) );
  XNOR2_X1 U10374 ( .A(n7893), .B(n7894), .ZN(n10589) );
  NAND2_X1 U10375 ( .A1(n7895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7897) );
  XNOR2_X1 U10376 ( .A(n7897), .B(n7896), .ZN(n14908) );
  OAI22_X1 U10377 ( .A1(n8182), .A2(n10623), .B1(n10638), .B2(n14908), .ZN(
        n7898) );
  INV_X1 U10378 ( .A(n7898), .ZN(n7899) );
  NAND2_X1 U10379 ( .A1(n7900), .A2(n7899), .ZN(n12538) );
  NAND2_X1 U10380 ( .A1(n12538), .A2(n8266), .ZN(n7908) );
  NAND2_X1 U10381 ( .A1(n10216), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10382 ( .A1(n7923), .A2(n7901), .ZN(n7902) );
  AND2_X1 U10383 ( .A1(n7951), .A2(n7902), .ZN(n15518) );
  NAND2_X1 U10384 ( .A1(n8396), .A2(n15518), .ZN(n7905) );
  NAND2_X1 U10385 ( .A1(n7976), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10386 ( .A1(n8442), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7903) );
  NAND4_X1 U10387 ( .A1(n7906), .A2(n7905), .A3(n7904), .A4(n7903), .ZN(n15667) );
  NAND2_X1 U10388 ( .A1(n15667), .A2(n8277), .ZN(n7907) );
  NAND2_X1 U10389 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  XNOR2_X1 U10390 ( .A(n7909), .B(n8448), .ZN(n11843) );
  NAND2_X1 U10391 ( .A1(n12538), .A2(n8277), .ZN(n7911) );
  OR2_X1 U10392 ( .A1(n11652), .A2(n8450), .ZN(n7910) );
  XNOR2_X1 U10393 ( .A(n7912), .B(n7913), .ZN(n10580) );
  NAND2_X1 U10394 ( .A1(n7914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7916) );
  XNOR2_X1 U10395 ( .A(n7915), .B(n7916), .ZN(n10847) );
  OAI22_X1 U10396 ( .A1(n8182), .A2(n10629), .B1(n10638), .B2(n10847), .ZN(
        n7917) );
  INV_X1 U10397 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10398 ( .A1(n12530), .A2(n8266), .ZN(n7929) );
  NAND2_X1 U10399 ( .A1(n10216), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7927) );
  INV_X1 U10400 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10401 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  AND2_X1 U10402 ( .A1(n7923), .A2(n7922), .ZN(n11505) );
  NAND2_X1 U10403 ( .A1(n8396), .A2(n11505), .ZN(n7926) );
  NAND2_X1 U10404 ( .A1(n7976), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10405 ( .A1(n8442), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7924) );
  NAND4_X2 U10406 ( .A1(n7927), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n15531) );
  NAND2_X1 U10407 ( .A1(n15531), .A2(n8277), .ZN(n7928) );
  NAND2_X1 U10408 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  XNOR2_X1 U10409 ( .A(n7930), .B(n8448), .ZN(n11645) );
  OR2_X1 U10410 ( .A1(n12338), .A2(n8450), .ZN(n7933) );
  NAND2_X1 U10411 ( .A1(n12530), .A2(n8277), .ZN(n7932) );
  AND2_X1 U10412 ( .A1(n7933), .A2(n7932), .ZN(n11646) );
  AOI22_X1 U10413 ( .A1(n11843), .A2(n11842), .B1(n11645), .B2(n11646), .ZN(
        n7934) );
  NAND2_X1 U10414 ( .A1(n11644), .A2(n7934), .ZN(n7941) );
  INV_X1 U10415 ( .A(n11843), .ZN(n7939) );
  INV_X1 U10416 ( .A(n11645), .ZN(n11839) );
  INV_X1 U10417 ( .A(n11646), .ZN(n11840) );
  NAND2_X1 U10418 ( .A1(n11839), .A2(n11840), .ZN(n7935) );
  NAND2_X1 U10419 ( .A1(n7935), .A2(n11842), .ZN(n7938) );
  INV_X1 U10420 ( .A(n11842), .ZN(n7936) );
  AND2_X1 U10421 ( .A1(n7936), .A2(n11840), .ZN(n7937) );
  AOI22_X1 U10422 ( .A1(n7939), .A2(n7938), .B1(n7937), .B2(n11839), .ZN(n7940) );
  XNOR2_X1 U10423 ( .A(n7943), .B(n7942), .ZN(n10618) );
  NAND2_X1 U10424 ( .A1(n7944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7946) );
  XNOR2_X1 U10425 ( .A(n7946), .B(n7945), .ZN(n10793) );
  OAI22_X1 U10426 ( .A1(n8182), .A2(n10619), .B1(n10638), .B2(n10793), .ZN(
        n7947) );
  INV_X1 U10427 ( .A(n7947), .ZN(n7948) );
  NAND2_X1 U10428 ( .A1(n12548), .A2(n8266), .ZN(n7959) );
  NAND2_X1 U10429 ( .A1(n10216), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10430 ( .A1(n7951), .A2(n7950), .ZN(n7952) );
  NAND2_X1 U10431 ( .A1(n7974), .A2(n7952), .ZN(n11614) );
  INV_X1 U10432 ( .A(n11614), .ZN(n7953) );
  NAND2_X1 U10433 ( .A1(n8396), .A2(n7953), .ZN(n7956) );
  NAND2_X1 U10434 ( .A1(n8121), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10435 ( .A1(n8442), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7954) );
  NAND4_X1 U10436 ( .A1(n7957), .A2(n7956), .A3(n7955), .A4(n7954), .ZN(n15514) );
  NAND2_X1 U10437 ( .A1(n15514), .A2(n8277), .ZN(n7958) );
  NAND2_X1 U10438 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  XNOR2_X1 U10439 ( .A(n7960), .B(n8448), .ZN(n7963) );
  INV_X1 U10440 ( .A(n15514), .ZN(n15385) );
  NOR2_X1 U10441 ( .A1(n8450), .A2(n15385), .ZN(n7961) );
  AOI21_X1 U10442 ( .B1(n12548), .B2(n8277), .A(n7961), .ZN(n7962) );
  XNOR2_X1 U10443 ( .A(n7963), .B(n7962), .ZN(n11596) );
  NAND2_X1 U10444 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  XNOR2_X1 U10445 ( .A(n7965), .B(n7966), .ZN(n10632) );
  NAND2_X1 U10446 ( .A1(n7967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7969) );
  OR2_X1 U10447 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U10448 ( .A1(n7969), .A2(n7968), .ZN(n7992) );
  AOI22_X1 U10449 ( .A1(n6604), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n14924), 
        .B2(n8064), .ZN(n7971) );
  NAND2_X1 U10450 ( .A1(n10216), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10451 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  AND2_X1 U10452 ( .A1(n7997), .A2(n7975), .ZN(n12133) );
  NAND2_X1 U10453 ( .A1(n8396), .A2(n12133), .ZN(n7979) );
  NAND2_X1 U10454 ( .A1(n8121), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U10455 ( .A1(n8442), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7977) );
  NAND4_X1 U10456 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n14821) );
  INV_X1 U10457 ( .A(n14821), .ZN(n15377) );
  NOR2_X1 U10458 ( .A1(n8450), .A2(n15377), .ZN(n7981) );
  AOI21_X1 U10459 ( .B1(n15389), .B2(n8277), .A(n7981), .ZN(n7986) );
  NAND2_X1 U10460 ( .A1(n15389), .A2(n8266), .ZN(n7983) );
  NAND2_X1 U10461 ( .A1(n14821), .A2(n8277), .ZN(n7982) );
  NAND2_X1 U10462 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U10463 ( .A(n7984), .B(n10208), .ZN(n12124) );
  NAND2_X2 U10464 ( .A1(n7987), .A2(n7585), .ZN(n12126) );
  INV_X1 U10465 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U10466 ( .A1(n7992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7993) );
  XNOR2_X1 U10467 ( .A(n7993), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U10468 ( .A1(n10854), .A2(n8064), .B1(n6604), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10469 ( .A1(n10216), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8002) );
  INV_X1 U10470 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10471 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  AND2_X1 U10472 ( .A1(n8012), .A2(n7998), .ZN(n12146) );
  NAND2_X1 U10473 ( .A1(n8396), .A2(n12146), .ZN(n8001) );
  NAND2_X1 U10474 ( .A1(n8121), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10475 ( .A1(n8442), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7999) );
  OAI22_X1 U10476 ( .A1(n15378), .A2(n6541), .B1(n15384), .B2(n6537), .ZN(
        n8003) );
  XNOR2_X1 U10477 ( .A(n8003), .B(n10208), .ZN(n8005) );
  OAI22_X1 U10478 ( .A1(n15378), .A2(n6537), .B1(n15384), .B2(n8450), .ZN(
        n8004) );
  AND2_X1 U10479 ( .A1(n8005), .A2(n8004), .ZN(n12065) );
  NAND2_X1 U10480 ( .A1(n10657), .A2(n6552), .ZN(n8011) );
  NAND2_X1 U10481 ( .A1(n8008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8009) );
  XNOR2_X1 U10482 ( .A(n8009), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U10483 ( .A1(n10818), .A2(n8064), .B1(n6604), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U10484 ( .A1(n10216), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10485 ( .A1(n8012), .A2(n10744), .ZN(n8013) );
  AND2_X1 U10486 ( .A1(n8040), .A2(n8013), .ZN(n12232) );
  NAND2_X1 U10487 ( .A1(n8396), .A2(n12232), .ZN(n8016) );
  NAND2_X1 U10488 ( .A1(n8145), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10489 ( .A1(n8442), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8014) );
  NAND4_X1 U10490 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n15362) );
  OAI22_X1 U10491 ( .A1(n12062), .A2(n6538), .B1(n12565), .B2(n8450), .ZN(
        n8019) );
  OAI22_X1 U10492 ( .A1(n12062), .A2(n6541), .B1(n12565), .B2(n6537), .ZN(
        n8018) );
  XNOR2_X1 U10493 ( .A(n8018), .B(n10208), .ZN(n8020) );
  XOR2_X1 U10494 ( .A(n8019), .B(n8020), .Z(n12229) );
  INV_X1 U10495 ( .A(n8019), .ZN(n8022) );
  INV_X1 U10496 ( .A(n8020), .ZN(n8021) );
  XOR2_X1 U10497 ( .A(n8024), .B(n8023), .Z(n12289) );
  MUX2_X1 U10498 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10575), .Z(n8051) );
  XNOR2_X1 U10499 ( .A(n8082), .B(n8076), .ZN(n10923) );
  NAND2_X1 U10500 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U10501 ( .A1(n8031), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10502 ( .A1(n8033), .A2(n8032), .ZN(n8062) );
  OR2_X1 U10503 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  AOI22_X1 U10504 ( .A1(n10981), .A2(n8064), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n6604), .ZN(n8035) );
  NAND2_X1 U10505 ( .A1(n10216), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8045) );
  AND2_X1 U10506 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8037) );
  INV_X1 U10507 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10824) );
  INV_X1 U10508 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8039) );
  OAI21_X1 U10509 ( .B1(n8040), .B2(n10824), .A(n8039), .ZN(n8041) );
  AND2_X1 U10510 ( .A1(n8067), .A2(n8041), .ZN(n14768) );
  NAND2_X1 U10511 ( .A1(n8396), .A2(n14768), .ZN(n8044) );
  NAND2_X1 U10512 ( .A1(n8121), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10513 ( .A1(n8442), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8042) );
  AOI22_X1 U10514 ( .A1(n15352), .A2(n8266), .B1(n8277), .B2(n15363), .ZN(
        n8046) );
  XNOR2_X1 U10515 ( .A(n8046), .B(n10208), .ZN(n8048) );
  AOI22_X1 U10516 ( .A1(n15352), .A2(n8277), .B1(n8404), .B2(n15363), .ZN(
        n8047) );
  XNOR2_X1 U10517 ( .A(n8048), .B(n8047), .ZN(n14763) );
  NAND2_X1 U10518 ( .A1(n8051), .A2(SI_13_), .ZN(n8079) );
  NAND2_X1 U10519 ( .A1(n8079), .A2(SI_14_), .ZN(n8059) );
  INV_X1 U10520 ( .A(n8051), .ZN(n8052) );
  AOI21_X1 U10521 ( .B1(n8052), .B2(n10815), .A(SI_14_), .ZN(n8049) );
  NAND3_X1 U10522 ( .A1(n8060), .A2(n8049), .A3(n8050), .ZN(n8058) );
  INV_X1 U10523 ( .A(n8059), .ZN(n8056) );
  INV_X1 U10524 ( .A(n8050), .ZN(n8055) );
  OAI21_X1 U10525 ( .B1(SI_14_), .B2(n10815), .A(n8051), .ZN(n8054) );
  INV_X1 U10526 ( .A(SI_14_), .ZN(n10921) );
  OAI21_X1 U10527 ( .B1(SI_13_), .B2(n10921), .A(n8052), .ZN(n8053) );
  AOI22_X1 U10528 ( .A1(n8056), .A2(n8055), .B1(n8054), .B2(n8053), .ZN(n8057)
         );
  OAI211_X1 U10529 ( .C1(n8060), .C2(n8059), .A(n8058), .B(n8057), .ZN(n8061)
         );
  MUX2_X1 U10530 ( .A(n10937), .B(n10939), .S(n10581), .Z(n8083) );
  XNOR2_X1 U10531 ( .A(n8061), .B(n8083), .ZN(n10935) );
  NAND2_X1 U10532 ( .A1(n10935), .A2(n6552), .ZN(n8066) );
  NAND2_X1 U10533 ( .A1(n8062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8063) );
  XNOR2_X1 U10534 ( .A(n8063), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U10535 ( .A1(n11630), .A2(n8064), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n6604), .ZN(n8065) );
  NAND2_X1 U10536 ( .A1(n10216), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8072) );
  INV_X1 U10537 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10974) );
  OR2_X2 U10538 ( .A1(n8067), .A2(n10974), .ZN(n8118) );
  NAND2_X1 U10539 ( .A1(n8067), .A2(n10974), .ZN(n8068) );
  AND2_X1 U10540 ( .A1(n8118), .A2(n8068), .ZN(n15193) );
  NAND2_X1 U10541 ( .A1(n8396), .A2(n15193), .ZN(n8071) );
  NAND2_X1 U10542 ( .A1(n8121), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10543 ( .A1(n8442), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8069) );
  OAI22_X1 U10544 ( .A1(n15346), .A2(n6541), .B1(n14766), .B2(n6537), .ZN(
        n8073) );
  XNOR2_X1 U10545 ( .A(n8073), .B(n10208), .ZN(n8075) );
  OAI22_X1 U10546 ( .A1(n15346), .A2(n6537), .B1(n14766), .B2(n8450), .ZN(
        n8074) );
  XNOR2_X1 U10547 ( .A(n8075), .B(n8074), .ZN(n14669) );
  INV_X1 U10548 ( .A(n8083), .ZN(n8077) );
  NAND2_X1 U10549 ( .A1(n8083), .A2(n10921), .ZN(n8084) );
  MUX2_X1 U10550 ( .A(n11038), .B(n11037), .S(n10575), .Z(n8086) );
  INV_X1 U10551 ( .A(SI_15_), .ZN(n10813) );
  INV_X1 U10552 ( .A(n8086), .ZN(n8087) );
  NAND2_X1 U10553 ( .A1(n8087), .A2(SI_15_), .ZN(n8088) );
  MUX2_X1 U10554 ( .A(n11178), .B(n11177), .S(n10575), .Z(n8090) );
  INV_X1 U10555 ( .A(SI_16_), .ZN(n10967) );
  NAND2_X1 U10556 ( .A1(n8090), .A2(n10967), .ZN(n8138) );
  INV_X1 U10557 ( .A(n8090), .ZN(n8091) );
  NAND2_X1 U10558 ( .A1(n8091), .A2(SI_16_), .ZN(n8092) );
  NAND2_X1 U10559 ( .A1(n8094), .A2(n8093), .ZN(n8110) );
  OR2_X1 U10560 ( .A1(n8110), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10561 ( .A1(n8112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8095) );
  MUX2_X1 U10562 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8095), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8098) );
  INV_X1 U10563 ( .A(n8112), .ZN(n8097) );
  NAND2_X1 U10564 ( .A1(n8097), .A2(n8096), .ZN(n8139) );
  NAND2_X1 U10565 ( .A1(n8098), .A2(n8139), .ZN(n11627) );
  OAI22_X1 U10566 ( .A1(n8182), .A2(n11178), .B1(n10638), .B2(n11627), .ZN(
        n8099) );
  INV_X1 U10567 ( .A(n8099), .ZN(n8100) );
  AND2_X2 U10568 ( .A1(n8101), .A2(n8100), .ZN(n15332) );
  INV_X1 U10569 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8117) );
  OR2_X2 U10570 ( .A1(n8118), .A2(n8117), .ZN(n8120) );
  INV_X1 U10571 ( .A(n8120), .ZN(n8102) );
  INV_X1 U10572 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10573 ( .A1(n8120), .A2(n8103), .ZN(n8104) );
  NAND2_X1 U10574 ( .A1(n8168), .A2(n8104), .ZN(n15176) );
  OR2_X1 U10575 ( .A1(n15176), .A2(n8464), .ZN(n8107) );
  AOI22_X1 U10576 ( .A1(n10216), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n7976), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10577 ( .A1(n8442), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8105) );
  OAI22_X1 U10578 ( .A1(n15332), .A2(n6541), .B1(n15321), .B2(n6538), .ZN(
        n8108) );
  XNOR2_X1 U10579 ( .A(n8108), .B(n10208), .ZN(n14723) );
  OAI22_X1 U10580 ( .A1(n15332), .A2(n6537), .B1(n15321), .B2(n8450), .ZN(
        n8132) );
  NAND2_X1 U10581 ( .A1(n14723), .A2(n8132), .ZN(n8131) );
  XNOR2_X1 U10582 ( .A(n8109), .B(n7648), .ZN(n11036) );
  NAND2_X1 U10583 ( .A1(n8110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8111) );
  MUX2_X1 U10584 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8111), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n8113) );
  NAND2_X1 U10585 ( .A1(n8113), .A2(n8112), .ZN(n11621) );
  OAI22_X1 U10586 ( .A1(n8182), .A2(n11038), .B1(n10638), .B2(n11621), .ZN(
        n8114) );
  INV_X1 U10587 ( .A(n8114), .ZN(n8115) );
  NAND2_X1 U10588 ( .A1(n12585), .A2(n8266), .ZN(n8127) );
  NAND2_X1 U10589 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  AND2_X1 U10590 ( .A1(n8120), .A2(n8119), .ZN(n14812) );
  NAND2_X1 U10591 ( .A1(n14812), .A2(n8396), .ZN(n8125) );
  NAND2_X1 U10592 ( .A1(n8121), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10593 ( .A1(n10216), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10594 ( .A1(n8442), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8122) );
  NAND4_X1 U10595 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n15344) );
  NAND2_X1 U10596 ( .A1(n15344), .A2(n8277), .ZN(n8126) );
  NAND2_X1 U10597 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  XNOR2_X1 U10598 ( .A(n8128), .B(n8448), .ZN(n14721) );
  INV_X1 U10599 ( .A(n15344), .ZN(n15197) );
  NOR2_X1 U10600 ( .A1(n8450), .A2(n15197), .ZN(n8129) );
  AOI21_X1 U10601 ( .B1(n12585), .B2(n8277), .A(n8129), .ZN(n14719) );
  OR2_X1 U10602 ( .A1(n14721), .A2(n14719), .ZN(n8130) );
  INV_X1 U10603 ( .A(n8132), .ZN(n14722) );
  AOI21_X1 U10604 ( .B1(n14721), .B2(n14719), .A(n14722), .ZN(n8133) );
  NAND3_X1 U10605 ( .A1(n14722), .A2(n14719), .A3(n14721), .ZN(n8134) );
  NAND2_X1 U10606 ( .A1(n8136), .A2(n7635), .ZN(n14732) );
  MUX2_X1 U10607 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10575), .Z(n8157) );
  INV_X1 U10608 ( .A(SI_17_), .ZN(n11009) );
  INV_X1 U10609 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U10610 ( .A1(n8139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8141) );
  XNOR2_X1 U10611 ( .A(n8141), .B(n8140), .ZN(n14939) );
  OAI22_X1 U10612 ( .A1(n8182), .A2(n11199), .B1(n14939), .B2(n10638), .ZN(
        n8142) );
  INV_X1 U10613 ( .A(n8142), .ZN(n8143) );
  XNOR2_X1 U10614 ( .A(n8168), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n15159) );
  NAND2_X1 U10615 ( .A1(n15159), .A2(n8396), .ZN(n8150) );
  INV_X1 U10616 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U10617 ( .A1(n10216), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U10618 ( .A1(n8145), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U10619 ( .C1(n12104), .C2(n12429), .A(n8147), .B(n8146), .ZN(n8148) );
  INV_X1 U10620 ( .A(n8148), .ZN(n8149) );
  NAND2_X1 U10621 ( .A1(n8150), .A2(n8149), .ZN(n15329) );
  OAI22_X1 U10622 ( .A1(n12592), .A2(n6541), .B1(n15181), .B2(n6537), .ZN(
        n8151) );
  XOR2_X1 U10623 ( .A(n10208), .B(n8151), .Z(n14734) );
  AOI22_X1 U10624 ( .A1(n15325), .A2(n8277), .B1(n8404), .B2(n15329), .ZN(
        n14733) );
  INV_X1 U10625 ( .A(n14734), .ZN(n8154) );
  INV_X1 U10626 ( .A(n14733), .ZN(n8153) );
  NAND2_X1 U10627 ( .A1(n8157), .A2(SI_17_), .ZN(n8175) );
  NAND2_X1 U10628 ( .A1(n8178), .A2(n8175), .ZN(n8159) );
  MUX2_X1 U10629 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10575), .Z(n8174) );
  XNOR2_X1 U10630 ( .A(n8174), .B(SI_18_), .ZN(n8158) );
  NAND2_X1 U10631 ( .A1(n11402), .A2(n6552), .ZN(n8165) );
  INV_X1 U10632 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11403) );
  NAND2_X1 U10633 ( .A1(n8160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8162) );
  XNOR2_X1 U10634 ( .A(n8162), .B(n8161), .ZN(n12113) );
  OAI22_X1 U10635 ( .A1(n8182), .A2(n11403), .B1(n10638), .B2(n12113), .ZN(
        n8163) );
  INV_X1 U10636 ( .A(n8163), .ZN(n8164) );
  INV_X1 U10637 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n14736) );
  INV_X1 U10638 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8166) );
  OAI21_X1 U10639 ( .B1(n8168), .B2(n14736), .A(n8166), .ZN(n8169) );
  NAND2_X1 U10640 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n8167) );
  AND2_X1 U10641 ( .A1(n8169), .A2(n8187), .ZN(n15144) );
  NAND2_X1 U10642 ( .A1(n15144), .A2(n8396), .ZN(n8172) );
  AOI22_X1 U10643 ( .A1(n10216), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8145), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10644 ( .A1(n8442), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8170) );
  OAI22_X1 U10645 ( .A1(n15315), .A2(n6538), .B1(n15322), .B2(n8450), .ZN(
        n8198) );
  OAI22_X1 U10646 ( .A1(n15315), .A2(n6541), .B1(n15322), .B2(n6537), .ZN(
        n8173) );
  XNOR2_X1 U10647 ( .A(n8173), .B(n10208), .ZN(n8197) );
  XOR2_X1 U10648 ( .A(n8198), .B(n8197), .Z(n14786) );
  INV_X1 U10649 ( .A(SI_18_), .ZN(n11196) );
  OAI21_X1 U10650 ( .B1(n8179), .B2(n11196), .A(n8175), .ZN(n8176) );
  INV_X1 U10651 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U10652 ( .A1(n8179), .A2(n11196), .ZN(n8207) );
  NAND2_X1 U10653 ( .A1(n8209), .A2(n8207), .ZN(n8181) );
  INV_X1 U10654 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11538) );
  MUX2_X1 U10655 ( .A(n11481), .B(n11538), .S(n10575), .Z(n8206) );
  XNOR2_X1 U10656 ( .A(n8206), .B(SI_19_), .ZN(n8180) );
  OAI22_X1 U10657 ( .A1(n8182), .A2(n11481), .B1(n15207), .B2(n10638), .ZN(
        n8183) );
  INV_X1 U10658 ( .A(n8183), .ZN(n8184) );
  INV_X1 U10659 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10660 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  NAND2_X1 U10661 ( .A1(n8214), .A2(n8188), .ZN(n15125) );
  OR2_X1 U10662 ( .A1(n15125), .A2(n8464), .ZN(n8194) );
  INV_X1 U10663 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10664 ( .A1(n8145), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10665 ( .A1(n8442), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8189) );
  OAI211_X1 U10666 ( .C1(n8219), .C2(n8191), .A(n8190), .B(n8189), .ZN(n8192)
         );
  INV_X1 U10667 ( .A(n8192), .ZN(n8193) );
  OAI22_X1 U10668 ( .A1(n15309), .A2(n6541), .B1(n15314), .B2(n6538), .ZN(
        n8195) );
  XNOR2_X1 U10669 ( .A(n8195), .B(n10208), .ZN(n8202) );
  NOR2_X1 U10670 ( .A1(n15314), .A2(n8450), .ZN(n8196) );
  AOI21_X1 U10671 ( .B1(n15131), .B2(n8277), .A(n8196), .ZN(n8203) );
  XNOR2_X1 U10672 ( .A(n8202), .B(n8203), .ZN(n14695) );
  INV_X1 U10673 ( .A(n8197), .ZN(n8200) );
  INV_X1 U10674 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10675 ( .A1(n8200), .A2(n8199), .ZN(n14693) );
  INV_X1 U10676 ( .A(n8203), .ZN(n8204) );
  OAI21_X1 U10677 ( .B1(n8210), .B2(SI_19_), .A(n8207), .ZN(n8208) );
  NAND2_X1 U10678 ( .A1(n8210), .A2(SI_19_), .ZN(n8211) );
  MUX2_X1 U10679 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10575), .Z(n8253) );
  NAND2_X1 U10680 ( .A1(n6604), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8212) );
  INV_X1 U10681 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14755) );
  NAND2_X1 U10682 ( .A1(n8214), .A2(n14755), .ZN(n8215) );
  NAND2_X1 U10683 ( .A1(n8238), .A2(n8215), .ZN(n15104) );
  INV_X1 U10684 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U10685 ( .A1(n8442), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10686 ( .A1(n8145), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8217) );
  OAI211_X1 U10687 ( .C1(n8219), .C2(n10475), .A(n8218), .B(n8217), .ZN(n8220)
         );
  INV_X1 U10688 ( .A(n8220), .ZN(n8221) );
  AND2_X1 U10689 ( .A1(n15306), .A2(n8404), .ZN(n8223) );
  AOI21_X1 U10690 ( .B1(n10129), .B2(n8277), .A(n8223), .ZN(n8226) );
  AOI22_X1 U10691 ( .A1(n10129), .A2(n8266), .B1(n8277), .B2(n15306), .ZN(
        n8224) );
  XNOR2_X1 U10692 ( .A(n8224), .B(n10208), .ZN(n8225) );
  XOR2_X1 U10693 ( .A(n8226), .B(n8225), .Z(n14753) );
  INV_X1 U10694 ( .A(n8225), .ZN(n8228) );
  INV_X1 U10695 ( .A(n8226), .ZN(n8227) );
  NAND2_X1 U10696 ( .A1(n8230), .A2(n8253), .ZN(n8233) );
  NAND2_X1 U10697 ( .A1(n8231), .A2(SI_20_), .ZN(n8232) );
  MUX2_X1 U10698 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10575), .Z(n8255) );
  XNOR2_X1 U10699 ( .A(n8255), .B(SI_21_), .ZN(n8234) );
  NAND2_X1 U10700 ( .A1(n6604), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10701 ( .A1(n15091), .A2(n8266), .ZN(n8246) );
  INV_X1 U10702 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U10703 ( .A1(n8238), .A2(n14703), .ZN(n8239) );
  NAND2_X1 U10704 ( .A1(n8286), .A2(n8239), .ZN(n15085) );
  INV_X1 U10705 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U10706 ( .A1(n10216), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10707 ( .A1(n8145), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8240) );
  OAI211_X1 U10708 ( .C1(n8242), .C2(n12429), .A(n8241), .B(n8240), .ZN(n8243)
         );
  INV_X1 U10709 ( .A(n8243), .ZN(n8244) );
  NAND2_X1 U10710 ( .A1(n14818), .A2(n8277), .ZN(n8245) );
  NAND2_X1 U10711 ( .A1(n8246), .A2(n8245), .ZN(n8247) );
  NAND2_X1 U10712 ( .A1(n15091), .A2(n8277), .ZN(n8249) );
  NAND2_X1 U10713 ( .A1(n14818), .A2(n8404), .ZN(n8248) );
  NAND2_X1 U10714 ( .A1(n8249), .A2(n8248), .ZN(n8299) );
  NAND2_X1 U10715 ( .A1(n14678), .A2(n8299), .ZN(n8298) );
  INV_X1 U10716 ( .A(n8255), .ZN(n8250) );
  INV_X1 U10717 ( .A(SI_21_), .ZN(n11536) );
  NAND2_X1 U10718 ( .A1(n8250), .A2(n11536), .ZN(n8256) );
  OAI21_X1 U10719 ( .B1(SI_20_), .B2(n8253), .A(n8256), .ZN(n8251) );
  INV_X1 U10720 ( .A(n8251), .ZN(n8252) );
  INV_X1 U10721 ( .A(n8253), .ZN(n8254) );
  INV_X1 U10722 ( .A(SI_20_), .ZN(n11484) );
  NOR2_X1 U10723 ( .A1(n8254), .A2(n11484), .ZN(n8257) );
  MUX2_X1 U10724 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10575), .Z(n8260) );
  NAND2_X1 U10725 ( .A1(n8260), .A2(SI_22_), .ZN(n8258) );
  INV_X1 U10726 ( .A(n8260), .ZN(n8804) );
  INV_X1 U10727 ( .A(SI_22_), .ZN(n8282) );
  NAND2_X1 U10728 ( .A1(n8804), .A2(n8282), .ZN(n8261) );
  MUX2_X1 U10729 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10575), .Z(n8312) );
  XNOR2_X1 U10730 ( .A(n8312), .B(SI_23_), .ZN(n8310) );
  INV_X1 U10731 ( .A(n8310), .ZN(n8263) );
  NAND2_X1 U10732 ( .A1(n11546), .A2(n6552), .ZN(n8265) );
  NAND2_X1 U10733 ( .A1(n6604), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8264) );
  NAND2_X2 U10734 ( .A1(n8265), .A2(n8264), .ZN(n15062) );
  NAND2_X1 U10735 ( .A1(n15062), .A2(n8266), .ZN(n8275) );
  INV_X1 U10736 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U10737 ( .A1(n8288), .A2(n14687), .ZN(n8268) );
  NAND2_X1 U10738 ( .A1(n8318), .A2(n8268), .ZN(n15058) );
  INV_X1 U10739 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U10740 ( .A1(n10216), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10741 ( .A1(n8145), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8269) );
  OAI211_X1 U10742 ( .C1(n15059), .C2(n12429), .A(n8270), .B(n8269), .ZN(n8271) );
  INV_X1 U10743 ( .A(n8271), .ZN(n8272) );
  NAND2_X1 U10744 ( .A1(n15045), .A2(n8277), .ZN(n8274) );
  NAND2_X1 U10745 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  XNOR2_X1 U10746 ( .A(n8276), .B(n10208), .ZN(n8302) );
  NAND2_X1 U10747 ( .A1(n15062), .A2(n8277), .ZN(n8279) );
  NAND2_X1 U10748 ( .A1(n15045), .A2(n8404), .ZN(n8278) );
  NAND2_X1 U10749 ( .A1(n8279), .A2(n8278), .ZN(n8303) );
  NAND2_X1 U10750 ( .A1(n8302), .A2(n8303), .ZN(n14683) );
  INV_X1 U10751 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10752 ( .A1(n8286), .A2(n8285), .ZN(n8287) );
  NAND2_X1 U10753 ( .A1(n8288), .A2(n8287), .ZN(n14778) );
  INV_X1 U10754 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U10755 ( .A1(n10216), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10756 ( .A1(n8145), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8289) );
  OAI211_X1 U10757 ( .C1(n12429), .C2(n8291), .A(n8290), .B(n8289), .ZN(n8292)
         );
  INV_X1 U10758 ( .A(n8292), .ZN(n8293) );
  OAI22_X1 U10759 ( .A1(n15076), .A2(n6541), .B1(n15089), .B2(n6537), .ZN(
        n8295) );
  XNOR2_X1 U10760 ( .A(n8295), .B(n10208), .ZN(n14680) );
  NAND2_X1 U10761 ( .A1(n15294), .A2(n8404), .ZN(n8296) );
  NAND2_X1 U10762 ( .A1(n8297), .A2(n8296), .ZN(n8300) );
  NAND2_X1 U10763 ( .A1(n14680), .A2(n8300), .ZN(n14685) );
  NAND4_X1 U10764 ( .A1(n14685), .A2(n14681), .A3(n14682), .A4(n14683), .ZN(
        n8308) );
  INV_X1 U10765 ( .A(n14680), .ZN(n8301) );
  INV_X1 U10766 ( .A(n8300), .ZN(n14679) );
  NAND3_X1 U10767 ( .A1(n8301), .A2(n14679), .A3(n14683), .ZN(n8306) );
  INV_X1 U10768 ( .A(n8302), .ZN(n8305) );
  INV_X1 U10769 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U10770 ( .A1(n8305), .A2(n8304), .ZN(n14742) );
  NAND2_X1 U10771 ( .A1(n8312), .A2(SI_23_), .ZN(n8334) );
  MUX2_X1 U10772 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10575), .Z(n8338) );
  XNOR2_X1 U10773 ( .A(n8338), .B(SI_24_), .ZN(n8313) );
  NAND2_X1 U10774 ( .A1(n11903), .A2(n6552), .ZN(n8316) );
  NAND2_X1 U10775 ( .A1(n6604), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8315) );
  INV_X1 U10776 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10777 ( .A1(n8318), .A2(n8317), .ZN(n8319) );
  NAND2_X1 U10778 ( .A1(n15044), .A2(n8396), .ZN(n8325) );
  INV_X1 U10779 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U10780 ( .A1(n10216), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10781 ( .A1(n8145), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8320) );
  OAI211_X1 U10782 ( .C1(n12429), .C2(n8322), .A(n8321), .B(n8320), .ZN(n8323)
         );
  INV_X1 U10783 ( .A(n8323), .ZN(n8324) );
  AND2_X2 U10784 ( .A1(n8325), .A2(n8324), .ZN(n14688) );
  OAI22_X1 U10785 ( .A1(n14752), .A2(n6541), .B1(n14688), .B2(n6538), .ZN(
        n8326) );
  XNOR2_X1 U10786 ( .A(n8326), .B(n8448), .ZN(n8329) );
  NAND2_X1 U10787 ( .A1(n15057), .A2(n8404), .ZN(n8327) );
  NAND2_X1 U10788 ( .A1(n8329), .A2(n8330), .ZN(n14709) );
  INV_X1 U10789 ( .A(n8329), .ZN(n8332) );
  INV_X1 U10790 ( .A(n8330), .ZN(n8331) );
  NAND2_X1 U10791 ( .A1(n8332), .A2(n8331), .ZN(n8333) );
  NAND2_X1 U10792 ( .A1(n14708), .A2(n14709), .ZN(n8364) );
  NAND2_X1 U10793 ( .A1(n8338), .A2(SI_24_), .ZN(n8335) );
  INV_X1 U10794 ( .A(n8338), .ZN(n8339) );
  INV_X1 U10795 ( .A(SI_24_), .ZN(n12273) );
  NAND2_X1 U10796 ( .A1(n8339), .A2(n12273), .ZN(n8340) );
  INV_X1 U10797 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9454) );
  INV_X1 U10798 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12121) );
  MUX2_X1 U10799 ( .A(n9454), .B(n12121), .S(n10575), .Z(n8342) );
  INV_X1 U10800 ( .A(SI_25_), .ZN(n12299) );
  NAND2_X1 U10801 ( .A1(n8342), .A2(n12299), .ZN(n8368) );
  INV_X1 U10802 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U10803 ( .A1(n8343), .A2(SI_25_), .ZN(n8344) );
  XNOR2_X1 U10804 ( .A(n8367), .B(n8366), .ZN(n12025) );
  NAND2_X1 U10805 ( .A1(n12025), .A2(n6552), .ZN(n8346) );
  NAND2_X1 U10806 ( .A1(n6604), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8345) );
  INV_X1 U10807 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10808 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  NAND2_X1 U10809 ( .A1(n8392), .A2(n8349), .ZN(n15029) );
  INV_X1 U10810 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10811 ( .A1(n10216), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8351) );
  NAND2_X1 U10812 ( .A1(n8145), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8350) );
  OAI211_X1 U10813 ( .C1(n8352), .C2(n12429), .A(n8351), .B(n8350), .ZN(n8353)
         );
  INV_X1 U10814 ( .A(n8353), .ZN(n8354) );
  AND2_X2 U10815 ( .A1(n8355), .A2(n8354), .ZN(n15274) );
  OAI22_X1 U10816 ( .A1(n15267), .A2(n6541), .B1(n15274), .B2(n6537), .ZN(
        n8356) );
  XNOR2_X1 U10817 ( .A(n8356), .B(n8448), .ZN(n8359) );
  NAND2_X1 U10818 ( .A1(n15015), .A2(n8404), .ZN(n8357) );
  NAND2_X1 U10819 ( .A1(n8359), .A2(n8360), .ZN(n8365) );
  INV_X1 U10820 ( .A(n8359), .ZN(n8362) );
  INV_X1 U10821 ( .A(n8360), .ZN(n8361) );
  NAND2_X1 U10822 ( .A1(n8362), .A2(n8361), .ZN(n8363) );
  NAND2_X1 U10823 ( .A1(n8364), .A2(n14710), .ZN(n14712) );
  NAND2_X1 U10824 ( .A1(n14712), .A2(n8365), .ZN(n14794) );
  MUX2_X1 U10825 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10575), .Z(n8384) );
  XNOR2_X1 U10826 ( .A(n8384), .B(SI_26_), .ZN(n8386) );
  INV_X1 U10827 ( .A(n8386), .ZN(n8370) );
  NAND2_X1 U10828 ( .A1(n12157), .A2(n6552), .ZN(n8372) );
  NAND2_X1 U10829 ( .A1(n6604), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10830 ( .A1(n15017), .A2(n8396), .ZN(n8378) );
  INV_X1 U10831 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10832 ( .A1(n10216), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U10833 ( .A1(n8145), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8373) );
  OAI211_X1 U10834 ( .C1(n8375), .C2(n12429), .A(n8374), .B(n8373), .ZN(n8376)
         );
  INV_X1 U10835 ( .A(n8376), .ZN(n8377) );
  OAI22_X1 U10836 ( .A1(n15261), .A2(n6541), .B1(n15251), .B2(n6538), .ZN(
        n8379) );
  XNOR2_X1 U10837 ( .A(n8379), .B(n10208), .ZN(n8381) );
  OAI22_X1 U10838 ( .A1(n15261), .A2(n6537), .B1(n15251), .B2(n8450), .ZN(
        n8380) );
  NOR2_X1 U10839 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  AOI21_X1 U10840 ( .B1(n8381), .B2(n8380), .A(n8382), .ZN(n14795) );
  NAND2_X1 U10841 ( .A1(n14794), .A2(n14795), .ZN(n14793) );
  INV_X1 U10842 ( .A(n8382), .ZN(n8383) );
  NAND2_X1 U10843 ( .A1(n14793), .A2(n8383), .ZN(n10256) );
  NAND2_X1 U10844 ( .A1(n8384), .A2(SI_26_), .ZN(n8385) );
  INV_X1 U10845 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12302) );
  INV_X1 U10846 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12401) );
  MUX2_X1 U10847 ( .A(n12302), .B(n12401), .S(n10581), .Z(n8435) );
  XNOR2_X1 U10848 ( .A(n8435), .B(SI_27_), .ZN(n8433) );
  INV_X1 U10849 ( .A(n8433), .ZN(n8388) );
  XNOR2_X1 U10850 ( .A(n8434), .B(n8388), .ZN(n12301) );
  NAND2_X1 U10851 ( .A1(n6604), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8389) );
  INV_X1 U10852 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14797) );
  INV_X1 U10853 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8391) );
  OAI21_X1 U10854 ( .B1(n8392), .B2(n14797), .A(n8391), .ZN(n8395) );
  AND2_X1 U10855 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n8393) );
  NAND2_X1 U10856 ( .A1(n14999), .A2(n8396), .ZN(n8401) );
  INV_X1 U10857 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U10858 ( .A1(n10216), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10859 ( .A1(n8145), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8397) );
  OAI211_X1 U10860 ( .C1(n10472), .C2(n12429), .A(n8398), .B(n8397), .ZN(n8399) );
  INV_X1 U10861 ( .A(n8399), .ZN(n8400) );
  AND2_X2 U10862 ( .A1(n8401), .A2(n8400), .ZN(n15242) );
  OAI22_X1 U10863 ( .A1(n15003), .A2(n6541), .B1(n15242), .B2(n6538), .ZN(
        n8402) );
  XNOR2_X1 U10864 ( .A(n8402), .B(n8448), .ZN(n8408) );
  INV_X1 U10865 ( .A(n8408), .ZN(n8410) );
  OR2_X1 U10866 ( .A1(n15003), .A2(n6538), .ZN(n8406) );
  NAND2_X1 U10867 ( .A1(n15016), .A2(n8404), .ZN(n8405) );
  INV_X1 U10868 ( .A(n8407), .ZN(n8409) );
  AOI21_X1 U10869 ( .B1(n8410), .B2(n8409), .A(n8456), .ZN(n10257) );
  NAND2_X1 U10870 ( .A1(n10256), .A2(n10257), .ZN(n10261) );
  INV_X1 U10871 ( .A(n10261), .ZN(n8453) );
  INV_X1 U10872 ( .A(P1_B_REG_SCAN_IN), .ZN(n10214) );
  OR2_X1 U10873 ( .A1(n12026), .A2(n10214), .ZN(n8411) );
  MUX2_X1 U10874 ( .A(n8411), .B(P1_B_REG_SCAN_IN), .S(n11904), .Z(n8412) );
  NAND2_X1 U10875 ( .A1(n8412), .A2(n10646), .ZN(n10644) );
  OAI22_X1 U10876 ( .A1(n10644), .A2(P1_D_REG_1__SCAN_IN), .B1(n12026), .B2(
        n10646), .ZN(n11005) );
  INV_X1 U10877 ( .A(n11005), .ZN(n10148) );
  INV_X1 U10878 ( .A(n10644), .ZN(n8415) );
  INV_X1 U10879 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8414) );
  NOR2_X1 U10880 ( .A1(n10646), .A2(n11904), .ZN(n8413) );
  AOI21_X1 U10881 ( .B1(n8415), .B2(n8414), .A(n8413), .ZN(n11006) );
  NOR4_X1 U10882 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n8423) );
  NOR4_X1 U10883 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n8422) );
  INV_X1 U10884 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15594) );
  INV_X1 U10885 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15602) );
  INV_X1 U10886 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15593) );
  INV_X1 U10887 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15595) );
  NAND4_X1 U10888 ( .A1(n15594), .A2(n15602), .A3(n15593), .A4(n15595), .ZN(
        n10294) );
  NOR4_X1 U10889 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8419) );
  NOR4_X1 U10890 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8418) );
  NOR4_X1 U10891 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n8417) );
  NOR4_X1 U10892 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8416) );
  NAND4_X1 U10893 ( .A1(n8419), .A2(n8418), .A3(n8417), .A4(n8416), .ZN(n8420)
         );
  NOR4_X1 U10894 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n10294), .A4(n8420), .ZN(n8421) );
  AND3_X1 U10895 ( .A1(n8423), .A2(n8422), .A3(n8421), .ZN(n8424) );
  NOR2_X1 U10896 ( .A1(n10644), .A2(n8424), .ZN(n10146) );
  INV_X1 U10897 ( .A(n10146), .ZN(n8425) );
  NAND3_X1 U10898 ( .A1(n10148), .A2(n11006), .A3(n8425), .ZN(n8462) );
  INV_X1 U10899 ( .A(n8462), .ZN(n8432) );
  OAI21_X1 U10900 ( .B1(n6660), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8426) );
  MUX2_X1 U10901 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8426), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8428) );
  NAND2_X1 U10902 ( .A1(n8428), .A2(n8427), .ZN(n10636) );
  AND2_X1 U10903 ( .A1(n10636), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10647) );
  NAND2_X1 U10904 ( .A1(n6608), .A2(n7760), .ZN(n12643) );
  NAND2_X1 U10905 ( .A1(n10645), .A2(n12643), .ZN(n8430) );
  NAND2_X1 U10906 ( .A1(n6755), .A2(n12645), .ZN(n15563) );
  NAND2_X1 U10907 ( .A1(n6755), .A2(n10213), .ZN(n8429) );
  NOR2_X1 U10908 ( .A1(n8430), .A2(n15388), .ZN(n8431) );
  INV_X1 U10909 ( .A(n8435), .ZN(n8436) );
  MUX2_X1 U10910 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10575), .Z(n9883) );
  NAND2_X1 U10911 ( .A1(n14664), .A2(n6552), .ZN(n8438) );
  NAND2_X1 U10912 ( .A1(n6604), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10913 ( .A1(n8439), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n10222) );
  INV_X1 U10914 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U10915 ( .A1(n8440), .A2(n10484), .ZN(n8441) );
  NAND2_X1 U10916 ( .A1(n10222), .A2(n8441), .ZN(n14986) );
  INV_X1 U10917 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U10918 ( .A1(n10216), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U10919 ( .A1(n8442), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8443) );
  OAI211_X1 U10920 ( .C1(n10331), .C2(n8216), .A(n8444), .B(n8443), .ZN(n8445)
         );
  INV_X1 U10921 ( .A(n8445), .ZN(n8446) );
  AND2_X2 U10922 ( .A1(n8447), .A2(n8446), .ZN(n15252) );
  OAI22_X1 U10923 ( .A1(n15224), .A2(n6541), .B1(n15252), .B2(n6538), .ZN(
        n8449) );
  XNOR2_X1 U10924 ( .A(n8449), .B(n8448), .ZN(n8452) );
  OAI22_X1 U10925 ( .A1(n15224), .A2(n6537), .B1(n15252), .B2(n8450), .ZN(
        n8451) );
  XNOR2_X1 U10926 ( .A(n8452), .B(n8451), .ZN(n8457) );
  INV_X1 U10927 ( .A(n8457), .ZN(n8455) );
  INV_X1 U10928 ( .A(n8456), .ZN(n8454) );
  NAND3_X1 U10929 ( .A1(n8457), .A2(n15491), .A3(n8456), .ZN(n8475) );
  NAND2_X1 U10930 ( .A1(n15540), .A2(n10213), .ZN(n11004) );
  NAND2_X1 U10931 ( .A1(n8462), .A2(n11004), .ZN(n10932) );
  NAND2_X1 U10932 ( .A1(n10932), .A2(n10645), .ZN(n11647) );
  INV_X1 U10933 ( .A(n14809), .ZN(n14769) );
  OAI21_X1 U10934 ( .B1(n12645), .B2(n10213), .A(n10637), .ZN(n8459) );
  AND2_X1 U10935 ( .A1(n10636), .A2(n10565), .ZN(n8458) );
  NAND2_X1 U10936 ( .A1(n10932), .A2(n12698), .ZN(n8460) );
  NAND2_X1 U10937 ( .A1(n8460), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15495) );
  OAI22_X1 U10938 ( .A1(n14986), .A2(n15495), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10484), .ZN(n8473) );
  NAND3_X1 U10939 ( .A1(n12698), .A2(n10637), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n8461) );
  NOR2_X2 U10940 ( .A1(n8471), .A2(n15430), .ZN(n14806) );
  OR2_X1 U10941 ( .A1(n10222), .A2(n8464), .ZN(n8470) );
  INV_X1 U10942 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10943 ( .A1(n10216), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10944 ( .A1(n8145), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8465) );
  OAI211_X1 U10945 ( .C1(n8467), .C2(n12429), .A(n8466), .B(n8465), .ZN(n8468)
         );
  INV_X1 U10946 ( .A(n8468), .ZN(n8469) );
  INV_X1 U10947 ( .A(n8471), .ZN(n15490) );
  NAND2_X1 U10948 ( .A1(n15490), .A2(n15430), .ZN(n14808) );
  OAI22_X1 U10949 ( .A1(n15242), .A2(n14798), .B1(n15241), .B2(n14808), .ZN(
        n8472) );
  AOI211_X1 U10950 ( .C1(n15244), .C2(n14769), .A(n8473), .B(n8472), .ZN(n8474) );
  NAND2_X1 U10951 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  AOI21_X1 U10952 ( .B1(n10261), .B2(n7641), .A(n8476), .ZN(n8477) );
  INV_X1 U10953 ( .A(n8887), .ZN(n8478) );
  INV_X1 U10954 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8488) );
  INV_X1 U10955 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10956 ( .A1(n8490), .A2(n8512), .ZN(n8974) );
  NAND2_X1 U10957 ( .A1(n8492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8494) );
  NAND2_X2 U10958 ( .A1(n8974), .A2(n12399), .ZN(n8542) );
  NAND2_X1 U10959 ( .A1(n8542), .A2(n10575), .ZN(n9939) );
  NAND2_X1 U10960 ( .A1(n12025), .A2(n9902), .ZN(n8496) );
  NAND2_X1 U10961 ( .A1(n8846), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8495) );
  INV_X1 U10962 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n14154) );
  INV_X1 U10963 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n13820) );
  INV_X1 U10964 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n14008) );
  INV_X1 U10965 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n14170) );
  INV_X1 U10966 ( .A(n8779), .ZN(n8503) );
  AND2_X1 U10967 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n8502) );
  INV_X1 U10968 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13949) );
  AND2_X1 U10969 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8504) );
  INV_X1 U10970 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13830) );
  OR2_X2 U10971 ( .A1(n8818), .A2(n13830), .ZN(n8830) );
  AND2_X1 U10972 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8506) );
  INV_X1 U10973 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13927) );
  INV_X1 U10974 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8508) );
  OAI21_X1 U10975 ( .B1(n8830), .B2(n13927), .A(n8508), .ZN(n8509) );
  NAND2_X1 U10976 ( .A1(n8838), .A2(n8509), .ZN(n14257) );
  INV_X1 U10977 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8510) );
  INV_X1 U10978 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14658) );
  XNOR2_X2 U10979 ( .A(n8511), .B(n14658), .ZN(n12703) );
  INV_X1 U10980 ( .A(n8849), .ZN(n8975) );
  BUF_X4 U10981 ( .A(n8557), .Z(n9945) );
  INV_X1 U10982 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8519) );
  CLKBUF_X3 U10983 ( .A(n8569), .Z(n9946) );
  NAND2_X1 U10984 ( .A1(n9946), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10985 ( .A1(n6597), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8517) );
  OAI211_X1 U10986 ( .C1(n8866), .C2(n8519), .A(n8518), .B(n8517), .ZN(n8520)
         );
  INV_X1 U10987 ( .A(n8520), .ZN(n8521) );
  INV_X1 U10988 ( .A(n8523), .ZN(n10615) );
  NAND2_X1 U10989 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8524) );
  MUX2_X1 U10990 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8524), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8525) );
  NAND2_X1 U10991 ( .A1(n8525), .A2(n6645), .ZN(n10867) );
  INV_X1 U10992 ( .A(n8530), .ZN(n8537) );
  NAND2_X1 U10993 ( .A1(n8569), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8532) );
  NAND4_X2 U10994 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n8543)
         );
  NAND2_X1 U10995 ( .A1(n8536), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10996 ( .A1(n8569), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10997 ( .A1(n8557), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10998 ( .A1(n8537), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8538) );
  XNOR2_X1 U10999 ( .A(n10572), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14668) );
  NAND2_X1 U11000 ( .A1(n9670), .A2(n11301), .ZN(n11333) );
  NAND2_X1 U11001 ( .A1(n11158), .A2(n8535), .ZN(n8544) );
  NAND2_X1 U11002 ( .A1(n8536), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U11003 ( .A1(n8569), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U11004 ( .A1(n8557), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U11005 ( .A1(n8594), .A2(n10592), .ZN(n8554) );
  NAND2_X1 U11006 ( .A1(n6645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8550) );
  INV_X1 U11007 ( .A(n14049), .ZN(n8551) );
  OR2_X1 U11008 ( .A1(n9940), .A2(n10593), .ZN(n8552) );
  XNOR2_X1 U11009 ( .A(n14041), .B(n15793), .ZN(n15762) );
  NAND2_X1 U11010 ( .A1(n15761), .A2(n15762), .ZN(n8556) );
  INV_X1 U11011 ( .A(n14041), .ZN(n10996) );
  NAND2_X1 U11012 ( .A1(n10996), .A2(n15793), .ZN(n8555) );
  NAND2_X1 U11013 ( .A1(n8556), .A2(n8555), .ZN(n11367) );
  NAND2_X1 U11014 ( .A1(n8569), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U11015 ( .A1(n6597), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U11016 ( .A1(n9945), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8559) );
  INV_X1 U11017 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U11018 ( .A1(n8849), .A2(n11371), .ZN(n8558) );
  NAND4_X1 U11019 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n14040) );
  NAND2_X1 U11020 ( .A1(n8594), .A2(n10576), .ZN(n8566) );
  INV_X1 U11021 ( .A(n8673), .ZN(n8563) );
  NAND2_X1 U11022 ( .A1(n8563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8562) );
  MUX2_X1 U11023 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8562), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8564) );
  AND2_X1 U11024 ( .A1(n8564), .A2(n8585), .ZN(n14058) );
  OR2_X1 U11025 ( .A1(n9940), .A2(n10585), .ZN(n8565) );
  NAND2_X1 U11026 ( .A1(n11367), .A2(n11368), .ZN(n8568) );
  INV_X1 U11027 ( .A(n14040), .ZN(n11327) );
  NAND2_X1 U11028 ( .A1(n11327), .A2(n15804), .ZN(n8567) );
  NAND2_X1 U11029 ( .A1(n8568), .A2(n8567), .ZN(n11318) );
  NAND2_X1 U11030 ( .A1(n8569), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11031 ( .A1(n6598), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8572) );
  OAI21_X1 U11032 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8579), .ZN(n11319) );
  INV_X1 U11033 ( .A(n11319), .ZN(n11238) );
  NAND2_X1 U11034 ( .A1(n8849), .A2(n11238), .ZN(n8571) );
  NAND2_X1 U11035 ( .A1(n9945), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8570) );
  NAND4_X1 U11036 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n14039) );
  NAND2_X1 U11037 ( .A1(n8585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U11038 ( .A(n8574), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U11039 ( .A1(n8846), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10798), 
        .B2(n14072), .ZN(n8576) );
  NAND2_X1 U11040 ( .A1(n10594), .A2(n8594), .ZN(n8575) );
  XNOR2_X1 U11041 ( .A(n14039), .B(n15811), .ZN(n8928) );
  INV_X1 U11042 ( .A(n14039), .ZN(n8929) );
  NAND2_X1 U11043 ( .A1(n8929), .A2(n15811), .ZN(n8577) );
  NAND2_X1 U11044 ( .A1(n9946), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11045 ( .A1(n6598), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8583) );
  INV_X1 U11046 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11047 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  AND2_X1 U11048 ( .A1(n8611), .A2(n8580), .ZN(n11391) );
  NAND2_X1 U11049 ( .A1(n8849), .A2(n11391), .ZN(n8582) );
  NAND2_X1 U11050 ( .A1(n9945), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8581) );
  NAND4_X1 U11051 ( .A1(n8584), .A2(n8583), .A3(n8582), .A4(n8581), .ZN(n14038) );
  INV_X1 U11052 ( .A(n8585), .ZN(n8587) );
  NAND2_X1 U11053 ( .A1(n8587), .A2(n8586), .ZN(n8589) );
  NAND2_X1 U11054 ( .A1(n8589), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8588) );
  MUX2_X1 U11055 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8588), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8590) );
  AND2_X1 U11056 ( .A1(n8590), .A2(n8603), .ZN(n14087) );
  AOI22_X1 U11057 ( .A1(n8846), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10798), 
        .B2(n14087), .ZN(n8592) );
  NAND2_X1 U11058 ( .A1(n10586), .A2(n9902), .ZN(n8591) );
  XNOR2_X1 U11059 ( .A(n14038), .B(n11520), .ZN(n11513) );
  INV_X1 U11060 ( .A(n14038), .ZN(n11436) );
  NAND2_X1 U11061 ( .A1(n11436), .A2(n11520), .ZN(n8593) );
  NAND2_X1 U11062 ( .A1(n10580), .A2(n8594), .ZN(n8597) );
  NAND2_X1 U11063 ( .A1(n8603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8595) );
  XNOR2_X1 U11064 ( .A(n8595), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14102) );
  AOI22_X1 U11065 ( .A1(n8846), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10798), 
        .B2(n14102), .ZN(n8596) );
  NAND2_X1 U11066 ( .A1(n6597), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U11067 ( .A1(n9946), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8600) );
  XNOR2_X1 U11068 ( .A(n8611), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U11069 ( .A1(n8849), .A2(n11559), .ZN(n8599) );
  NAND2_X1 U11070 ( .A1(n9945), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8598) );
  NAND4_X1 U11071 ( .A1(n8601), .A2(n8600), .A3(n8599), .A4(n8598), .ZN(n14037) );
  XNOR2_X1 U11072 ( .A(n11561), .B(n14037), .ZN(n11552) );
  INV_X1 U11073 ( .A(n14037), .ZN(n11734) );
  NAND2_X1 U11074 ( .A1(n11734), .A2(n11561), .ZN(n8602) );
  NAND2_X1 U11075 ( .A1(n10589), .A2(n9902), .ZN(n8608) );
  INV_X1 U11076 ( .A(n8603), .ZN(n8605) );
  INV_X1 U11077 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11078 ( .A1(n8605), .A2(n8604), .ZN(n8617) );
  NAND2_X1 U11079 ( .A1(n8617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U11080 ( .A(n8606), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U11081 ( .A1(n8846), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10798), 
        .B2(n14115), .ZN(n8607) );
  NAND2_X1 U11082 ( .A1(n6598), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U11083 ( .A1(n9946), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8615) );
  INV_X1 U11084 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8610) );
  INV_X1 U11085 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8609) );
  OAI21_X1 U11086 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8612) );
  AND2_X1 U11087 ( .A1(n8624), .A2(n8612), .ZN(n11529) );
  NAND2_X1 U11088 ( .A1(n8849), .A2(n11529), .ZN(n8614) );
  NAND2_X1 U11089 ( .A1(n9945), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8613) );
  OR2_X1 U11090 ( .A1(n15834), .A2(n11873), .ZN(n8936) );
  NAND2_X1 U11091 ( .A1(n15834), .A2(n11873), .ZN(n8935) );
  NAND2_X1 U11092 ( .A1(n8936), .A2(n8935), .ZN(n11733) );
  INV_X1 U11093 ( .A(n11873), .ZN(n14036) );
  NAND2_X1 U11094 ( .A1(n10618), .A2(n8594), .ZN(n8622) );
  NAND2_X1 U11095 ( .A1(n8619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8618) );
  MUX2_X1 U11096 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8618), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8620) );
  INV_X1 U11097 ( .A(n14129), .ZN(n10882) );
  AOI22_X1 U11098 ( .A1(n8846), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10882), 
        .B2(n10798), .ZN(n8621) );
  NAND2_X1 U11099 ( .A1(n6597), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11100 ( .A1(n9946), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8628) );
  INV_X1 U11101 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11102 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  AND2_X1 U11103 ( .A1(n8640), .A2(n8625), .ZN(n11590) );
  NAND2_X1 U11104 ( .A1(n8849), .A2(n11590), .ZN(n8627) );
  NAND2_X1 U11105 ( .A1(n9945), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8626) );
  NAND4_X1 U11106 ( .A1(n8629), .A2(n8628), .A3(n8627), .A4(n8626), .ZN(n14035) );
  XNOR2_X1 U11107 ( .A(n6607), .B(n14035), .ZN(n9982) );
  NAND2_X1 U11108 ( .A1(n6607), .A2(n14035), .ZN(n8630) );
  OAI21_X1 U11109 ( .B1(n11581), .B2(n9982), .A(n8630), .ZN(n11980) );
  NAND2_X1 U11110 ( .A1(n10632), .A2(n9902), .ZN(n8638) );
  NAND2_X1 U11111 ( .A1(n8632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8631) );
  MUX2_X1 U11112 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8631), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8635) );
  INV_X1 U11113 ( .A(n8632), .ZN(n8634) );
  INV_X1 U11114 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U11115 ( .A1(n8634), .A2(n8633), .ZN(n8660) );
  INV_X1 U11116 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10633) );
  INV_X1 U11117 ( .A(n8636), .ZN(n8637) );
  NAND2_X1 U11118 ( .A1(n9946), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11119 ( .A1(n6597), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U11120 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  AND2_X1 U11121 ( .A1(n8651), .A2(n8641), .ZN(n13937) );
  NAND2_X1 U11122 ( .A1(n8849), .A2(n13937), .ZN(n8643) );
  NAND2_X1 U11123 ( .A1(n9945), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11124 ( .A(n14604), .B(n13839), .ZN(n11984) );
  INV_X1 U11125 ( .A(n13839), .ZN(n14034) );
  NAND2_X1 U11126 ( .A1(n14604), .A2(n14034), .ZN(n8646) );
  NAND2_X1 U11127 ( .A1(n10653), .A2(n9902), .ZN(n8649) );
  NAND2_X1 U11128 ( .A1(n8660), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8647) );
  XNOR2_X1 U11129 ( .A(n8647), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U11130 ( .A1(n10908), .A2(n10798), .B1(n8846), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U11131 ( .A1(n6597), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11132 ( .A1(n9946), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8655) );
  INV_X1 U11133 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11134 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  AND2_X1 U11135 ( .A1(n8664), .A2(n8652), .ZN(n12008) );
  NAND2_X1 U11136 ( .A1(n8849), .A2(n12008), .ZN(n8654) );
  NAND2_X1 U11137 ( .A1(n9945), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11138 ( .A1(n13842), .A2(n13977), .ZN(n14467) );
  OR2_X1 U11139 ( .A1(n13842), .A2(n13977), .ZN(n8657) );
  INV_X1 U11140 ( .A(n12014), .ZN(n8658) );
  INV_X1 U11141 ( .A(n13977), .ZN(n14497) );
  OR2_X1 U11142 ( .A1(n13842), .A2(n14497), .ZN(n8659) );
  NAND2_X1 U11143 ( .A1(n12005), .A2(n8659), .ZN(n14504) );
  NAND2_X1 U11144 ( .A1(n10657), .A2(n9902), .ZN(n8663) );
  OAI21_X1 U11145 ( .B1(n8660), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8661) );
  AOI22_X1 U11146 ( .A1(n11352), .A2(n10798), .B1(n8846), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11147 ( .A1(n6598), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11148 ( .A1(n9946), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8668) );
  NAND2_X1 U11149 ( .A1(n8664), .A2(n10890), .ZN(n8665) );
  AND2_X1 U11150 ( .A1(n8678), .A2(n8665), .ZN(n14501) );
  NAND2_X1 U11151 ( .A1(n8849), .A2(n14501), .ZN(n8667) );
  NAND2_X1 U11152 ( .A1(n9945), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8666) );
  NAND4_X1 U11153 ( .A1(n8669), .A2(n8668), .A3(n8667), .A4(n8666), .ZN(n14033) );
  XNOR2_X1 U11154 ( .A(n14598), .B(n14033), .ZN(n14503) );
  NAND2_X1 U11155 ( .A1(n14598), .A2(n14033), .ZN(n8672) );
  NAND2_X1 U11156 ( .A1(n10683), .A2(n9902), .ZN(n8950) );
  OR2_X1 U11157 ( .A1(n9940), .A2(n10751), .ZN(n8676) );
  NAND2_X1 U11158 ( .A1(n8684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8674) );
  XNOR2_X1 U11159 ( .A(n8674), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15746) );
  NAND2_X1 U11160 ( .A1(n10798), .A2(n15746), .ZN(n8675) );
  NAND2_X1 U11161 ( .A1(n6597), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U11162 ( .A1(n9946), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8682) );
  INV_X1 U11163 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11164 ( .A1(n8678), .A2(n8677), .ZN(n8679) );
  AND2_X1 U11165 ( .A1(n8726), .A2(n8679), .ZN(n14483) );
  NAND2_X1 U11166 ( .A1(n8849), .A2(n14483), .ZN(n8681) );
  NAND2_X1 U11167 ( .A1(n9945), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8680) );
  XNOR2_X1 U11168 ( .A(n14593), .B(n13958), .ZN(n14475) );
  INV_X1 U11169 ( .A(n8684), .ZN(n8686) );
  INV_X1 U11170 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8687) );
  INV_X1 U11171 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8688) );
  INV_X1 U11172 ( .A(n8749), .ZN(n8689) );
  NAND2_X1 U11173 ( .A1(n8689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8690) );
  XNOR2_X1 U11174 ( .A(n8690), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U11175 ( .A1(n8846), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6606), 
        .B2(n14173), .ZN(n8691) );
  INV_X1 U11176 ( .A(n6598), .ZN(n8853) );
  INV_X1 U11177 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11968) );
  INV_X1 U11178 ( .A(n8693), .ZN(n8705) );
  INV_X1 U11179 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U11180 ( .A1(n8705), .A2(n13909), .ZN(n8694) );
  NAND2_X1 U11181 ( .A1(n8753), .A2(n8694), .ZN(n14407) );
  OR2_X1 U11182 ( .A1(n14407), .A2(n8975), .ZN(n8698) );
  NAND2_X1 U11183 ( .A1(n9946), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11184 ( .A1(n9945), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8695) );
  AND2_X1 U11185 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  OAI211_X1 U11186 ( .C1(n8853), .C2(n11968), .A(n8698), .B(n8697), .ZN(n14029) );
  NAND2_X1 U11187 ( .A1(n11036), .A2(n9902), .ZN(n8703) );
  INV_X1 U11188 ( .A(n8699), .ZN(n8700) );
  NAND2_X1 U11189 ( .A1(n8700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U11190 ( .A(n8701), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U11191 ( .A1(n8846), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10798), 
        .B2(n11964), .ZN(n8702) );
  NAND2_X1 U11192 ( .A1(n8715), .A2(n14008), .ZN(n8704) );
  AND2_X1 U11193 ( .A1(n8705), .A2(n8704), .ZN(n14423) );
  NAND2_X1 U11194 ( .A1(n14423), .A2(n8849), .ZN(n8709) );
  NAND2_X1 U11195 ( .A1(n6598), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11196 ( .A1(n9946), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U11197 ( .A1(n9945), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8706) );
  NAND4_X1 U11198 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n14030) );
  OR2_X1 U11199 ( .A1(n14578), .A2(n14030), .ZN(n14403) );
  NAND2_X1 U11200 ( .A1(n10935), .A2(n9902), .ZN(n8713) );
  INV_X1 U11201 ( .A(n8873), .ZN(n8722) );
  NAND2_X1 U11202 ( .A1(n8722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8711) );
  XNOR2_X1 U11203 ( .A(n8711), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U11204 ( .A1(n8846), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10798), 
        .B2(n11568), .ZN(n8712) );
  NAND2_X1 U11205 ( .A1(n9946), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11206 ( .A1(n6597), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11207 ( .A1(n8728), .A2(n13820), .ZN(n8714) );
  AND2_X1 U11208 ( .A1(n8715), .A2(n8714), .ZN(n14442) );
  NAND2_X1 U11209 ( .A1(n8849), .A2(n14442), .ZN(n8717) );
  NAND2_X1 U11210 ( .A1(n9945), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8716) );
  NAND4_X1 U11211 ( .A1(n8719), .A2(n8718), .A3(n8717), .A4(n8716), .ZN(n14031) );
  OR2_X1 U11212 ( .A1(n14583), .A2(n14031), .ZN(n8733) );
  NAND2_X1 U11213 ( .A1(n10923), .A2(n9902), .ZN(n8725) );
  NAND2_X1 U11214 ( .A1(n8720), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8721) );
  MUX2_X1 U11215 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8721), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8723) );
  NAND2_X1 U11216 ( .A1(n8723), .A2(n8722), .ZN(n14155) );
  INV_X1 U11217 ( .A(n14155), .ZN(n11357) );
  AOI22_X1 U11218 ( .A1(n8846), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10798), 
        .B2(n11357), .ZN(n8724) );
  NAND2_X1 U11219 ( .A1(n9946), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11220 ( .A1(n6597), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11221 ( .A1(n8726), .A2(n14154), .ZN(n8727) );
  AND2_X1 U11222 ( .A1(n8728), .A2(n8727), .ZN(n14453) );
  NAND2_X1 U11223 ( .A1(n8849), .A2(n14453), .ZN(n8730) );
  NAND2_X1 U11224 ( .A1(n9945), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8729) );
  NAND4_X1 U11225 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n14032) );
  OR2_X1 U11226 ( .A1(n14589), .A2(n14032), .ZN(n14435) );
  NAND2_X1 U11227 ( .A1(n8733), .A2(n14435), .ZN(n14400) );
  NOR2_X1 U11228 ( .A1(n8735), .A2(n14400), .ZN(n8734) );
  INV_X1 U11229 ( .A(n8735), .ZN(n8745) );
  NAND2_X1 U11230 ( .A1(n14589), .A2(n14032), .ZN(n8736) );
  INV_X1 U11231 ( .A(n14031), .ZN(n9783) );
  NAND2_X1 U11232 ( .A1(n8736), .A2(n9783), .ZN(n8737) );
  NAND2_X1 U11233 ( .A1(n8737), .A2(n14583), .ZN(n8739) );
  NAND3_X1 U11234 ( .A1(n14589), .A2(n14031), .A3(n14032), .ZN(n8738) );
  NAND2_X1 U11235 ( .A1(n8739), .A2(n8738), .ZN(n14401) );
  NAND2_X1 U11236 ( .A1(n14578), .A2(n14030), .ZN(n8740) );
  INV_X1 U11237 ( .A(n14029), .ZN(n9799) );
  NAND2_X1 U11238 ( .A1(n8740), .A2(n9799), .ZN(n8741) );
  NAND2_X1 U11239 ( .A1(n14573), .A2(n8741), .ZN(n8743) );
  NAND3_X1 U11240 ( .A1(n14578), .A2(n14029), .A3(n14030), .ZN(n8742) );
  NAND2_X1 U11241 ( .A1(n8743), .A2(n8742), .ZN(n8744) );
  AOI21_X1 U11242 ( .B1(n8745), .B2(n14401), .A(n8744), .ZN(n8746) );
  NAND2_X1 U11243 ( .A1(n11198), .A2(n9902), .ZN(n8752) );
  INV_X1 U11244 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11245 ( .A1(n8757), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11246 ( .A(n8750), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U11247 ( .A1(n14186), .A2(n10798), .B1(n8846), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11248 ( .A1(n8753), .A2(n14170), .ZN(n8754) );
  NAND2_X1 U11249 ( .A1(n8779), .A2(n8754), .ZN(n14390) );
  AOI22_X1 U11250 ( .A1(n6597), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9946), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11251 ( .A1(n9945), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8755) );
  OAI211_X1 U11252 ( .C1(n14390), .C2(n8975), .A(n8756), .B(n8755), .ZN(n14028) );
  AND2_X1 U11253 ( .A1(n14568), .A2(n14028), .ZN(n14374) );
  NAND2_X1 U11254 ( .A1(n11402), .A2(n9902), .ZN(n8762) );
  NAND2_X1 U11255 ( .A1(n8773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8760) );
  XNOR2_X1 U11256 ( .A(n8760), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U11257 ( .A1(n14189), .A2(n10798), .B1(n8846), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8761) );
  XNOR2_X1 U11258 ( .A(n8779), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U11259 ( .A1(n14369), .A2(n8849), .ZN(n8768) );
  INV_X1 U11260 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11261 ( .A1(n6598), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11262 ( .A1(n9946), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8763) );
  OAI211_X1 U11263 ( .C1(n8765), .C2(n8866), .A(n8764), .B(n8763), .ZN(n8766)
         );
  INV_X1 U11264 ( .A(n8766), .ZN(n8767) );
  NAND2_X1 U11265 ( .A1(n8768), .A2(n8767), .ZN(n14027) );
  AND2_X1 U11266 ( .A1(n14562), .A2(n14027), .ZN(n8769) );
  INV_X1 U11267 ( .A(n14562), .ZN(n14371) );
  OAI21_X1 U11268 ( .B1(n14568), .B2(n14028), .A(n14027), .ZN(n8771) );
  INV_X1 U11269 ( .A(n14568), .ZN(n13924) );
  NOR2_X1 U11270 ( .A1(n14027), .A2(n14028), .ZN(n8770) );
  AOI22_X1 U11271 ( .A1(n14371), .A2(n8771), .B1(n13924), .B2(n8770), .ZN(
        n8772) );
  NAND2_X1 U11272 ( .A1(n11480), .A2(n9902), .ZN(n8777) );
  INV_X1 U11273 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8774) );
  AOI22_X1 U11274 ( .A1(n14214), .A2(n6606), .B1(n8846), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8776) );
  INV_X1 U11275 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13988) );
  INV_X1 U11276 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8778) );
  OAI21_X1 U11277 ( .B1(n8779), .B2(n13988), .A(n8778), .ZN(n8780) );
  NAND2_X1 U11278 ( .A1(n8788), .A2(n8780), .ZN(n14358) );
  OR2_X1 U11279 ( .A1(n14358), .A2(n8975), .ZN(n8785) );
  INV_X1 U11280 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U11281 ( .A1(n9945), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U11282 ( .A1(n9946), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8781) );
  OAI211_X1 U11283 ( .C1(n8853), .C2(n14204), .A(n8782), .B(n8781), .ZN(n8783)
         );
  INV_X1 U11284 ( .A(n8783), .ZN(n8784) );
  INV_X1 U11285 ( .A(n14337), .ZN(n14026) );
  NAND2_X1 U11286 ( .A1(n14557), .A2(n14026), .ZN(n8786) );
  NAND2_X1 U11287 ( .A1(n8846), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11288 ( .A1(n8788), .A2(n13949), .ZN(n8789) );
  AND2_X1 U11289 ( .A1(n8809), .A2(n8789), .ZN(n14339) );
  NAND2_X1 U11290 ( .A1(n14339), .A2(n8849), .ZN(n8795) );
  INV_X1 U11291 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U11292 ( .A1(n6598), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U11293 ( .A1(n9946), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8790) );
  OAI211_X1 U11294 ( .C1(n8792), .C2(n8866), .A(n8791), .B(n8790), .ZN(n8793)
         );
  INV_X1 U11295 ( .A(n8793), .ZN(n8794) );
  INV_X1 U11296 ( .A(n14349), .ZN(n14025) );
  NAND2_X1 U11297 ( .A1(n14553), .A2(n14025), .ZN(n8796) );
  NAND2_X1 U11298 ( .A1(n8846), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8797) );
  XNOR2_X1 U11299 ( .A(n8809), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n14323) );
  NAND2_X1 U11300 ( .A1(n14323), .A2(n8849), .ZN(n8803) );
  INV_X1 U11301 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U11302 ( .A1(n9945), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U11303 ( .A1(n9946), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8799) );
  OAI211_X1 U11304 ( .C1(n8853), .C2(n14549), .A(n8800), .B(n8799), .ZN(n8801)
         );
  INV_X1 U11305 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U11306 ( .A1(n8803), .A2(n8802), .ZN(n14024) );
  XNOR2_X1 U11307 ( .A(n14548), .B(n14024), .ZN(n14316) );
  XNOR2_X1 U11308 ( .A(n8805), .B(n8804), .ZN(n11771) );
  NAND2_X1 U11309 ( .A1(n11771), .A2(n9902), .ZN(n8807) );
  NAND2_X1 U11310 ( .A1(n8846), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8806) );
  INV_X1 U11311 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13875) );
  INV_X1 U11312 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8808) );
  OAI21_X1 U11313 ( .B1(n8809), .B2(n13875), .A(n8808), .ZN(n8810) );
  NAND2_X1 U11314 ( .A1(n8810), .A2(n8818), .ZN(n14307) );
  OR2_X1 U11315 ( .A1(n14307), .A2(n8975), .ZN(n8815) );
  INV_X1 U11316 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U11317 ( .A1(n9945), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8812) );
  NAND2_X1 U11318 ( .A1(n9946), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8811) );
  OAI211_X1 U11319 ( .C1(n8853), .C2(n14544), .A(n8812), .B(n8811), .ZN(n8813)
         );
  INV_X1 U11320 ( .A(n8813), .ZN(n8814) );
  INV_X1 U11321 ( .A(n14287), .ZN(n14023) );
  NAND2_X1 U11322 ( .A1(n11546), .A2(n8594), .ZN(n8817) );
  NAND2_X1 U11323 ( .A1(n8846), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U11324 ( .A1(n8818), .A2(n13830), .ZN(n8819) );
  AND2_X1 U11325 ( .A1(n8830), .A2(n8819), .ZN(n14291) );
  NAND2_X1 U11326 ( .A1(n14291), .A2(n8849), .ZN(n8825) );
  INV_X1 U11327 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11328 ( .A1(n9946), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11329 ( .A1(n6598), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8820) );
  OAI211_X1 U11330 ( .C1(n8822), .C2(n8866), .A(n8821), .B(n8820), .ZN(n8823)
         );
  INV_X1 U11331 ( .A(n8823), .ZN(n8824) );
  NAND2_X1 U11332 ( .A1(n14538), .A2(n14268), .ZN(n8967) );
  INV_X1 U11333 ( .A(n14268), .ZN(n14022) );
  INV_X1 U11334 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11979) );
  OR2_X1 U11335 ( .A1(n9940), .A2(n11979), .ZN(n8828) );
  XNOR2_X1 U11336 ( .A(n8830), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n14269) );
  NAND2_X1 U11337 ( .A1(n14269), .A2(n8849), .ZN(n8835) );
  INV_X1 U11338 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U11339 ( .A1(n9946), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11340 ( .A1(n6597), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8831) );
  OAI211_X1 U11341 ( .C1(n8866), .C2(n14271), .A(n8832), .B(n8831), .ZN(n8833)
         );
  INV_X1 U11342 ( .A(n8833), .ZN(n8834) );
  NAND2_X2 U11343 ( .A1(n8835), .A2(n8834), .ZN(n14021) );
  NAND2_X1 U11344 ( .A1(n8846), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8836) );
  INV_X1 U11345 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10380) );
  NAND2_X1 U11346 ( .A1(n8838), .A2(n10380), .ZN(n8839) );
  INV_X1 U11347 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11348 ( .A1(n6598), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11349 ( .A1(n9946), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8840) );
  OAI211_X1 U11350 ( .C1(n8842), .C2(n8866), .A(n8841), .B(n8840), .ZN(n8843)
         );
  AOI21_X1 U11351 ( .B1(n14238), .B2(n8849), .A(n8843), .ZN(n13801) );
  NAND2_X1 U11352 ( .A1(n8844), .A2(n13801), .ZN(n8845) );
  NAND2_X1 U11353 ( .A1(n8846), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8847) );
  XNOR2_X1 U11354 ( .A(n8860), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U11355 ( .A1(n14224), .A2(n8849), .ZN(n8856) );
  INV_X1 U11356 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8852) );
  NAND2_X1 U11357 ( .A1(n9945), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11358 ( .A1(n9946), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8850) );
  OAI211_X1 U11359 ( .C1(n8853), .C2(n8852), .A(n8851), .B(n8850), .ZN(n8854)
         );
  INV_X1 U11360 ( .A(n8854), .ZN(n8855) );
  INV_X1 U11361 ( .A(n14018), .ZN(n8857) );
  INV_X1 U11362 ( .A(n10519), .ZN(n10522) );
  NAND2_X1 U11363 ( .A1(n14222), .A2(n10522), .ZN(n8871) );
  INV_X1 U11364 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9508) );
  OR2_X1 U11365 ( .A1(n9940), .A2(n9508), .ZN(n8858) );
  INV_X1 U11366 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13805) );
  INV_X1 U11367 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13866) );
  OAI21_X1 U11368 ( .B1(n8860), .B2(n13805), .A(n13866), .ZN(n8863) );
  INV_X1 U11369 ( .A(n8860), .ZN(n8862) );
  AND2_X1 U11370 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8861) );
  NAND2_X1 U11371 ( .A1(n8862), .A2(n8861), .ZN(n10542) );
  NAND2_X1 U11372 ( .A1(n8863), .A2(n10542), .ZN(n14213) );
  OR2_X1 U11373 ( .A1(n14213), .A2(n8975), .ZN(n8870) );
  INV_X1 U11374 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U11375 ( .A1(n6598), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U11376 ( .A1(n9946), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8864) );
  OAI211_X1 U11377 ( .C1(n8867), .C2(n8866), .A(n8865), .B(n8864), .ZN(n8868)
         );
  INV_X1 U11378 ( .A(n8868), .ZN(n8869) );
  NAND2_X1 U11379 ( .A1(n14218), .A2(n14017), .ZN(n10521) );
  INV_X1 U11380 ( .A(n14221), .ZN(n8921) );
  NOR2_X1 U11381 ( .A1(n8887), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11382 ( .A1(n8875), .A2(n8874), .ZN(n8879) );
  NAND2_X1 U11383 ( .A1(n8881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8876) );
  MUX2_X1 U11384 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8876), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8878) );
  NAND2_X1 U11385 ( .A1(n8878), .A2(n8877), .ZN(n12123) );
  INV_X1 U11386 ( .A(n12123), .ZN(n8885) );
  NAND2_X1 U11387 ( .A1(n8879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8880) );
  MUX2_X1 U11388 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8880), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8882) );
  NAND2_X1 U11389 ( .A1(n8882), .A2(n8881), .ZN(n11976) );
  NAND2_X1 U11390 ( .A1(n8877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11391 ( .A(n8883), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8914) );
  INV_X1 U11392 ( .A(n8914), .ZN(n12159) );
  NOR2_X1 U11393 ( .A1(n11976), .A2(n12159), .ZN(n8884) );
  NAND2_X1 U11394 ( .A1(n8885), .A2(n8884), .ZN(n10563) );
  NAND2_X1 U11395 ( .A1(n8887), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11396 ( .A1(n8911), .A2(n8888), .ZN(n8889) );
  XNOR2_X1 U11397 ( .A(n8889), .B(P2_IR_REG_23__SCAN_IN), .ZN(n10799) );
  XNOR2_X1 U11398 ( .A(n11976), .B(P2_B_REG_SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11399 ( .A1(n8890), .A2(n12123), .ZN(n8891) );
  INV_X1 U11400 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15784) );
  NAND2_X1 U11401 ( .A1(n15771), .A2(n15784), .ZN(n8893) );
  NAND2_X1 U11402 ( .A1(n12123), .A2(n12159), .ZN(n8892) );
  NAND2_X1 U11403 ( .A1(n8893), .A2(n8892), .ZN(n10941) );
  AND2_X1 U11404 ( .A1(n15781), .A2(n10941), .ZN(n15782) );
  NOR2_X1 U11405 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8897) );
  NOR4_X1 U11406 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8896) );
  NOR4_X1 U11407 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8895) );
  NOR4_X1 U11408 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8894) );
  AND4_X1 U11409 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n8903)
         );
  NOR4_X1 U11410 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8901) );
  NOR4_X1 U11411 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8900) );
  NOR4_X1 U11412 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8899) );
  NOR4_X1 U11413 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8898) );
  AND4_X1 U11414 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n8902)
         );
  NAND2_X1 U11415 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  NAND2_X1 U11416 ( .A1(n15771), .A2(n8904), .ZN(n10940) );
  NAND2_X1 U11417 ( .A1(n8905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11418 ( .A1(n6547), .A2(n11605), .ZN(n9996) );
  NAND2_X1 U11419 ( .A1(n8911), .A2(n8908), .ZN(n8909) );
  NAND2_X1 U11420 ( .A1(n9996), .A2(n10954), .ZN(n10947) );
  NAND2_X1 U11421 ( .A1(n10940), .A2(n10947), .ZN(n10532) );
  INV_X1 U11422 ( .A(n10005), .ZN(n11880) );
  NOR2_X1 U11423 ( .A1(n10532), .A2(n10945), .ZN(n8912) );
  INV_X1 U11424 ( .A(n11976), .ZN(n8915) );
  INV_X1 U11425 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15779) );
  NAND2_X1 U11426 ( .A1(n15771), .A2(n15779), .ZN(n8913) );
  OAI21_X1 U11427 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n15780) );
  INV_X1 U11428 ( .A(n15780), .ZN(n10943) );
  NAND2_X1 U11429 ( .A1(n14214), .A2(n11772), .ZN(n9943) );
  OR2_X1 U11430 ( .A1(n9943), .A2(n6553), .ZN(n15808) );
  INV_X1 U11431 ( .A(n10991), .ZN(n9671) );
  NAND2_X1 U11432 ( .A1(n15808), .A2(n8920), .ZN(n15797) );
  NAND2_X1 U11433 ( .A1(n15864), .A2(n15797), .ZN(n14586) );
  NAND2_X1 U11434 ( .A1(n8921), .A2(n14590), .ZN(n8999) );
  NOR2_X1 U11435 ( .A1(n9670), .A2(n11335), .ZN(n11338) );
  NAND2_X1 U11436 ( .A1(n11338), .A2(n11334), .ZN(n11340) );
  NAND2_X1 U11437 ( .A1(n11340), .A2(n8922), .ZN(n15754) );
  NAND2_X1 U11438 ( .A1(n14041), .A2(n15793), .ZN(n8923) );
  NAND2_X1 U11439 ( .A1(n15754), .A2(n8923), .ZN(n8925) );
  NAND2_X1 U11440 ( .A1(n10996), .A2(n15764), .ZN(n8924) );
  NAND2_X1 U11441 ( .A1(n8925), .A2(n8924), .ZN(n11375) );
  INV_X1 U11442 ( .A(n11368), .ZN(n11376) );
  NAND2_X1 U11443 ( .A1(n11375), .A2(n11376), .ZN(n8927) );
  NAND2_X1 U11444 ( .A1(n11327), .A2(n11370), .ZN(n8926) );
  NAND2_X1 U11445 ( .A1(n8927), .A2(n8926), .ZN(n11325) );
  NAND2_X1 U11446 ( .A1(n11325), .A2(n11326), .ZN(n8931) );
  NAND2_X1 U11447 ( .A1(n8929), .A2(n11324), .ZN(n8930) );
  NOR2_X1 U11448 ( .A1(n14038), .A2(n11520), .ZN(n8932) );
  NAND2_X1 U11449 ( .A1(n14038), .A2(n11520), .ZN(n11550) );
  OAI211_X1 U11450 ( .C1(n11734), .C2(n15827), .A(n8936), .B(n11550), .ZN(
        n8933) );
  INV_X1 U11451 ( .A(n8933), .ZN(n8934) );
  NAND2_X1 U11452 ( .A1(n11551), .A2(n8934), .ZN(n8939) );
  NAND2_X1 U11453 ( .A1(n11734), .A2(n15827), .ZN(n11728) );
  NAND2_X1 U11454 ( .A1(n8935), .A2(n11728), .ZN(n8937) );
  NAND2_X1 U11455 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  INV_X1 U11456 ( .A(n9982), .ZN(n11582) );
  INV_X1 U11457 ( .A(n14035), .ZN(n13939) );
  OR2_X1 U11458 ( .A1(n6607), .A2(n13939), .ZN(n8940) );
  NAND2_X1 U11459 ( .A1(n14604), .A2(n13839), .ZN(n12012) );
  NAND2_X1 U11460 ( .A1(n11983), .A2(n12012), .ZN(n8942) );
  NAND2_X1 U11461 ( .A1(n8942), .A2(n7627), .ZN(n8946) );
  NAND3_X1 U11462 ( .A1(n8950), .A2(n8949), .A3(n14467), .ZN(n8944) );
  NAND2_X1 U11463 ( .A1(n14467), .A2(n14495), .ZN(n8943) );
  NAND2_X1 U11464 ( .A1(n8944), .A2(n8943), .ZN(n8945) );
  INV_X1 U11465 ( .A(n14033), .ZN(n14472) );
  NAND2_X1 U11466 ( .A1(n14598), .A2(n14472), .ZN(n14469) );
  NAND2_X1 U11467 ( .A1(n8946), .A2(n6687), .ZN(n8954) );
  NAND3_X1 U11468 ( .A1(n8950), .A2(n8949), .A3(n14033), .ZN(n8948) );
  NAND2_X1 U11469 ( .A1(n14495), .A2(n14033), .ZN(n8947) );
  NAND2_X1 U11470 ( .A1(n8948), .A2(n8947), .ZN(n8952) );
  INV_X1 U11471 ( .A(n14598), .ZN(n14505) );
  AND2_X1 U11472 ( .A1(n14495), .A2(n8949), .ZN(n8951) );
  AOI22_X1 U11473 ( .A1(n8952), .A2(n14505), .B1(n8951), .B2(n8950), .ZN(n8953) );
  NAND2_X1 U11474 ( .A1(n8954), .A2(n8953), .ZN(n14458) );
  INV_X1 U11475 ( .A(n14032), .ZN(n14474) );
  NOR2_X1 U11476 ( .A1(n14589), .A2(n14474), .ZN(n8956) );
  NAND2_X1 U11477 ( .A1(n14589), .A2(n14474), .ZN(n8955) );
  XNOR2_X1 U11478 ( .A(n14583), .B(n9783), .ZN(n14438) );
  OAI22_X1 U11479 ( .A1(n14437), .A2(n14438), .B1(n9783), .B2(n14583), .ZN(
        n14427) );
  INV_X1 U11480 ( .A(n14030), .ZN(n9791) );
  XNOR2_X1 U11481 ( .A(n14578), .B(n9791), .ZN(n14430) );
  NAND2_X1 U11482 ( .A1(n14578), .A2(n9791), .ZN(n8957) );
  OR2_X1 U11483 ( .A1(n14573), .A2(n9799), .ZN(n14382) );
  XNOR2_X1 U11484 ( .A(n14568), .B(n14028), .ZN(n14373) );
  INV_X1 U11485 ( .A(n14028), .ZN(n13987) );
  OR2_X1 U11486 ( .A1(n14568), .A2(n13987), .ZN(n8959) );
  INV_X1 U11487 ( .A(n14027), .ZN(n14348) );
  NAND2_X1 U11488 ( .A1(n14562), .A2(n14348), .ZN(n8960) );
  OR2_X1 U11489 ( .A1(n14562), .A2(n14348), .ZN(n14345) );
  OR2_X1 U11490 ( .A1(n14557), .A2(n14337), .ZN(n8961) );
  AND2_X1 U11491 ( .A1(n14345), .A2(n8961), .ZN(n8962) );
  NAND2_X1 U11492 ( .A1(n14553), .A2(n14349), .ZN(n8963) );
  INV_X1 U11493 ( .A(n14024), .ZN(n14336) );
  OR2_X1 U11494 ( .A1(n14548), .A2(n14336), .ZN(n8964) );
  NAND2_X1 U11495 ( .A1(n14548), .A2(n14336), .ZN(n8965) );
  INV_X1 U11496 ( .A(n14021), .ZN(n14286) );
  NAND2_X1 U11497 ( .A1(n14532), .A2(n14286), .ZN(n8968) );
  INV_X1 U11498 ( .A(n14020), .ZN(n14267) );
  AND2_X1 U11499 ( .A1(n14527), .A2(n14267), .ZN(n8969) );
  NAND2_X1 U11500 ( .A1(n14214), .A2(n8917), .ZN(n8972) );
  NAND2_X1 U11501 ( .A1(n10005), .A2(n6553), .ZN(n8971) );
  INV_X1 U11502 ( .A(n10954), .ZN(n8982) );
  OR2_X1 U11503 ( .A1(n8982), .A2(n8974), .ZN(n14471) );
  NAND2_X1 U11504 ( .A1(n14018), .A2(n14496), .ZN(n8984) );
  OR2_X1 U11505 ( .A1(n10542), .A2(n8975), .ZN(n8980) );
  NAND2_X1 U11506 ( .A1(n6597), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11507 ( .A1(n9946), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11508 ( .A1(n9945), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8976) );
  AND3_X1 U11509 ( .A1(n8978), .A2(n8977), .A3(n8976), .ZN(n8979) );
  INV_X1 U11510 ( .A(n8974), .ZN(n8981) );
  OR2_X1 U11511 ( .A1(n11213), .A2(n14473), .ZN(n8983) );
  NAND2_X1 U11512 ( .A1(n8984), .A2(n8983), .ZN(n13870) );
  INV_X1 U11513 ( .A(n11520), .ZN(n15819) );
  INV_X1 U11514 ( .A(n15834), .ZN(n11741) );
  INV_X1 U11515 ( .A(n13842), .ZN(n12009) );
  INV_X1 U11516 ( .A(n14583), .ZN(n14445) );
  INV_X1 U11517 ( .A(n14578), .ZN(n14425) );
  INV_X1 U11518 ( .A(n14557), .ZN(n14361) );
  INV_X1 U11519 ( .A(n14543), .ZN(n14310) );
  INV_X1 U11520 ( .A(n14538), .ZN(n14293) );
  INV_X1 U11521 ( .A(n10275), .ZN(n8991) );
  INV_X1 U11522 ( .A(n14218), .ZN(n13867) );
  OAI211_X1 U11523 ( .C1(n8991), .C2(n13867), .A(n10957), .B(n10537), .ZN(
        n14215) );
  AND2_X2 U11524 ( .A1(n9996), .A2(n6591), .ZN(n15835) );
  INV_X1 U11525 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U11526 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  NAND2_X1 U11527 ( .A1(n8997), .A2(n8996), .ZN(n8998) );
  NAND2_X1 U11528 ( .A1(n8999), .A2(n8998), .ZN(P2_U3527) );
  AND2_X2 U11529 ( .A1(n9000), .A2(n15780), .ZN(n15850) );
  NAND2_X1 U11530 ( .A1(n15850), .A2(n15797), .ZN(n14649) );
  NAND2_X1 U11531 ( .A1(n8921), .A2(n9001), .ZN(n9007) );
  INV_X1 U11532 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11533 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  NAND2_X1 U11534 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U11535 ( .A1(n9007), .A2(n9006), .ZN(P2_U3495) );
  NAND4_X1 U11536 ( .A1(n9009), .A2(n9148), .A3(n9150), .A4(n9112), .ZN(n9010)
         );
  NOR2_X1 U11537 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), 
        .ZN(n9012) );
  NAND4_X1 U11538 ( .A1(n9012), .A2(n9011), .A3(n9294), .A4(n9212), .ZN(n9336)
         );
  NAND3_X1 U11539 ( .A1(n9176), .A2(n9198), .A3(n9338), .ZN(n9013) );
  NOR2_X1 U11540 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n9015) );
  NOR2_X1 U11541 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), 
        .ZN(n9014) );
  NAND4_X1 U11542 ( .A1(n9015), .A2(n9014), .A3(n9640), .A4(n9357), .ZN(n9615)
         );
  NAND3_X1 U11543 ( .A1(n9322), .A2(n9016), .A3(n9623), .ZN(n9017) );
  INV_X1 U11544 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11545 ( .A1(n9030), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U11546 ( .A1(n9065), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9029) );
  INV_X1 U11548 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9023) );
  OR2_X1 U11549 ( .A1(n9396), .A2(n9023), .ZN(n9028) );
  NAND2_X1 U11550 ( .A1(n6542), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9027) );
  INV_X1 U11551 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15912) );
  OR2_X1 U11552 ( .A1(n9437), .A2(n15912), .ZN(n9026) );
  NAND2_X1 U11553 ( .A1(n9034), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9031) );
  MUX2_X1 U11554 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9031), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n9032) );
  NAND2_X1 U11555 ( .A1(n9625), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9033) );
  NAND2_X4 U11556 ( .A1(n12424), .A2(n6545), .ZN(n9603) );
  INV_X1 U11557 ( .A(n9166), .ZN(n9119) );
  XNOR2_X1 U11558 ( .A(n7665), .B(P1_DATAO_REG_2__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U11559 ( .A(n9071), .B(n9037), .ZN(n10613) );
  INV_X1 U11560 ( .A(n10613), .ZN(n9038) );
  NAND2_X1 U11561 ( .A1(n9040), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9042) );
  XNOR2_X2 U11562 ( .A(n9042), .B(n9041), .ZN(n11088) );
  NAND2_X1 U11563 ( .A1(n9359), .A2(n11088), .ZN(n9043) );
  INV_X1 U11564 ( .A(n9556), .ZN(n9063) );
  NAND2_X1 U11565 ( .A1(n9065), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11566 ( .A1(n9345), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11567 ( .A1(n9166), .A2(SI_1_), .ZN(n9051) );
  XNOR2_X1 U11568 ( .A(n9047), .B(n9057), .ZN(n10568) );
  NAND2_X1 U11569 ( .A1(n9335), .A2(n10568), .ZN(n9050) );
  NAND2_X1 U11570 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9048) );
  XNOR2_X2 U11571 ( .A(n9048), .B(P3_IR_REG_1__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U11572 ( .A1(n9359), .A2(n11085), .ZN(n9049) );
  INV_X1 U11573 ( .A(n11665), .ZN(n9553) );
  NAND2_X1 U11574 ( .A1(n9345), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11575 ( .A1(n9065), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11576 ( .A1(n6542), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U11577 ( .A1(n9066), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9053) );
  INV_X1 U11578 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n13152) );
  MUX2_X1 U11579 ( .A(n13152), .B(n10572), .S(n9603), .Z(n9062) );
  INV_X1 U11580 ( .A(n9057), .ZN(n9060) );
  NAND2_X1 U11581 ( .A1(n9058), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11582 ( .A1(n9060), .A2(n9059), .ZN(n10571) );
  NAND2_X1 U11583 ( .A1(n9335), .A2(n10571), .ZN(n9061) );
  NAND2_X1 U11584 ( .A1(n9062), .A2(n9061), .ZN(n15869) );
  INV_X1 U11585 ( .A(n15869), .ZN(n11401) );
  NAND2_X1 U11586 ( .A1(n15866), .A2(n9554), .ZN(n9552) );
  NAND2_X1 U11587 ( .A1(n9553), .A2(n11667), .ZN(n11775) );
  NAND2_X1 U11588 ( .A1(n9063), .A2(n11775), .ZN(n9064) );
  NAND2_X1 U11589 ( .A1(n11671), .A2(n12809), .ZN(n12808) );
  NAND2_X1 U11590 ( .A1(n9064), .A2(n12808), .ZN(n11785) );
  NAND2_X1 U11591 ( .A1(n9065), .A2(n9082), .ZN(n9070) );
  NAND2_X1 U11592 ( .A1(n9066), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U11593 ( .A1(n9345), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9067) );
  INV_X1 U11594 ( .A(n13150), .ZN(n9080) );
  NAND2_X1 U11595 ( .A1(n10593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11596 ( .A1(n7665), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11597 ( .A1(n9074), .A2(n9073), .ZN(n9090) );
  XNOR2_X1 U11598 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9075) );
  XNOR2_X1 U11599 ( .A(n9090), .B(n9075), .ZN(n10611) );
  NAND2_X1 U11600 ( .A1(n9335), .A2(n10611), .ZN(n9079) );
  NAND2_X1 U11601 ( .A1(n9076), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9077) );
  XNOR2_X1 U11602 ( .A(n9077), .B(n9008), .ZN(n11152) );
  NAND2_X1 U11603 ( .A1(n9359), .A2(n11152), .ZN(n9078) );
  OAI211_X1 U11604 ( .C1(n9119), .C2(SI_3_), .A(n9079), .B(n9078), .ZN(n15913)
         );
  INV_X1 U11605 ( .A(n15913), .ZN(n12985) );
  NAND2_X1 U11606 ( .A1(n13150), .A2(n15913), .ZN(n12813) );
  NAND2_X1 U11607 ( .A1(n11785), .A2(n11790), .ZN(n11787) );
  NAND2_X1 U11608 ( .A1(n11787), .A2(n12812), .ZN(n11828) );
  NAND2_X1 U11609 ( .A1(n9345), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9087) );
  INV_X2 U11610 ( .A(n9437), .ZN(n9497) );
  NAND2_X1 U11611 ( .A1(n9497), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U11612 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9083) );
  NAND2_X1 U11613 ( .A1(n9101), .A2(n9083), .ZN(n13063) );
  NAND2_X1 U11614 ( .A1(n9065), .A2(n13063), .ZN(n9085) );
  NAND2_X1 U11615 ( .A1(n6542), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11616 ( .A1(n10596), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9091) );
  NAND2_X1 U11617 ( .A1(n9093), .A2(n9092), .ZN(n9094) );
  NAND2_X1 U11618 ( .A1(n9108), .A2(n9094), .ZN(n10607) );
  NAND2_X1 U11619 ( .A1(n9490), .A2(n10607), .ZN(n9098) );
  NAND2_X1 U11620 ( .A1(n9095), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9096) );
  XNOR2_X1 U11621 ( .A(n9096), .B(n9112), .ZN(n11094) );
  NAND2_X1 U11622 ( .A1(n9359), .A2(n11094), .ZN(n9097) );
  OAI211_X1 U11623 ( .C1(n9119), .C2(SI_4_), .A(n9098), .B(n9097), .ZN(n15918)
         );
  INV_X1 U11624 ( .A(n15918), .ZN(n13062) );
  OR2_X1 U11625 ( .A1(n11803), .A2(n13062), .ZN(n12818) );
  NAND2_X1 U11626 ( .A1(n11803), .A2(n13062), .ZN(n12819) );
  NAND2_X1 U11627 ( .A1(n12818), .A2(n12819), .ZN(n12762) );
  NAND2_X1 U11628 ( .A1(n11828), .A2(n12815), .ZN(n9099) );
  NAND2_X1 U11629 ( .A1(n9099), .A2(n12819), .ZN(n11802) );
  NAND2_X1 U11630 ( .A1(n9497), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U11631 ( .A1(n9345), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11632 ( .A1(n9101), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U11633 ( .A1(n9121), .A2(n9102), .ZN(n11808) );
  NAND2_X1 U11634 ( .A1(n9065), .A2(n11808), .ZN(n9104) );
  NAND2_X1 U11635 ( .A1(n6542), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11636 ( .A1(n10588), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9109) );
  OAI21_X1 U11637 ( .B1(n9111), .B2(n9110), .A(n9128), .ZN(n10609) );
  NAND2_X1 U11638 ( .A1(n9490), .A2(n10609), .ZN(n9118) );
  INV_X1 U11639 ( .A(n9095), .ZN(n9113) );
  NAND2_X1 U11640 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  NAND2_X1 U11641 ( .A1(n9115), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U11642 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9114), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9116) );
  NAND2_X1 U11643 ( .A1(n9116), .A2(n9147), .ZN(n11248) );
  NAND2_X1 U11644 ( .A1(n9359), .A2(n11248), .ZN(n9117) );
  OAI211_X1 U11645 ( .C1(n9119), .C2(SI_5_), .A(n9118), .B(n9117), .ZN(n11682)
         );
  INV_X1 U11646 ( .A(n11682), .ZN(n15923) );
  OR2_X1 U11647 ( .A1(n12180), .A2(n15923), .ZN(n12825) );
  NAND2_X1 U11648 ( .A1(n12180), .A2(n15923), .ZN(n12796) );
  NAND2_X1 U11649 ( .A1(n12825), .A2(n12796), .ZN(n12763) );
  NAND2_X1 U11650 ( .A1(n11802), .A2(n12821), .ZN(n9120) );
  NAND2_X1 U11651 ( .A1(n9497), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U11652 ( .A1(n9345), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U11653 ( .A1(n9121), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U11654 ( .A1(n9134), .A2(n9122), .ZN(n13112) );
  NAND2_X1 U11655 ( .A1(n9524), .A2(n13112), .ZN(n9124) );
  NAND2_X1 U11656 ( .A1(n6542), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9123) );
  XNOR2_X1 U11657 ( .A(n9142), .B(n9140), .ZN(n10601) );
  NAND2_X1 U11658 ( .A1(n12751), .A2(SI_6_), .ZN(n9131) );
  NAND2_X1 U11659 ( .A1(n9147), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U11660 ( .A1(n9359), .A2(n11283), .ZN(n9130) );
  OAI211_X1 U11661 ( .C1(n9516), .C2(n10601), .A(n9131), .B(n9130), .ZN(n13109) );
  OR2_X1 U11662 ( .A1(n12183), .A2(n13109), .ZN(n12827) );
  NAND2_X1 U11663 ( .A1(n12183), .A2(n13109), .ZN(n12830) );
  NAND2_X1 U11664 ( .A1(n12827), .A2(n12830), .ZN(n11817) );
  INV_X1 U11665 ( .A(n11817), .ZN(n12765) );
  NAND2_X1 U11666 ( .A1(n9497), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9139) );
  NAND2_X1 U11667 ( .A1(n12028), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11668 ( .A1(n9134), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11669 ( .A1(n9155), .A2(n9135), .ZN(n12953) );
  NAND2_X1 U11670 ( .A1(n9524), .A2(n12953), .ZN(n9137) );
  NAND2_X1 U11671 ( .A1(n6542), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9136) );
  INV_X1 U11672 ( .A(n9140), .ZN(n9141) );
  NAND2_X1 U11673 ( .A1(n10591), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U11674 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U11675 ( .A1(n9162), .A2(n9146), .ZN(n10603) );
  NAND2_X1 U11676 ( .A1(n10603), .A2(n9490), .ZN(n9154) );
  INV_X1 U11677 ( .A(SI_7_), .ZN(n10602) );
  NAND2_X1 U11678 ( .A1(n12751), .A2(n10602), .ZN(n9153) );
  INV_X1 U11679 ( .A(n9147), .ZN(n9149) );
  NAND2_X1 U11680 ( .A1(n9149), .A2(n9148), .ZN(n9167) );
  NAND2_X1 U11681 ( .A1(n9167), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9151) );
  XNOR2_X1 U11682 ( .A(n9151), .B(n9150), .ZN(n11266) );
  NAND2_X1 U11683 ( .A1(n9359), .A2(n11266), .ZN(n9152) );
  INV_X1 U11684 ( .A(n13147), .ZN(n11897) );
  NAND2_X1 U11685 ( .A1(n11897), .A2(n15935), .ZN(n12832) );
  NAND2_X1 U11686 ( .A1(n9497), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11687 ( .A1(n12028), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U11688 ( .A1(n9155), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11689 ( .A1(n9181), .A2(n9156), .ZN(n13004) );
  NAND2_X1 U11690 ( .A1(n9065), .A2(n13004), .ZN(n9158) );
  NAND2_X1 U11691 ( .A1(n6542), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U11692 ( .A1(n10619), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9172) );
  INV_X1 U11693 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U11694 ( .A1(n10621), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9163) );
  OAI21_X1 U11695 ( .B1(n9165), .B2(n9164), .A(n9173), .ZN(n10598) );
  OR2_X1 U11696 ( .A1(n10598), .A2(n9516), .ZN(n9170) );
  OAI21_X1 U11697 ( .B1(n9167), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9168) );
  XNOR2_X1 U11698 ( .A(n9168), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U11699 ( .A1(n12751), .A2(SI_8_), .B1(n9359), .B2(n11471), .ZN(
        n9169) );
  NAND2_X1 U11700 ( .A1(n9170), .A2(n9169), .ZN(n13003) );
  OR2_X1 U11701 ( .A1(n12193), .A2(n13003), .ZN(n12846) );
  NAND2_X1 U11702 ( .A1(n12193), .A2(n13003), .ZN(n12841) );
  NAND2_X1 U11703 ( .A1(n12846), .A2(n12841), .ZN(n12769) );
  INV_X1 U11704 ( .A(n12769), .ZN(n12835) );
  NAND2_X1 U11705 ( .A1(n11894), .A2(n12835), .ZN(n9171) );
  XNOR2_X1 U11706 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .ZN(n9188) );
  XNOR2_X1 U11707 ( .A(n9191), .B(n9188), .ZN(n10605) );
  NAND2_X1 U11708 ( .A1(n10605), .A2(n9490), .ZN(n9179) );
  INV_X1 U11709 ( .A(SI_9_), .ZN(n10604) );
  INV_X1 U11710 ( .A(n9174), .ZN(n9195) );
  NAND2_X1 U11711 ( .A1(n9195), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9177) );
  XNOR2_X1 U11712 ( .A(n9177), .B(n9176), .ZN(n11472) );
  AOI22_X1 U11713 ( .A1(n12751), .A2(n10604), .B1(n9359), .B2(n11472), .ZN(
        n9178) );
  NAND2_X1 U11714 ( .A1(n12028), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U11715 ( .A1(n6542), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11716 ( .A1(n9181), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11717 ( .A1(n9203), .A2(n9182), .ZN(n12209) );
  NAND2_X1 U11718 ( .A1(n9065), .A2(n12209), .ZN(n9184) );
  NAND2_X1 U11719 ( .A1(n9497), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9183) );
  NAND4_X1 U11720 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(n13145) );
  NAND2_X1 U11721 ( .A1(n12192), .A2(n12251), .ZN(n12851) );
  INV_X1 U11722 ( .A(n12851), .ZN(n9187) );
  INV_X1 U11723 ( .A(n9188), .ZN(n9190) );
  NAND2_X1 U11724 ( .A1(n10633), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9189) );
  INV_X1 U11725 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U11726 ( .A1(n10656), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9209) );
  INV_X1 U11727 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U11728 ( .A1(n10654), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U11729 ( .A1(n9192), .A2(n6759), .ZN(n9194) );
  NAND2_X1 U11730 ( .A1(n9210), .A2(n9194), .ZN(n10631) );
  NAND2_X1 U11731 ( .A1(n10631), .A2(n9490), .ZN(n9202) );
  NAND2_X1 U11732 ( .A1(n9197), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9196) );
  MUX2_X1 U11733 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9196), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n9200) );
  INV_X1 U11734 ( .A(n9197), .ZN(n9199) );
  NAND2_X1 U11735 ( .A1(n9199), .A2(n9198), .ZN(n9337) );
  NAND2_X1 U11736 ( .A1(n9200), .A2(n9337), .ZN(n11756) );
  AOI22_X1 U11737 ( .A1(n12751), .A2(n10630), .B1(n9359), .B2(n11756), .ZN(
        n9201) );
  NAND2_X1 U11738 ( .A1(n9497), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11739 ( .A1(n12028), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U11740 ( .A1(n9203), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U11741 ( .A1(n9216), .A2(n9204), .ZN(n12264) );
  NAND2_X1 U11742 ( .A1(n9065), .A2(n12264), .ZN(n9206) );
  NAND2_X1 U11743 ( .A1(n6542), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11744 ( .A1(n12847), .A2(n13087), .ZN(n12843) );
  XNOR2_X1 U11745 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9211) );
  XNOR2_X1 U11746 ( .A(n9223), .B(n9211), .ZN(n10652) );
  NAND2_X1 U11747 ( .A1(n10652), .A2(n9490), .ZN(n9215) );
  NAND2_X1 U11748 ( .A1(n9337), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U11749 ( .A(n9213), .B(n9212), .ZN(n11765) );
  AOI22_X1 U11750 ( .A1(n12751), .A2(n10651), .B1(n9359), .B2(n11765), .ZN(
        n9214) );
  NAND2_X1 U11751 ( .A1(n9497), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11752 ( .A1(n12028), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9220) );
  INV_X1 U11753 ( .A(n9230), .ZN(n9231) );
  NAND2_X1 U11754 ( .A1(n9216), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11755 ( .A1(n9231), .A2(n9217), .ZN(n13092) );
  NAND2_X1 U11756 ( .A1(n9065), .A2(n13092), .ZN(n9219) );
  NAND2_X1 U11757 ( .A1(n6542), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11758 ( .A1(n13095), .A2(n13144), .ZN(n12857) );
  NAND2_X1 U11759 ( .A1(n12856), .A2(n12857), .ZN(n12854) );
  NAND2_X1 U11760 ( .A1(n10659), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11761 ( .A1(n9223), .A2(n9222), .ZN(n9225) );
  NAND2_X1 U11762 ( .A1(n10661), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9224) );
  XNOR2_X1 U11763 ( .A(n9240), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n9237) );
  XNOR2_X1 U11764 ( .A(n9239), .B(n9237), .ZN(n10662) );
  NAND2_X1 U11765 ( .A1(n10662), .A2(n9490), .ZN(n9228) );
  NAND2_X1 U11766 ( .A1(n9243), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9226) );
  XNOR2_X1 U11767 ( .A(n9226), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U11768 ( .A1(n12751), .A2(SI_12_), .B1(n9359), .B2(n11938), .ZN(
        n9227) );
  NAND2_X1 U11769 ( .A1(n9228), .A2(n9227), .ZN(n13030) );
  NAND2_X1 U11770 ( .A1(n9497), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U11771 ( .A1(n12028), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9235) );
  INV_X2 U11772 ( .A(n9531), .ZN(n9524) );
  INV_X1 U11773 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11774 ( .A1(n9231), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11775 ( .A1(n9247), .A2(n9232), .ZN(n13029) );
  NAND2_X1 U11776 ( .A1(n9524), .A2(n13029), .ZN(n9234) );
  NAND2_X1 U11777 ( .A1(n6542), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9233) );
  NAND4_X1 U11778 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n13143) );
  OR2_X1 U11779 ( .A1(n13030), .A2(n13090), .ZN(n12861) );
  NAND2_X1 U11780 ( .A1(n13030), .A2(n13090), .ZN(n12860) );
  INV_X1 U11781 ( .A(n9237), .ZN(n9238) );
  NAND2_X1 U11782 ( .A1(n9240), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9241) );
  XNOR2_X1 U11783 ( .A(n9254), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U11784 ( .A1(n10816), .A2(n9490), .ZN(n9246) );
  NAND2_X1 U11785 ( .A1(n9259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9244) );
  INV_X1 U11786 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9260) );
  XNOR2_X1 U11787 ( .A(n9244), .B(n9260), .ZN(n13185) );
  AOI22_X1 U11788 ( .A1(n12751), .A2(n10815), .B1(n9359), .B2(n13185), .ZN(
        n9245) );
  NAND2_X1 U11789 ( .A1(n9497), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U11790 ( .A1(n12028), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11791 ( .A1(n9247), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U11792 ( .A1(n9269), .A2(n9248), .ZN(n13578) );
  NAND2_X1 U11793 ( .A1(n9524), .A2(n13578), .ZN(n9250) );
  NAND2_X1 U11794 ( .A1(n6542), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9249) );
  INV_X1 U11795 ( .A(n12866), .ZN(n9253) );
  NAND2_X1 U11796 ( .A1(n9254), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9256) );
  INV_X1 U11797 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U11798 ( .A1(n9276), .A2(n10925), .ZN(n9255) );
  NAND2_X1 U11799 ( .A1(n9256), .A2(n9255), .ZN(n9258) );
  XNOR2_X1 U11800 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9257) );
  XNOR2_X1 U11801 ( .A(n9258), .B(n9257), .ZN(n10922) );
  NAND2_X1 U11802 ( .A1(n10922), .A2(n9490), .ZN(n9268) );
  INV_X1 U11803 ( .A(n9259), .ZN(n9261) );
  NAND2_X1 U11804 ( .A1(n9261), .A2(n9260), .ZN(n9263) );
  NAND2_X1 U11805 ( .A1(n9263), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9262) );
  MUX2_X1 U11806 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9262), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n9266) );
  INV_X1 U11807 ( .A(n9263), .ZN(n9265) );
  INV_X1 U11808 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11809 ( .A1(n9265), .A2(n9264), .ZN(n9293) );
  NAND2_X1 U11810 ( .A1(n9266), .A2(n9293), .ZN(n13195) );
  AOI22_X1 U11811 ( .A1(n13195), .A2(n9359), .B1(n12751), .B2(n10921), .ZN(
        n9267) );
  NAND2_X1 U11812 ( .A1(n9497), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9274) );
  INV_X2 U11813 ( .A(n9396), .ZN(n12028) );
  NAND2_X1 U11814 ( .A1(n12028), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11815 ( .A1(n9269), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11816 ( .A1(n9298), .A2(n9270), .ZN(n13571) );
  NAND2_X1 U11817 ( .A1(n9524), .A2(n13571), .ZN(n9272) );
  NAND2_X1 U11818 ( .A1(n6542), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9271) );
  NAND4_X1 U11819 ( .A1(n9274), .A2(n9273), .A3(n9272), .A4(n9271), .ZN(n13545) );
  NAND2_X1 U11820 ( .A1(n13707), .A2(n13545), .ZN(n12870) );
  INV_X1 U11821 ( .A(n12870), .ZN(n13530) );
  INV_X1 U11822 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U11823 ( .A1(n10924), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9275) );
  AOI22_X1 U11824 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n10925), .B1(n10937), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11825 ( .A1(n11038), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11826 ( .A1(n11037), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11827 ( .A1(n9279), .A2(n9278), .ZN(n9291) );
  NAND2_X1 U11828 ( .A1(n11178), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11829 ( .A1(n11177), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11830 ( .A1(n9315), .A2(n9280), .ZN(n9312) );
  XNOR2_X1 U11831 ( .A(n9314), .B(n9312), .ZN(n10966) );
  NAND2_X1 U11832 ( .A1(n10966), .A2(n9490), .ZN(n9283) );
  OAI21_X1 U11833 ( .B1(n9293), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9281) );
  XNOR2_X1 U11834 ( .A(n9281), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U11835 ( .A1(n13272), .A2(n9359), .B1(SI_16_), .B2(n12751), .ZN(
        n9282) );
  INV_X1 U11836 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13539) );
  INV_X1 U11837 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11838 ( .A1(n9300), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11839 ( .A1(n9342), .A2(n9286), .ZN(n13537) );
  NAND2_X1 U11840 ( .A1(n13537), .A2(n9524), .ZN(n9290) );
  NAND2_X1 U11841 ( .A1(n12028), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11842 ( .A1(n9066), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9287) );
  AND2_X1 U11843 ( .A1(n9288), .A2(n9287), .ZN(n9289) );
  OAI211_X1 U11844 ( .C1(n9467), .C2(n13539), .A(n9290), .B(n9289), .ZN(n13546) );
  INV_X1 U11845 ( .A(n13546), .ZN(n13510) );
  OR2_X1 U11846 ( .A1(n13541), .A2(n13510), .ZN(n12876) );
  NAND2_X1 U11847 ( .A1(n13541), .A2(n13510), .ZN(n12877) );
  XNOR2_X1 U11848 ( .A(n9292), .B(n9291), .ZN(n10814) );
  NAND2_X1 U11849 ( .A1(n10814), .A2(n9490), .ZN(n9297) );
  NAND2_X1 U11850 ( .A1(n9293), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9295) );
  XNOR2_X1 U11851 ( .A(n9295), .B(n9294), .ZN(n13226) );
  AOI22_X1 U11852 ( .A1(n13226), .A2(n9359), .B1(n12751), .B2(n10813), .ZN(
        n9296) );
  NAND2_X1 U11853 ( .A1(n9298), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11854 ( .A1(n9300), .A2(n9299), .ZN(n13552) );
  NAND2_X1 U11855 ( .A1(n13552), .A2(n9524), .ZN(n9304) );
  NAND2_X1 U11856 ( .A1(n9497), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11857 ( .A1(n12028), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11858 ( .A1(n6542), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9301) );
  NAND4_X1 U11859 ( .A1(n9304), .A2(n9303), .A3(n9302), .A4(n9301), .ZN(n13565) );
  INV_X1 U11860 ( .A(n9308), .ZN(n9306) );
  NAND2_X1 U11861 ( .A1(n13651), .A2(n13565), .ZN(n12873) );
  AND2_X1 U11862 ( .A1(n13549), .A2(n13535), .ZN(n9305) );
  NOR2_X1 U11863 ( .A1(n9306), .A2(n9305), .ZN(n9310) );
  OR2_X1 U11864 ( .A1(n13530), .A2(n9310), .ZN(n9307) );
  AND2_X1 U11865 ( .A1(n13531), .A2(n9308), .ZN(n9309) );
  OR2_X1 U11866 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  INV_X1 U11867 ( .A(n9312), .ZN(n9313) );
  NAND2_X1 U11868 ( .A1(n9314), .A2(n9313), .ZN(n9316) );
  INV_X1 U11869 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U11870 ( .A1(n11201), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11871 ( .A1(n9333), .A2(n9317), .ZN(n9319) );
  NAND2_X1 U11872 ( .A1(n11199), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11873 ( .A1(n9319), .A2(n9318), .ZN(n9354) );
  XNOR2_X1 U11874 ( .A(n11403), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U11875 ( .A(n9354), .B(n9352), .ZN(n11195) );
  NAND2_X1 U11876 ( .A1(n11195), .A2(n9490), .ZN(n9326) );
  INV_X1 U11877 ( .A(n9323), .ZN(n9320) );
  NAND2_X1 U11878 ( .A1(n9320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9321) );
  MUX2_X1 U11879 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9321), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9324) );
  NAND2_X1 U11880 ( .A1(n9324), .A2(n9614), .ZN(n13311) );
  INV_X1 U11881 ( .A(n13311), .ZN(n13323) );
  AOI22_X1 U11882 ( .A1(n12751), .A2(SI_18_), .B1(n9359), .B2(n13323), .ZN(
        n9325) );
  INV_X1 U11883 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U11884 ( .A1(n9344), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11885 ( .A1(n9364), .A2(n9327), .ZN(n13502) );
  NAND2_X1 U11886 ( .A1(n13502), .A2(n9524), .ZN(n9332) );
  INV_X1 U11887 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U11888 ( .A1(n6542), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U11889 ( .A1(n12028), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9328) );
  OAI211_X1 U11890 ( .C1(n9437), .C2(n13698), .A(n9329), .B(n9328), .ZN(n9330)
         );
  INV_X1 U11891 ( .A(n9330), .ZN(n9331) );
  NAND2_X1 U11892 ( .A1(n9332), .A2(n9331), .ZN(n13141) );
  NAND2_X1 U11893 ( .A1(n13492), .A2(n13512), .ZN(n12880) );
  INV_X1 U11894 ( .A(n12880), .ZN(n9349) );
  XNOR2_X1 U11895 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n9334) );
  XNOR2_X1 U11896 ( .A(n9333), .B(n9334), .ZN(n11010) );
  NAND2_X1 U11897 ( .A1(n11010), .A2(n9490), .ZN(n9341) );
  OAI21_X1 U11898 ( .B1(n9337), .B2(n9336), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9339) );
  XNOR2_X1 U11899 ( .A(n9339), .B(n9338), .ZN(n13294) );
  AOI22_X1 U11900 ( .A1(n12751), .A2(n11009), .B1(n9359), .B2(n13294), .ZN(
        n9340) );
  INV_X1 U11901 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U11902 ( .A1(n9342), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11903 ( .A1(n9344), .A2(n9343), .ZN(n13519) );
  NAND2_X1 U11904 ( .A1(n13519), .A2(n9524), .ZN(n9347) );
  AOI22_X1 U11905 ( .A1(n9066), .A2(P3_REG0_REG_17__SCAN_IN), .B1(n9345), .B2(
        P3_REG1_REG_17__SCAN_IN), .ZN(n9346) );
  OAI211_X1 U11906 ( .C1(n9467), .C2(n13521), .A(n9347), .B(n9346), .ZN(n13527) );
  INV_X1 U11907 ( .A(n13489), .ZN(n9348) );
  NAND2_X1 U11908 ( .A1(n13643), .A2(n13527), .ZN(n9577) );
  INV_X1 U11909 ( .A(n9577), .ZN(n9350) );
  NAND2_X1 U11910 ( .A1(n12880), .A2(n9350), .ZN(n9351) );
  AND2_X1 U11911 ( .A1(n9351), .A2(n13477), .ZN(n9371) );
  INV_X1 U11912 ( .A(n9352), .ZN(n9353) );
  NAND2_X1 U11913 ( .A1(n11403), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9355) );
  XNOR2_X1 U11914 ( .A(n11481), .B(P1_DATAO_REG_19__SCAN_IN), .ZN(n9373) );
  XNOR2_X1 U11915 ( .A(n9375), .B(n9373), .ZN(n11364) );
  NAND2_X1 U11916 ( .A1(n11364), .A2(n9490), .ZN(n9361) );
  NAND2_X1 U11917 ( .A1(n9614), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9358) );
  INV_X1 U11918 ( .A(n13316), .ZN(n12754) );
  AOI22_X1 U11919 ( .A1(n12751), .A2(SI_19_), .B1(n12754), .B2(n9359), .ZN(
        n9360) );
  INV_X1 U11920 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11921 ( .A1(n9364), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U11922 ( .A1(n9380), .A2(n9365), .ZN(n13483) );
  NAND2_X1 U11923 ( .A1(n13483), .A2(n9524), .ZN(n9370) );
  INV_X1 U11924 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13309) );
  NAND2_X1 U11925 ( .A1(n9066), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11926 ( .A1(n12028), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9366) );
  OAI211_X1 U11927 ( .C1(n13309), .C2(n9467), .A(n9367), .B(n9366), .ZN(n9368)
         );
  INV_X1 U11928 ( .A(n9368), .ZN(n9369) );
  INV_X1 U11929 ( .A(n13499), .ZN(n13473) );
  OR2_X1 U11930 ( .A1(n12990), .A2(n13473), .ZN(n12886) );
  NAND2_X1 U11931 ( .A1(n12990), .A2(n13473), .ZN(n12885) );
  INV_X1 U11932 ( .A(n9373), .ZN(n9374) );
  NAND2_X1 U11933 ( .A1(n11481), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9376) );
  INV_X1 U11934 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11606) );
  XNOR2_X1 U11935 ( .A(n11606), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n9377) );
  XNOR2_X1 U11936 ( .A(n9388), .B(n9377), .ZN(n11482) );
  NAND2_X1 U11937 ( .A1(n11482), .A2(n9490), .ZN(n9379) );
  NAND2_X1 U11938 ( .A1(n12751), .A2(SI_20_), .ZN(n9378) );
  NAND2_X1 U11939 ( .A1(n9380), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U11940 ( .A1(n9392), .A2(n9381), .ZN(n13466) );
  NAND2_X1 U11941 ( .A1(n13466), .A2(n9524), .ZN(n9386) );
  INV_X1 U11942 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U11943 ( .A1(n12028), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U11944 ( .A1(n6542), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9382) );
  OAI211_X1 U11945 ( .C1(n9437), .C2(n10330), .A(n9383), .B(n9382), .ZN(n9384)
         );
  INV_X1 U11946 ( .A(n9384), .ZN(n9385) );
  OR2_X1 U11947 ( .A1(n13628), .A2(n13482), .ZN(n12889) );
  INV_X1 U11948 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11608) );
  AND2_X1 U11949 ( .A1(n11608), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9387) );
  INV_X1 U11950 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11883) );
  NAND2_X1 U11951 ( .A1(n11883), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9401) );
  INV_X1 U11952 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11881) );
  NAND2_X1 U11953 ( .A1(n11881), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9389) );
  AND2_X1 U11954 ( .A1(n9401), .A2(n9389), .ZN(n9400) );
  XNOR2_X1 U11955 ( .A(n9402), .B(n9400), .ZN(n11534) );
  NAND2_X1 U11956 ( .A1(n11534), .A2(n9490), .ZN(n9391) );
  NAND2_X1 U11957 ( .A1(n12751), .A2(SI_21_), .ZN(n9390) );
  NAND2_X1 U11958 ( .A1(n9392), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U11959 ( .A1(n9410), .A2(n9393), .ZN(n13460) );
  NAND2_X1 U11960 ( .A1(n13460), .A2(n9524), .ZN(n9399) );
  INV_X1 U11961 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U11962 ( .A1(n9066), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U11963 ( .A1(n6542), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9394) );
  OAI211_X1 U11964 ( .C1(n9396), .C2(n13625), .A(n9395), .B(n9394), .ZN(n9397)
         );
  INV_X1 U11965 ( .A(n9397), .ZN(n9398) );
  NAND2_X1 U11966 ( .A1(n13459), .A2(n13474), .ZN(n13439) );
  INV_X1 U11967 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U11968 ( .A1(n9403), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9423) );
  INV_X1 U11969 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U11970 ( .A1(n11774), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9404) );
  AND2_X1 U11971 ( .A1(n9423), .A2(n9404), .ZN(n9405) );
  NAND2_X1 U11972 ( .A1(n9406), .A2(n9405), .ZN(n9424) );
  OR2_X1 U11973 ( .A1(n9406), .A2(n9405), .ZN(n9407) );
  AND2_X1 U11974 ( .A1(n9424), .A2(n9407), .ZN(n11542) );
  NAND2_X1 U11975 ( .A1(n11542), .A2(n9490), .ZN(n9409) );
  NAND2_X1 U11976 ( .A1(n12751), .A2(SI_22_), .ZN(n9408) );
  NAND2_X1 U11977 ( .A1(n9410), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11978 ( .A1(n9445), .A2(n9411), .ZN(n13448) );
  NAND2_X1 U11979 ( .A1(n13448), .A2(n9524), .ZN(n9417) );
  INV_X1 U11980 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11981 ( .A1(n12028), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11982 ( .A1(n9497), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9412) );
  OAI211_X1 U11983 ( .C1(n9414), .C2(n9467), .A(n9413), .B(n9412), .ZN(n9415)
         );
  INV_X1 U11984 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11985 ( .A1(n13080), .A2(n13458), .ZN(n12896) );
  AND2_X1 U11986 ( .A1(n13439), .A2(n12896), .ZN(n9418) );
  NAND2_X1 U11987 ( .A1(n13438), .A2(n9418), .ZN(n9422) );
  INV_X1 U11988 ( .A(n12896), .ZN(n9420) );
  NAND2_X1 U11989 ( .A1(n13687), .A2(n13427), .ZN(n12895) );
  AND2_X1 U11990 ( .A1(n13440), .A2(n12895), .ZN(n9419) );
  NAND2_X1 U11991 ( .A1(n9422), .A2(n9421), .ZN(n13380) );
  INV_X1 U11992 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9425) );
  XNOR2_X1 U11993 ( .A(n9425), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11994 ( .A1(n9425), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9426) );
  INV_X1 U11995 ( .A(n9429), .ZN(n9428) );
  INV_X1 U11996 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9427) );
  XNOR2_X1 U11997 ( .A(n9453), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12271) );
  NAND2_X1 U11998 ( .A1(n12271), .A2(n9490), .ZN(n9432) );
  NAND2_X1 U11999 ( .A1(n12751), .A2(SI_24_), .ZN(n9431) );
  NAND2_X2 U12000 ( .A1(n9432), .A2(n9431), .ZN(n13610) );
  INV_X1 U12001 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U12002 ( .A1(n9447), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U12003 ( .A1(n9463), .A2(n9434), .ZN(n13414) );
  NAND2_X1 U12004 ( .A1(n13414), .A2(n9524), .ZN(n9440) );
  INV_X1 U12005 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n10378) );
  NAND2_X1 U12006 ( .A1(n6542), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U12007 ( .A1(n12028), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9435) );
  OAI211_X1 U12008 ( .C1(n9437), .C2(n10378), .A(n9436), .B(n9435), .ZN(n9438)
         );
  INV_X1 U12009 ( .A(n9438), .ZN(n9439) );
  XNOR2_X1 U12010 ( .A(n9442), .B(n9441), .ZN(n11852) );
  NAND2_X1 U12011 ( .A1(n11852), .A2(n9490), .ZN(n9444) );
  NAND2_X1 U12012 ( .A1(n12751), .A2(SI_23_), .ZN(n9443) );
  NAND2_X1 U12013 ( .A1(n9445), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U12014 ( .A1(n9447), .A2(n9446), .ZN(n13423) );
  NAND2_X1 U12015 ( .A1(n13423), .A2(n9524), .ZN(n9452) );
  INV_X1 U12016 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13424) );
  NAND2_X1 U12017 ( .A1(n9497), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U12018 ( .A1(n12028), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9448) );
  OAI211_X1 U12019 ( .C1(n13424), .C2(n9467), .A(n9449), .B(n9448), .ZN(n9450)
         );
  INV_X1 U12020 ( .A(n9450), .ZN(n9451) );
  OR3_X2 U12021 ( .A1(n13380), .A2(n12899), .A3(n13404), .ZN(n9473) );
  NAND2_X1 U12022 ( .A1(n13614), .A2(n13447), .ZN(n9588) );
  NAND2_X1 U12023 ( .A1(n9454), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12024 ( .A1(n12121), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9455) );
  AND2_X1 U12025 ( .A1(n9475), .A2(n9455), .ZN(n9456) );
  NAND2_X1 U12026 ( .A1(n12751), .A2(SI_25_), .ZN(n9459) );
  INV_X1 U12027 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U12028 ( .A1(n9463), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U12029 ( .A1(n9481), .A2(n9464), .ZN(n13395) );
  NAND2_X1 U12030 ( .A1(n13395), .A2(n9524), .ZN(n9470) );
  INV_X1 U12031 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U12032 ( .A1(n9066), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U12033 ( .A1(n12028), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9465) );
  OAI211_X1 U12034 ( .C1(n13396), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9468)
         );
  INV_X1 U12035 ( .A(n9468), .ZN(n9469) );
  NAND2_X1 U12036 ( .A1(n13399), .A2(n13410), .ZN(n12905) );
  OAI211_X1 U12037 ( .C1(n12899), .C2(n9588), .A(n12905), .B(n13383), .ZN(
        n9471) );
  INV_X1 U12038 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U12039 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  INV_X1 U12040 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U12041 ( .A1(n12160), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9487) );
  INV_X1 U12042 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U12043 ( .A1(n12158), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9477) );
  AND2_X1 U12044 ( .A1(n9487), .A2(n9477), .ZN(n9478) );
  NAND2_X1 U12045 ( .A1(n9479), .A2(n9478), .ZN(n9488) );
  NAND2_X1 U12046 ( .A1(n12751), .A2(SI_26_), .ZN(n9480) );
  NAND2_X1 U12047 ( .A1(n9481), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U12048 ( .A1(n9495), .A2(n9482), .ZN(n13375) );
  NAND2_X1 U12049 ( .A1(n6542), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U12050 ( .A1(n9066), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U12051 ( .A1(n12028), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9483) );
  AND3_X1 U12052 ( .A1(n9485), .A2(n9484), .A3(n9483), .ZN(n9486) );
  NAND2_X1 U12053 ( .A1(n9594), .A2(n13357), .ZN(n12761) );
  NAND2_X1 U12054 ( .A1(n12302), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U12055 ( .A1(n12401), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U12056 ( .A1(n9506), .A2(n9489), .ZN(n9503) );
  XNOR2_X1 U12057 ( .A(n9505), .B(n9503), .ZN(n13726) );
  NAND2_X1 U12058 ( .A1(n13726), .A2(n9490), .ZN(n9492) );
  NAND2_X1 U12059 ( .A1(n12751), .A2(SI_27_), .ZN(n9491) );
  INV_X1 U12060 ( .A(n9495), .ZN(n9494) );
  INV_X1 U12061 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U12062 ( .A1(n9495), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U12063 ( .A1(n9518), .A2(n9496), .ZN(n13361) );
  NAND2_X1 U12064 ( .A1(n13361), .A2(n9524), .ZN(n9502) );
  NAND2_X1 U12065 ( .A1(n6542), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U12066 ( .A1(n9497), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U12067 ( .A1(n12028), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9498) );
  AND3_X1 U12068 ( .A1(n9500), .A2(n9499), .A3(n9498), .ZN(n9501) );
  INV_X1 U12069 ( .A(n13343), .ZN(n13370) );
  INV_X1 U12070 ( .A(n9503), .ZN(n9504) );
  NAND2_X1 U12071 ( .A1(n9505), .A2(n9504), .ZN(n9507) );
  INV_X1 U12072 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15432) );
  NAND2_X1 U12073 ( .A1(n15432), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12074 ( .A1(n9508), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9509) );
  AND2_X1 U12075 ( .A1(n9526), .A2(n9509), .ZN(n9511) );
  INV_X1 U12076 ( .A(n9510), .ZN(n9513) );
  INV_X1 U12077 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U12078 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  NAND2_X1 U12079 ( .A1(n9527), .A2(n9514), .ZN(n12425) );
  NAND2_X1 U12080 ( .A1(n12751), .A2(SI_28_), .ZN(n9515) );
  OAI21_X2 U12081 ( .B1(n12425), .B2(n9516), .A(n9515), .ZN(n9525) );
  NAND2_X1 U12082 ( .A1(n9518), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U12083 ( .A1(n12716), .A2(n9519), .ZN(n13349) );
  NAND2_X1 U12084 ( .A1(n6542), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U12085 ( .A1(n12028), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U12086 ( .A1(n9066), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9520) );
  NAND3_X1 U12087 ( .A1(n9522), .A2(n9521), .A3(n9520), .ZN(n9523) );
  INV_X1 U12088 ( .A(n12916), .ZN(n12920) );
  NAND2_X1 U12089 ( .A1(n9525), .A2(n13358), .ZN(n12918) );
  INV_X1 U12090 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12734) );
  XNOR2_X1 U12091 ( .A(n12734), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n9528) );
  XNOR2_X1 U12092 ( .A(n12736), .B(n9528), .ZN(n13721) );
  NAND2_X1 U12093 ( .A1(n13721), .A2(n9490), .ZN(n9530) );
  NAND2_X1 U12094 ( .A1(n12751), .A2(SI_29_), .ZN(n9529) );
  NAND2_X1 U12095 ( .A1(n9066), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9534) );
  NAND2_X1 U12096 ( .A1(n12028), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U12097 ( .A1(n6542), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9532) );
  AND3_X1 U12098 ( .A1(n9534), .A2(n9533), .A3(n9532), .ZN(n9535) );
  NAND2_X1 U12099 ( .A1(n9664), .A2(n13345), .ZN(n12925) );
  XNOR2_X1 U12100 ( .A(n12757), .B(n12914), .ZN(n12720) );
  INV_X1 U12101 ( .A(n9540), .ZN(n9537) );
  NAND2_X1 U12102 ( .A1(n9537), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9538) );
  INV_X1 U12103 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U12104 ( .A1(n9540), .A2(n9539), .ZN(n9631) );
  INV_X1 U12105 ( .A(n9541), .ZN(n9542) );
  NAND2_X1 U12106 ( .A1(n9542), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9543) );
  OAI21_X1 U12107 ( .B1(n12800), .B2(n12790), .A(n12754), .ZN(n9546) );
  NAND2_X1 U12108 ( .A1(n9544), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U12109 ( .A1(n9546), .A2(n12801), .ZN(n9548) );
  OAI21_X1 U12110 ( .B1(n12790), .B2(n12755), .A(n12800), .ZN(n9547) );
  NAND2_X1 U12111 ( .A1(n9548), .A2(n9547), .ZN(n11687) );
  AND2_X1 U12112 ( .A1(n15928), .A2(n12937), .ZN(n9549) );
  NAND2_X1 U12113 ( .A1(n11687), .A2(n9549), .ZN(n9551) );
  AND2_X1 U12114 ( .A1(n12790), .A2(n13316), .ZN(n9550) );
  NAND2_X1 U12115 ( .A1(n12946), .A2(n9550), .ZN(n9656) );
  NAND2_X1 U12116 ( .A1(n11659), .A2(n12754), .ZN(n11417) );
  OR2_X1 U12117 ( .A1(n12946), .A2(n11417), .ZN(n15930) );
  OR2_X1 U12118 ( .A1(n12720), .A2(n13630), .ZN(n9613) );
  INV_X1 U12119 ( .A(n13358), .ZN(n13138) );
  INV_X1 U12120 ( .A(n9552), .ZN(n12803) );
  INV_X1 U12121 ( .A(n11668), .ZN(n12403) );
  INV_X1 U12122 ( .A(n11663), .ZN(n9555) );
  NAND2_X1 U12123 ( .A1(n11777), .A2(n12804), .ZN(n11793) );
  INV_X1 U12124 ( .A(n11790), .ZN(n12764) );
  NAND2_X1 U12125 ( .A1(n11671), .A2(n11670), .ZN(n11789) );
  AND2_X1 U12126 ( .A1(n12764), .A2(n11789), .ZN(n11792) );
  OR2_X1 U12127 ( .A1(n11803), .A2(n15918), .ZN(n9559) );
  INV_X1 U12128 ( .A(n9559), .ZN(n9557) );
  OR2_X1 U12129 ( .A1(n9557), .A2(n12762), .ZN(n9558) );
  NAND2_X1 U12130 ( .A1(n13150), .A2(n12985), .ZN(n11829) );
  INV_X1 U12131 ( .A(n13109), .ZN(n15929) );
  OR2_X1 U12132 ( .A1(n12183), .A2(n15929), .ZN(n11949) );
  NAND2_X1 U12133 ( .A1(n12763), .A2(n11949), .ZN(n9561) );
  NAND2_X1 U12134 ( .A1(n12180), .A2(n11682), .ZN(n11818) );
  NAND2_X1 U12135 ( .A1(n11817), .A2(n11818), .ZN(n11815) );
  AOI21_X1 U12136 ( .B1(n11815), .B2(n11949), .A(n12829), .ZN(n9560) );
  NAND2_X1 U12137 ( .A1(n13147), .A2(n15935), .ZN(n9562) );
  NAND2_X1 U12138 ( .A1(n9563), .A2(n9562), .ZN(n11895) );
  NAND2_X1 U12139 ( .A1(n12192), .A2(n13145), .ZN(n11998) );
  NAND2_X1 U12140 ( .A1(n11998), .A2(n12769), .ZN(n9566) );
  NAND2_X1 U12141 ( .A1(n12845), .A2(n12851), .ZN(n12042) );
  INV_X1 U12142 ( .A(n13003), .ZN(n12038) );
  NAND2_X1 U12143 ( .A1(n12193), .A2(n12038), .ZN(n11996) );
  NAND2_X1 U12144 ( .A1(n12042), .A2(n11996), .ZN(n9564) );
  NAND2_X1 U12145 ( .A1(n9564), .A2(n11998), .ZN(n9565) );
  OAI211_X1 U12146 ( .C1(n11895), .C2(n9566), .A(n12850), .B(n9565), .ZN(n9568) );
  INV_X1 U12147 ( .A(n13087), .ZN(n12207) );
  OR2_X1 U12148 ( .A1(n12847), .A2(n12207), .ZN(n9567) );
  NAND2_X1 U12149 ( .A1(n9568), .A2(n9567), .ZN(n12241) );
  NOR2_X1 U12150 ( .A1(n13095), .A2(n13085), .ZN(n12240) );
  NAND2_X1 U12151 ( .A1(n13095), .A2(n13085), .ZN(n12242) );
  OAI21_X1 U12152 ( .B1(n12241), .B2(n12240), .A(n7643), .ZN(n9572) );
  INV_X1 U12153 ( .A(n9569), .ZN(n9570) );
  AND2_X1 U12154 ( .A1(n13030), .A2(n13143), .ZN(n12325) );
  NAND2_X1 U12155 ( .A1(n9570), .A2(n12325), .ZN(n9571) );
  OAI211_X1 U12156 ( .C1(n13027), .C2(n13583), .A(n9572), .B(n9571), .ZN(
        n13561) );
  INV_X1 U12157 ( .A(n13545), .ZN(n12313) );
  OR2_X1 U12158 ( .A1(n13707), .A2(n12313), .ZN(n9573) );
  INV_X1 U12159 ( .A(n13565), .ZN(n12968) );
  NAND2_X1 U12160 ( .A1(n13651), .A2(n12968), .ZN(n9574) );
  OR2_X1 U12161 ( .A1(n13651), .A2(n12968), .ZN(n9575) );
  OR2_X1 U12162 ( .A1(n13541), .A2(n13546), .ZN(n9576) );
  NAND2_X1 U12163 ( .A1(n13477), .A2(n12880), .ZN(n12881) );
  INV_X1 U12164 ( .A(n13527), .ZN(n13046) );
  OR2_X1 U12165 ( .A1(n13643), .A2(n13046), .ZN(n13495) );
  AND2_X1 U12166 ( .A1(n12881), .A2(n13495), .ZN(n9580) );
  NAND3_X1 U12167 ( .A1(n12881), .A2(n13517), .A3(n13495), .ZN(n9578) );
  OAI21_X1 U12168 ( .B1(n13492), .B2(n13141), .A(n9578), .ZN(n9579) );
  OR2_X1 U12169 ( .A1(n12990), .A2(n13499), .ZN(n12778) );
  NAND2_X1 U12170 ( .A1(n12990), .A2(n13499), .ZN(n12777) );
  NAND2_X1 U12171 ( .A1(n13628), .A2(n13013), .ZN(n9581) );
  OR2_X1 U12172 ( .A1(n13459), .A2(n13140), .ZN(n9584) );
  NAND2_X1 U12173 ( .A1(n13080), .A2(n13427), .ZN(n9585) );
  NAND2_X1 U12174 ( .A1(n13687), .A2(n13458), .ZN(n9586) );
  NAND2_X1 U12175 ( .A1(n13614), .A2(n13139), .ZN(n9589) );
  AND2_X1 U12176 ( .A1(n13399), .A2(n13119), .ZN(n9591) );
  OR2_X1 U12177 ( .A1(n13407), .A2(n9591), .ZN(n9593) );
  INV_X1 U12178 ( .A(n9591), .ZN(n9592) );
  OR2_X1 U12179 ( .A1(n13610), .A2(n13428), .ZN(n13387) );
  OR2_X1 U12180 ( .A1(n9594), .A2(n13385), .ZN(n9595) );
  NAND2_X1 U12181 ( .A1(n13369), .A2(n9595), .ZN(n9597) );
  NAND2_X1 U12182 ( .A1(n9594), .A2(n13385), .ZN(n9596) );
  OR2_X1 U12183 ( .A1(n13674), .A2(n13343), .ZN(n9599) );
  INV_X2 U12184 ( .A(n13338), .ZN(n13340) );
  XNOR2_X1 U12185 ( .A(n12914), .B(n9600), .ZN(n9612) );
  OR2_X1 U12186 ( .A1(n12800), .A2(n13316), .ZN(n10231) );
  NAND2_X1 U12187 ( .A1(n12755), .A2(n12790), .ZN(n9601) );
  INV_X1 U12188 ( .A(n12424), .ZN(n12942) );
  NAND2_X1 U12189 ( .A1(n12942), .A2(n6821), .ZN(n11082) );
  NAND2_X1 U12190 ( .A1(n11082), .A2(n9603), .ZN(n11700) );
  INV_X1 U12191 ( .A(n11700), .ZN(n9604) );
  NAND2_X1 U12192 ( .A1(n9602), .A2(n9604), .ZN(n13509) );
  NAND2_X1 U12193 ( .A1(n6542), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9607) );
  NAND2_X1 U12194 ( .A1(n9066), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U12195 ( .A1(n12028), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9605) );
  AND3_X1 U12196 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(n9608) );
  NAND2_X1 U12197 ( .A1(n9602), .A2(n11700), .ZN(n13511) );
  INV_X1 U12198 ( .A(P3_B_REG_SCAN_IN), .ZN(n9609) );
  NOR2_X1 U12199 ( .A1(n12424), .A2(n9609), .ZN(n9610) );
  OR2_X1 U12200 ( .A1(n13511), .A2(n9610), .ZN(n13332) );
  OAI22_X1 U12201 ( .A1(n13358), .A2(n13509), .B1(n12930), .B2(n13332), .ZN(
        n9611) );
  NAND2_X1 U12202 ( .A1(n9613), .A2(n12714), .ZN(n10238) );
  INV_X1 U12203 ( .A(n9615), .ZN(n9616) );
  NAND2_X1 U12204 ( .A1(n9618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9617) );
  MUX2_X1 U12205 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9617), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9619) );
  XNOR2_X1 U12206 ( .A(P3_IR_REG_24__SCAN_IN), .B(P3_IR_REG_23__SCAN_IN), .ZN(
        n9620) );
  XNOR2_X1 U12207 ( .A(n9620), .B(P3_B_REG_SCAN_IN), .ZN(n9621) );
  NAND2_X1 U12208 ( .A1(n9622), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9624) );
  INV_X1 U12209 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9632) );
  XNOR2_X1 U12210 ( .A(n9633), .B(n9632), .ZN(n9637) );
  NAND2_X1 U12211 ( .A1(n9637), .A2(n12323), .ZN(n9634) );
  INV_X1 U12212 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U12213 ( .A1(n10752), .A2(n10617), .ZN(n9636) );
  NAND2_X1 U12214 ( .A1(n12323), .A2(n12300), .ZN(n9635) );
  NAND2_X1 U12215 ( .A1(n9636), .A2(n9635), .ZN(n11406) );
  XNOR2_X1 U12216 ( .A(n11658), .B(n11410), .ZN(n9653) );
  INV_X1 U12217 ( .A(n9637), .ZN(n9639) );
  NOR2_X1 U12218 ( .A1(n12323), .A2(n12300), .ZN(n9638) );
  NAND2_X1 U12219 ( .A1(n9639), .A2(n9638), .ZN(n11692) );
  NAND2_X1 U12220 ( .A1(n9631), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9641) );
  XNOR2_X1 U12221 ( .A(n9641), .B(n9640), .ZN(n11069) );
  NOR2_X1 U12222 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .ZN(
        n9645) );
  NOR4_X1 U12223 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9644) );
  NOR4_X1 U12224 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9643) );
  NOR4_X1 U12225 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9642) );
  NAND4_X1 U12226 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(n9651)
         );
  NOR4_X1 U12227 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9649) );
  NOR4_X1 U12228 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9648) );
  NOR4_X1 U12229 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9647) );
  NOR4_X1 U12230 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9646) );
  NAND4_X1 U12231 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(n9650)
         );
  OAI21_X1 U12232 ( .B1(n9651), .B2(n9650), .A(n10752), .ZN(n10233) );
  INV_X1 U12233 ( .A(n10233), .ZN(n10229) );
  NOR2_X1 U12234 ( .A1(n11702), .A2(n10229), .ZN(n9652) );
  NAND2_X1 U12235 ( .A1(n12946), .A2(n13316), .ZN(n9654) );
  OAI21_X1 U12236 ( .B1(n15928), .B2(n12790), .A(n9654), .ZN(n9655) );
  AOI21_X1 U12237 ( .B1(n9655), .B2(n11661), .A(n9602), .ZN(n9660) );
  INV_X1 U12238 ( .A(n9656), .ZN(n9657) );
  NAND2_X1 U12239 ( .A1(n9602), .A2(n11661), .ZN(n11690) );
  NAND2_X1 U12240 ( .A1(n11409), .A2(n11690), .ZN(n9658) );
  NAND2_X1 U12241 ( .A1(n9658), .A2(n11410), .ZN(n9659) );
  OAI21_X1 U12242 ( .B1(n9660), .B2(n11410), .A(n9659), .ZN(n9661) );
  INV_X1 U12243 ( .A(n9661), .ZN(n9662) );
  INV_X1 U12244 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9663) );
  NOR2_X1 U12245 ( .A1(n15954), .A2(n9663), .ZN(n9665) );
  INV_X1 U12246 ( .A(n15928), .ZN(n15936) );
  NAND2_X1 U12247 ( .A1(n9667), .A2(n9666), .ZN(P3_U3488) );
  NAND2_X1 U12248 ( .A1(n6596), .A2(n9722), .ZN(n9669) );
  NOR2_X1 U12249 ( .A1(n11301), .A2(n9671), .ZN(n9673) );
  NAND2_X1 U12250 ( .A1(n11301), .A2(n9671), .ZN(n9672) );
  OAI211_X1 U12251 ( .C1(n9670), .C2(n9673), .A(n9722), .B(n9672), .ZN(n9675)
         );
  NAND2_X1 U12252 ( .A1(n9670), .A2(n11335), .ZN(n10958) );
  NAND2_X1 U12253 ( .A1(n9675), .A2(n9674), .ZN(n9680) );
  NAND2_X1 U12254 ( .A1(n9680), .A2(n9681), .ZN(n9678) );
  NAND2_X1 U12255 ( .A1(n9787), .A2(n6596), .ZN(n9676) );
  OAI21_X1 U12256 ( .B1(n9787), .B2(n8535), .A(n9676), .ZN(n9677) );
  NAND2_X1 U12257 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  NAND2_X1 U12258 ( .A1(n9787), .A2(n14041), .ZN(n9683) );
  NAND2_X1 U12259 ( .A1(n9914), .A2(n15764), .ZN(n9682) );
  NAND2_X1 U12260 ( .A1(n9683), .A2(n9682), .ZN(n9688) );
  NAND2_X1 U12261 ( .A1(n14041), .A2(n6595), .ZN(n9684) );
  OAI21_X1 U12262 ( .B1(n15793), .B2(n6550), .A(n9684), .ZN(n9685) );
  NAND2_X1 U12263 ( .A1(n9686), .A2(n9685), .ZN(n9692) );
  INV_X1 U12264 ( .A(n9687), .ZN(n9690) );
  INV_X1 U12265 ( .A(n9688), .ZN(n9689) );
  CLKBUF_X1 U12266 ( .A(n9722), .Z(n9815) );
  NAND2_X1 U12267 ( .A1(n14040), .A2(n9914), .ZN(n9693) );
  OAI21_X1 U12268 ( .B1(n6550), .B2(n15804), .A(n9693), .ZN(n9696) );
  NAND2_X1 U12269 ( .A1(n9787), .A2(n14040), .ZN(n9694) );
  OAI21_X1 U12270 ( .B1(n9787), .B2(n15804), .A(n9694), .ZN(n9695) );
  INV_X1 U12271 ( .A(n9696), .ZN(n9697) );
  NAND2_X1 U12272 ( .A1(n9787), .A2(n14039), .ZN(n9699) );
  NAND2_X1 U12273 ( .A1(n11324), .A2(n6550), .ZN(n9698) );
  NAND2_X1 U12274 ( .A1(n9699), .A2(n9698), .ZN(n9704) );
  NAND2_X1 U12275 ( .A1(n9703), .A2(n9704), .ZN(n9702) );
  NAND2_X1 U12276 ( .A1(n14039), .A2(n6600), .ZN(n9700) );
  OAI21_X1 U12277 ( .B1(n15811), .B2(n6550), .A(n9700), .ZN(n9701) );
  NAND2_X1 U12278 ( .A1(n9702), .A2(n9701), .ZN(n9708) );
  INV_X1 U12279 ( .A(n9703), .ZN(n9706) );
  INV_X1 U12280 ( .A(n9704), .ZN(n9705) );
  NAND2_X1 U12281 ( .A1(n9706), .A2(n9705), .ZN(n9707) );
  NAND2_X1 U12282 ( .A1(n14038), .A2(n6550), .ZN(n9709) );
  OAI21_X1 U12283 ( .B1(n9914), .B2(n11520), .A(n9709), .ZN(n9712) );
  NAND2_X1 U12284 ( .A1(n9787), .A2(n14038), .ZN(n9710) );
  OAI21_X1 U12285 ( .B1(n9787), .B2(n11520), .A(n9710), .ZN(n9711) );
  NAND2_X1 U12286 ( .A1(n6546), .A2(n14037), .ZN(n9713) );
  OAI21_X1 U12287 ( .B1(n6546), .B2(n11561), .A(n9713), .ZN(n9718) );
  NAND2_X1 U12288 ( .A1(n14037), .A2(n6550), .ZN(n9714) );
  OAI21_X1 U12289 ( .B1(n11561), .B2(n6550), .A(n9714), .ZN(n9715) );
  NAND2_X1 U12290 ( .A1(n9716), .A2(n9715), .ZN(n9721) );
  INV_X1 U12291 ( .A(n9718), .ZN(n9719) );
  NAND2_X1 U12292 ( .A1(n15834), .A2(n6546), .ZN(n9723) );
  OAI21_X1 U12293 ( .B1(n11873), .B2(n6546), .A(n9723), .ZN(n9725) );
  MUX2_X1 U12294 ( .A(n11873), .B(n11741), .S(n6600), .Z(n9724) );
  NAND2_X1 U12295 ( .A1(n6607), .A2(n6600), .ZN(n9729) );
  NAND2_X1 U12296 ( .A1(n6546), .A2(n14035), .ZN(n9728) );
  NAND2_X1 U12297 ( .A1(n6607), .A2(n6546), .ZN(n9730) );
  OAI21_X1 U12298 ( .B1(n13939), .B2(n6546), .A(n9730), .ZN(n9731) );
  NAND2_X1 U12299 ( .A1(n14604), .A2(n6546), .ZN(n9733) );
  NAND2_X1 U12300 ( .A1(n14034), .A2(n9914), .ZN(n9732) );
  NAND2_X1 U12301 ( .A1(n9733), .A2(n9732), .ZN(n9738) );
  NAND2_X1 U12302 ( .A1(n9737), .A2(n9738), .ZN(n9736) );
  NAND2_X1 U12303 ( .A1(n14604), .A2(n6600), .ZN(n9734) );
  OAI21_X1 U12304 ( .B1(n13839), .B2(n6595), .A(n9734), .ZN(n9735) );
  NAND2_X1 U12305 ( .A1(n9736), .A2(n9735), .ZN(n9742) );
  INV_X1 U12306 ( .A(n9737), .ZN(n9740) );
  INV_X1 U12307 ( .A(n9738), .ZN(n9739) );
  NAND2_X1 U12308 ( .A1(n9740), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U12309 ( .A1(n13842), .A2(n9914), .ZN(n9744) );
  NAND2_X1 U12310 ( .A1(n14497), .A2(n6546), .ZN(n9743) );
  NAND2_X1 U12311 ( .A1(n9744), .A2(n9743), .ZN(n9749) );
  NAND2_X1 U12312 ( .A1(n9748), .A2(n9749), .ZN(n9747) );
  NAND2_X1 U12313 ( .A1(n13842), .A2(n6546), .ZN(n9745) );
  OAI21_X1 U12314 ( .B1(n13977), .B2(n6546), .A(n9745), .ZN(n9746) );
  NAND2_X1 U12315 ( .A1(n9747), .A2(n9746), .ZN(n9753) );
  INV_X1 U12316 ( .A(n9748), .ZN(n9751) );
  INV_X1 U12317 ( .A(n9749), .ZN(n9750) );
  NAND2_X1 U12318 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U12319 ( .A1(n14598), .A2(n6546), .ZN(n9755) );
  NAND2_X1 U12320 ( .A1(n14033), .A2(n6600), .ZN(n9754) );
  NAND2_X1 U12321 ( .A1(n9755), .A2(n9754), .ZN(n9758) );
  NAND2_X1 U12322 ( .A1(n14598), .A2(n6595), .ZN(n9756) );
  OAI21_X1 U12323 ( .B1(n14472), .B2(n6595), .A(n9756), .ZN(n9757) );
  INV_X1 U12324 ( .A(n9758), .ZN(n9759) );
  NAND2_X1 U12325 ( .A1(n14593), .A2(n9914), .ZN(n9761) );
  NAND2_X1 U12326 ( .A1(n14495), .A2(n6546), .ZN(n9760) );
  NAND2_X1 U12327 ( .A1(n9761), .A2(n9760), .ZN(n9765) );
  NAND2_X1 U12328 ( .A1(n9764), .A2(n9765), .ZN(n9763) );
  MUX2_X1 U12329 ( .A(n14495), .B(n14593), .S(n6546), .Z(n9762) );
  NAND2_X1 U12330 ( .A1(n9763), .A2(n9762), .ZN(n9769) );
  INV_X1 U12331 ( .A(n9764), .ZN(n9767) );
  INV_X1 U12332 ( .A(n9765), .ZN(n9766) );
  NAND2_X1 U12333 ( .A1(n9767), .A2(n9766), .ZN(n9768) );
  NAND2_X1 U12334 ( .A1(n9769), .A2(n9768), .ZN(n9774) );
  NAND2_X1 U12335 ( .A1(n14589), .A2(n6546), .ZN(n9771) );
  NAND2_X1 U12336 ( .A1(n14032), .A2(n6550), .ZN(n9770) );
  NAND2_X1 U12337 ( .A1(n9771), .A2(n9770), .ZN(n9775) );
  NAND2_X1 U12338 ( .A1(n9774), .A2(n9775), .ZN(n9773) );
  MUX2_X1 U12339 ( .A(n14032), .B(n14589), .S(n9914), .Z(n9772) );
  NAND2_X1 U12340 ( .A1(n9773), .A2(n9772), .ZN(n9779) );
  INV_X1 U12341 ( .A(n9774), .ZN(n9777) );
  INV_X1 U12342 ( .A(n9775), .ZN(n9776) );
  NAND2_X1 U12343 ( .A1(n9777), .A2(n9776), .ZN(n9778) );
  NAND2_X1 U12344 ( .A1(n14583), .A2(n9914), .ZN(n9781) );
  NAND2_X1 U12345 ( .A1(n6546), .A2(n14031), .ZN(n9780) );
  NAND2_X1 U12346 ( .A1(n9781), .A2(n9780), .ZN(n9786) );
  NAND2_X1 U12347 ( .A1(n14583), .A2(n6546), .ZN(n9782) );
  OAI21_X1 U12348 ( .B1(n9783), .B2(n6546), .A(n9782), .ZN(n9784) );
  NAND2_X1 U12349 ( .A1(n14578), .A2(n6546), .ZN(n9789) );
  NAND2_X1 U12350 ( .A1(n14030), .A2(n6595), .ZN(n9788) );
  NAND2_X1 U12351 ( .A1(n9789), .A2(n9788), .ZN(n9794) );
  NAND2_X1 U12352 ( .A1(n14578), .A2(n9914), .ZN(n9790) );
  OAI21_X1 U12353 ( .B1(n9791), .B2(n6550), .A(n9790), .ZN(n9792) );
  NAND2_X1 U12354 ( .A1(n14573), .A2(n6600), .ZN(n9797) );
  NAND2_X1 U12355 ( .A1(n14029), .A2(n6546), .ZN(n9796) );
  NAND2_X1 U12356 ( .A1(n9797), .A2(n9796), .ZN(n9803) );
  NAND2_X1 U12357 ( .A1(n14573), .A2(n6546), .ZN(n9798) );
  OAI21_X1 U12358 ( .B1(n9799), .B2(n6546), .A(n9798), .ZN(n9800) );
  NAND2_X1 U12359 ( .A1(n9801), .A2(n9800), .ZN(n9807) );
  INV_X1 U12360 ( .A(n9802), .ZN(n9805) );
  INV_X1 U12361 ( .A(n9803), .ZN(n9804) );
  NAND2_X1 U12362 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  NAND2_X1 U12363 ( .A1(n9807), .A2(n9806), .ZN(n9812) );
  NAND2_X1 U12364 ( .A1(n14568), .A2(n6546), .ZN(n9809) );
  NAND2_X1 U12365 ( .A1(n14028), .A2(n6595), .ZN(n9808) );
  NAND2_X1 U12366 ( .A1(n9809), .A2(n9808), .ZN(n9813) );
  NAND2_X1 U12367 ( .A1(n14568), .A2(n6595), .ZN(n9810) );
  OAI21_X1 U12368 ( .B1(n13987), .B2(n6595), .A(n9810), .ZN(n9811) );
  AND2_X1 U12369 ( .A1(n14021), .A2(n6600), .ZN(n9814) );
  AOI21_X1 U12370 ( .B1(n14532), .B2(n6546), .A(n9814), .ZN(n9862) );
  NAND2_X1 U12371 ( .A1(n14532), .A2(n6600), .ZN(n9817) );
  NAND2_X1 U12372 ( .A1(n14021), .A2(n6546), .ZN(n9816) );
  NAND2_X1 U12373 ( .A1(n9817), .A2(n9816), .ZN(n9861) );
  NAND2_X1 U12374 ( .A1(n9862), .A2(n9861), .ZN(n9866) );
  NOR2_X1 U12375 ( .A1(n14268), .A2(n6546), .ZN(n9818) );
  AOI21_X1 U12376 ( .B1(n14538), .B2(n6546), .A(n9818), .ZN(n9858) );
  NAND2_X1 U12377 ( .A1(n14538), .A2(n9914), .ZN(n9820) );
  OR2_X1 U12378 ( .A1(n14268), .A2(n9914), .ZN(n9819) );
  NAND2_X1 U12379 ( .A1(n9820), .A2(n9819), .ZN(n9857) );
  NAND2_X1 U12380 ( .A1(n9858), .A2(n9857), .ZN(n9821) );
  NAND2_X1 U12381 ( .A1(n9866), .A2(n9821), .ZN(n9869) );
  NOR2_X1 U12382 ( .A1(n14287), .A2(n6546), .ZN(n9822) );
  AOI21_X1 U12383 ( .B1(n14543), .B2(n6546), .A(n9822), .ZN(n9868) );
  NAND2_X1 U12384 ( .A1(n14543), .A2(n9914), .ZN(n9824) );
  NAND2_X1 U12385 ( .A1(n14023), .A2(n6546), .ZN(n9823) );
  NAND2_X1 U12386 ( .A1(n9824), .A2(n9823), .ZN(n9867) );
  AND2_X1 U12387 ( .A1(n9868), .A2(n9867), .ZN(n9825) );
  AND2_X1 U12388 ( .A1(n14024), .A2(n9914), .ZN(n9826) );
  AOI21_X1 U12389 ( .B1(n14548), .B2(n6546), .A(n9826), .ZN(n9874) );
  NAND2_X1 U12390 ( .A1(n14548), .A2(n6550), .ZN(n9828) );
  NAND2_X1 U12391 ( .A1(n14024), .A2(n6546), .ZN(n9827) );
  NAND2_X1 U12392 ( .A1(n9828), .A2(n9827), .ZN(n9873) );
  AND2_X1 U12393 ( .A1(n9874), .A2(n9873), .ZN(n9829) );
  NOR2_X1 U12394 ( .A1(n14349), .A2(n6546), .ZN(n9830) );
  AOI21_X1 U12395 ( .B1(n14553), .B2(n6546), .A(n9830), .ZN(n9852) );
  NAND2_X1 U12396 ( .A1(n14553), .A2(n6550), .ZN(n9832) );
  NAND2_X1 U12397 ( .A1(n14025), .A2(n6546), .ZN(n9831) );
  NAND2_X1 U12398 ( .A1(n9832), .A2(n9831), .ZN(n9851) );
  AND2_X1 U12399 ( .A1(n9852), .A2(n9851), .ZN(n9833) );
  NOR2_X1 U12400 ( .A1(n14337), .A2(n6546), .ZN(n9834) );
  AOI21_X1 U12401 ( .B1(n14557), .B2(n6546), .A(n9834), .ZN(n9844) );
  NAND2_X1 U12402 ( .A1(n14557), .A2(n6600), .ZN(n9836) );
  NAND2_X1 U12403 ( .A1(n14026), .A2(n6546), .ZN(n9835) );
  NAND2_X1 U12404 ( .A1(n9836), .A2(n9835), .ZN(n9843) );
  AND2_X1 U12405 ( .A1(n9844), .A2(n9843), .ZN(n9837) );
  AND2_X1 U12406 ( .A1(n14027), .A2(n6595), .ZN(n9838) );
  AOI21_X1 U12407 ( .B1(n14562), .B2(n6546), .A(n9838), .ZN(n9847) );
  NAND2_X1 U12408 ( .A1(n14562), .A2(n9914), .ZN(n9840) );
  NAND2_X1 U12409 ( .A1(n14027), .A2(n6546), .ZN(n9839) );
  NAND2_X1 U12410 ( .A1(n9840), .A2(n9839), .ZN(n9846) );
  NAND2_X1 U12411 ( .A1(n9847), .A2(n9846), .ZN(n9841) );
  INV_X1 U12412 ( .A(n9846), .ZN(n9849) );
  INV_X1 U12413 ( .A(n9847), .ZN(n9848) );
  NAND3_X1 U12414 ( .A1(n9850), .A2(n9849), .A3(n9848), .ZN(n9882) );
  OR3_X1 U12415 ( .A1(n9853), .A2(n9852), .A3(n9851), .ZN(n9881) );
  AND2_X1 U12416 ( .A1(n14020), .A2(n6595), .ZN(n9854) );
  AOI21_X1 U12417 ( .B1(n14527), .B2(n6546), .A(n9854), .ZN(n9918) );
  NAND2_X1 U12418 ( .A1(n14527), .A2(n6600), .ZN(n9856) );
  NAND2_X1 U12419 ( .A1(n14020), .A2(n6546), .ZN(n9855) );
  NAND2_X1 U12420 ( .A1(n9856), .A2(n9855), .ZN(n9917) );
  INV_X1 U12421 ( .A(n9857), .ZN(n9860) );
  INV_X1 U12422 ( .A(n9858), .ZN(n9859) );
  AND2_X1 U12423 ( .A1(n9860), .A2(n9859), .ZN(n9865) );
  INV_X1 U12424 ( .A(n9861), .ZN(n9864) );
  INV_X1 U12425 ( .A(n9862), .ZN(n9863) );
  AOI22_X1 U12426 ( .A1(n9866), .A2(n9865), .B1(n9864), .B2(n9863), .ZN(n9871)
         );
  OR3_X1 U12427 ( .A1(n9869), .A2(n9868), .A3(n9867), .ZN(n9870) );
  OAI211_X1 U12428 ( .C1(n9918), .C2(n9917), .A(n9871), .B(n9870), .ZN(n9872)
         );
  INV_X1 U12429 ( .A(n9872), .ZN(n9880) );
  OR3_X1 U12430 ( .A1(n9875), .A2(n9874), .A3(n9873), .ZN(n9879) );
  NOR2_X1 U12431 ( .A1(n13801), .A2(n6595), .ZN(n9876) );
  AOI21_X1 U12432 ( .B1(n14519), .B2(n6600), .A(n9876), .ZN(n9920) );
  NAND2_X1 U12433 ( .A1(n14519), .A2(n6546), .ZN(n9878) );
  OR2_X1 U12434 ( .A1(n13801), .A2(n6546), .ZN(n9877) );
  NAND2_X1 U12435 ( .A1(n9878), .A2(n9877), .ZN(n9919) );
  NAND2_X1 U12436 ( .A1(n9920), .A2(n9919), .ZN(n9924) );
  INV_X1 U12437 ( .A(n9883), .ZN(n9884) );
  INV_X1 U12438 ( .A(SI_28_), .ZN(n12423) );
  NAND2_X1 U12439 ( .A1(n9884), .A2(n12423), .ZN(n9885) );
  INV_X1 U12440 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15427) );
  MUX2_X1 U12441 ( .A(n15427), .B(n12734), .S(n10581), .Z(n9888) );
  XNOR2_X1 U12442 ( .A(n9888), .B(SI_29_), .ZN(n9900) );
  NAND2_X1 U12443 ( .A1(n9901), .A2(n9900), .ZN(n9890) );
  INV_X1 U12444 ( .A(SI_29_), .ZN(n13722) );
  NAND2_X1 U12445 ( .A1(n9888), .A2(n13722), .ZN(n9889) );
  NAND2_X1 U12446 ( .A1(n9890), .A2(n9889), .ZN(n9936) );
  MUX2_X1 U12447 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10575), .Z(n9891) );
  NAND2_X1 U12448 ( .A1(n9891), .A2(SI_30_), .ZN(n9892) );
  OAI21_X1 U12449 ( .B1(SI_30_), .B2(n9891), .A(n9892), .ZN(n9935) );
  MUX2_X1 U12450 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10575), .Z(n9893) );
  XNOR2_X1 U12451 ( .A(n9893), .B(SI_31_), .ZN(n9894) );
  INV_X1 U12452 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14660) );
  OR2_X1 U12453 ( .A1(n9940), .A2(n14660), .ZN(n9896) );
  NAND2_X1 U12454 ( .A1(n6598), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U12455 ( .A1(n9945), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12456 ( .A1(n9946), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9897) );
  NAND3_X1 U12457 ( .A1(n9899), .A2(n9898), .A3(n9897), .ZN(n14015) );
  NAND2_X1 U12458 ( .A1(n12318), .A2(n9902), .ZN(n9904) );
  OR2_X1 U12459 ( .A1(n9940), .A2(n12734), .ZN(n9903) );
  NOR2_X1 U12460 ( .A1(n11213), .A2(n6546), .ZN(n9905) );
  AOI21_X1 U12461 ( .B1(n12722), .B2(n6546), .A(n9905), .ZN(n9956) );
  NAND2_X1 U12462 ( .A1(n12722), .A2(n9914), .ZN(n9907) );
  OR2_X1 U12463 ( .A1(n11213), .A2(n6595), .ZN(n9906) );
  NAND2_X1 U12464 ( .A1(n9907), .A2(n9906), .ZN(n9955) );
  NAND2_X1 U12465 ( .A1(n9956), .A2(n9955), .ZN(n9961) );
  NOR2_X1 U12466 ( .A1(n10551), .A2(n6546), .ZN(n9908) );
  AOI21_X1 U12467 ( .B1(n14218), .B2(n6546), .A(n9908), .ZN(n9959) );
  NAND2_X1 U12468 ( .A1(n14218), .A2(n9914), .ZN(n9910) );
  NAND2_X1 U12469 ( .A1(n14017), .A2(n6546), .ZN(n9909) );
  NAND2_X1 U12470 ( .A1(n9910), .A2(n9909), .ZN(n9958) );
  NAND2_X1 U12471 ( .A1(n9959), .A2(n9958), .ZN(n9911) );
  AND2_X1 U12472 ( .A1(n9961), .A2(n9911), .ZN(n9912) );
  AND2_X1 U12473 ( .A1(n14018), .A2(n6600), .ZN(n9913) );
  AOI21_X1 U12474 ( .B1(n14225), .B2(n6546), .A(n9913), .ZN(n9929) );
  NAND2_X1 U12475 ( .A1(n14225), .A2(n9914), .ZN(n9916) );
  NAND2_X1 U12476 ( .A1(n14018), .A2(n6546), .ZN(n9915) );
  NAND2_X1 U12477 ( .A1(n9916), .A2(n9915), .ZN(n9930) );
  NAND2_X1 U12478 ( .A1(n9929), .A2(n9930), .ZN(n9926) );
  AND2_X1 U12479 ( .A1(n9918), .A2(n9917), .ZN(n9923) );
  INV_X1 U12480 ( .A(n9919), .ZN(n9922) );
  INV_X1 U12481 ( .A(n9920), .ZN(n9921) );
  AOI22_X1 U12482 ( .A1(n9924), .A2(n9923), .B1(n9922), .B2(n9921), .ZN(n9925)
         );
  NAND2_X1 U12483 ( .A1(n9928), .A2(n9927), .ZN(n9967) );
  INV_X1 U12484 ( .A(n9929), .ZN(n9932) );
  INV_X1 U12485 ( .A(n9930), .ZN(n9931) );
  MUX2_X1 U12486 ( .A(n14015), .B(n6546), .S(n12395), .Z(n9934) );
  NAND2_X1 U12487 ( .A1(n6546), .A2(n14015), .ZN(n9972) );
  NAND2_X1 U12488 ( .A1(n9934), .A2(n9972), .ZN(n9957) );
  NAND2_X1 U12489 ( .A1(n9936), .A2(n9935), .ZN(n9937) );
  INV_X1 U12490 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12739) );
  OR2_X1 U12491 ( .A1(n9940), .A2(n12739), .ZN(n9941) );
  MUX2_X1 U12492 ( .A(n14015), .B(n9943), .S(n11605), .Z(n9944) );
  INV_X1 U12493 ( .A(n9944), .ZN(n9951) );
  NAND2_X1 U12494 ( .A1(n6597), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U12495 ( .A1(n9945), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12496 ( .A1(n9946), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9947) );
  NAND3_X1 U12497 ( .A1(n9949), .A2(n9948), .A3(n9947), .ZN(n14016) );
  INV_X1 U12498 ( .A(n14016), .ZN(n9950) );
  AOI21_X1 U12499 ( .B1(n9951), .B2(n10005), .A(n9950), .ZN(n9952) );
  AOI21_X1 U12500 ( .B1(n12705), .B2(n6546), .A(n9952), .ZN(n9969) );
  NAND2_X1 U12501 ( .A1(n12705), .A2(n6595), .ZN(n9954) );
  NAND2_X1 U12502 ( .A1(n6546), .A2(n14016), .ZN(n9953) );
  NAND2_X1 U12503 ( .A1(n9954), .A2(n9953), .ZN(n9968) );
  INV_X1 U12504 ( .A(n9958), .ZN(n9962) );
  INV_X1 U12505 ( .A(n9959), .ZN(n9960) );
  NAND4_X1 U12506 ( .A1(n9994), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9963)
         );
  NAND2_X1 U12507 ( .A1(n9967), .A2(n9966), .ZN(n9975) );
  NAND2_X1 U12508 ( .A1(n9969), .A2(n9968), .ZN(n9974) );
  INV_X1 U12509 ( .A(n14015), .ZN(n9970) );
  NAND3_X1 U12510 ( .A1(n12395), .A2(n9970), .A3(n6595), .ZN(n9971) );
  OAI21_X1 U12511 ( .B1(n12395), .B2(n9972), .A(n9971), .ZN(n9973) );
  MUX2_X1 U12512 ( .A(n11772), .B(n11880), .S(n6553), .Z(n9976) );
  OR2_X1 U12513 ( .A1(n10799), .A2(n6531), .ZN(n11540) );
  NOR3_X1 U12514 ( .A1(n6547), .A2(n9976), .A3(n11540), .ZN(n10000) );
  INV_X1 U12515 ( .A(n14316), .ZN(n14318) );
  XNOR2_X1 U12516 ( .A(n14562), .B(n14348), .ZN(n14376) );
  XNOR2_X1 U12517 ( .A(n14589), .B(n14474), .ZN(n14459) );
  OAI21_X1 U12518 ( .B1(n9670), .B2(n11301), .A(n11333), .ZN(n11304) );
  NAND2_X1 U12519 ( .A1(n11304), .A2(n6553), .ZN(n9978) );
  NOR2_X1 U12520 ( .A1(n9978), .A2(n9977), .ZN(n9979) );
  INV_X1 U12521 ( .A(n15762), .ZN(n15755) );
  NAND4_X1 U12522 ( .A1(n9979), .A2(n11376), .A3(n11326), .A4(n15755), .ZN(
        n9980) );
  NOR4_X1 U12523 ( .A1(n9980), .A2(n11733), .A3(n11552), .A4(n11513), .ZN(
        n9983) );
  INV_X1 U12524 ( .A(n11984), .ZN(n9981) );
  NOR2_X1 U12525 ( .A1(n14438), .A2(n9984), .ZN(n9985) );
  NOR2_X1 U12526 ( .A1(n14289), .A2(n9986), .ZN(n9988) );
  NOR2_X1 U12527 ( .A1(n9990), .A2(n9989), .ZN(n9992) );
  XNOR2_X1 U12528 ( .A(n12705), .B(n14016), .ZN(n9991) );
  AND4_X1 U12529 ( .A1(n10552), .A2(n9992), .A3(n10271), .A4(n9991), .ZN(n9993) );
  NAND2_X1 U12530 ( .A1(n9994), .A2(n9993), .ZN(n10003) );
  INV_X1 U12531 ( .A(n10003), .ZN(n9995) );
  NOR2_X1 U12532 ( .A1(n11540), .A2(n10005), .ZN(n10002) );
  INV_X1 U12533 ( .A(n12399), .ZN(n10802) );
  INV_X1 U12534 ( .A(n9996), .ZN(n10961) );
  NAND4_X1 U12535 ( .A1(n15781), .A2(n14496), .A3(n10802), .A4(n10961), .ZN(
        n9997) );
  OAI211_X1 U12536 ( .C1(n8917), .C2(n11540), .A(n9997), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9998) );
  NAND3_X1 U12537 ( .A1(n10003), .A2(n14214), .A3(n10002), .ZN(n10004) );
  OR2_X1 U12538 ( .A1(n10005), .A2(n11605), .ZN(n10540) );
  NAND2_X1 U12539 ( .A1(n6547), .A2(n10540), .ZN(n10007) );
  AOI21_X1 U12540 ( .B1(n10007), .B2(n10006), .A(n11540), .ZN(n10008) );
  INV_X1 U12541 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n10098) );
  INV_X1 U12542 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n13253) );
  NAND2_X1 U12543 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n13253), .ZN(n10036) );
  INV_X1 U12544 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U12545 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n10012), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n13253), .ZN(n10038) );
  INV_X1 U12546 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13230) );
  NOR2_X1 U12547 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n13230), .ZN(n10034) );
  INV_X1 U12548 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U12549 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .B1(n15510), .B2(n13230), .ZN(n10092) );
  INV_X1 U12550 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10975) );
  INV_X1 U12551 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10032) );
  INV_X1 U12552 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10825) );
  INV_X1 U12553 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10029) );
  XOR2_X1 U12554 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n10029), .Z(n10040) );
  INV_X1 U12555 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10853) );
  INV_X1 U12556 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15899) );
  INV_X1 U12557 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U12558 ( .A1(n11151), .A2(n10014), .ZN(n10015) );
  XNOR2_X1 U12559 ( .A(n10016), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n10047) );
  INV_X1 U12560 ( .A(n10047), .ZN(n10018) );
  AOI21_X1 U12561 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  INV_X1 U12562 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U12563 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n10840), .ZN(n10022) );
  OAI21_X1 U12564 ( .B1(P3_ADDR_REG_6__SCAN_IN), .B2(n10840), .A(n10022), .ZN(
        n10065) );
  NOR2_X1 U12565 ( .A1(n10066), .A2(n10065), .ZN(n10023) );
  INV_X1 U12566 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11309) );
  NAND2_X1 U12567 ( .A1(n10024), .A2(n11309), .ZN(n10026) );
  INV_X1 U12568 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10481) );
  XNOR2_X1 U12569 ( .A(n15899), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n10041) );
  INV_X1 U12570 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11456) );
  XNOR2_X1 U12571 ( .A(n11456), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U12572 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n10825), .ZN(n10030) );
  OAI21_X1 U12573 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n10825), .A(n10030), 
        .ZN(n10083) );
  INV_X1 U12574 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n13177) );
  XOR2_X1 U12575 ( .A(n13177), .B(n10032), .Z(n10085) );
  XOR2_X1 U12576 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n10975), .Z(n10088) );
  NAND2_X1 U12577 ( .A1(n10038), .A2(n10037), .ZN(n10035) );
  XNOR2_X1 U12578 ( .A(n10038), .B(n10037), .ZN(n15480) );
  XNOR2_X1 U12579 ( .A(n10040), .B(n10039), .ZN(n10080) );
  XOR2_X1 U12580 ( .A(n10042), .B(n10041), .Z(n10073) );
  XNOR2_X1 U12581 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n10043) );
  XNOR2_X1 U12582 ( .A(n10046), .B(n10045), .ZN(n10061) );
  XNOR2_X1 U12583 ( .A(n10048), .B(n10047), .ZN(n10049) );
  XOR2_X1 U12584 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n10050), .Z(n15966) );
  XOR2_X1 U12585 ( .A(n10052), .B(n10051), .Z(n15440) );
  OAI21_X1 U12586 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10053), .A(n10054), .ZN(
        n15961) );
  NAND2_X1 U12587 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15961), .ZN(n15971) );
  NOR2_X1 U12588 ( .A1(n15971), .A2(n15970), .ZN(n15969) );
  NOR2_X1 U12589 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NAND2_X1 U12590 ( .A1(n15440), .A2(n15439), .ZN(n15438) );
  NAND2_X1 U12591 ( .A1(n15966), .A2(n15967), .ZN(n15965) );
  INV_X1 U12592 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15959) );
  NAND2_X1 U12593 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  XOR2_X1 U12594 ( .A(n10066), .B(n10065), .Z(n15445) );
  NOR2_X1 U12595 ( .A1(n10067), .A2(n10064), .ZN(n10068) );
  INV_X1 U12596 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10390) );
  XNOR2_X1 U12597 ( .A(n10070), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15964) );
  INV_X1 U12598 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14900) );
  XOR2_X1 U12599 ( .A(n14900), .B(n10069), .Z(n15963) );
  NAND2_X1 U12600 ( .A1(n15964), .A2(n15963), .ZN(n15962) );
  NAND2_X1 U12601 ( .A1(n10070), .A2(n10390), .ZN(n10071) );
  NAND2_X1 U12602 ( .A1(n15448), .A2(n15447), .ZN(n10072) );
  NOR2_X1 U12603 ( .A1(n15448), .A2(n15447), .ZN(n15446) );
  AOI21_X2 U12604 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n10072), .A(n15446), .ZN(
        n10074) );
  XNOR2_X1 U12605 ( .A(n10074), .B(n10073), .ZN(n15450) );
  INV_X1 U12606 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15730) );
  XOR2_X1 U12607 ( .A(n10077), .B(n10076), .Z(n15453) );
  INV_X1 U12608 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15459) );
  NAND2_X1 U12609 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  XOR2_X1 U12610 ( .A(n10084), .B(n10083), .Z(n15463) );
  XOR2_X1 U12611 ( .A(n10086), .B(n10085), .Z(n15466) );
  INV_X1 U12612 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10087) );
  XNOR2_X1 U12613 ( .A(n10089), .B(n10088), .ZN(n15471) );
  NOR2_X1 U12614 ( .A1(n15470), .A2(n15471), .ZN(n10090) );
  NAND2_X1 U12615 ( .A1(n15471), .A2(n15470), .ZN(n15469) );
  XNOR2_X1 U12616 ( .A(n10092), .B(n10091), .ZN(n10093) );
  NOR2_X2 U12617 ( .A1(n10094), .A2(n10093), .ZN(n15474) );
  INV_X1 U12618 ( .A(n15474), .ZN(n15475) );
  INV_X1 U12619 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15477) );
  NAND2_X1 U12620 ( .A1(n10094), .A2(n10093), .ZN(n15476) );
  NAND2_X1 U12621 ( .A1(n15477), .A2(n15476), .ZN(n15473) );
  INV_X1 U12622 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10341) );
  INV_X1 U12623 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10360) );
  NOR2_X1 U12624 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n10360), .ZN(n10096) );
  AOI21_X1 U12625 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n10360), .A(n10096), 
        .ZN(n10248) );
  NAND2_X1 U12626 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n10097), .ZN(n10101) );
  NAND2_X1 U12627 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  NAND2_X1 U12628 ( .A1(n10101), .A2(n10100), .ZN(n10247) );
  XNOR2_X1 U12629 ( .A(n10248), .B(n10247), .ZN(n10244) );
  INV_X1 U12630 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U12631 ( .A1(n15564), .A2(n12490), .ZN(n12501) );
  NAND2_X1 U12632 ( .A1(n12495), .A2(n12497), .ZN(n12649) );
  NAND2_X1 U12633 ( .A1(n12501), .A2(n12649), .ZN(n10105) );
  NAND2_X1 U12634 ( .A1(n15566), .A2(n6593), .ZN(n12648) );
  NAND2_X1 U12635 ( .A1(n10105), .A2(n12648), .ZN(n11487) );
  NAND2_X1 U12636 ( .A1(n15647), .A2(n10156), .ZN(n12515) );
  NAND2_X1 U12637 ( .A1(n15629), .A2(n15557), .ZN(n12514) );
  AND2_X1 U12638 ( .A1(n12515), .A2(n12514), .ZN(n12511) );
  NAND2_X1 U12639 ( .A1(n15547), .A2(n12511), .ZN(n10106) );
  NAND2_X1 U12640 ( .A1(n10106), .A2(n12514), .ZN(n11884) );
  NAND2_X1 U12641 ( .A1(n15487), .A2(n12520), .ZN(n10107) );
  NAND2_X1 U12642 ( .A1(n15659), .A2(n15666), .ZN(n10109) );
  NAND2_X1 U12643 ( .A1(n12338), .A2(n12530), .ZN(n10110) );
  XNOR2_X1 U12644 ( .A(n12538), .B(n11652), .ZN(n15512) );
  INV_X1 U12645 ( .A(n15512), .ZN(n10111) );
  NAND2_X1 U12646 ( .A1(n12538), .A2(n11652), .ZN(n10112) );
  XNOR2_X1 U12647 ( .A(n12548), .B(n15514), .ZN(n12658) );
  INV_X1 U12648 ( .A(n12658), .ZN(n10115) );
  OR2_X1 U12649 ( .A1(n12548), .A2(n15385), .ZN(n10114) );
  OAI21_X1 U12650 ( .B1(n11610), .B2(n10115), .A(n10114), .ZN(n11909) );
  INV_X1 U12651 ( .A(n15384), .ZN(n14820) );
  NAND2_X1 U12652 ( .A1(n15389), .A2(n15377), .ZN(n12050) );
  OAI21_X1 U12653 ( .B1(n15378), .B2(n14820), .A(n12050), .ZN(n10116) );
  INV_X1 U12654 ( .A(n10116), .ZN(n10117) );
  NAND2_X1 U12655 ( .A1(n11909), .A2(n10117), .ZN(n10122) );
  OAI21_X1 U12656 ( .B1(n15389), .B2(n15377), .A(n15384), .ZN(n10120) );
  NAND2_X1 U12657 ( .A1(n14820), .A2(n14821), .ZN(n10118) );
  NOR2_X1 U12658 ( .A1(n15389), .A2(n10118), .ZN(n10119) );
  AOI21_X1 U12659 ( .B1(n15378), .B2(n10120), .A(n10119), .ZN(n10121) );
  NAND2_X1 U12660 ( .A1(n10122), .A2(n10121), .ZN(n12053) );
  XNOR2_X1 U12661 ( .A(n15372), .B(n12565), .ZN(n12662) );
  INV_X1 U12662 ( .A(n12662), .ZN(n12052) );
  XNOR2_X1 U12663 ( .A(n12098), .B(n15353), .ZN(n12569) );
  AND2_X1 U12664 ( .A1(n12052), .A2(n12569), .ZN(n10123) );
  NAND2_X1 U12665 ( .A1(n12053), .A2(n10123), .ZN(n12091) );
  INV_X1 U12666 ( .A(n12569), .ZN(n10124) );
  OR2_X1 U12667 ( .A1(n15372), .A2(n12565), .ZN(n12088) );
  OR2_X1 U12668 ( .A1(n15352), .A2(n14673), .ZN(n15202) );
  OR2_X1 U12669 ( .A1(n12098), .A2(n12217), .ZN(n12222) );
  NAND2_X1 U12670 ( .A1(n15202), .A2(n12222), .ZN(n12578) );
  INV_X1 U12671 ( .A(n12578), .ZN(n10125) );
  AND2_X1 U12672 ( .A1(n12090), .A2(n10125), .ZN(n10126) );
  NAND2_X1 U12673 ( .A1(n15352), .A2(n14673), .ZN(n12580) );
  XNOR2_X1 U12674 ( .A(n12585), .B(n15344), .ZN(n12664) );
  INV_X1 U12675 ( .A(n12664), .ZN(n12274) );
  INV_X1 U12676 ( .A(n15321), .ZN(n14819) );
  XNOR2_X1 U12677 ( .A(n15183), .B(n14819), .ZN(n15170) );
  INV_X1 U12678 ( .A(n15170), .ZN(n15172) );
  XOR2_X1 U12679 ( .A(n15329), .B(n15325), .Z(n15156) );
  NOR2_X1 U12680 ( .A1(n15325), .A2(n15181), .ZN(n12597) );
  NAND2_X1 U12681 ( .A1(n15315), .A2(n15305), .ZN(n15096) );
  XNOR2_X1 U12682 ( .A(n10129), .B(n15306), .ZN(n15108) );
  NOR2_X1 U12683 ( .A1(n15315), .A2(n15305), .ZN(n10131) );
  OAI21_X1 U12684 ( .B1(n10131), .B2(n15314), .A(n15131), .ZN(n10130) );
  INV_X1 U12685 ( .A(n15306), .ZN(n15129) );
  XNOR2_X1 U12686 ( .A(n15062), .B(n15045), .ZN(n15055) );
  NAND2_X1 U12687 ( .A1(n15062), .A2(n15273), .ZN(n10137) );
  NAND2_X1 U12688 ( .A1(n15276), .A2(n14688), .ZN(n10138) );
  XNOR2_X1 U12689 ( .A(n15034), .B(n15274), .ZN(n12669) );
  NAND2_X1 U12690 ( .A1(n15261), .A2(n15028), .ZN(n10140) );
  NAND2_X1 U12691 ( .A1(n15255), .A2(n15242), .ZN(n10142) );
  XNOR2_X2 U12692 ( .A(n15244), .B(n15223), .ZN(n14983) );
  NOR2_X1 U12693 ( .A1(n15224), .A2(n15223), .ZN(n15227) );
  AOI21_X1 U12694 ( .B1(n15232), .B2(n14983), .A(n15227), .ZN(n10145) );
  NAND2_X1 U12695 ( .A1(n12318), .A2(n6552), .ZN(n10144) );
  NAND2_X1 U12696 ( .A1(n6604), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n10143) );
  INV_X1 U12697 ( .A(n15228), .ZN(n15222) );
  XNOR2_X1 U12698 ( .A(n10145), .B(n15222), .ZN(n10228) );
  NAND2_X1 U12699 ( .A1(n12698), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10930) );
  NOR2_X1 U12700 ( .A1(n10930), .A2(n10146), .ZN(n11007) );
  INV_X1 U12701 ( .A(n11006), .ZN(n10147) );
  NAND2_X1 U12702 ( .A1(n15395), .A2(n10148), .ZN(n10219) );
  INV_X1 U12703 ( .A(n11004), .ZN(n10149) );
  NAND2_X1 U12704 ( .A1(n6608), .A2(n10213), .ZN(n10151) );
  INV_X1 U12705 ( .A(n7760), .ZN(n12646) );
  OR2_X1 U12706 ( .A1(n12646), .A2(n12430), .ZN(n10150) );
  OR2_X1 U12707 ( .A1(n15564), .A2(n12492), .ZN(n15577) );
  NAND2_X1 U12708 ( .A1(n15566), .A2(n12497), .ZN(n10152) );
  NAND2_X1 U12709 ( .A1(n15577), .A2(n10152), .ZN(n15579) );
  NAND2_X1 U12710 ( .A1(n10153), .A2(n6593), .ZN(n15576) );
  NAND2_X1 U12711 ( .A1(n15579), .A2(n15576), .ZN(n11486) );
  NAND2_X1 U12712 ( .A1(n15486), .A2(n12508), .ZN(n10154) );
  NAND2_X1 U12713 ( .A1(n15629), .A2(n10156), .ZN(n10157) );
  NAND2_X1 U12714 ( .A1(n15487), .A2(n12519), .ZN(n10158) );
  NAND2_X1 U12715 ( .A1(n10159), .A2(n10158), .ZN(n15527) );
  XNOR2_X1 U12716 ( .A(n15666), .B(n12526), .ZN(n12651) );
  NAND2_X1 U12717 ( .A1(n11506), .A2(n15659), .ZN(n11498) );
  OR2_X1 U12718 ( .A1(n15531), .A2(n12530), .ZN(n10160) );
  AND2_X1 U12719 ( .A1(n11498), .A2(n10160), .ZN(n10162) );
  INV_X1 U12720 ( .A(n10160), .ZN(n10161) );
  XNOR2_X2 U12721 ( .A(n12338), .B(n12530), .ZN(n12655) );
  OR2_X1 U12722 ( .A1(n12538), .A2(n15667), .ZN(n10163) );
  XNOR2_X1 U12723 ( .A(n15389), .B(n14821), .ZN(n12657) );
  OR2_X1 U12724 ( .A1(n15389), .A2(n14821), .ZN(n10166) );
  OR2_X1 U12725 ( .A1(n15378), .A2(n15384), .ZN(n10167) );
  OR2_X1 U12726 ( .A1(n12098), .A2(n15353), .ZN(n10168) );
  OR2_X1 U12727 ( .A1(n15352), .A2(n15363), .ZN(n15189) );
  NAND2_X1 U12728 ( .A1(n15189), .A2(n15354), .ZN(n10169) );
  NAND2_X1 U12729 ( .A1(n10169), .A2(n15346), .ZN(n10171) );
  OR2_X1 U12730 ( .A1(n15189), .A2(n15354), .ZN(n10170) );
  NAND2_X1 U12731 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  INV_X1 U12732 ( .A(n10172), .ZN(n12276) );
  OR2_X1 U12733 ( .A1(n15346), .A2(n14766), .ZN(n10173) );
  NAND2_X1 U12734 ( .A1(n15202), .A2(n12580), .ZN(n12663) );
  NAND2_X1 U12735 ( .A1(n10173), .A2(n12663), .ZN(n12277) );
  AND2_X1 U12736 ( .A1(n12276), .A2(n12277), .ZN(n10174) );
  NOR2_X1 U12737 ( .A1(n10174), .A2(n12664), .ZN(n10175) );
  OR2_X1 U12738 ( .A1(n12585), .A2(n15344), .ZN(n10177) );
  OR2_X1 U12739 ( .A1(n15332), .A2(n15321), .ZN(n10179) );
  AND2_X1 U12740 ( .A1(n15332), .A2(n15321), .ZN(n10178) );
  NAND2_X1 U12741 ( .A1(n12592), .A2(n15181), .ZN(n10180) );
  NAND2_X1 U12742 ( .A1(n15153), .A2(n10180), .ZN(n10182) );
  OR2_X1 U12743 ( .A1(n12592), .A2(n15181), .ZN(n10181) );
  NAND2_X1 U12744 ( .A1(n10182), .A2(n10181), .ZN(n15115) );
  INV_X1 U12745 ( .A(n15115), .ZN(n10184) );
  OR2_X1 U12746 ( .A1(n15315), .A2(n15322), .ZN(n15116) );
  INV_X1 U12747 ( .A(n15314), .ZN(n15145) );
  NAND2_X1 U12748 ( .A1(n15131), .A2(n15145), .ZN(n10183) );
  AOI21_X1 U12749 ( .B1(n15131), .B2(n15145), .A(n15305), .ZN(n10185) );
  AOI22_X1 U12750 ( .A1(n10185), .A2(n15315), .B1(n15309), .B2(n15314), .ZN(
        n10186) );
  NAND2_X1 U12751 ( .A1(n10129), .A2(n15306), .ZN(n10189) );
  NAND2_X1 U12752 ( .A1(n15076), .A2(n15089), .ZN(n10193) );
  INV_X1 U12753 ( .A(n10193), .ZN(n10190) );
  AND2_X1 U12754 ( .A1(n15082), .A2(n10192), .ZN(n10191) );
  INV_X1 U12755 ( .A(n10192), .ZN(n10195) );
  OR2_X1 U12756 ( .A1(n15091), .A2(n14818), .ZN(n15067) );
  AND2_X1 U12757 ( .A1(n15067), .A2(n10193), .ZN(n10194) );
  NOR2_X1 U12758 ( .A1(n15062), .A2(n15045), .ZN(n10198) );
  NAND2_X1 U12759 ( .A1(n15267), .A2(n15274), .ZN(n10199) );
  NAND2_X1 U12760 ( .A1(n14752), .A2(n14688), .ZN(n15024) );
  NOR2_X1 U12761 ( .A1(n14752), .A2(n14688), .ZN(n10200) );
  AOI22_X1 U12762 ( .A1(n10200), .A2(n10199), .B1(n15034), .B2(n15015), .ZN(
        n10201) );
  OR2_X1 U12763 ( .A1(n15261), .A2(n15251), .ZN(n10202) );
  NAND2_X1 U12764 ( .A1(n15003), .A2(n15242), .ZN(n10204) );
  XOR2_X1 U12765 ( .A(n15228), .B(n10206), .Z(n15239) );
  AOI21_X1 U12766 ( .B1(n12491), .B2(n6608), .A(n10213), .ZN(n10207) );
  NAND2_X1 U12767 ( .A1(n10208), .A2(n10207), .ZN(n15137) );
  OR2_X1 U12768 ( .A1(n10209), .A2(n15207), .ZN(n15149) );
  AND2_X1 U12769 ( .A1(n15137), .A2(n15149), .ZN(n10210) );
  NAND2_X1 U12770 ( .A1(n15554), .A2(n10156), .ZN(n15555) );
  INV_X1 U12771 ( .A(n15555), .ZN(n10211) );
  INV_X1 U12772 ( .A(n12530), .ZN(n11507) );
  INV_X1 U12773 ( .A(n12538), .ZN(n15683) );
  INV_X1 U12774 ( .A(n12585), .ZN(n15339) );
  NOR2_X4 U12775 ( .A1(n15083), .A2(n7418), .ZN(n15073) );
  OR2_X2 U12776 ( .A1(n14984), .A2(n12448), .ZN(n14976) );
  AOI21_X1 U12777 ( .B1(n14984), .B2(n12448), .A(n15574), .ZN(n10212) );
  INV_X1 U12778 ( .A(n15430), .ZN(n10710) );
  OR2_X1 U12779 ( .A1(n15584), .A2(n15630), .ZN(n15162) );
  NAND2_X1 U12780 ( .A1(n15584), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12781 ( .A1(n12696), .A2(n10214), .ZN(n10215) );
  NOR2_X1 U12782 ( .A1(n15628), .A2(n10215), .ZN(n14972) );
  INV_X1 U12783 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U12784 ( .A1(n10216), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12785 ( .A1(n8442), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n10217) );
  OAI211_X1 U12786 ( .C1(n8216), .C2(n10504), .A(n10218), .B(n10217), .ZN(
        n14817) );
  NAND2_X1 U12787 ( .A1(n14972), .A2(n14817), .ZN(n15233) );
  OR2_X1 U12788 ( .A1(n10219), .A2(n15233), .ZN(n10220) );
  OAI211_X1 U12789 ( .C1(n10222), .C2(n15549), .A(n10221), .B(n10220), .ZN(
        n10223) );
  AOI21_X1 U12790 ( .B1(n15223), .B2(n15192), .A(n10223), .ZN(n10224) );
  OAI21_X1 U12791 ( .B1(n15237), .B2(n15552), .A(n10224), .ZN(n10225) );
  INV_X1 U12792 ( .A(n11658), .ZN(n13714) );
  NOR2_X1 U12793 ( .A1(n11406), .A2(n10229), .ZN(n10230) );
  NAND2_X1 U12794 ( .A1(n13714), .A2(n10230), .ZN(n11688) );
  INV_X1 U12795 ( .A(n11688), .ZN(n11704) );
  NAND2_X1 U12796 ( .A1(n12801), .A2(n12790), .ZN(n11657) );
  NOR2_X1 U12797 ( .A1(n10231), .A2(n11657), .ZN(n11689) );
  INV_X1 U12798 ( .A(n11689), .ZN(n11683) );
  NAND2_X1 U12799 ( .A1(n9602), .A2(n12937), .ZN(n11048) );
  OAI21_X1 U12800 ( .B1(n11683), .B2(n11702), .A(n11698), .ZN(n10232) );
  NAND2_X1 U12801 ( .A1(n11704), .A2(n10232), .ZN(n10237) );
  AND2_X1 U12802 ( .A1(n11406), .A2(n10233), .ZN(n10234) );
  NAND2_X1 U12803 ( .A1(n11658), .A2(n10234), .ZN(n11697) );
  INV_X1 U12804 ( .A(n11697), .ZN(n10235) );
  INV_X1 U12805 ( .A(n11702), .ZN(n11685) );
  NAND3_X1 U12806 ( .A1(n10235), .A2(n11685), .A3(n11687), .ZN(n10236) );
  INV_X2 U12807 ( .A(n15941), .ZN(n15943) );
  NAND2_X1 U12808 ( .A1(n10238), .A2(n15943), .ZN(n10243) );
  INV_X1 U12809 ( .A(n9664), .ZN(n10240) );
  INV_X1 U12810 ( .A(n10241), .ZN(n10242) );
  NAND2_X1 U12811 ( .A1(n10243), .A2(n10242), .ZN(P3_U3456) );
  NAND2_X1 U12812 ( .A1(n10248), .A2(n10247), .ZN(n10249) );
  OAI21_X1 U12813 ( .B1(n10360), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n10249), 
        .ZN(n10251) );
  XNOR2_X1 U12814 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10250) );
  XNOR2_X1 U12815 ( .A(n10251), .B(n10250), .ZN(n10253) );
  XNOR2_X1 U12816 ( .A(n10255), .B(n10254), .ZN(SUB_1596_U4) );
  INV_X1 U12817 ( .A(n10256), .ZN(n10259) );
  INV_X1 U12818 ( .A(n10257), .ZN(n10258) );
  NAND2_X1 U12819 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  NAND2_X1 U12820 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  NAND2_X1 U12821 ( .A1(n10262), .A2(n15491), .ZN(n10268) );
  AOI22_X1 U12822 ( .A1(n14999), .A2(n14813), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10263) );
  OAI21_X1 U12823 ( .B1(n15252), .B2(n14808), .A(n10263), .ZN(n10264) );
  AOI21_X1 U12824 ( .B1(n14806), .B2(n15028), .A(n10264), .ZN(n10265) );
  INV_X1 U12825 ( .A(n10266), .ZN(n10267) );
  NAND2_X1 U12826 ( .A1(n10268), .A2(n10267), .ZN(P1_U3214) );
  XNOR2_X1 U12827 ( .A(n10270), .B(n10271), .ZN(n10272) );
  OAI22_X1 U12828 ( .A1(n10551), .A2(n14473), .B1(n13801), .B2(n14471), .ZN(
        n13810) );
  INV_X1 U12829 ( .A(n14236), .ZN(n10273) );
  AOI21_X1 U12830 ( .B1(n10273), .B2(n14225), .A(n14482), .ZN(n10274) );
  NAND2_X1 U12831 ( .A1(n10275), .A2(n10274), .ZN(n14228) );
  NAND2_X1 U12832 ( .A1(n14225), .A2(n15835), .ZN(n10276) );
  NAND2_X1 U12833 ( .A1(n10277), .A2(n7631), .ZN(n14610) );
  NAND2_X1 U12834 ( .A1(n14610), .A2(n15864), .ZN(n10279) );
  NAND2_X1 U12835 ( .A1(n10279), .A2(n10278), .ZN(n10518) );
  NOR4_X1 U12836 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), .A3(SI_13_), .A4(SI_11_), .ZN(n10291) );
  INV_X1 U12837 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13667) );
  NAND4_X1 U12838 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_REG0_REG_0__SCAN_IN), 
        .A3(n11484), .A4(n13667), .ZN(n10281) );
  NAND4_X1 U12839 ( .A1(P3_D_REG_0__SCAN_IN), .A2(SI_25_), .A3(
        P1_REG2_REG_24__SCAN_IN), .A4(P2_REG2_REG_4__SCAN_IN), .ZN(n10280) );
  NOR2_X1 U12840 ( .A1(n10281), .A2(n10280), .ZN(n10285) );
  NAND2_X1 U12841 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10806) );
  NOR2_X1 U12842 ( .A1(n11349), .A2(n10806), .ZN(n10284) );
  INV_X1 U12843 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n14088) );
  NOR4_X1 U12844 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(P2_REG2_REG_24__SCAN_IN), 
        .A3(n14204), .A4(n14088), .ZN(n10283) );
  NOR4_X1 U12845 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .A3(P2_REG0_REG_4__SCAN_IN), .A4(n11199), .ZN(n10282) );
  NAND4_X1 U12846 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  NOR2_X1 U12847 ( .A1(n14687), .A2(n10286), .ZN(n10290) );
  INV_X1 U12848 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10738) );
  NAND4_X1 U12849 ( .A1(n10738), .A2(P1_REG0_REG_28__SCAN_IN), .A3(SI_2_), 
        .A4(P2_DATAO_REG_9__SCAN_IN), .ZN(n10288) );
  NAND4_X1 U12850 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .A3(P3_IR_REG_28__SCAN_IN), .A4(P3_REG3_REG_22__SCAN_IN), .ZN(n10287)
         );
  NOR2_X1 U12851 ( .A1(n10288), .A2(n10287), .ZN(n10289) );
  NAND4_X1 U12852 ( .A1(n10291), .A2(P1_ADDR_REG_3__SCAN_IN), .A3(n10290), 
        .A4(n10289), .ZN(n10295) );
  NAND4_X1 U12853 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .A3(P2_ADDR_REG_7__SCAN_IN), .A4(P2_ADDR_REG_5__SCAN_IN), .ZN(n10293)
         );
  OR4_X1 U12854 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(P3_ADDR_REG_8__SCAN_IN), 
        .A3(P1_ADDR_REG_8__SCAN_IN), .A4(P2_ADDR_REG_17__SCAN_IN), .ZN(n10292)
         );
  NOR4_X1 U12855 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10303) );
  INV_X1 U12856 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11783) );
  INV_X1 U12857 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U12858 ( .A1(n10330), .A2(n11783), .A3(n10362), .A4(
        P3_REG3_REG_3__SCAN_IN), .ZN(n10301) );
  INV_X1 U12859 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10297) );
  INV_X1 U12860 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10296) );
  NAND4_X1 U12861 ( .A1(n10297), .A2(n10296), .A3(P2_REG2_REG_7__SCAN_IN), 
        .A4(P2_REG0_REG_8__SCAN_IN), .ZN(n10300) );
  INV_X1 U12862 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U12863 ( .A1(n10904), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_18__SCAN_IN), .A4(P2_REG1_REG_21__SCAN_IN), .ZN(n10299) );
  INV_X1 U12864 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n12727) );
  OR4_X1 U12865 ( .A1(P3_DATAO_REG_18__SCAN_IN), .A2(n12727), .A3(keyinput74), 
        .A4(P3_DATAO_REG_13__SCAN_IN), .ZN(n10298) );
  NOR4_X1 U12866 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10302) );
  NAND4_X1 U12867 ( .A1(n10303), .A2(n10302), .A3(P2_D_REG_27__SCAN_IN), .A4(
        P2_D_REG_20__SCAN_IN), .ZN(n10321) );
  NOR4_X1 U12868 ( .A1(n11979), .A2(n13625), .A3(n10472), .A4(n10475), .ZN(
        n10307) );
  NOR4_X1 U12869 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(P3_DATAO_REG_20__SCAN_IN), .A4(n10974), .ZN(n10306) );
  INV_X1 U12870 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10778) );
  INV_X1 U12871 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10781) );
  NOR4_X1 U12872 ( .A1(P3_REG0_REG_7__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(n10778), .A4(n10781), .ZN(n10305) );
  NOR4_X1 U12873 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P2_DATAO_REG_27__SCAN_IN), 
        .A3(P3_REG0_REG_24__SCAN_IN), .A4(P2_REG3_REG_0__SCAN_IN), .ZN(n10304)
         );
  AND4_X1 U12874 ( .A1(n10307), .A2(n10306), .A3(n10305), .A4(n10304), .ZN(
        n10311) );
  NOR4_X1 U12875 ( .A1(P3_D_REG_14__SCAN_IN), .A2(SI_10_), .A3(
        P1_IR_REG_29__SCAN_IN), .A4(P3_DATAO_REG_29__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U12876 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), 
        .A3(P2_REG3_REG_8__SCAN_IN), .A4(P2_REG1_REG_22__SCAN_IN), .ZN(n10308)
         );
  NOR3_X1 U12877 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P3_DATAO_REG_6__SCAN_IN), 
        .A3(n10308), .ZN(n10309) );
  NAND3_X1 U12878 ( .A1(n10311), .A2(n10310), .A3(n10309), .ZN(n10320) );
  INV_X1 U12879 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10312) );
  NOR4_X1 U12880 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_REG0_REG_28__SCAN_IN), 
        .A3(P2_REG1_REG_12__SCAN_IN), .A4(n10312), .ZN(n10316) );
  NOR4_X1 U12881 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .A3(P1_B_REG_SCAN_IN), .A4(P1_ADDR_REG_18__SCAN_IN), .ZN(n10315) );
  NOR4_X1 U12882 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P1_REG2_REG_22__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(n13253), .ZN(n10314) );
  INV_X1 U12883 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15776) );
  INV_X1 U12884 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15772) );
  NOR4_X1 U12885 ( .A1(SI_8_), .A2(P1_REG3_REG_1__SCAN_IN), .A3(n15776), .A4(
        n15772), .ZN(n10313) );
  NAND4_X1 U12886 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10319) );
  NOR4_X1 U12887 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(P2_REG3_REG_20__SCAN_IN), .A4(P2_ADDR_REG_15__SCAN_IN), .ZN(n10317) );
  NAND3_X1 U12888 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(P3_DATAO_REG_25__SCAN_IN), .A3(n10317), .ZN(n10318) );
  NOR4_X1 U12889 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10327) );
  NAND4_X1 U12890 ( .A1(P3_REG0_REG_18__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), 
        .A3(P1_REG2_REG_13__SCAN_IN), .A4(P1_REG1_REG_3__SCAN_IN), .ZN(n10325)
         );
  INV_X1 U12891 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15856) );
  NAND4_X1 U12892 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P3_REG2_REG_1__SCAN_IN), 
        .A3(P1_D_REG_31__SCAN_IN), .A4(n15856), .ZN(n10324) );
  INV_X1 U12893 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U12894 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), 
        .A3(P1_REG0_REG_30__SCAN_IN), .A4(n11548), .ZN(n10323) );
  INV_X1 U12895 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n10496) );
  INV_X1 U12896 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15799) );
  NAND4_X1 U12897 ( .A1(n10496), .A2(n11251), .A3(n13830), .A4(n15799), .ZN(
        n10322) );
  NOR4_X1 U12898 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  AOI21_X1 U12899 ( .B1(n10327), .B2(n10326), .A(keyinput82), .ZN(n10516) );
  INV_X1 U12900 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15441) );
  INV_X1 U12901 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n10666) );
  INV_X1 U12902 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15773) );
  AOI22_X1 U12903 ( .A1(n10666), .A2(keyinput59), .B1(n15773), .B2(keyinput86), 
        .ZN(n10328) );
  OAI221_X1 U12904 ( .B1(n10666), .B2(keyinput59), .C1(n15773), .C2(keyinput86), .A(n10328), .ZN(n10335) );
  AOI22_X1 U12905 ( .A1(n10331), .A2(keyinput8), .B1(n10330), .B2(keyinput69), 
        .ZN(n10329) );
  OAI221_X1 U12906 ( .B1(n10331), .B2(keyinput8), .C1(n10330), .C2(keyinput69), 
        .A(n10329), .ZN(n10334) );
  XNOR2_X1 U12907 ( .A(keyinput33), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n10332)
         );
  OAI21_X1 U12908 ( .B1(n15441), .B2(keyinput82), .A(n10332), .ZN(n10333) );
  NOR3_X1 U12909 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10353) );
  INV_X1 U12910 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U12911 ( .A1(n14703), .A2(keyinput112), .B1(keyinput9), .B2(n11714), 
        .ZN(n10336) );
  OAI221_X1 U12912 ( .B1(n14703), .B2(keyinput112), .C1(n11714), .C2(keyinput9), .A(n10336), .ZN(n10339) );
  INV_X1 U12913 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U12914 ( .A1(n10825), .A2(keyinput115), .B1(keyinput30), .B2(n10670), .ZN(n10337) );
  OAI221_X1 U12915 ( .B1(n10825), .B2(keyinput115), .C1(n10670), .C2(
        keyinput30), .A(n10337), .ZN(n10338) );
  NOR2_X1 U12916 ( .A1(n10339), .A2(n10338), .ZN(n10352) );
  INV_X1 U12917 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U12918 ( .A1(n10342), .A2(keyinput62), .B1(keyinput56), .B2(n10341), 
        .ZN(n10340) );
  OAI221_X1 U12919 ( .B1(n10342), .B2(keyinput62), .C1(n10341), .C2(keyinput56), .A(n10340), .ZN(n10345) );
  INV_X1 U12920 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U12921 ( .A1(n9082), .A2(keyinput31), .B1(keyinput49), .B2(n15849), 
        .ZN(n10343) );
  OAI221_X1 U12922 ( .B1(n9082), .B2(keyinput31), .C1(n15849), .C2(keyinput49), 
        .A(n10343), .ZN(n10344) );
  NOR2_X1 U12923 ( .A1(n10345), .A2(n10344), .ZN(n10351) );
  INV_X1 U12924 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n12156) );
  INV_X1 U12925 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U12926 ( .A1(n12156), .A2(keyinput95), .B1(n10759), .B2(keyinput40), 
        .ZN(n10346) );
  OAI221_X1 U12927 ( .B1(n12156), .B2(keyinput95), .C1(n10759), .C2(keyinput40), .A(n10346), .ZN(n10349) );
  INV_X1 U12928 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13668) );
  INV_X1 U12929 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U12930 ( .A1(n13668), .A2(keyinput3), .B1(n10775), .B2(keyinput99), 
        .ZN(n10347) );
  OAI221_X1 U12931 ( .B1(n13668), .B2(keyinput3), .C1(n10775), .C2(keyinput99), 
        .A(n10347), .ZN(n10348) );
  NOR2_X1 U12932 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  AND4_X1 U12933 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10374) );
  INV_X1 U12934 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U12935 ( .A1(n15772), .A2(keyinput72), .B1(n10355), .B2(keyinput57), 
        .ZN(n10354) );
  OAI221_X1 U12936 ( .B1(n15772), .B2(keyinput72), .C1(n10355), .C2(keyinput57), .A(n10354), .ZN(n10358) );
  AOI22_X1 U12937 ( .A1(n15593), .A2(keyinput123), .B1(keyinput88), .B2(n12727), .ZN(n10356) );
  OAI221_X1 U12938 ( .B1(n15593), .B2(keyinput123), .C1(n12727), .C2(
        keyinput88), .A(n10356), .ZN(n10357) );
  NOR2_X1 U12939 ( .A1(n10358), .A2(n10357), .ZN(n10373) );
  INV_X1 U12940 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U12941 ( .A1(n10360), .A2(keyinput87), .B1(n12036), .B2(keyinput106), .ZN(n10359) );
  OAI221_X1 U12942 ( .B1(n10360), .B2(keyinput87), .C1(n12036), .C2(
        keyinput106), .A(n10359), .ZN(n10364) );
  INV_X1 U12943 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15774) );
  AOI22_X1 U12944 ( .A1(n15774), .A2(keyinput29), .B1(n10362), .B2(keyinput77), 
        .ZN(n10361) );
  OAI221_X1 U12945 ( .B1(n15774), .B2(keyinput29), .C1(n10362), .C2(keyinput77), .A(n10361), .ZN(n10363) );
  NOR2_X1 U12946 ( .A1(n10364), .A2(n10363), .ZN(n10372) );
  INV_X1 U12947 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U12948 ( .A1(n14544), .A2(keyinput85), .B1(n15603), .B2(keyinput121), .ZN(n10365) );
  OAI221_X1 U12949 ( .B1(n14544), .B2(keyinput85), .C1(n15603), .C2(
        keyinput121), .A(n10365), .ZN(n10370) );
  INV_X1 U12950 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n14116) );
  INV_X1 U12951 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U12952 ( .A1(n14116), .A2(keyinput6), .B1(n10367), .B2(keyinput127), 
        .ZN(n10366) );
  OAI221_X1 U12953 ( .B1(n14116), .B2(keyinput6), .C1(n10367), .C2(keyinput127), .A(n10366), .ZN(n10369) );
  INV_X1 U12954 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15586) );
  XNOR2_X1 U12955 ( .A(n15586), .B(keyinput120), .ZN(n10368) );
  NOR3_X1 U12956 ( .A1(n10370), .A2(n10369), .A3(n10368), .ZN(n10371) );
  NAND4_X1 U12957 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10468) );
  INV_X1 U12958 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U12959 ( .A1(n15477), .A2(keyinput25), .B1(n10855), .B2(keyinput26), 
        .ZN(n10375) );
  OAI221_X1 U12960 ( .B1(n15477), .B2(keyinput25), .C1(n10855), .C2(keyinput26), .A(n10375), .ZN(n10383) );
  INV_X1 U12961 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U12962 ( .A1(n10378), .A2(keyinput124), .B1(keyinput71), .B2(n10377), .ZN(n10376) );
  OAI221_X1 U12963 ( .B1(n10378), .B2(keyinput124), .C1(n10377), .C2(
        keyinput71), .A(n10376), .ZN(n10382) );
  AOI22_X1 U12964 ( .A1(n10380), .A2(keyinput42), .B1(keyinput32), .B2(n13949), 
        .ZN(n10379) );
  OAI221_X1 U12965 ( .B1(n10380), .B2(keyinput42), .C1(n13949), .C2(keyinput32), .A(n10379), .ZN(n10381) );
  NOR3_X1 U12966 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n10400) );
  AOI22_X1 U12967 ( .A1(n14687), .A2(keyinput90), .B1(keyinput102), .B2(n10904), .ZN(n10384) );
  OAI221_X1 U12968 ( .B1(n14687), .B2(keyinput90), .C1(n10904), .C2(
        keyinput102), .A(n10384), .ZN(n10387) );
  AOI22_X1 U12969 ( .A1(n10781), .A2(keyinput50), .B1(keyinput11), .B2(n10778), 
        .ZN(n10385) );
  OAI221_X1 U12970 ( .B1(n10781), .B2(keyinput50), .C1(n10778), .C2(keyinput11), .A(n10385), .ZN(n10386) );
  NOR2_X1 U12971 ( .A1(n10387), .A2(n10386), .ZN(n10399) );
  AOI22_X1 U12972 ( .A1(n11349), .A2(keyinput114), .B1(keyinput83), .B2(n11281), .ZN(n10388) );
  OAI221_X1 U12973 ( .B1(n11349), .B2(keyinput114), .C1(n11281), .C2(
        keyinput83), .A(n10388), .ZN(n10392) );
  INV_X1 U12974 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14822) );
  AOI22_X1 U12975 ( .A1(n14822), .A2(keyinput79), .B1(keyinput28), .B2(n10390), 
        .ZN(n10389) );
  OAI221_X1 U12976 ( .B1(n14822), .B2(keyinput79), .C1(n10390), .C2(keyinput28), .A(n10389), .ZN(n10391) );
  NOR2_X1 U12977 ( .A1(n10392), .A2(n10391), .ZN(n10398) );
  INV_X1 U12978 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U12979 ( .A1(n8322), .A2(keyinput13), .B1(keyinput61), .B2(n14073), 
        .ZN(n10393) );
  OAI221_X1 U12980 ( .B1(n8322), .B2(keyinput13), .C1(n14073), .C2(keyinput61), 
        .A(n10393), .ZN(n10396) );
  AOI22_X1 U12981 ( .A1(n15776), .A2(keyinput19), .B1(keyinput73), .B2(n10840), 
        .ZN(n10394) );
  OAI221_X1 U12982 ( .B1(n15776), .B2(keyinput19), .C1(n10840), .C2(keyinput73), .A(n10394), .ZN(n10395) );
  NOR2_X1 U12983 ( .A1(n10396), .A2(n10395), .ZN(n10397) );
  NAND4_X1 U12984 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10467) );
  AOI22_X1 U12985 ( .A1(n14271), .A2(keyinput68), .B1(keyinput64), .B2(n14088), 
        .ZN(n10401) );
  OAI221_X1 U12986 ( .B1(n14271), .B2(keyinput68), .C1(n14088), .C2(keyinput64), .A(n10401), .ZN(n10409) );
  INV_X1 U12987 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U12988 ( .A1(n11296), .A2(keyinput80), .B1(n12302), .B2(keyinput45), 
        .ZN(n10402) );
  OAI221_X1 U12989 ( .B1(n11296), .B2(keyinput80), .C1(n12302), .C2(keyinput45), .A(n10402), .ZN(n10408) );
  XNOR2_X1 U12990 ( .A(SI_25_), .B(keyinput119), .ZN(n10406) );
  XNOR2_X1 U12991 ( .A(SI_10_), .B(keyinput98), .ZN(n10405) );
  XNOR2_X1 U12992 ( .A(SI_20_), .B(keyinput5), .ZN(n10404) );
  XNOR2_X1 U12993 ( .A(SI_8_), .B(keyinput96), .ZN(n10403) );
  NAND4_X1 U12994 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10407) );
  NOR3_X1 U12995 ( .A1(n10409), .A2(n10408), .A3(n10407), .ZN(n10465) );
  XNOR2_X1 U12996 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput39), .ZN(n10413) );
  XNOR2_X1 U12997 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput0), .ZN(n10412) );
  XNOR2_X1 U12998 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput54), .ZN(n10411) );
  XNOR2_X1 U12999 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput27), .ZN(n10410) );
  NAND4_X1 U13000 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10419) );
  XNOR2_X1 U13001 ( .A(P1_REG2_REG_22__SCAN_IN), .B(keyinput104), .ZN(n10417)
         );
  XNOR2_X1 U13002 ( .A(P1_B_REG_SCAN_IN), .B(keyinput34), .ZN(n10416) );
  XNOR2_X1 U13003 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput4), .ZN(n10415) );
  XNOR2_X1 U13004 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput92), .ZN(n10414) );
  NAND4_X1 U13005 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  NOR2_X1 U13006 ( .A1(n10419), .A2(n10418), .ZN(n10431) );
  XNOR2_X1 U13007 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput101), .ZN(n10423) );
  XNOR2_X1 U13008 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput35), .ZN(n10422) );
  XNOR2_X1 U13009 ( .A(P2_REG1_REG_12__SCAN_IN), .B(keyinput66), .ZN(n10421)
         );
  XNOR2_X1 U13010 ( .A(P3_REG0_REG_30__SCAN_IN), .B(keyinput23), .ZN(n10420)
         );
  NAND4_X1 U13011 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10429) );
  XNOR2_X1 U13012 ( .A(P3_D_REG_0__SCAN_IN), .B(keyinput20), .ZN(n10427) );
  XNOR2_X1 U13013 ( .A(P3_REG2_REG_1__SCAN_IN), .B(keyinput14), .ZN(n10426) );
  XNOR2_X1 U13014 ( .A(SI_13_), .B(keyinput107), .ZN(n10425) );
  XNOR2_X1 U13015 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput111), .ZN(n10424) );
  NAND4_X1 U13016 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10428) );
  NOR2_X1 U13017 ( .A1(n10429), .A2(n10428), .ZN(n10430) );
  AND2_X1 U13018 ( .A1(n10431), .A2(n10430), .ZN(n10464) );
  XNOR2_X1 U13019 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput91), .ZN(n10435) );
  XNOR2_X1 U13020 ( .A(SI_2_), .B(keyinput100), .ZN(n10434) );
  XNOR2_X1 U13021 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput84), .ZN(n10433)
         );
  XNOR2_X1 U13022 ( .A(P3_REG2_REG_2__SCAN_IN), .B(keyinput89), .ZN(n10432) );
  NAND4_X1 U13023 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10441) );
  XNOR2_X1 U13024 ( .A(SI_11_), .B(keyinput47), .ZN(n10439) );
  XNOR2_X1 U13025 ( .A(keyinput74), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10438) );
  XNOR2_X1 U13026 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput43), .ZN(n10437) );
  XNOR2_X1 U13027 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput24), .ZN(n10436)
         );
  NAND4_X1 U13028 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10440) );
  NOR2_X1 U13029 ( .A1(n10441), .A2(n10440), .ZN(n10453) );
  XNOR2_X1 U13030 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput37), .ZN(n10445) );
  XNOR2_X1 U13031 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput17), .ZN(n10444) );
  XNOR2_X1 U13032 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput18), .ZN(n10443)
         );
  XNOR2_X1 U13033 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput2), .ZN(n10442)
         );
  NAND4_X1 U13034 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10451) );
  XNOR2_X1 U13035 ( .A(keyinput117), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10449)
         );
  XNOR2_X1 U13036 ( .A(P2_REG1_REG_15__SCAN_IN), .B(keyinput15), .ZN(n10448)
         );
  XNOR2_X1 U13037 ( .A(keyinput109), .B(P3_REG0_REG_7__SCAN_IN), .ZN(n10447)
         );
  XNOR2_X1 U13038 ( .A(keyinput110), .B(P3_DATAO_REG_18__SCAN_IN), .ZN(n10446)
         );
  NAND4_X1 U13039 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10450) );
  NOR2_X1 U13040 ( .A1(n10451), .A2(n10450), .ZN(n10452) );
  AND2_X1 U13041 ( .A1(n10453), .A2(n10452), .ZN(n10463) );
  AOI22_X1 U13042 ( .A1(n15602), .A2(keyinput16), .B1(keyinput113), .B2(n13253), .ZN(n10454) );
  OAI221_X1 U13043 ( .B1(n15602), .B2(keyinput16), .C1(n13253), .C2(
        keyinput113), .A(n10454), .ZN(n10461) );
  XNOR2_X1 U13044 ( .A(n15594), .B(keyinput78), .ZN(n10460) );
  XNOR2_X1 U13045 ( .A(keyinput81), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U13046 ( .A(keyinput97), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n10457)
         );
  XNOR2_X1 U13047 ( .A(keyinput38), .B(P2_REG1_REG_0__SCAN_IN), .ZN(n10456) );
  XNOR2_X1 U13048 ( .A(keyinput67), .B(P2_REG0_REG_0__SCAN_IN), .ZN(n10455) );
  NAND4_X1 U13049 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10459) );
  NOR3_X1 U13050 ( .A1(n10461), .A2(n10460), .A3(n10459), .ZN(n10462) );
  NAND4_X1 U13051 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10466) );
  NOR3_X1 U13052 ( .A1(n10468), .A2(n10467), .A3(n10466), .ZN(n10514) );
  AOI22_X1 U13053 ( .A1(n13625), .A2(keyinput75), .B1(n11979), .B2(keyinput70), 
        .ZN(n10469) );
  OAI221_X1 U13054 ( .B1(n13625), .B2(keyinput75), .C1(n11979), .C2(keyinput70), .A(n10469), .ZN(n10479) );
  INV_X1 U13055 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U13056 ( .A1(n11035), .A2(keyinput93), .B1(n10974), .B2(keyinput52), 
        .ZN(n10470) );
  OAI221_X1 U13057 ( .B1(n11035), .B2(keyinput93), .C1(n10974), .C2(keyinput52), .A(n10470), .ZN(n10478) );
  AOI22_X1 U13058 ( .A1(n10472), .A2(keyinput7), .B1(n15595), .B2(keyinput108), 
        .ZN(n10471) );
  OAI221_X1 U13059 ( .B1(n10472), .B2(keyinput7), .C1(n15595), .C2(keyinput108), .A(n10471), .ZN(n10477) );
  AOI22_X1 U13060 ( .A1(n10475), .A2(keyinput22), .B1(n10474), .B2(keyinput12), 
        .ZN(n10473) );
  OAI221_X1 U13061 ( .B1(n10475), .B2(keyinput22), .C1(n10474), .C2(keyinput12), .A(n10473), .ZN(n10476) );
  NOR4_X1 U13062 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10491) );
  AOI22_X1 U13063 ( .A1(n10481), .A2(keyinput21), .B1(n11201), .B2(keyinput105), .ZN(n10480) );
  OAI221_X1 U13064 ( .B1(n10481), .B2(keyinput21), .C1(n11201), .C2(
        keyinput105), .A(n10480), .ZN(n10489) );
  INV_X1 U13065 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13066 ( .A1(n10668), .A2(keyinput63), .B1(n11199), .B2(keyinput36), 
        .ZN(n10482) );
  OAI221_X1 U13067 ( .B1(n10668), .B2(keyinput63), .C1(n11199), .C2(keyinput36), .A(n10482), .ZN(n10488) );
  INV_X1 U13068 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15815) );
  AOI22_X1 U13069 ( .A1(n15815), .A2(keyinput46), .B1(n10484), .B2(keyinput65), 
        .ZN(n10483) );
  OAI221_X1 U13070 ( .B1(n15815), .B2(keyinput46), .C1(n10484), .C2(keyinput65), .A(n10483), .ZN(n10487) );
  INV_X1 U13071 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U13072 ( .A1(n11427), .A2(keyinput125), .B1(keyinput48), .B2(n14204), .ZN(n10485) );
  OAI221_X1 U13073 ( .B1(n11427), .B2(keyinput125), .C1(n14204), .C2(
        keyinput48), .A(n10485), .ZN(n10486) );
  NOR4_X1 U13074 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10490) );
  AND2_X1 U13075 ( .A1(n10491), .A2(n10490), .ZN(n10513) );
  AOI22_X1 U13076 ( .A1(n14900), .A2(keyinput103), .B1(n15856), .B2(keyinput94), .ZN(n10492) );
  OAI221_X1 U13077 ( .B1(n14900), .B2(keyinput103), .C1(n15856), .C2(
        keyinput94), .A(n10492), .ZN(n10500) );
  INV_X1 U13078 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15605) );
  AOI22_X1 U13079 ( .A1(n15605), .A2(keyinput1), .B1(n13698), .B2(keyinput44), 
        .ZN(n10493) );
  OAI221_X1 U13080 ( .B1(n15605), .B2(keyinput1), .C1(n13698), .C2(keyinput44), 
        .A(n10493), .ZN(n10499) );
  INV_X1 U13081 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15703) );
  INV_X1 U13082 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13083 ( .A1(n15703), .A2(keyinput55), .B1(n10980), .B2(keyinput10), 
        .ZN(n10494) );
  OAI221_X1 U13084 ( .B1(n15703), .B2(keyinput55), .C1(n10980), .C2(keyinput10), .A(n10494), .ZN(n10498) );
  AOI22_X1 U13085 ( .A1(n10496), .A2(keyinput58), .B1(keyinput60), .B2(n13830), 
        .ZN(n10495) );
  OAI221_X1 U13086 ( .B1(n10496), .B2(keyinput58), .C1(n13830), .C2(keyinput60), .A(n10495), .ZN(n10497) );
  NOR4_X1 U13087 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10512) );
  AOI22_X1 U13088 ( .A1(n11251), .A2(keyinput118), .B1(keyinput116), .B2(
        n15799), .ZN(n10501) );
  OAI221_X1 U13089 ( .B1(n11251), .B2(keyinput118), .C1(n15799), .C2(
        keyinput116), .A(n10501), .ZN(n10510) );
  INV_X1 U13090 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15775) );
  INV_X1 U13091 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U13092 ( .A1(n15775), .A2(keyinput122), .B1(n12408), .B2(keyinput76), .ZN(n10502) );
  OAI221_X1 U13093 ( .B1(n15775), .B2(keyinput122), .C1(n12408), .C2(
        keyinput76), .A(n10502), .ZN(n10509) );
  AOI22_X1 U13094 ( .A1(n10504), .A2(keyinput51), .B1(n11548), .B2(keyinput41), 
        .ZN(n10503) );
  OAI221_X1 U13095 ( .B1(n10504), .B2(keyinput51), .C1(n11548), .C2(keyinput41), .A(n10503), .ZN(n10508) );
  INV_X1 U13096 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10827) );
  INV_X1 U13097 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13098 ( .A1(n10827), .A2(keyinput126), .B1(keyinput53), .B2(n10506), .ZN(n10505) );
  OAI221_X1 U13099 ( .B1(n10827), .B2(keyinput126), .C1(n10506), .C2(
        keyinput53), .A(n10505), .ZN(n10507) );
  NOR4_X1 U13100 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10511) );
  AND4_X1 U13101 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n10515) );
  OAI21_X1 U13102 ( .B1(n10516), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n10515), .ZN(
        n10517) );
  XNOR2_X1 U13103 ( .A(n10518), .B(n10517), .ZN(P2_U3526) );
  INV_X1 U13104 ( .A(n10524), .ZN(n10523) );
  NOR3_X1 U13105 ( .A1(n14222), .A2(n10546), .A3(n10523), .ZN(n10531) );
  INV_X1 U13106 ( .A(n14222), .ZN(n10529) );
  INV_X1 U13107 ( .A(n10521), .ZN(n10520) );
  NAND2_X1 U13108 ( .A1(n10546), .A2(n6670), .ZN(n10528) );
  OAI211_X1 U13109 ( .C1(n10523), .C2(n10522), .A(n10552), .B(n10521), .ZN(
        n10526) );
  NAND2_X1 U13110 ( .A1(n10546), .A2(n10524), .ZN(n10525) );
  NAND2_X1 U13111 ( .A1(n10526), .A2(n10525), .ZN(n10527) );
  INV_X1 U13112 ( .A(n10532), .ZN(n10534) );
  INV_X1 U13113 ( .A(n10941), .ZN(n10533) );
  NAND4_X1 U13114 ( .A1(n10534), .A2(n10533), .A3(n15781), .A4(n15780), .ZN(
        n10539) );
  NAND2_X2 U13115 ( .A1(n10539), .A2(n14406), .ZN(n14499) );
  NOR2_X1 U13116 ( .A1(n6547), .A2(n10991), .ZN(n10535) );
  NAND2_X1 U13117 ( .A1(n14499), .A2(n10535), .ZN(n14488) );
  INV_X1 U13118 ( .A(n8920), .ZN(n15818) );
  NAND2_X1 U13119 ( .A1(n14499), .A2(n15818), .ZN(n10536) );
  NOR2_X1 U13120 ( .A1(n10539), .A2(n14214), .ZN(n14457) );
  INV_X1 U13121 ( .A(n14507), .ZN(n15767) );
  NOR2_X1 U13122 ( .A1(n8917), .A2(n10540), .ZN(n10951) );
  INV_X1 U13123 ( .A(n10951), .ZN(n10541) );
  INV_X1 U13124 ( .A(n10542), .ZN(n10543) );
  INV_X1 U13125 ( .A(n14406), .ZN(n15760) );
  AOI22_X1 U13126 ( .A1(n10543), .A2(n15760), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14484), .ZN(n10544) );
  OAI21_X1 U13127 ( .B1(n7524), .B2(n14486), .A(n10544), .ZN(n10545) );
  AOI21_X1 U13128 ( .B1(n12721), .B2(n15767), .A(n10545), .ZN(n10560) );
  NAND3_X1 U13129 ( .A1(n10548), .A2(n10546), .A3(n15757), .ZN(n10558) );
  OAI211_X1 U13130 ( .C1(n10551), .C2(n14218), .A(n10552), .B(n15757), .ZN(
        n10547) );
  NOR2_X1 U13131 ( .A1(n10548), .A2(n10547), .ZN(n10557) );
  INV_X1 U13132 ( .A(P2_B_REG_SCAN_IN), .ZN(n10549) );
  NOR2_X1 U13133 ( .A1(n12399), .A2(n10549), .ZN(n10550) );
  NOR2_X1 U13134 ( .A1(n14473), .A2(n10550), .ZN(n12394) );
  NOR2_X1 U13135 ( .A1(n10551), .A2(n14471), .ZN(n10554) );
  NOR4_X1 U13136 ( .A1(n10552), .A2(n10551), .A3(n14461), .A4(n14218), .ZN(
        n10553) );
  AOI211_X1 U13137 ( .C1(n12394), .C2(n14016), .A(n10554), .B(n10553), .ZN(
        n10555) );
  NAND2_X1 U13138 ( .A1(n12726), .A2(n14499), .ZN(n10559) );
  OAI21_X1 U13139 ( .B1(n12733), .B2(n14465), .A(n10561), .ZN(P2_U3236) );
  INV_X1 U13140 ( .A(n10799), .ZN(n10562) );
  NOR2_X1 U13141 ( .A1(n10563), .A2(n10562), .ZN(n10801) );
  AND2_X1 U13142 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10801), .ZN(P2_U3947) );
  INV_X1 U13143 ( .A(n11692), .ZN(n10564) );
  AND2_X2 U13144 ( .A1(n10564), .A2(n13713), .ZN(P3_U3897) );
  NOR2_X1 U13145 ( .A1(n10565), .A2(P1_U3086), .ZN(n10566) );
  AND2_X2 U13146 ( .A1(n10566), .A2(n10636), .ZN(P1_U4016) );
  INV_X1 U13147 ( .A(n11085), .ZN(n11194) );
  NAND2_X1 U13148 ( .A1(n10581), .A2(P3_U3151), .ZN(n13731) );
  INV_X1 U13149 ( .A(SI_1_), .ZN(n10570) );
  NAND2_X1 U13150 ( .A1(n10567), .A2(P3_U3151), .ZN(n13729) );
  INV_X1 U13151 ( .A(n10568), .ZN(n10569) );
  OAI222_X1 U13152 ( .A1(P3_U3151), .A2(n11194), .B1(n13731), .B2(n10570), 
        .C1(n13729), .C2(n10569), .ZN(P3_U3294) );
  INV_X1 U13153 ( .A(n10571), .ZN(n10574) );
  INV_X1 U13154 ( .A(n13729), .ZN(n11851) );
  INV_X1 U13155 ( .A(n11851), .ZN(n13725) );
  MUX2_X1 U13156 ( .A(n10572), .B(n13152), .S(P3_STATE_REG_SCAN_IN), .Z(n10573) );
  OAI21_X1 U13157 ( .B1(n10574), .B2(n13725), .A(n10573), .ZN(P3_U3295) );
  AND2_X1 U13158 ( .A1(n10567), .A2(P1_U3086), .ZN(n11545) );
  INV_X1 U13159 ( .A(n10576), .ZN(n10584) );
  OAI222_X1 U13160 ( .A1(n15433), .A2(n10577), .B1(n6554), .B2(n10584), .C1(
        P1_U3086), .C2(n14859), .ZN(P1_U3352) );
  INV_X1 U13161 ( .A(n14825), .ZN(n10579) );
  OAI222_X1 U13162 ( .A1(n10579), .A2(P1_U3086), .B1(n6554), .B2(n10615), .C1(
        n10578), .C2(n15433), .ZN(P1_U3354) );
  INV_X1 U13163 ( .A(n10580), .ZN(n10628) );
  NAND2_X1 U13164 ( .A1(n10567), .A2(n6531), .ZN(n12702) );
  INV_X1 U13165 ( .A(n12702), .ZN(n14666) );
  AOI22_X1 U13166 ( .A1(n14102), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n14666), .ZN(n10582) );
  OAI21_X1 U13167 ( .B1(n10628), .B2(n11978), .A(n10582), .ZN(P2_U3321) );
  INV_X1 U13168 ( .A(n14666), .ZN(n14659) );
  INV_X1 U13169 ( .A(n14058), .ZN(n10583) );
  OAI222_X1 U13170 ( .A1(n14659), .A2(n10585), .B1(n11978), .B2(n10584), .C1(
        P2_U3088), .C2(n10583), .ZN(P2_U3324) );
  INV_X1 U13171 ( .A(n10586), .ZN(n10624) );
  INV_X1 U13172 ( .A(n14087), .ZN(n10587) );
  OAI222_X1 U13173 ( .A1(n14659), .A2(n10588), .B1(n11978), .B2(n10624), .C1(
        P2_U3088), .C2(n10587), .ZN(P2_U3322) );
  INV_X1 U13174 ( .A(n10589), .ZN(n10622) );
  INV_X1 U13175 ( .A(n14115), .ZN(n10590) );
  OAI222_X1 U13176 ( .A1(n14659), .A2(n10591), .B1(n11978), .B2(n10622), .C1(
        P2_U3088), .C2(n10590), .ZN(P2_U3320) );
  INV_X1 U13177 ( .A(n10592), .ZN(n10642) );
  OAI222_X1 U13178 ( .A1(n14659), .A2(n10593), .B1(n11978), .B2(n10642), .C1(
        P2_U3088), .C2(n8551), .ZN(P2_U3325) );
  INV_X1 U13179 ( .A(n10594), .ZN(n10626) );
  INV_X1 U13180 ( .A(n14072), .ZN(n10595) );
  OAI222_X1 U13181 ( .A1(n14659), .A2(n10596), .B1(n11978), .B2(n10626), .C1(
        P2_U3088), .C2(n10595), .ZN(P2_U3323) );
  INV_X1 U13182 ( .A(n13731), .ZN(n13718) );
  INV_X1 U13183 ( .A(n13718), .ZN(n11854) );
  INV_X1 U13184 ( .A(SI_8_), .ZN(n10597) );
  INV_X1 U13185 ( .A(n11471), .ZN(n11457) );
  OAI222_X1 U13186 ( .A1(n13729), .A2(n10598), .B1(n11854), .B2(n10597), .C1(
        n11457), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U13187 ( .A(SI_6_), .ZN(n10600) );
  INV_X1 U13188 ( .A(n11283), .ZN(n10599) );
  OAI222_X1 U13189 ( .A1(n13725), .A2(n10601), .B1(n11854), .B2(n10600), .C1(
        n10599), .C2(P3_U3151), .ZN(P3_U3289) );
  OAI222_X1 U13190 ( .A1(n13729), .A2(n10603), .B1(n11854), .B2(n10602), .C1(
        n11266), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U13191 ( .A1(n13729), .A2(n10605), .B1(n11854), .B2(n10604), .C1(
        n11472), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U13192 ( .A(SI_4_), .ZN(n10606) );
  OAI222_X1 U13193 ( .A1(n13729), .A2(n10607), .B1(n11854), .B2(n10606), .C1(
        n11094), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U13194 ( .A(SI_5_), .ZN(n10608) );
  OAI222_X1 U13195 ( .A1(n13729), .A2(n10609), .B1(n11854), .B2(n10608), .C1(
        n11248), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U13196 ( .A(SI_3_), .ZN(n10610) );
  OAI222_X1 U13197 ( .A1(n13729), .A2(n10611), .B1(n11854), .B2(n10610), .C1(
        n11152), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U13198 ( .A(SI_2_), .ZN(n10612) );
  OAI222_X1 U13199 ( .A1(n11088), .A2(P3_U3151), .B1(n13729), .B2(n10613), 
        .C1(n10612), .C2(n11854), .ZN(P3_U3293) );
  OAI222_X1 U13200 ( .A1(n10867), .A2(P2_U3088), .B1(n11978), .B2(n10615), 
        .C1(n10614), .C2(n12702), .ZN(P2_U3326) );
  NAND2_X1 U13201 ( .A1(n11410), .A2(n13713), .ZN(n10616) );
  OAI21_X1 U13202 ( .B1(n13713), .B2(n10617), .A(n10616), .ZN(P3_U3377) );
  INV_X1 U13203 ( .A(n10618), .ZN(n10620) );
  OAI222_X1 U13204 ( .A1(n15433), .A2(n10619), .B1(n6554), .B2(n10620), .C1(
        P1_U3086), .C2(n10793), .ZN(P1_U3347) );
  OAI222_X1 U13205 ( .A1(n12702), .A2(n10621), .B1(n11978), .B2(n10620), .C1(
        P2_U3088), .C2(n14129), .ZN(P2_U3319) );
  OAI222_X1 U13206 ( .A1(n15433), .A2(n10623), .B1(n6554), .B2(n10622), .C1(
        P1_U3086), .C2(n14908), .ZN(P1_U3348) );
  OAI222_X1 U13207 ( .A1(n15433), .A2(n10625), .B1(n6554), .B2(n10624), .C1(
        P1_U3086), .C2(n14886), .ZN(P1_U3350) );
  OAI222_X1 U13208 ( .A1(n15433), .A2(n10627), .B1(n6554), .B2(n10626), .C1(
        P1_U3086), .C2(n14873), .ZN(P1_U3351) );
  OAI222_X1 U13209 ( .A1(n15433), .A2(n10629), .B1(n6554), .B2(n10628), .C1(
        P1_U3086), .C2(n10847), .ZN(P1_U3349) );
  OAI222_X1 U13210 ( .A1(n13729), .A2(n10631), .B1(n11854), .B2(n10630), .C1(
        n11756), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U13211 ( .A(n10632), .ZN(n10641) );
  OAI222_X1 U13212 ( .A1(n14659), .A2(n10633), .B1(n11978), .B2(n10641), .C1(
        P2_U3088), .C2(n15718), .ZN(P2_U3318) );
  INV_X1 U13213 ( .A(n10645), .ZN(n10635) );
  INV_X1 U13214 ( .A(n10636), .ZN(n10634) );
  NAND2_X1 U13215 ( .A1(n10634), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12701) );
  NAND2_X1 U13216 ( .A1(n10635), .A2(n12701), .ZN(n10673) );
  NAND2_X1 U13217 ( .A1(n10637), .A2(n10636), .ZN(n10639) );
  NAND2_X1 U13218 ( .A1(n10639), .A2(n10638), .ZN(n10671) );
  NAND2_X1 U13219 ( .A1(n10673), .A2(n10671), .ZN(n15509) );
  INV_X1 U13220 ( .A(n15509), .ZN(n14938) );
  NOR2_X1 U13221 ( .A1(n14938), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13222 ( .A(n14924), .ZN(n10702) );
  INV_X1 U13223 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10640) );
  OAI222_X1 U13224 ( .A1(n10702), .A2(P1_U3086), .B1(n6554), .B2(n10641), .C1(
        n10640), .C2(n15433), .ZN(P1_U3346) );
  INV_X1 U13225 ( .A(n14844), .ZN(n10643) );
  OAI222_X1 U13226 ( .A1(n10643), .A2(P1_U3086), .B1(n6554), .B2(n10642), .C1(
        n7665), .C2(n15433), .ZN(P1_U3353) );
  AND2_X2 U13227 ( .A1(n10645), .A2(n10644), .ZN(n15616) );
  INV_X1 U13228 ( .A(n10646), .ZN(n12162) );
  NAND2_X1 U13229 ( .A1(n10647), .A2(n12162), .ZN(n10649) );
  OAI22_X1 U13230 ( .A1(n15616), .A2(P1_D_REG_0__SCAN_IN), .B1(n11904), .B2(
        n10649), .ZN(n10648) );
  INV_X1 U13231 ( .A(n10648), .ZN(P1_U3445) );
  OAI22_X1 U13232 ( .A1(n15616), .A2(P1_D_REG_1__SCAN_IN), .B1(n12026), .B2(
        n10649), .ZN(n10650) );
  INV_X1 U13233 ( .A(n10650), .ZN(P1_U3446) );
  OAI222_X1 U13234 ( .A1(n13729), .A2(n10652), .B1(n11854), .B2(n10651), .C1(
        n11765), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U13235 ( .A(n10653), .ZN(n10655) );
  INV_X1 U13236 ( .A(n10908), .ZN(n14143) );
  OAI222_X1 U13237 ( .A1(n14659), .A2(n10654), .B1(n11978), .B2(n10655), .C1(
        P2_U3088), .C2(n14143), .ZN(P2_U3317) );
  INV_X1 U13238 ( .A(n10854), .ZN(n10861) );
  OAI222_X1 U13239 ( .A1(n15433), .A2(n10656), .B1(n6554), .B2(n10655), .C1(
        P1_U3086), .C2(n10861), .ZN(P1_U3345) );
  INV_X1 U13240 ( .A(n10657), .ZN(n10660) );
  INV_X1 U13241 ( .A(n11352), .ZN(n10658) );
  OAI222_X1 U13242 ( .A1(n14659), .A2(n10659), .B1(n11978), .B2(n10660), .C1(
        P2_U3088), .C2(n10658), .ZN(P2_U3316) );
  INV_X1 U13243 ( .A(n10818), .ZN(n10747) );
  OAI222_X1 U13244 ( .A1(n15433), .A2(n10661), .B1(n6554), .B2(n10660), .C1(
        P1_U3086), .C2(n10747), .ZN(P1_U3344) );
  INV_X1 U13245 ( .A(n10662), .ZN(n10664) );
  INV_X1 U13246 ( .A(n11938), .ZN(n13167) );
  OAI222_X1 U13247 ( .A1(n13725), .A2(n10664), .B1(n11854), .B2(n10663), .C1(
        n13167), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U13248 ( .A1(P3_U3897), .A2(n13087), .ZN(n10665) );
  OAI21_X1 U13249 ( .B1(P3_U3897), .B2(n10666), .A(n10665), .ZN(P3_U3501) );
  NAND2_X1 U13250 ( .A1(n13568), .A2(P3_U3897), .ZN(n10667) );
  OAI21_X1 U13251 ( .B1(P3_U3897), .B2(n10668), .A(n10667), .ZN(P3_U3504) );
  INV_X1 U13252 ( .A(n12183), .ZN(n12952) );
  NAND2_X1 U13253 ( .A1(n12952), .A2(P3_U3897), .ZN(n10669) );
  OAI21_X1 U13254 ( .B1(P3_U3897), .B2(n10670), .A(n10669), .ZN(P3_U3497) );
  INV_X1 U13255 ( .A(n10671), .ZN(n10672) );
  NAND2_X1 U13256 ( .A1(n10673), .A2(n10672), .ZN(n10712) );
  INV_X1 U13257 ( .A(n12696), .ZN(n14832) );
  INV_X1 U13258 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13259 ( .A1(n14832), .A2(n10674), .ZN(n10675) );
  NAND2_X1 U13260 ( .A1(n10710), .A2(n10675), .ZN(n14835) );
  INV_X1 U13261 ( .A(n14835), .ZN(n10676) );
  OAI21_X1 U13262 ( .B1(n14832), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10676), .ZN(
        n10677) );
  MUX2_X1 U13263 ( .A(n10677), .B(n10676), .S(P1_IR_REG_0__SCAN_IN), .Z(n10679) );
  INV_X1 U13264 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10678) );
  OAI22_X1 U13265 ( .A1(n10712), .A2(n10679), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10678), .ZN(n10681) );
  OR2_X1 U13266 ( .A1(n10712), .A2(n14832), .ZN(n14962) );
  NOR3_X1 U13267 ( .A1(n14962), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n7559), .ZN(
        n10680) );
  AOI211_X1 U13268 ( .C1(n14938), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10681), .B(
        n10680), .ZN(n10682) );
  INV_X1 U13269 ( .A(n10682), .ZN(P1_U3243) );
  INV_X1 U13270 ( .A(n10683), .ZN(n10750) );
  INV_X1 U13271 ( .A(n15433), .ZN(n15422) );
  AOI22_X1 U13272 ( .A1(n10977), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15422), .ZN(n10684) );
  OAI21_X1 U13273 ( .B1(n10750), .B2(n6554), .A(n10684), .ZN(P1_U3343) );
  INV_X1 U13274 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10685) );
  MUX2_X1 U13275 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10685), .S(n14844), .Z(
        n10688) );
  INV_X1 U13276 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10686) );
  MUX2_X1 U13277 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10686), .S(n14825), .Z(
        n14827) );
  AND2_X1 U13278 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14828) );
  NAND2_X1 U13279 ( .A1(n14827), .A2(n14828), .ZN(n14841) );
  NAND2_X1 U13280 ( .A1(n14825), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14840) );
  NAND2_X1 U13281 ( .A1(n14841), .A2(n14840), .ZN(n10687) );
  NAND2_X1 U13282 ( .A1(n10688), .A2(n10687), .ZN(n14861) );
  NAND2_X1 U13283 ( .A1(n14844), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U13284 ( .A1(n14861), .A2(n14860), .ZN(n10690) );
  MUX2_X1 U13285 ( .A(n15703), .B(P1_REG1_REG_3__SCAN_IN), .S(n14859), .Z(
        n10689) );
  OR2_X1 U13286 ( .A1(n14859), .A2(n15703), .ZN(n14875) );
  NAND2_X1 U13287 ( .A1(n14876), .A2(n14875), .ZN(n10693) );
  INV_X1 U13288 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10691) );
  MUX2_X1 U13289 ( .A(n10691), .B(P1_REG1_REG_4__SCAN_IN), .S(n14873), .Z(
        n10692) );
  NAND2_X1 U13290 ( .A1(n10693), .A2(n10692), .ZN(n14878) );
  OR2_X1 U13291 ( .A1(n14873), .A2(n10691), .ZN(n10694) );
  INV_X1 U13292 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15706) );
  MUX2_X1 U13293 ( .A(n15706), .B(P1_REG1_REG_5__SCAN_IN), .S(n14886), .Z(
        n14894) );
  NAND2_X1 U13294 ( .A1(n14893), .A2(n14894), .ZN(n14892) );
  NAND2_X1 U13295 ( .A1(n14886), .A2(n15706), .ZN(n10695) );
  NAND2_X1 U13296 ( .A1(n14892), .A2(n10695), .ZN(n10837) );
  INV_X1 U13297 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15708) );
  MUX2_X1 U13298 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15708), .S(n10847), .Z(
        n10836) );
  OR2_X1 U13299 ( .A1(n10847), .A2(n15708), .ZN(n14910) );
  NAND2_X1 U13300 ( .A1(n14911), .A2(n14910), .ZN(n10698) );
  INV_X1 U13301 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10696) );
  MUX2_X1 U13302 ( .A(n10696), .B(P1_REG1_REG_7__SCAN_IN), .S(n14908), .Z(
        n10697) );
  NAND2_X1 U13303 ( .A1(n10698), .A2(n10697), .ZN(n14913) );
  OR2_X1 U13304 ( .A1(n14908), .A2(n10696), .ZN(n10699) );
  INV_X1 U13305 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15712) );
  MUX2_X1 U13306 ( .A(n15712), .B(P1_REG1_REG_8__SCAN_IN), .S(n10793), .Z(
        n10786) );
  NAND2_X1 U13307 ( .A1(n10787), .A2(n10786), .ZN(n10785) );
  NAND2_X1 U13308 ( .A1(n10793), .A2(n15712), .ZN(n10700) );
  NAND2_X1 U13309 ( .A1(n10785), .A2(n10700), .ZN(n14921) );
  INV_X1 U13310 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10701) );
  XNOR2_X1 U13311 ( .A(n14924), .B(n10701), .ZN(n14922) );
  NAND2_X1 U13312 ( .A1(n14921), .A2(n14922), .ZN(n14920) );
  NAND2_X1 U13313 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  NAND2_X1 U13314 ( .A1(n14920), .A2(n10703), .ZN(n10849) );
  XNOR2_X1 U13315 ( .A(n10854), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n10850) );
  INV_X1 U13316 ( .A(n10708), .ZN(n10848) );
  AND2_X1 U13317 ( .A1(n10854), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10705) );
  OR2_X1 U13318 ( .A1(n10818), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10828) );
  NAND2_X1 U13319 ( .A1(n10818), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13320 ( .A1(n10828), .A2(n10704), .ZN(n10706) );
  OAI21_X1 U13321 ( .B1(n10848), .B2(n10705), .A(n10706), .ZN(n10709) );
  NOR2_X1 U13322 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  NAND2_X1 U13323 ( .A1(n10708), .A2(n10707), .ZN(n10829) );
  AOI21_X1 U13324 ( .B1(n10709), .B2(n10829), .A(n14962), .ZN(n10749) );
  OR2_X1 U13325 ( .A1(n10712), .A2(n10710), .ZN(n14957) );
  NAND2_X1 U13326 ( .A1(n10710), .A2(n14832), .ZN(n10711) );
  OR2_X1 U13327 ( .A1(n10712), .A2(n10711), .ZN(n14960) );
  INV_X1 U13328 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14845) );
  MUX2_X1 U13329 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14845), .S(n14844), .Z(
        n10716) );
  INV_X1 U13330 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10713) );
  MUX2_X1 U13331 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10713), .S(n14825), .Z(
        n14826) );
  AND2_X1 U13332 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10714) );
  NAND2_X1 U13333 ( .A1(n14826), .A2(n10714), .ZN(n14847) );
  NAND2_X1 U13334 ( .A1(n14825), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U13335 ( .A1(n14847), .A2(n14846), .ZN(n10715) );
  NAND2_X1 U13336 ( .A1(n10716), .A2(n10715), .ZN(n14856) );
  NAND2_X1 U13337 ( .A1(n14844), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U13338 ( .A1(n14856), .A2(n14855), .ZN(n10719) );
  INV_X1 U13339 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10717) );
  MUX2_X1 U13340 ( .A(n10717), .B(P1_REG2_REG_3__SCAN_IN), .S(n14859), .Z(
        n10718) );
  NAND2_X1 U13341 ( .A1(n10719), .A2(n10718), .ZN(n14871) );
  OR2_X1 U13342 ( .A1(n14859), .A2(n10717), .ZN(n14870) );
  NAND2_X1 U13343 ( .A1(n14871), .A2(n14870), .ZN(n10722) );
  INV_X1 U13344 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10720) );
  MUX2_X1 U13345 ( .A(n10720), .B(P1_REG2_REG_4__SCAN_IN), .S(n14873), .Z(
        n10721) );
  NAND2_X1 U13346 ( .A1(n10722), .A2(n10721), .ZN(n14889) );
  OR2_X1 U13347 ( .A1(n14873), .A2(n10720), .ZN(n14888) );
  NAND2_X1 U13348 ( .A1(n14889), .A2(n14888), .ZN(n10725) );
  INV_X1 U13349 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10723) );
  MUX2_X1 U13350 ( .A(n10723), .B(P1_REG2_REG_5__SCAN_IN), .S(n14886), .Z(
        n10724) );
  NAND2_X1 U13351 ( .A1(n10725), .A2(n10724), .ZN(n14891) );
  INV_X1 U13352 ( .A(n14886), .ZN(n14885) );
  NAND2_X1 U13353 ( .A1(n14885), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U13354 ( .A1(n14891), .A2(n10843), .ZN(n10727) );
  INV_X1 U13355 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11503) );
  MUX2_X1 U13356 ( .A(n11503), .B(P1_REG2_REG_6__SCAN_IN), .S(n10847), .Z(
        n10726) );
  NAND2_X1 U13357 ( .A1(n10727), .A2(n10726), .ZN(n14905) );
  OR2_X1 U13358 ( .A1(n10847), .A2(n11503), .ZN(n14904) );
  NAND2_X1 U13359 ( .A1(n14905), .A2(n14904), .ZN(n10729) );
  INV_X1 U13360 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10730) );
  MUX2_X1 U13361 ( .A(n10730), .B(P1_REG2_REG_7__SCAN_IN), .S(n14908), .Z(
        n10728) );
  NAND2_X1 U13362 ( .A1(n10729), .A2(n10728), .ZN(n14907) );
  OR2_X1 U13363 ( .A1(n14908), .A2(n10730), .ZN(n10789) );
  NAND2_X1 U13364 ( .A1(n14907), .A2(n10789), .ZN(n10732) );
  INV_X1 U13365 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11612) );
  MUX2_X1 U13366 ( .A(n11612), .B(P1_REG2_REG_8__SCAN_IN), .S(n10793), .Z(
        n10731) );
  NAND2_X1 U13367 ( .A1(n10732), .A2(n10731), .ZN(n14927) );
  OR2_X1 U13368 ( .A1(n10793), .A2(n11612), .ZN(n14926) );
  NAND2_X1 U13369 ( .A1(n14927), .A2(n14926), .ZN(n10735) );
  INV_X1 U13370 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10733) );
  MUX2_X1 U13371 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10733), .S(n14924), .Z(
        n10734) );
  NAND2_X1 U13372 ( .A1(n10735), .A2(n10734), .ZN(n14929) );
  NAND2_X1 U13373 ( .A1(n14924), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10857) );
  NAND2_X1 U13374 ( .A1(n14929), .A2(n10857), .ZN(n10737) );
  MUX2_X1 U13375 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10855), .S(n10854), .Z(
        n10736) );
  NAND2_X1 U13376 ( .A1(n10737), .A2(n10736), .ZN(n10859) );
  NAND2_X1 U13377 ( .A1(n10854), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13378 ( .A1(n10859), .A2(n10742), .ZN(n10740) );
  MUX2_X1 U13379 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10738), .S(n10818), .Z(
        n10739) );
  NAND2_X1 U13380 ( .A1(n10740), .A2(n10739), .ZN(n10820) );
  MUX2_X1 U13381 ( .A(n10738), .B(P1_REG2_REG_11__SCAN_IN), .S(n10818), .Z(
        n10741) );
  NAND3_X1 U13382 ( .A1(n10859), .A2(n10742), .A3(n10741), .ZN(n10743) );
  NAND3_X1 U13383 ( .A1(n15505), .A2(n10820), .A3(n10743), .ZN(n10746) );
  NOR2_X1 U13384 ( .A1(n10744), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12231) );
  AOI21_X1 U13385 ( .B1(n14938), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n12231), 
        .ZN(n10745) );
  OAI211_X1 U13386 ( .C1(n14957), .C2(n10747), .A(n10746), .B(n10745), .ZN(
        n10748) );
  OR2_X1 U13387 ( .A1(n10749), .A2(n10748), .ZN(P1_U3254) );
  INV_X1 U13388 ( .A(n15746), .ZN(n11347) );
  OAI222_X1 U13389 ( .A1(n12702), .A2(n10751), .B1(n11978), .B2(n10750), .C1(
        n11347), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13390 ( .A(n13713), .ZN(n11718) );
  NOR2_X1 U13391 ( .A1(n11718), .A2(n10752), .ZN(n10754) );
  INV_X1 U13392 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10753) );
  NOR2_X1 U13393 ( .A1(n10779), .A2(n10753), .ZN(P3_U3245) );
  CLKBUF_X1 U13394 ( .A(n10754), .Z(n10779) );
  INV_X1 U13395 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10755) );
  NOR2_X1 U13396 ( .A1(n10779), .A2(n10755), .ZN(P3_U3246) );
  INV_X1 U13397 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10756) );
  NOR2_X1 U13398 ( .A1(n10779), .A2(n10756), .ZN(P3_U3248) );
  INV_X1 U13399 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10757) );
  NOR2_X1 U13400 ( .A1(n10779), .A2(n10757), .ZN(P3_U3249) );
  INV_X1 U13401 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10758) );
  NOR2_X1 U13402 ( .A1(n10779), .A2(n10758), .ZN(P3_U3250) );
  NOR2_X1 U13403 ( .A1(n10779), .A2(n10759), .ZN(P3_U3251) );
  INV_X1 U13404 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10760) );
  NOR2_X1 U13405 ( .A1(n10779), .A2(n10760), .ZN(P3_U3252) );
  INV_X1 U13406 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10761) );
  NOR2_X1 U13407 ( .A1(n10779), .A2(n10761), .ZN(P3_U3253) );
  INV_X1 U13408 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10762) );
  NOR2_X1 U13409 ( .A1(n10779), .A2(n10762), .ZN(P3_U3254) );
  INV_X1 U13410 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10763) );
  NOR2_X1 U13411 ( .A1(n10779), .A2(n10763), .ZN(P3_U3255) );
  INV_X1 U13412 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10764) );
  NOR2_X1 U13413 ( .A1(n10779), .A2(n10764), .ZN(P3_U3256) );
  INV_X1 U13414 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10765) );
  NOR2_X1 U13415 ( .A1(n10779), .A2(n10765), .ZN(P3_U3257) );
  INV_X1 U13416 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10766) );
  NOR2_X1 U13417 ( .A1(n10754), .A2(n10766), .ZN(P3_U3258) );
  INV_X1 U13418 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10767) );
  NOR2_X1 U13419 ( .A1(n10779), .A2(n10767), .ZN(P3_U3259) );
  INV_X1 U13420 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10768) );
  NOR2_X1 U13421 ( .A1(n10754), .A2(n10768), .ZN(P3_U3260) );
  INV_X1 U13422 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10769) );
  NOR2_X1 U13423 ( .A1(n10779), .A2(n10769), .ZN(P3_U3261) );
  INV_X1 U13424 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10770) );
  NOR2_X1 U13425 ( .A1(n10754), .A2(n10770), .ZN(P3_U3262) );
  INV_X1 U13426 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10771) );
  NOR2_X1 U13427 ( .A1(n10779), .A2(n10771), .ZN(P3_U3263) );
  INV_X1 U13428 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10772) );
  NOR2_X1 U13429 ( .A1(n10754), .A2(n10772), .ZN(P3_U3244) );
  INV_X1 U13430 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10773) );
  NOR2_X1 U13431 ( .A1(n10754), .A2(n10773), .ZN(P3_U3243) );
  INV_X1 U13432 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10774) );
  NOR2_X1 U13433 ( .A1(n10754), .A2(n10774), .ZN(P3_U3242) );
  NOR2_X1 U13434 ( .A1(n10754), .A2(n10775), .ZN(P3_U3241) );
  INV_X1 U13435 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10776) );
  NOR2_X1 U13436 ( .A1(n10754), .A2(n10776), .ZN(P3_U3240) );
  INV_X1 U13437 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10777) );
  NOR2_X1 U13438 ( .A1(n10754), .A2(n10777), .ZN(P3_U3239) );
  NOR2_X1 U13439 ( .A1(n10779), .A2(n10778), .ZN(P3_U3247) );
  INV_X1 U13440 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10780) );
  NOR2_X1 U13441 ( .A1(n10754), .A2(n10780), .ZN(P3_U3237) );
  NOR2_X1 U13442 ( .A1(n10754), .A2(n10781), .ZN(P3_U3236) );
  INV_X1 U13443 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10782) );
  NOR2_X1 U13444 ( .A1(n10779), .A2(n10782), .ZN(P3_U3235) );
  INV_X1 U13445 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10783) );
  NOR2_X1 U13446 ( .A1(n10779), .A2(n10783), .ZN(P3_U3234) );
  INV_X1 U13447 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10784) );
  NOR2_X1 U13448 ( .A1(n10779), .A2(n10784), .ZN(P3_U3238) );
  OAI21_X1 U13449 ( .B1(n10787), .B2(n10786), .A(n10785), .ZN(n10795) );
  MUX2_X1 U13450 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11612), .S(n10793), .Z(
        n10788) );
  NAND3_X1 U13451 ( .A1(n14907), .A2(n10789), .A3(n10788), .ZN(n10790) );
  NAND3_X1 U13452 ( .A1(n15505), .A2(n14927), .A3(n10790), .ZN(n10792) );
  AND2_X1 U13453 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11597) );
  AOI21_X1 U13454 ( .B1(n14938), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11597), .ZN(
        n10791) );
  OAI211_X1 U13455 ( .C1(n14957), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI21_X1 U13456 ( .B1(n15504), .B2(n10795), .A(n10794), .ZN(n10796) );
  INV_X1 U13457 ( .A(n10796), .ZN(P1_U3251) );
  AND2_X1 U13458 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10865) );
  INV_X1 U13459 ( .A(n10865), .ZN(n10797) );
  XNOR2_X1 U13460 ( .A(n10867), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n10866) );
  MUX2_X1 U13461 ( .A(n10797), .B(n10865), .S(n10866), .Z(n10812) );
  AOI21_X1 U13462 ( .B1(n10954), .B2(n10799), .A(n10798), .ZN(n10800) );
  OR2_X1 U13463 ( .A1(n10801), .A2(n10800), .ZN(n10804) );
  NOR2_X1 U13464 ( .A1(n8974), .A2(n6531), .ZN(n14665) );
  AND2_X1 U13465 ( .A1(n10804), .A2(n14665), .ZN(n10807) );
  INV_X1 U13466 ( .A(n15734), .ZN(n14197) );
  NOR2_X2 U13467 ( .A1(n10804), .A2(n6531), .ZN(n15715) );
  AND2_X1 U13468 ( .A1(n8974), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10803) );
  NAND2_X1 U13469 ( .A1(n10804), .A2(n10803), .ZN(n14206) );
  INV_X1 U13470 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11336) );
  OAI22_X1 U13471 ( .A1(n14206), .A2(n10867), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11336), .ZN(n10805) );
  AOI21_X1 U13472 ( .B1(n15715), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n10805), .ZN(
        n10811) );
  XNOR2_X1 U13473 ( .A(n10867), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n10809) );
  INV_X1 U13474 ( .A(n10806), .ZN(n10808) );
  NAND2_X1 U13475 ( .A1(n10807), .A2(n12399), .ZN(n14207) );
  NAND2_X1 U13476 ( .A1(n10809), .A2(n10808), .ZN(n10895) );
  OAI211_X1 U13477 ( .C1(n10809), .C2(n10808), .A(n15744), .B(n10895), .ZN(
        n10810) );
  OAI211_X1 U13478 ( .C1(n10812), .C2(n14197), .A(n10811), .B(n10810), .ZN(
        P2_U3215) );
  OAI222_X1 U13479 ( .A1(n13725), .A2(n10814), .B1(n13731), .B2(n10813), .C1(
        n13226), .C2(P3_U3151), .ZN(P3_U3280) );
  OAI222_X1 U13480 ( .A1(n13725), .A2(n10816), .B1(n13731), .B2(n10815), .C1(
        n13185), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U13481 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10817) );
  MUX2_X1 U13482 ( .A(n10817), .B(P1_REG2_REG_12__SCAN_IN), .S(n10977), .Z(
        n10823) );
  NAND2_X1 U13483 ( .A1(n10818), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13484 ( .A1(n10820), .A2(n10819), .ZN(n10822) );
  INV_X1 U13485 ( .A(n10979), .ZN(n10821) );
  AOI21_X1 U13486 ( .B1(n10823), .B2(n10822), .A(n10821), .ZN(n10835) );
  INV_X1 U13487 ( .A(n14957), .ZN(n15501) );
  NOR2_X1 U13488 ( .A1(n10824), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12291) );
  NOR2_X1 U13489 ( .A1(n15509), .A2(n10825), .ZN(n10826) );
  AOI211_X1 U13490 ( .C1(n15501), .C2(n10977), .A(n12291), .B(n10826), .ZN(
        n10834) );
  XNOR2_X1 U13491 ( .A(n10977), .B(n10827), .ZN(n10831) );
  NAND2_X1 U13492 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  NAND2_X1 U13493 ( .A1(n10830), .A2(n10831), .ZN(n11012) );
  OAI21_X1 U13494 ( .B1(n10831), .B2(n10830), .A(n11012), .ZN(n10832) );
  NAND2_X1 U13495 ( .A1(n10832), .A2(n15504), .ZN(n10833) );
  OAI211_X1 U13496 ( .C1(n10835), .C2(n14960), .A(n10834), .B(n10833), .ZN(
        P1_U3255) );
  AND2_X1 U13497 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U13498 ( .A1(n10837), .A2(n10836), .ZN(n10838) );
  NAND3_X1 U13499 ( .A1(n15504), .A2(n14911), .A3(n10838), .ZN(n10839) );
  OAI21_X1 U13500 ( .B1(n10840), .B2(n15509), .A(n10839), .ZN(n10841) );
  NOR2_X1 U13501 ( .A1(n11648), .A2(n10841), .ZN(n10846) );
  MUX2_X1 U13502 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11503), .S(n10847), .Z(
        n10842) );
  NAND3_X1 U13503 ( .A1(n14891), .A2(n10843), .A3(n10842), .ZN(n10844) );
  NAND3_X1 U13504 ( .A1(n15505), .A2(n14905), .A3(n10844), .ZN(n10845) );
  OAI211_X1 U13505 ( .C1(n14957), .C2(n10847), .A(n10846), .B(n10845), .ZN(
        P1_U3249) );
  AOI211_X1 U13506 ( .C1(n10850), .C2(n10849), .A(n14962), .B(n10848), .ZN(
        n10851) );
  INV_X1 U13507 ( .A(n10851), .ZN(n10852) );
  OAI21_X1 U13508 ( .B1(n10853), .B2(n15509), .A(n10852), .ZN(n10863) );
  MUX2_X1 U13509 ( .A(n10855), .B(P1_REG2_REG_10__SCAN_IN), .S(n10854), .Z(
        n10856) );
  NAND3_X1 U13510 ( .A1(n14929), .A2(n10857), .A3(n10856), .ZN(n10858) );
  NAND3_X1 U13511 ( .A1(n15505), .A2(n10859), .A3(n10858), .ZN(n10860) );
  NAND2_X1 U13512 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12068)
         );
  OAI211_X1 U13513 ( .C1(n14957), .C2(n10861), .A(n10860), .B(n12068), .ZN(
        n10862) );
  OR2_X1 U13514 ( .A1(n10863), .A2(n10862), .ZN(P1_U3253) );
  INV_X1 U13515 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11379) );
  MUX2_X1 U13516 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11379), .S(n14058), .Z(
        n10871) );
  INV_X1 U13517 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13518 ( .A1(n10866), .A2(n10865), .ZN(n10869) );
  INV_X1 U13519 ( .A(n10867), .ZN(n10893) );
  NAND2_X1 U13520 ( .A1(n10893), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U13521 ( .A1(n10869), .A2(n10868), .ZN(n14047) );
  NAND2_X1 U13522 ( .A1(n14049), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U13523 ( .A1(n10871), .A2(n10870), .ZN(n14076) );
  NAND2_X1 U13524 ( .A1(n14058), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14075) );
  NAND2_X1 U13525 ( .A1(n14076), .A2(n14075), .ZN(n10873) );
  MUX2_X1 U13526 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n14073), .S(n14072), .Z(
        n10872) );
  NAND2_X1 U13527 ( .A1(n10873), .A2(n10872), .ZN(n14090) );
  NAND2_X1 U13528 ( .A1(n14072), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n14089) );
  NAND2_X1 U13529 ( .A1(n14090), .A2(n14089), .ZN(n10875) );
  MUX2_X1 U13530 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n14088), .S(n14087), .Z(
        n10874) );
  NAND2_X1 U13531 ( .A1(n10875), .A2(n10874), .ZN(n14105) );
  NAND2_X1 U13532 ( .A1(n14087), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14104) );
  NAND2_X1 U13533 ( .A1(n14105), .A2(n14104), .ZN(n10877) );
  INV_X1 U13534 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11557) );
  MUX2_X1 U13535 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11557), .S(n14102), .Z(
        n10876) );
  NAND2_X1 U13536 ( .A1(n10877), .A2(n10876), .ZN(n14119) );
  NAND2_X1 U13537 ( .A1(n14102), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U13538 ( .A1(n14119), .A2(n14118), .ZN(n10879) );
  MUX2_X1 U13539 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n14116), .S(n14115), .Z(
        n10878) );
  NAND2_X1 U13540 ( .A1(n10879), .A2(n10878), .ZN(n14132) );
  NAND2_X1 U13541 ( .A1(n14115), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U13542 ( .A1(n14132), .A2(n14131), .ZN(n10881) );
  INV_X1 U13543 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11588) );
  MUX2_X1 U13544 ( .A(n11588), .B(P2_REG2_REG_8__SCAN_IN), .S(n14129), .Z(
        n10880) );
  NAND2_X1 U13545 ( .A1(n10882), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10883) );
  INV_X1 U13546 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10884) );
  MUX2_X1 U13547 ( .A(n10884), .B(P2_REG2_REG_9__SCAN_IN), .S(n15718), .Z(
        n15717) );
  NAND2_X1 U13548 ( .A1(n15718), .A2(n10884), .ZN(n10885) );
  INV_X1 U13549 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n12021) );
  MUX2_X1 U13550 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n12021), .S(n10908), .Z(
        n14146) );
  NAND2_X1 U13551 ( .A1(n14147), .A2(n14146), .ZN(n14145) );
  NAND2_X1 U13552 ( .A1(n10908), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13553 ( .A1(n14145), .A2(n10886), .ZN(n10889) );
  INV_X1 U13554 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n14500) );
  MUX2_X1 U13555 ( .A(n14500), .B(P2_REG2_REG_11__SCAN_IN), .S(n11352), .Z(
        n10888) );
  INV_X1 U13556 ( .A(n15733), .ZN(n10887) );
  AOI21_X1 U13557 ( .B1(n10889), .B2(n10888), .A(n10887), .ZN(n10914) );
  INV_X1 U13558 ( .A(n14206), .ZN(n15747) );
  NOR2_X1 U13559 ( .A1(n10890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13980) );
  INV_X1 U13560 ( .A(n15715), .ZN(n15753) );
  NOR2_X1 U13561 ( .A1(n15753), .A2(n15459), .ZN(n10891) );
  AOI211_X1 U13562 ( .C1(n15747), .C2(n11352), .A(n13980), .B(n10891), .ZN(
        n10913) );
  INV_X1 U13563 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10892) );
  XNOR2_X1 U13564 ( .A(n11352), .B(n10892), .ZN(n10911) );
  INV_X1 U13565 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n15853) );
  MUX2_X1 U13566 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n15853), .S(n14049), .Z(
        n14045) );
  NAND2_X1 U13567 ( .A1(n10893), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13568 ( .A1(n10895), .A2(n10894), .ZN(n14044) );
  NAND2_X1 U13569 ( .A1(n14045), .A2(n14044), .ZN(n14043) );
  NAND2_X1 U13570 ( .A1(n14049), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10896) );
  NAND2_X1 U13571 ( .A1(n14043), .A2(n10896), .ZN(n14055) );
  INV_X1 U13572 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10897) );
  XNOR2_X1 U13573 ( .A(n14058), .B(n10897), .ZN(n14056) );
  NAND2_X1 U13574 ( .A1(n14055), .A2(n14056), .ZN(n14054) );
  NAND2_X1 U13575 ( .A1(n14058), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U13576 ( .A1(n14054), .A2(n10898), .ZN(n14068) );
  MUX2_X1 U13577 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15856), .S(n14072), .Z(
        n14069) );
  NAND2_X1 U13578 ( .A1(n14068), .A2(n14069), .ZN(n14067) );
  NAND2_X1 U13579 ( .A1(n14072), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13580 ( .A1(n14067), .A2(n10899), .ZN(n14083) );
  INV_X1 U13581 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10900) );
  XNOR2_X1 U13582 ( .A(n14087), .B(n10900), .ZN(n14084) );
  NAND2_X1 U13583 ( .A1(n14083), .A2(n14084), .ZN(n14082) );
  NAND2_X1 U13584 ( .A1(n14087), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U13585 ( .A1(n14082), .A2(n10901), .ZN(n14098) );
  INV_X1 U13586 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15859) );
  MUX2_X1 U13587 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15859), .S(n14102), .Z(
        n14099) );
  NAND2_X1 U13588 ( .A1(n14098), .A2(n14099), .ZN(n14097) );
  NAND2_X1 U13589 ( .A1(n14102), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U13590 ( .A1(n14097), .A2(n10902), .ZN(n14112) );
  INV_X1 U13591 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15861) );
  MUX2_X1 U13592 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15861), .S(n14115), .Z(
        n14113) );
  NAND2_X1 U13593 ( .A1(n14112), .A2(n14113), .ZN(n14111) );
  NAND2_X1 U13594 ( .A1(n14115), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U13595 ( .A1(n14111), .A2(n10903), .ZN(n14127) );
  MUX2_X1 U13596 ( .A(n10904), .B(P2_REG1_REG_8__SCAN_IN), .S(n14129), .Z(
        n14128) );
  NAND2_X1 U13597 ( .A1(n14127), .A2(n14128), .ZN(n15719) );
  INV_X1 U13598 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10906) );
  XNOR2_X1 U13599 ( .A(n15718), .B(n10906), .ZN(n15720) );
  NOR2_X1 U13600 ( .A1(n14129), .A2(n10904), .ZN(n15721) );
  NOR2_X1 U13601 ( .A1(n15720), .A2(n15721), .ZN(n10905) );
  NAND2_X1 U13602 ( .A1(n15719), .A2(n10905), .ZN(n15723) );
  NAND2_X1 U13603 ( .A1(n15718), .A2(n10906), .ZN(n10907) );
  NAND2_X1 U13604 ( .A1(n15723), .A2(n10907), .ZN(n14138) );
  XNOR2_X1 U13605 ( .A(n10908), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U13606 ( .A1(n10908), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10909) );
  NAND2_X1 U13607 ( .A1(n14140), .A2(n10909), .ZN(n10910) );
  NAND2_X1 U13608 ( .A1(n10910), .A2(n10911), .ZN(n15738) );
  OAI211_X1 U13609 ( .C1(n10911), .C2(n10910), .A(n15738), .B(n15744), .ZN(
        n10912) );
  OAI211_X1 U13610 ( .C1(n10914), .C2(n14197), .A(n10913), .B(n10912), .ZN(
        P2_U3225) );
  AOI22_X1 U13611 ( .A1(n15744), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15734), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10918) );
  INV_X1 U13612 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11299) );
  NAND2_X1 U13613 ( .A1(n15734), .A2(n11299), .ZN(n10915) );
  OAI211_X1 U13614 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14207), .A(n10915), .B(
        n14206), .ZN(n10916) );
  INV_X1 U13615 ( .A(n10916), .ZN(n10917) );
  MUX2_X1 U13616 ( .A(n10918), .B(n10917), .S(P2_IR_REG_0__SCAN_IN), .Z(n10920) );
  AOI22_X1 U13617 ( .A1(n15715), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n6531), .ZN(n10919) );
  NAND2_X1 U13618 ( .A1(n10920), .A2(n10919), .ZN(P2_U3214) );
  OAI222_X1 U13619 ( .A1(n13725), .A2(n10922), .B1(n13731), .B2(n10921), .C1(
        n13195), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U13620 ( .A(n10923), .ZN(n10926) );
  OAI222_X1 U13621 ( .A1(n12702), .A2(n10924), .B1(n11978), .B2(n10926), .C1(
        n14155), .C2(n6531), .ZN(P2_U3314) );
  INV_X1 U13622 ( .A(n10981), .ZN(n11024) );
  OAI222_X1 U13623 ( .A1(P1_U3086), .A2(n11024), .B1(n6554), .B2(n10926), .C1(
        n10925), .C2(n15433), .ZN(P1_U3342) );
  OAI21_X1 U13624 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(n14834) );
  INV_X1 U13625 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U13626 ( .A1(n10932), .A2(n10931), .ZN(n11042) );
  AOI22_X1 U13627 ( .A1(n14834), .A2(n15491), .B1(n11042), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U13628 ( .A1(n14779), .A2(n15566), .ZN(n10933) );
  OAI211_X1 U13629 ( .C1(n14809), .C2(n12492), .A(n10934), .B(n10933), .ZN(
        P1_U3232) );
  INV_X1 U13630 ( .A(n10935), .ZN(n10938) );
  INV_X1 U13631 ( .A(n11630), .ZN(n10936) );
  OAI222_X1 U13632 ( .A1(n15433), .A2(n10937), .B1(n6554), .B2(n10938), .C1(
        P1_U3086), .C2(n10936), .ZN(P1_U3341) );
  OAI222_X1 U13633 ( .A1(n12702), .A2(n10939), .B1(n11978), .B2(n10938), .C1(
        P2_U3088), .C2(n7051), .ZN(P2_U3313) );
  INV_X1 U13634 ( .A(n10940), .ZN(n10942) );
  NOR2_X1 U13635 ( .A1(n10942), .A2(n10941), .ZN(n10944) );
  NAND2_X1 U13636 ( .A1(n10944), .A2(n10943), .ZN(n10960) );
  INV_X1 U13637 ( .A(n10945), .ZN(n10946) );
  NAND2_X1 U13638 ( .A1(n10960), .A2(n10946), .ZN(n10950) );
  AND2_X1 U13639 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  NAND2_X1 U13640 ( .A1(n10950), .A2(n10949), .ZN(n11204) );
  NOR2_X1 U13641 ( .A1(n11204), .A2(n6531), .ZN(n11175) );
  NAND2_X1 U13642 ( .A1(n15781), .A2(n10951), .ZN(n10952) );
  OR2_X1 U13643 ( .A1(n10960), .A2(n10952), .ZN(n10953) );
  NOR2_X1 U13644 ( .A1(n15835), .A2(n10954), .ZN(n10955) );
  NAND2_X1 U13645 ( .A1(n15781), .A2(n10955), .ZN(n10956) );
  OAI21_X1 U13646 ( .B1(n13800), .B2(n10958), .A(n7647), .ZN(n10959) );
  AOI22_X1 U13647 ( .A1(n14000), .A2(n11301), .B1(n14004), .B2(n10959), .ZN(
        n10965) );
  INV_X1 U13648 ( .A(n10960), .ZN(n10963) );
  AND2_X1 U13649 ( .A1(n15781), .A2(n10961), .ZN(n10962) );
  NAND2_X1 U13650 ( .A1(n13992), .A2(n14494), .ZN(n13950) );
  INV_X1 U13651 ( .A(n13950), .ZN(n13981) );
  NAND2_X1 U13652 ( .A1(n13981), .A2(n6596), .ZN(n10964) );
  OAI211_X1 U13653 ( .C1(n11175), .C2(n11296), .A(n10965), .B(n10964), .ZN(
        P2_U3204) );
  INV_X1 U13654 ( .A(n13272), .ZN(n10969) );
  INV_X1 U13655 ( .A(n10966), .ZN(n10968) );
  OAI222_X1 U13656 ( .A1(n10969), .A2(P3_U3151), .B1(n13729), .B2(n10968), 
        .C1(n10967), .C2(n11854), .ZN(P3_U3279) );
  INV_X1 U13657 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10970) );
  XNOR2_X1 U13658 ( .A(n10981), .B(n10970), .ZN(n11014) );
  OR2_X1 U13659 ( .A1(n10977), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11011) );
  AND2_X1 U13660 ( .A1(n11014), .A2(n11011), .ZN(n10971) );
  NAND2_X1 U13661 ( .A1(n11012), .A2(n10971), .ZN(n11013) );
  NAND2_X1 U13662 ( .A1(n10981), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U13663 ( .A1(n11013), .A2(n10972), .ZN(n11629) );
  XOR2_X1 U13664 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11630), .Z(n10973) );
  XNOR2_X1 U13665 ( .A(n11629), .B(n10973), .ZN(n10990) );
  NOR2_X1 U13666 ( .A1(n10974), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14670) );
  NOR2_X1 U13667 ( .A1(n15509), .A2(n10975), .ZN(n10976) );
  AOI211_X1 U13668 ( .C1(n15501), .C2(n11630), .A(n14670), .B(n10976), .ZN(
        n10989) );
  OR2_X1 U13669 ( .A1(n10977), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13670 ( .A1(n10979), .A2(n10978), .ZN(n11016) );
  MUX2_X1 U13671 ( .A(n10980), .B(P1_REG2_REG_13__SCAN_IN), .S(n10981), .Z(
        n11017) );
  NAND2_X1 U13672 ( .A1(n10981), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10986) );
  NAND2_X1 U13673 ( .A1(n11018), .A2(n10986), .ZN(n10984) );
  INV_X1 U13674 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10982) );
  MUX2_X1 U13675 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10982), .S(n11630), .Z(
        n10983) );
  NAND2_X1 U13676 ( .A1(n10984), .A2(n10983), .ZN(n11620) );
  MUX2_X1 U13677 ( .A(n10982), .B(P1_REG2_REG_14__SCAN_IN), .S(n11630), .Z(
        n10985) );
  NAND3_X1 U13678 ( .A1(n11018), .A2(n10986), .A3(n10985), .ZN(n10987) );
  NAND3_X1 U13679 ( .A1(n11620), .A2(n15505), .A3(n10987), .ZN(n10988) );
  OAI211_X1 U13680 ( .C1(n10990), .C2(n14962), .A(n10989), .B(n10988), .ZN(
        P1_U3257) );
  XNOR2_X1 U13681 ( .A(n11164), .B(n11165), .ZN(n10995) );
  NAND2_X1 U13682 ( .A1(n13864), .A2(n11335), .ZN(n10993) );
  OAI21_X1 U13683 ( .B1(n10995), .B2(n10994), .A(n11168), .ZN(n11000) );
  OAI22_X1 U13684 ( .A1(n13950), .A2(n10996), .B1(n14014), .B2(n8535), .ZN(
        n10999) );
  NAND2_X1 U13685 ( .A1(n13992), .A2(n14496), .ZN(n13978) );
  INV_X1 U13686 ( .A(n9670), .ZN(n10997) );
  OAI22_X1 U13687 ( .A1(n11175), .A2(n11336), .B1(n13978), .B2(n10997), .ZN(
        n10998) );
  AOI211_X1 U13688 ( .C1(n14004), .C2(n11000), .A(n10999), .B(n10998), .ZN(
        n11001) );
  INV_X1 U13689 ( .A(n11001), .ZN(P2_U3194) );
  OR2_X1 U13690 ( .A1(n11002), .A2(n15207), .ZN(n15674) );
  NAND2_X1 U13691 ( .A1(n15694), .A2(n15651), .ZN(n11003) );
  INV_X1 U13692 ( .A(n15564), .ZN(n15567) );
  XNOR2_X1 U13693 ( .A(n15567), .B(n12492), .ZN(n12650) );
  AOI222_X1 U13694 ( .A1(n11003), .A2(n12650), .B1(n12490), .B2(n6755), .C1(
        n15566), .C2(n15668), .ZN(n15618) );
  AND2_X1 U13695 ( .A1(n11005), .A2(n11004), .ZN(n15394) );
  AND3_X2 U13696 ( .A1(n11007), .A2(n15394), .A3(n11006), .ZN(n15714) );
  NAND2_X1 U13697 ( .A1(n15711), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n11008) );
  OAI21_X1 U13698 ( .B1(n15618), .B2(n15711), .A(n11008), .ZN(P1_U3528) );
  OAI222_X1 U13699 ( .A1(n13725), .A2(n11010), .B1(n13731), .B2(n11009), .C1(
        n13294), .C2(P3_U3151), .ZN(P3_U3278) );
  AND2_X1 U13700 ( .A1(n11012), .A2(n11011), .ZN(n11015) );
  OAI211_X1 U13701 ( .C1(n11015), .C2(n11014), .A(n15504), .B(n11013), .ZN(
        n11023) );
  NAND2_X1 U13702 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14764)
         );
  AOI21_X1 U13703 ( .B1(n11017), .B2(n11016), .A(n14960), .ZN(n11019) );
  NAND2_X1 U13704 ( .A1(n11019), .A2(n11018), .ZN(n11020) );
  NAND2_X1 U13705 ( .A1(n14764), .A2(n11020), .ZN(n11021) );
  AOI21_X1 U13706 ( .B1(n14938), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11021), 
        .ZN(n11022) );
  OAI211_X1 U13707 ( .C1(n14957), .C2(n11024), .A(n11023), .B(n11022), .ZN(
        P1_U3256) );
  NOR2_X1 U13708 ( .A1(n10269), .A2(n11304), .ZN(n11025) );
  OAI22_X1 U13709 ( .A1(n11304), .A2(n14461), .B1(n11158), .B2(n14473), .ZN(
        n11297) );
  AOI211_X1 U13710 ( .C1(n6591), .C2(n11301), .A(n11025), .B(n11297), .ZN(
        n11028) );
  NAND2_X1 U13711 ( .A1(n8995), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n11026) );
  OAI21_X1 U13712 ( .B1(n11028), .B2(n8995), .A(n11026), .ZN(P2_U3499) );
  NAND2_X1 U13713 ( .A1(n9003), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n11027) );
  OAI21_X1 U13714 ( .B1(n11028), .B2(n9003), .A(n11027), .ZN(P2_U3430) );
  XOR2_X1 U13715 ( .A(n11030), .B(n11029), .Z(n11033) );
  INV_X1 U13716 ( .A(n15491), .ZN(n14815) );
  AOI22_X1 U13717 ( .A1(n14806), .A2(n15566), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n11042), .ZN(n11032) );
  NOR2_X1 U13718 ( .A1(n15682), .A2(n12508), .ZN(n15633) );
  INV_X1 U13719 ( .A(n11647), .ZN(n15483) );
  AOI22_X1 U13720 ( .A1(n14779), .A2(n15647), .B1(n15633), .B2(n15483), .ZN(
        n11031) );
  OAI211_X1 U13721 ( .C1(n11033), .C2(n14815), .A(n11032), .B(n11031), .ZN(
        P1_U3237) );
  NAND2_X1 U13722 ( .A1(n13013), .A2(P3_U3897), .ZN(n11034) );
  OAI21_X1 U13723 ( .B1(P3_U3897), .B2(n11035), .A(n11034), .ZN(P3_U3511) );
  INV_X1 U13724 ( .A(n11964), .ZN(n11571) );
  INV_X1 U13725 ( .A(n11036), .ZN(n11039) );
  OAI222_X1 U13726 ( .A1(P2_U3088), .A2(n11571), .B1(n11978), .B2(n11039), 
        .C1(n11037), .C2(n14659), .ZN(P2_U3312) );
  OAI222_X1 U13727 ( .A1(P1_U3086), .A2(n11621), .B1(n6554), .B2(n11039), .C1(
        n11038), .C2(n15433), .ZN(P1_U3340) );
  XOR2_X1 U13728 ( .A(n11041), .B(n11040), .Z(n11046) );
  AOI22_X1 U13729 ( .A1(n14779), .A2(n15562), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n11042), .ZN(n11043) );
  OAI21_X1 U13730 ( .B1(n15564), .B2(n14798), .A(n11043), .ZN(n11044) );
  AOI21_X1 U13731 ( .B1(n14769), .B2(n12497), .A(n11044), .ZN(n11045) );
  OAI21_X1 U13732 ( .B1(n14815), .B2(n11046), .A(n11045), .ZN(P1_U3222) );
  AND2_X1 U13733 ( .A1(n11047), .A2(n11401), .ZN(n12799) );
  NOR2_X1 U13734 ( .A1(n12802), .A2(n12799), .ZN(n15868) );
  NAND2_X1 U13735 ( .A1(n11048), .A2(n15928), .ZN(n11049) );
  OR2_X1 U13736 ( .A1(n15868), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U13737 ( .A1(n15866), .A2(n13566), .ZN(n11050) );
  AND2_X1 U13738 ( .A1(n11051), .A2(n11050), .ZN(n11416) );
  INV_X1 U13739 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11052) );
  MUX2_X1 U13740 ( .A(n11416), .B(n11052), .S(n15941), .Z(n11053) );
  OAI21_X1 U13741 ( .B1(n11401), .B2(n13711), .A(n11053), .ZN(P3_U3390) );
  MUX2_X1 U13742 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13285), .Z(n11243) );
  INV_X1 U13743 ( .A(n11248), .ZN(n11244) );
  XNOR2_X1 U13744 ( .A(n11243), .B(n11244), .ZN(n11241) );
  XNOR2_X1 U13745 ( .A(n11054), .B(n11085), .ZN(n11180) );
  INV_X1 U13746 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11415) );
  INV_X1 U13747 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11399) );
  INV_X1 U13748 ( .A(n11054), .ZN(n11055) );
  NAND2_X1 U13749 ( .A1(n11055), .A2(n11085), .ZN(n11056) );
  NAND2_X1 U13750 ( .A1(n11057), .A2(n11056), .ZN(n11108) );
  MUX2_X1 U13751 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13727), .Z(n11058) );
  INV_X1 U13752 ( .A(n11088), .ZN(n11122) );
  XNOR2_X1 U13753 ( .A(n11058), .B(n11122), .ZN(n11109) );
  INV_X1 U13754 ( .A(n11058), .ZN(n11059) );
  NAND2_X1 U13755 ( .A1(n11059), .A2(n11122), .ZN(n11060) );
  MUX2_X1 U13756 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13727), .Z(n11061) );
  INV_X1 U13757 ( .A(n11152), .ZN(n11076) );
  XNOR2_X1 U13758 ( .A(n11061), .B(n11076), .ZN(n11145) );
  NAND2_X1 U13759 ( .A1(n11144), .A2(n11145), .ZN(n11064) );
  INV_X1 U13760 ( .A(n11061), .ZN(n11062) );
  NAND2_X1 U13761 ( .A1(n11062), .A2(n11076), .ZN(n11063) );
  MUX2_X1 U13762 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13727), .Z(n11065) );
  INV_X1 U13763 ( .A(n11094), .ZN(n11141) );
  XNOR2_X1 U13764 ( .A(n11065), .B(n11141), .ZN(n11126) );
  INV_X1 U13765 ( .A(n11065), .ZN(n11066) );
  NAND2_X1 U13766 ( .A1(n11066), .A2(n11141), .ZN(n11067) );
  XOR2_X1 U13767 ( .A(n11242), .B(n11241), .Z(n11107) );
  NAND2_X1 U13768 ( .A1(P3_U3897), .A2(n12424), .ZN(n15892) );
  INV_X1 U13769 ( .A(n11069), .ZN(n11068) );
  AND2_X1 U13770 ( .A1(n11068), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12941) );
  INV_X1 U13771 ( .A(n12941), .ZN(n12945) );
  NAND2_X1 U13772 ( .A1(n11702), .A2(n12945), .ZN(n11099) );
  NAND2_X1 U13773 ( .A1(n9602), .A2(n11069), .ZN(n11070) );
  NAND2_X1 U13774 ( .A1(n11070), .A2(n9603), .ZN(n11098) );
  INV_X1 U13775 ( .A(n11098), .ZN(n11071) );
  NAND2_X1 U13776 ( .A1(n11099), .A2(n11071), .ZN(n11083) );
  INV_X1 U13777 ( .A(n11083), .ZN(n11072) );
  NOR2_X1 U13778 ( .A1(n11399), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n13157) );
  INV_X1 U13779 ( .A(n13157), .ZN(n11073) );
  NAND2_X1 U13780 ( .A1(n11085), .A2(n11073), .ZN(n11074) );
  NAND2_X1 U13781 ( .A1(n11074), .A2(n6643), .ZN(n11186) );
  INV_X1 U13782 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n11187) );
  OR2_X1 U13783 ( .A1(n11186), .A2(n11187), .ZN(n11184) );
  NAND2_X1 U13784 ( .A1(n11088), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U13785 ( .A1(n11148), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U13786 ( .A1(n11077), .A2(n11152), .ZN(n11078) );
  NAND2_X1 U13787 ( .A1(n11079), .A2(n11078), .ZN(n11133) );
  INV_X1 U13788 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11080) );
  MUX2_X1 U13789 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n11080), .S(n11094), .Z(
        n11134) );
  NAND2_X1 U13790 ( .A1(n11133), .A2(n11134), .ZN(n11132) );
  NAND2_X1 U13791 ( .A1(n11094), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U13792 ( .A1(n11132), .A2(n11081), .ZN(n11249) );
  XNOR2_X1 U13793 ( .A(n11247), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n11105) );
  MUX2_X1 U13794 ( .A(n11083), .B(n13142), .S(n12942), .Z(n13317) );
  OR2_X1 U13795 ( .A1(n11083), .A2(n11082), .ZN(n13329) );
  XNOR2_X1 U13796 ( .A(n11088), .B(n11783), .ZN(n11112) );
  NAND2_X1 U13797 ( .A1(n13152), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U13798 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  NAND2_X1 U13799 ( .A1(n11086), .A2(n11087), .ZN(n11181) );
  INV_X1 U13800 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U13801 ( .A1(n11183), .A2(n11087), .ZN(n11111) );
  NAND2_X1 U13802 ( .A1(n11112), .A2(n11111), .ZN(n11110) );
  NAND2_X1 U13803 ( .A1(n11088), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11089) );
  NAND2_X1 U13804 ( .A1(n11110), .A2(n11089), .ZN(n11090) );
  NAND2_X1 U13805 ( .A1(n11090), .A2(n11152), .ZN(n11128) );
  NAND2_X1 U13806 ( .A1(n11146), .A2(n11128), .ZN(n11093) );
  INV_X1 U13807 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11092) );
  XNOR2_X1 U13808 ( .A(n11094), .B(n11092), .ZN(n11127) );
  NAND2_X1 U13809 ( .A1(n11094), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13810 ( .A1(n11131), .A2(n11095), .ZN(n11096) );
  NAND2_X1 U13811 ( .A1(n11096), .A2(n11248), .ZN(n11252) );
  OAI21_X1 U13812 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n6768), .A(n11253), .ZN(
        n11102) );
  NAND2_X1 U13813 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n11706) );
  OAI21_X1 U13814 ( .B1(n15898), .B2(n11100), .A(n11706), .ZN(n11101) );
  AOI21_X1 U13815 ( .B1(n15888), .B2(n11102), .A(n11101), .ZN(n11103) );
  OAI21_X1 U13816 ( .B1(n11248), .B2(n13317), .A(n11103), .ZN(n11104) );
  AOI21_X1 U13817 ( .B1(n15895), .B2(n11105), .A(n11104), .ZN(n11106) );
  OAI21_X1 U13818 ( .B1(n11107), .B2(n15892), .A(n11106), .ZN(P3_U3187) );
  XOR2_X1 U13819 ( .A(n11108), .B(n11109), .Z(n11124) );
  OAI21_X1 U13820 ( .B1(n11112), .B2(n11111), .A(n11110), .ZN(n11113) );
  NAND2_X1 U13821 ( .A1(n15888), .A2(n11113), .ZN(n11120) );
  OAI21_X1 U13822 ( .B1(n11116), .B2(n11115), .A(n11114), .ZN(n11117) );
  NAND2_X1 U13823 ( .A1(n15895), .A2(n11117), .ZN(n11119) );
  AOI22_X1 U13824 ( .A1(n15865), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11118) );
  NAND3_X1 U13825 ( .A1(n11120), .A2(n11119), .A3(n11118), .ZN(n11121) );
  AOI21_X1 U13826 ( .B1(n11122), .B2(n15886), .A(n11121), .ZN(n11123) );
  OAI21_X1 U13827 ( .B1(n11124), .B2(n15892), .A(n11123), .ZN(P3_U3184) );
  XOR2_X1 U13828 ( .A(n11125), .B(n11126), .Z(n11143) );
  INV_X1 U13829 ( .A(n11127), .ZN(n11129) );
  NAND3_X1 U13830 ( .A1(n11146), .A2(n11129), .A3(n11128), .ZN(n11130) );
  AOI21_X1 U13831 ( .B1(n11131), .B2(n11130), .A(n13329), .ZN(n11140) );
  INV_X1 U13832 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n11138) );
  OAI21_X1 U13833 ( .B1(n11134), .B2(n11133), .A(n11132), .ZN(n11135) );
  NAND2_X1 U13834 ( .A1(n15895), .A2(n11135), .ZN(n11137) );
  AND2_X1 U13835 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n13061) );
  INV_X1 U13836 ( .A(n13061), .ZN(n11136) );
  OAI211_X1 U13837 ( .C1(n15898), .C2(n11138), .A(n11137), .B(n11136), .ZN(
        n11139) );
  AOI211_X1 U13838 ( .C1(n15886), .C2(n11141), .A(n11140), .B(n11139), .ZN(
        n11142) );
  OAI21_X1 U13839 ( .B1(n11143), .B2(n15892), .A(n11142), .ZN(P3_U3186) );
  XOR2_X1 U13840 ( .A(n11144), .B(n11145), .Z(n11157) );
  OAI21_X1 U13841 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11147), .A(n11146), .ZN(
        n11155) );
  XNOR2_X1 U13842 ( .A(n11148), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U13843 ( .A1(n15895), .A2(n11149), .ZN(n11150) );
  NAND2_X1 U13844 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n12983) );
  OAI211_X1 U13845 ( .C1(n11151), .C2(n15898), .A(n11150), .B(n12983), .ZN(
        n11154) );
  NOR2_X1 U13846 ( .A1(n13317), .A2(n11152), .ZN(n11153) );
  AOI211_X1 U13847 ( .C1(n15888), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11156) );
  OAI21_X1 U13848 ( .B1(n11157), .B2(n15892), .A(n11156), .ZN(P3_U3185) );
  INV_X1 U13849 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11174) );
  OAI22_X1 U13850 ( .A1(n11158), .A2(n14471), .B1(n11327), .B2(n14473), .ZN(
        n15756) );
  AOI22_X1 U13851 ( .A1(n14000), .A2(n15764), .B1(n13992), .B2(n15756), .ZN(
        n11173) );
  XNOR2_X1 U13852 ( .A(n11225), .B(n15764), .ZN(n11159) );
  AND2_X1 U13853 ( .A1(n13862), .A2(n14041), .ZN(n11160) );
  NAND2_X1 U13854 ( .A1(n11159), .A2(n11160), .ZN(n11214) );
  INV_X1 U13855 ( .A(n11214), .ZN(n11220) );
  INV_X1 U13856 ( .A(n11159), .ZN(n11162) );
  INV_X1 U13857 ( .A(n11160), .ZN(n11161) );
  NAND2_X1 U13858 ( .A1(n11162), .A2(n11161), .ZN(n11216) );
  INV_X1 U13859 ( .A(n11216), .ZN(n11163) );
  NOR2_X1 U13860 ( .A1(n11220), .A2(n11163), .ZN(n11170) );
  INV_X1 U13861 ( .A(n11164), .ZN(n11166) );
  INV_X1 U13862 ( .A(n11215), .ZN(n11167) );
  NAND2_X1 U13863 ( .A1(n11168), .A2(n11167), .ZN(n11169) );
  NAND2_X1 U13864 ( .A1(n11169), .A2(n11170), .ZN(n11202) );
  OAI21_X1 U13865 ( .B1(n11170), .B2(n11169), .A(n11202), .ZN(n11171) );
  NAND2_X1 U13866 ( .A1(n11171), .A2(n14004), .ZN(n11172) );
  OAI211_X1 U13867 ( .C1(n11175), .C2(n11174), .A(n11173), .B(n11172), .ZN(
        P2_U3209) );
  INV_X1 U13868 ( .A(n11176), .ZN(n11179) );
  INV_X1 U13869 ( .A(n14173), .ZN(n14165) );
  OAI222_X1 U13870 ( .A1(n12702), .A2(n11177), .B1(n11978), .B2(n11179), .C1(
        n14165), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI222_X1 U13871 ( .A1(P1_U3086), .A2(n11627), .B1(n6554), .B2(n11179), .C1(
        n11178), .C2(n15433), .ZN(P1_U3339) );
  XNOR2_X1 U13872 ( .A(n11180), .B(n13155), .ZN(n11192) );
  INV_X1 U13873 ( .A(n15892), .ZN(n13154) );
  NAND2_X1 U13874 ( .A1(n11181), .A2(n12410), .ZN(n11182) );
  AOI21_X1 U13875 ( .B1(n11183), .B2(n11182), .A(n13329), .ZN(n11191) );
  INV_X1 U13876 ( .A(n11184), .ZN(n11185) );
  AOI21_X1 U13877 ( .B1(n11187), .B2(n11186), .A(n11185), .ZN(n11189) );
  AOI22_X1 U13878 ( .A1(n15865), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11188) );
  OAI21_X1 U13879 ( .B1(n13237), .B2(n11189), .A(n11188), .ZN(n11190) );
  AOI211_X1 U13880 ( .C1(n11192), .C2(n13154), .A(n11191), .B(n11190), .ZN(
        n11193) );
  OAI21_X1 U13881 ( .B1(n11194), .B2(n13317), .A(n11193), .ZN(P3_U3183) );
  INV_X1 U13882 ( .A(n11195), .ZN(n11197) );
  OAI222_X1 U13883 ( .A1(n13725), .A2(n11197), .B1(n13731), .B2(n11196), .C1(
        n13311), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13884 ( .A(n11198), .ZN(n11200) );
  OAI222_X1 U13885 ( .A1(P1_U3086), .A2(n14939), .B1(n6554), .B2(n11200), .C1(
        n11199), .C2(n15433), .ZN(P1_U3338) );
  INV_X1 U13886 ( .A(n14186), .ZN(n14182) );
  OAI222_X1 U13887 ( .A1(n12702), .A2(n11201), .B1(n11978), .B2(n11200), .C1(
        n14182), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13888 ( .A1(n11202), .A2(n11216), .ZN(n11203) );
  XNOR2_X1 U13889 ( .A(n11225), .B(n11370), .ZN(n11223) );
  NAND2_X1 U13890 ( .A1(n13862), .A2(n14040), .ZN(n11221) );
  XNOR2_X1 U13891 ( .A(n11223), .B(n11221), .ZN(n11218) );
  XNOR2_X1 U13892 ( .A(n11203), .B(n11218), .ZN(n11210) );
  NAND2_X1 U13893 ( .A1(n11204), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13990) );
  NAND2_X1 U13894 ( .A1(n14000), .A2(n11370), .ZN(n11208) );
  NAND2_X1 U13895 ( .A1(n14039), .A2(n14494), .ZN(n11206) );
  NAND2_X1 U13896 ( .A1(n14041), .A2(n14496), .ZN(n11205) );
  NAND2_X1 U13897 ( .A1(n11206), .A2(n11205), .ZN(n11377) );
  AOI22_X1 U13898 ( .A1(n13992), .A2(n11377), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n6531), .ZN(n11207) );
  OAI211_X1 U13899 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n13990), .A(n11208), .B(
        n11207), .ZN(n11209) );
  AOI21_X1 U13900 ( .B1(n11210), .B2(n14004), .A(n11209), .ZN(n11211) );
  INV_X1 U13901 ( .A(n11211), .ZN(P2_U3190) );
  INV_X2 U13902 ( .A(P2_U3947), .ZN(n14042) );
  NAND2_X1 U13903 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n14042), .ZN(n11212) );
  OAI21_X1 U13904 ( .B1(n11213), .B2(n14042), .A(n11212), .ZN(P2_U3560) );
  NAND2_X1 U13905 ( .A1(n11215), .A2(n11214), .ZN(n11217) );
  INV_X1 U13906 ( .A(n11221), .ZN(n11222) );
  NAND2_X1 U13907 ( .A1(n11223), .A2(n11222), .ZN(n11224) );
  XNOR2_X1 U13908 ( .A(n13864), .B(n15811), .ZN(n11226) );
  NAND2_X1 U13909 ( .A1(n13862), .A2(n14039), .ZN(n11227) );
  NAND2_X1 U13910 ( .A1(n11226), .A2(n11227), .ZN(n11387) );
  INV_X1 U13911 ( .A(n11226), .ZN(n11229) );
  INV_X1 U13912 ( .A(n11227), .ZN(n11228) );
  NAND2_X1 U13913 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  NAND2_X1 U13914 ( .A1(n11387), .A2(n11230), .ZN(n11234) );
  INV_X1 U13915 ( .A(n11388), .ZN(n11233) );
  AOI21_X1 U13916 ( .B1(n11235), .B2(n11234), .A(n11233), .ZN(n11240) );
  INV_X1 U13917 ( .A(n13990), .ZN(n14011) );
  NAND2_X1 U13918 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(n6531), .ZN(n14070) );
  OAI21_X1 U13919 ( .B1(n14014), .B2(n15811), .A(n14070), .ZN(n11237) );
  OAI22_X1 U13920 ( .A1(n11327), .A2(n13978), .B1(n13950), .B2(n11436), .ZN(
        n11236) );
  AOI211_X1 U13921 ( .C1(n11238), .C2(n14011), .A(n11237), .B(n11236), .ZN(
        n11239) );
  OAI21_X1 U13922 ( .B1(n11240), .B2(n14002), .A(n11239), .ZN(P2_U3202) );
  MUX2_X1 U13923 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13285), .Z(n11272) );
  XNOR2_X1 U13924 ( .A(n11272), .B(n11283), .ZN(n11270) );
  INV_X1 U13925 ( .A(n11243), .ZN(n11245) );
  NAND2_X1 U13926 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  XOR2_X1 U13927 ( .A(n11271), .B(n11270), .Z(n11261) );
  NAND2_X1 U13928 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  INV_X1 U13929 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11251) );
  MUX2_X1 U13930 ( .A(n11251), .B(P3_REG1_REG_6__SCAN_IN), .S(n11283), .Z(
        n11262) );
  XNOR2_X1 U13931 ( .A(n11263), .B(n11262), .ZN(n11259) );
  NAND3_X1 U13932 ( .A1(n11253), .A2(n6771), .A3(n11252), .ZN(n11254) );
  AND2_X1 U13933 ( .A1(n11285), .A2(n11254), .ZN(n11257) );
  NAND2_X1 U13934 ( .A1(n15886), .A2(n11283), .ZN(n11256) );
  AND2_X1 U13935 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n13108) );
  AOI21_X1 U13936 ( .B1(n15865), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n13108), .ZN(
        n11255) );
  OAI211_X1 U13937 ( .C1(n11257), .C2(n13329), .A(n11256), .B(n11255), .ZN(
        n11258) );
  AOI21_X1 U13938 ( .B1(n15895), .B2(n11259), .A(n11258), .ZN(n11260) );
  OAI21_X1 U13939 ( .B1(n11261), .B2(n15892), .A(n11260), .ZN(P3_U3188) );
  XNOR2_X1 U13940 ( .A(n11471), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11469) );
  OR2_X1 U13941 ( .A1(n11283), .A2(n11251), .ZN(n11264) );
  NAND2_X1 U13942 ( .A1(n11265), .A2(n11264), .ZN(n11267) );
  XNOR2_X1 U13943 ( .A(n11267), .B(n11307), .ZN(n11305) );
  NAND2_X1 U13944 ( .A1(n11305), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U13945 ( .A1(n11267), .A2(n11266), .ZN(n11268) );
  XOR2_X1 U13946 ( .A(n11469), .B(n11470), .Z(n11295) );
  NAND2_X1 U13947 ( .A1(n11271), .A2(n11270), .ZN(n11275) );
  INV_X1 U13948 ( .A(n11272), .ZN(n11273) );
  NAND2_X1 U13949 ( .A1(n11273), .A2(n11283), .ZN(n11274) );
  MUX2_X1 U13950 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13285), .Z(n11276) );
  XNOR2_X1 U13951 ( .A(n11276), .B(n11307), .ZN(n11311) );
  NAND2_X1 U13952 ( .A1(n11310), .A2(n11311), .ZN(n11279) );
  INV_X1 U13953 ( .A(n11276), .ZN(n11277) );
  NAND2_X1 U13954 ( .A1(n11277), .A2(n11307), .ZN(n11278) );
  NAND2_X1 U13955 ( .A1(n11279), .A2(n11278), .ZN(n11446) );
  MUX2_X1 U13956 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13285), .Z(n11447) );
  XNOR2_X1 U13957 ( .A(n11447), .B(n11471), .ZN(n11445) );
  XNOR2_X1 U13958 ( .A(n11446), .B(n11445), .ZN(n11293) );
  NAND2_X1 U13959 ( .A1(n15886), .A2(n11471), .ZN(n11280) );
  NAND2_X1 U13960 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n13001) );
  OAI211_X1 U13961 ( .C1(n11281), .C2(n15898), .A(n11280), .B(n13001), .ZN(
        n11292) );
  INV_X1 U13962 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11282) );
  OR2_X1 U13963 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  INV_X1 U13964 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11944) );
  XNOR2_X1 U13965 ( .A(n11471), .B(n11944), .ZN(n11288) );
  INV_X1 U13966 ( .A(n11459), .ZN(n11290) );
  NAND3_X1 U13967 ( .A1(n11287), .A2(n11288), .A3(n7316), .ZN(n11289) );
  AOI21_X1 U13968 ( .B1(n11290), .B2(n11289), .A(n13329), .ZN(n11291) );
  AOI211_X1 U13969 ( .C1(n13154), .C2(n11293), .A(n11292), .B(n11291), .ZN(
        n11294) );
  OAI21_X1 U13970 ( .B1(n11295), .B2(n13237), .A(n11294), .ZN(P3_U3190) );
  AOI211_X1 U13971 ( .C1(n15760), .C2(P2_REG3_REG_0__SCAN_IN), .A(n11298), .B(
        n11297), .ZN(n11300) );
  MUX2_X1 U13972 ( .A(n11300), .B(n11299), .S(n14484), .Z(n11303) );
  NAND2_X1 U13973 ( .A1(n15759), .A2(n11301), .ZN(n11302) );
  OAI211_X1 U13974 ( .C1(n14465), .C2(n11304), .A(n11303), .B(n11302), .ZN(
        P2_U3265) );
  XOR2_X1 U13975 ( .A(n11305), .B(P3_REG1_REG_7__SCAN_IN), .Z(n11317) );
  OAI21_X1 U13976 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n11306), .A(n11287), .ZN(
        n11315) );
  NAND2_X1 U13977 ( .A1(n15886), .A2(n11307), .ZN(n11308) );
  NAND2_X1 U13978 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n12950) );
  OAI211_X1 U13979 ( .C1(n11309), .C2(n15898), .A(n11308), .B(n12950), .ZN(
        n11314) );
  XOR2_X1 U13980 ( .A(n11310), .B(n11311), .Z(n11312) );
  NOR2_X1 U13981 ( .A1(n11312), .A2(n15892), .ZN(n11313) );
  AOI211_X1 U13982 ( .C1(n15888), .C2(n11315), .A(n11314), .B(n11313), .ZN(
        n11316) );
  OAI21_X1 U13983 ( .B1(n11317), .B2(n13237), .A(n11316), .ZN(P3_U3189) );
  XNOR2_X1 U13984 ( .A(n11318), .B(n11326), .ZN(n15809) );
  OAI22_X1 U13985 ( .A1(n14499), .A2(n14073), .B1(n11319), .B2(n14406), .ZN(
        n11323) );
  OAI211_X1 U13986 ( .C1(n8987), .C2(n15811), .A(n10957), .B(n11321), .ZN(
        n15810) );
  NOR2_X1 U13987 ( .A1(n14507), .A2(n15810), .ZN(n11322) );
  AOI211_X1 U13988 ( .C1(n15759), .C2(n11324), .A(n11323), .B(n11322), .ZN(
        n11332) );
  XNOR2_X1 U13989 ( .A(n11325), .B(n11326), .ZN(n11329) );
  OAI22_X1 U13990 ( .A1(n11436), .A2(n14473), .B1(n11327), .B2(n14471), .ZN(
        n11328) );
  AOI21_X1 U13991 ( .B1(n11329), .B2(n15757), .A(n11328), .ZN(n11330) );
  OAI21_X1 U13992 ( .B1(n15809), .B2(n8920), .A(n11330), .ZN(n15812) );
  NAND2_X1 U13993 ( .A1(n15812), .A2(n14499), .ZN(n11331) );
  OAI211_X1 U13994 ( .C1(n15809), .C2(n14488), .A(n11332), .B(n11331), .ZN(
        P2_U3261) );
  XNOR2_X1 U13995 ( .A(n11334), .B(n11333), .ZN(n15785) );
  OAI211_X1 U13996 ( .C1(n11335), .C2(n8535), .A(n10957), .B(n15763), .ZN(
        n15786) );
  OAI22_X1 U13997 ( .A1(n14507), .A2(n15786), .B1(n11336), .B2(n14406), .ZN(
        n11337) );
  AOI21_X1 U13998 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n14484), .A(n11337), .ZN(
        n11346) );
  INV_X1 U13999 ( .A(n11338), .ZN(n11339) );
  NAND2_X1 U14000 ( .A1(n11339), .A2(n9977), .ZN(n11341) );
  NAND2_X1 U14001 ( .A1(n11341), .A2(n11340), .ZN(n11342) );
  NAND2_X1 U14002 ( .A1(n11342), .A2(n15757), .ZN(n11344) );
  AOI22_X1 U14003 ( .A1(n14494), .A2(n14041), .B1(n9670), .B2(n14496), .ZN(
        n11343) );
  NAND2_X1 U14004 ( .A1(n11344), .A2(n11343), .ZN(n15787) );
  AOI22_X1 U14005 ( .A1(n15759), .A2(n8529), .B1(n14499), .B2(n15787), .ZN(
        n11345) );
  OAI211_X1 U14006 ( .C1(n14465), .C2(n15785), .A(n11346), .B(n11345), .ZN(
        P2_U3264) );
  INV_X1 U14007 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11348) );
  OR2_X1 U14008 ( .A1(n11352), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15731) );
  MUX2_X1 U14009 ( .A(n11348), .B(P2_REG2_REG_12__SCAN_IN), .S(n15746), .Z(
        n15732) );
  AOI21_X1 U14010 ( .B1(n15733), .B2(n15731), .A(n15732), .ZN(n15736) );
  AOI21_X1 U14011 ( .B1(n11348), .B2(n11347), .A(n15736), .ZN(n14153) );
  INV_X1 U14012 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11349) );
  MUX2_X1 U14013 ( .A(n11349), .B(P2_REG2_REG_13__SCAN_IN), .S(n14155), .Z(
        n14152) );
  XNOR2_X1 U14014 ( .A(n11565), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11363) );
  NOR2_X1 U14015 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13820), .ZN(n11351) );
  NOR2_X1 U14016 ( .A1(n14206), .A2(n7051), .ZN(n11350) );
  AOI211_X1 U14017 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n15715), .A(n11351), 
        .B(n11350), .ZN(n11362) );
  NAND2_X1 U14018 ( .A1(n11352), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n15737) );
  INV_X1 U14019 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11353) );
  XNOR2_X1 U14020 ( .A(n15746), .B(n11353), .ZN(n15739) );
  AND2_X1 U14021 ( .A1(n15737), .A2(n15739), .ZN(n11354) );
  NAND2_X1 U14022 ( .A1(n15738), .A2(n11354), .ZN(n15742) );
  OR2_X1 U14023 ( .A1(n15746), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14024 ( .A1(n15742), .A2(n11355), .ZN(n14159) );
  INV_X1 U14025 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11356) );
  XNOR2_X1 U14026 ( .A(n14155), .B(n11356), .ZN(n14158) );
  NAND2_X1 U14027 ( .A1(n11357), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11358) );
  NAND2_X1 U14028 ( .A1(n14160), .A2(n11358), .ZN(n11360) );
  INV_X1 U14029 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14584) );
  XNOR2_X1 U14030 ( .A(n11568), .B(n14584), .ZN(n11359) );
  NAND2_X1 U14031 ( .A1(n11360), .A2(n11359), .ZN(n11570) );
  OAI211_X1 U14032 ( .C1(n11360), .C2(n11359), .A(n11570), .B(n15744), .ZN(
        n11361) );
  OAI211_X1 U14033 ( .C1(n11363), .C2(n14197), .A(n11362), .B(n11361), .ZN(
        P2_U3228) );
  INV_X1 U14034 ( .A(SI_19_), .ZN(n11366) );
  INV_X1 U14035 ( .A(n11364), .ZN(n11365) );
  OAI222_X1 U14036 ( .A1(P3_U3151), .A2(n13316), .B1(n13731), .B2(n11366), 
        .C1(n13725), .C2(n11365), .ZN(P3_U3276) );
  INV_X1 U14037 ( .A(n14465), .ZN(n15768) );
  XNOR2_X1 U14038 ( .A(n11368), .B(n11367), .ZN(n15800) );
  OAI211_X1 U14039 ( .C1(n11369), .C2(n15804), .A(n10957), .B(n11320), .ZN(
        n15802) );
  NAND2_X1 U14040 ( .A1(n15759), .A2(n11370), .ZN(n11373) );
  NAND2_X1 U14041 ( .A1(n15760), .A2(n11371), .ZN(n11372) );
  OAI211_X1 U14042 ( .C1(n14507), .C2(n15802), .A(n11373), .B(n11372), .ZN(
        n11374) );
  AOI21_X1 U14043 ( .B1(n15768), .B2(n15800), .A(n11374), .ZN(n11381) );
  XNOR2_X1 U14044 ( .A(n11376), .B(n11375), .ZN(n11378) );
  AOI21_X1 U14045 ( .B1(n11378), .B2(n15757), .A(n11377), .ZN(n15803) );
  MUX2_X1 U14046 ( .A(n11379), .B(n15803), .S(n14499), .Z(n11380) );
  NAND2_X1 U14047 ( .A1(n11381), .A2(n11380), .ZN(P2_U3262) );
  XNOR2_X1 U14048 ( .A(n13864), .B(n11520), .ZN(n11382) );
  NAND2_X1 U14049 ( .A1(n13862), .A2(n14038), .ZN(n11383) );
  NAND2_X1 U14050 ( .A1(n11382), .A2(n11383), .ZN(n11434) );
  INV_X1 U14051 ( .A(n11382), .ZN(n11385) );
  INV_X1 U14052 ( .A(n11383), .ZN(n11384) );
  NAND2_X1 U14053 ( .A1(n11385), .A2(n11384), .ZN(n11386) );
  AND2_X1 U14054 ( .A1(n11434), .A2(n11386), .ZN(n11390) );
  OAI21_X1 U14055 ( .B1(n11390), .B2(n11389), .A(n11435), .ZN(n11397) );
  INV_X1 U14056 ( .A(n11391), .ZN(n11519) );
  NOR2_X1 U14057 ( .A1(n13990), .A2(n11519), .ZN(n11396) );
  NAND2_X1 U14058 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(n6531), .ZN(n14085) );
  NAND2_X1 U14059 ( .A1(n14037), .A2(n14494), .ZN(n11393) );
  NAND2_X1 U14060 ( .A1(n14039), .A2(n14496), .ZN(n11392) );
  NAND2_X1 U14061 ( .A1(n11393), .A2(n11392), .ZN(n11516) );
  NAND2_X1 U14062 ( .A1(n13992), .A2(n11516), .ZN(n11394) );
  OAI211_X1 U14063 ( .C1(n14014), .C2(n11520), .A(n14085), .B(n11394), .ZN(
        n11395) );
  AOI211_X1 U14064 ( .C1(n11397), .C2(n14004), .A(n11396), .B(n11395), .ZN(
        n11398) );
  INV_X1 U14065 ( .A(n11398), .ZN(P2_U3199) );
  MUX2_X1 U14066 ( .A(n11416), .B(n11399), .S(n15951), .Z(n11400) );
  OAI21_X1 U14067 ( .B1(n11401), .B2(n13660), .A(n11400), .ZN(P3_U3459) );
  INV_X1 U14068 ( .A(n11402), .ZN(n11404) );
  OAI222_X1 U14069 ( .A1(n15433), .A2(n11403), .B1(n6554), .B2(n11404), .C1(
        P1_U3086), .C2(n12113), .ZN(P1_U3337) );
  INV_X1 U14070 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11405) );
  OAI222_X1 U14071 ( .A1(n12702), .A2(n11405), .B1(n11978), .B2(n11404), .C1(
        P2_U3088), .C2(n7042), .ZN(P2_U3309) );
  NAND2_X1 U14072 ( .A1(n11690), .A2(n11406), .ZN(n11407) );
  NAND2_X1 U14073 ( .A1(n11407), .A2(n11409), .ZN(n11408) );
  OAI21_X1 U14074 ( .B1(n11410), .B2(n11409), .A(n11408), .ZN(n11411) );
  INV_X1 U14075 ( .A(n11411), .ZN(n11412) );
  NAND2_X1 U14076 ( .A1(n11413), .A2(n11412), .ZN(n11419) );
  OR2_X1 U14077 ( .A1(n15928), .A2(n11417), .ZN(n11414) );
  MUX2_X1 U14078 ( .A(n11416), .B(n11415), .S(n13580), .Z(n11421) );
  INV_X1 U14079 ( .A(n11417), .ZN(n12936) );
  OR2_X1 U14080 ( .A1(n15928), .A2(n12936), .ZN(n11418) );
  AOI22_X1 U14081 ( .A1(n13557), .A2(n15869), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n13579), .ZN(n11420) );
  NAND2_X1 U14082 ( .A1(n11421), .A2(n11420), .ZN(P3_U3233) );
  NAND2_X1 U14083 ( .A1(n11422), .A2(n11423), .ZN(n11425) );
  XNOR2_X1 U14084 ( .A(n11425), .B(n11424), .ZN(n11432) );
  NAND2_X1 U14085 ( .A1(n15388), .A2(n12520), .ZN(n15648) );
  OAI22_X1 U14086 ( .A1(n14808), .A2(n11506), .B1(n15648), .B2(n11647), .ZN(
        n11426) );
  INV_X1 U14087 ( .A(n11426), .ZN(n11429) );
  NOR2_X1 U14088 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11427), .ZN(n14868) );
  AOI21_X1 U14089 ( .B1(n14806), .B2(n15647), .A(n14868), .ZN(n11428) );
  OAI211_X1 U14090 ( .C1(n11430), .C2(n15495), .A(n11429), .B(n11428), .ZN(
        n11431) );
  AOI21_X1 U14091 ( .B1(n11432), .B2(n15491), .A(n11431), .ZN(n11433) );
  INV_X1 U14092 ( .A(n11433), .ZN(P1_U3230) );
  XNOR2_X1 U14093 ( .A(n13864), .B(n11561), .ZN(n11527) );
  NAND2_X1 U14094 ( .A1(n13862), .A2(n14037), .ZN(n11526) );
  XNOR2_X1 U14095 ( .A(n11527), .B(n11526), .ZN(n11525) );
  XNOR2_X1 U14096 ( .A(n11524), .B(n11525), .ZN(n11440) );
  NAND2_X1 U14097 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n6531), .ZN(n14100) );
  OAI21_X1 U14098 ( .B1(n14014), .B2(n11561), .A(n14100), .ZN(n11438) );
  OAI22_X1 U14099 ( .A1(n11436), .A2(n13978), .B1(n13950), .B2(n11873), .ZN(
        n11437) );
  AOI211_X1 U14100 ( .C1(n11559), .C2(n14011), .A(n11438), .B(n11437), .ZN(
        n11439) );
  OAI21_X1 U14101 ( .B1(n11440), .B2(n14002), .A(n11439), .ZN(P2_U3211) );
  INV_X1 U14102 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11441) );
  INV_X1 U14103 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12175) );
  MUX2_X1 U14104 ( .A(n11441), .B(n12175), .S(n13285), .Z(n11442) );
  INV_X1 U14105 ( .A(n11756), .ZN(n11468) );
  NAND2_X1 U14106 ( .A1(n11442), .A2(n11468), .ZN(n11760) );
  INV_X1 U14107 ( .A(n11442), .ZN(n11443) );
  NAND2_X1 U14108 ( .A1(n11443), .A2(n11756), .ZN(n11444) );
  NAND2_X1 U14109 ( .A1(n11760), .A2(n11444), .ZN(n11455) );
  NAND2_X1 U14110 ( .A1(n11446), .A2(n11445), .ZN(n11450) );
  INV_X1 U14111 ( .A(n11447), .ZN(n11448) );
  NAND2_X1 U14112 ( .A1(n11448), .A2(n11471), .ZN(n11449) );
  INV_X1 U14113 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12076) );
  INV_X1 U14114 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12172) );
  MUX2_X1 U14115 ( .A(n12076), .B(n12172), .S(n13285), .Z(n11451) );
  INV_X1 U14116 ( .A(n11472), .ZN(n15887) );
  AND2_X1 U14117 ( .A1(n11451), .A2(n15887), .ZN(n15880) );
  INV_X1 U14118 ( .A(n11451), .ZN(n11452) );
  NAND2_X1 U14119 ( .A1(n11452), .A2(n11472), .ZN(n15881) );
  INV_X1 U14120 ( .A(n11761), .ZN(n11453) );
  AOI21_X1 U14121 ( .B1(n11455), .B2(n11454), .A(n11453), .ZN(n11479) );
  NAND2_X1 U14122 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12259)
         );
  OAI21_X1 U14123 ( .B1(n15898), .B2(n11456), .A(n12259), .ZN(n11467) );
  INV_X1 U14124 ( .A(n11461), .ZN(n11463) );
  XNOR2_X1 U14125 ( .A(n11756), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11464) );
  NAND3_X1 U14126 ( .A1(n11462), .A2(n11464), .A3(n11463), .ZN(n11465) );
  AOI21_X1 U14127 ( .B1(n6635), .B2(n11465), .A(n13329), .ZN(n11466) );
  AOI211_X1 U14128 ( .C1(n15886), .C2(n11468), .A(n11467), .B(n11466), .ZN(
        n11478) );
  NAND2_X1 U14129 ( .A1(n15879), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11475) );
  NAND2_X1 U14130 ( .A1(n11473), .A2(n11472), .ZN(n11474) );
  NAND2_X1 U14131 ( .A1(n11475), .A2(n11474), .ZN(n11755) );
  XNOR2_X1 U14132 ( .A(n11756), .B(n12175), .ZN(n11754) );
  XNOR2_X1 U14133 ( .A(n11755), .B(n11754), .ZN(n11476) );
  NAND2_X1 U14134 ( .A1(n11476), .A2(n15895), .ZN(n11477) );
  OAI211_X1 U14135 ( .C1(n11479), .C2(n15892), .A(n11478), .B(n11477), .ZN(
        P3_U3192) );
  INV_X1 U14136 ( .A(n11480), .ZN(n11537) );
  OAI222_X1 U14137 ( .A1(n15433), .A2(n11481), .B1(n6554), .B2(n11537), .C1(
        n15207), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U14138 ( .A(n11482), .ZN(n11483) );
  OAI222_X1 U14139 ( .A1(P3_U3151), .A2(n11659), .B1(n13731), .B2(n11484), 
        .C1(n13725), .C2(n11483), .ZN(P3_U3275) );
  XNOR2_X1 U14140 ( .A(n11486), .B(n12652), .ZN(n15636) );
  XNOR2_X1 U14141 ( .A(n11487), .B(n12652), .ZN(n11488) );
  NOR2_X1 U14142 ( .A1(n11488), .A2(n15651), .ZN(n15634) );
  OR2_X1 U14143 ( .A1(n15584), .A2(n15628), .ZN(n15196) );
  NAND2_X1 U14144 ( .A1(n15565), .A2(n11489), .ZN(n11490) );
  NAND2_X1 U14145 ( .A1(n11490), .A2(n15540), .ZN(n11491) );
  OR2_X1 U14146 ( .A1(n11491), .A2(n15554), .ZN(n15627) );
  INV_X1 U14147 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14838) );
  OAI22_X1 U14148 ( .A1(n15185), .A2(n15627), .B1(n14838), .B2(n15549), .ZN(
        n11492) );
  INV_X1 U14149 ( .A(n11492), .ZN(n11494) );
  NAND2_X1 U14150 ( .A1(n15584), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n11493) );
  OAI211_X1 U14151 ( .C1(n15196), .C2(n15629), .A(n11494), .B(n11493), .ZN(
        n11496) );
  OAI22_X1 U14152 ( .A1(n6804), .A2(n15162), .B1(n15552), .B2(n12508), .ZN(
        n11495) );
  AOI211_X1 U14153 ( .C1(n15634), .C2(n15178), .A(n11496), .B(n11495), .ZN(
        n11497) );
  OAI21_X1 U14154 ( .B1(n15214), .B2(n15636), .A(n11497), .ZN(P1_U3291) );
  NAND2_X1 U14155 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  XOR2_X1 U14156 ( .A(n12655), .B(n11500), .Z(n15675) );
  XNOR2_X1 U14157 ( .A(n12655), .B(n11501), .ZN(n11502) );
  NAND2_X1 U14158 ( .A1(n11502), .A2(n15568), .ZN(n15673) );
  MUX2_X1 U14159 ( .A(n11503), .B(n15673), .S(n15178), .Z(n11511) );
  OAI21_X1 U14160 ( .B1(n6753), .B2(n11507), .A(n15540), .ZN(n11504) );
  NOR2_X1 U14161 ( .A1(n11504), .A2(n15523), .ZN(n15669) );
  INV_X1 U14162 ( .A(n11505), .ZN(n11649) );
  OAI22_X1 U14163 ( .A1(n15162), .A2(n11506), .B1(n11649), .B2(n15549), .ZN(
        n11509) );
  OAI22_X1 U14164 ( .A1(n11507), .A2(n15552), .B1(n15196), .B2(n11652), .ZN(
        n11508) );
  AOI211_X1 U14165 ( .C1(n15582), .C2(n15669), .A(n11509), .B(n11508), .ZN(
        n11510) );
  OAI211_X1 U14166 ( .C1(n15675), .C2(n15214), .A(n11511), .B(n11510), .ZN(
        P1_U3287) );
  INV_X1 U14167 ( .A(n11513), .ZN(n11514) );
  XNOR2_X1 U14168 ( .A(n11512), .B(n11514), .ZN(n15816) );
  XNOR2_X1 U14169 ( .A(n11515), .B(n11514), .ZN(n11517) );
  AOI21_X1 U14170 ( .B1(n11517), .B2(n15757), .A(n11516), .ZN(n15823) );
  MUX2_X1 U14171 ( .A(n14088), .B(n15823), .S(n14499), .Z(n11523) );
  AOI21_X1 U14172 ( .B1(n11321), .B2(n15819), .A(n14482), .ZN(n11518) );
  AND2_X1 U14173 ( .A1(n11558), .A2(n11518), .ZN(n15821) );
  OAI22_X1 U14174 ( .A1(n14486), .A2(n11520), .B1(n14406), .B2(n11519), .ZN(
        n11521) );
  AOI21_X1 U14175 ( .B1(n15767), .B2(n15821), .A(n11521), .ZN(n11522) );
  OAI211_X1 U14176 ( .C1(n14465), .C2(n15816), .A(n11523), .B(n11522), .ZN(
        P2_U3260) );
  OR2_X1 U14177 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  XNOR2_X1 U14178 ( .A(n15834), .B(n13799), .ZN(n11858) );
  NOR2_X1 U14179 ( .A1(n11873), .A2(n13800), .ZN(n11859) );
  XNOR2_X1 U14180 ( .A(n11858), .B(n11859), .ZN(n11856) );
  XNOR2_X1 U14181 ( .A(n11857), .B(n11856), .ZN(n11533) );
  OAI22_X1 U14182 ( .A1(n13950), .A2(n13939), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8609), .ZN(n11531) );
  INV_X1 U14183 ( .A(n11529), .ZN(n11740) );
  OAI22_X1 U14184 ( .A1(n13978), .A2(n11734), .B1(n13990), .B2(n11740), .ZN(
        n11530) );
  AOI211_X1 U14185 ( .C1(n15834), .C2(n14000), .A(n11531), .B(n11530), .ZN(
        n11532) );
  OAI21_X1 U14186 ( .B1(n11533), .B2(n14002), .A(n11532), .ZN(P2_U3185) );
  INV_X1 U14187 ( .A(n11534), .ZN(n11535) );
  OAI222_X1 U14188 ( .A1(P3_U3151), .A2(n12801), .B1(n13731), .B2(n11536), 
        .C1(n13725), .C2(n11535), .ZN(P3_U3274) );
  OAI222_X1 U14189 ( .A1(n14659), .A2(n11538), .B1(P2_U3088), .B2(n6547), .C1(
        n11978), .C2(n11537), .ZN(P2_U3308) );
  INV_X1 U14190 ( .A(n11546), .ZN(n11541) );
  NAND2_X1 U14191 ( .A1(n14666), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11539) );
  OAI211_X1 U14192 ( .C1(n11541), .C2(n11978), .A(n11540), .B(n11539), .ZN(
        P2_U3304) );
  INV_X1 U14193 ( .A(n11542), .ZN(n11544) );
  OAI22_X1 U14194 ( .A1(n12946), .A2(P3_U3151), .B1(SI_22_), .B2(n11854), .ZN(
        n11543) );
  AOI21_X1 U14195 ( .B1(n11544), .B2(n11851), .A(n11543), .ZN(P3_U3273) );
  NAND2_X1 U14196 ( .A1(n11546), .A2(n11545), .ZN(n11547) );
  OAI211_X1 U14197 ( .C1(n11548), .C2(n15433), .A(n11547), .B(n12701), .ZN(
        P1_U3332) );
  XOR2_X1 U14198 ( .A(n11549), .B(n11552), .Z(n15830) );
  NAND2_X1 U14199 ( .A1(n11551), .A2(n11550), .ZN(n11553) );
  INV_X1 U14200 ( .A(n11553), .ZN(n11555) );
  INV_X1 U14201 ( .A(n11552), .ZN(n11554) );
  NOR2_X1 U14202 ( .A1(n11553), .A2(n11552), .ZN(n11730) );
  INV_X1 U14203 ( .A(n11730), .ZN(n11727) );
  OAI21_X1 U14204 ( .B1(n11555), .B2(n11554), .A(n11727), .ZN(n11556) );
  AOI222_X1 U14205 ( .A1(n11556), .A2(n15757), .B1(n14038), .B2(n14496), .C1(
        n14036), .C2(n14494), .ZN(n15829) );
  MUX2_X1 U14206 ( .A(n11557), .B(n15829), .S(n14499), .Z(n11564) );
  AOI211_X1 U14207 ( .C1(n15827), .C2(n11558), .A(n14482), .B(n11737), .ZN(
        n15826) );
  INV_X1 U14208 ( .A(n11559), .ZN(n11560) );
  OAI22_X1 U14209 ( .A1(n14486), .A2(n11561), .B1(n14406), .B2(n11560), .ZN(
        n11562) );
  AOI21_X1 U14210 ( .B1(n15826), .B2(n14457), .A(n11562), .ZN(n11563) );
  OAI211_X1 U14211 ( .C1(n14465), .C2(n15830), .A(n11564), .B(n11563), .ZN(
        P2_U3259) );
  XNOR2_X1 U14212 ( .A(n11958), .B(n11964), .ZN(n11960) );
  XNOR2_X1 U14213 ( .A(n11960), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11575) );
  NOR2_X1 U14214 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14008), .ZN(n11567) );
  NOR2_X1 U14215 ( .A1(n14206), .A2(n11571), .ZN(n11566) );
  AOI211_X1 U14216 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n15715), .A(n11567), 
        .B(n11566), .ZN(n11574) );
  NAND2_X1 U14217 ( .A1(n11568), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14218 ( .A1(n11570), .A2(n11569), .ZN(n11965) );
  XNOR2_X1 U14219 ( .A(n11965), .B(n11571), .ZN(n11572) );
  NAND2_X1 U14220 ( .A1(n11572), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11967) );
  OAI211_X1 U14221 ( .C1(n11572), .C2(P2_REG1_REG_15__SCAN_IN), .A(n11967), 
        .B(n15744), .ZN(n11573) );
  OAI211_X1 U14222 ( .C1(n11575), .C2(n14197), .A(n11574), .B(n11573), .ZN(
        P2_U3229) );
  OAI21_X1 U14223 ( .B1(n15584), .B2(n11576), .A(n15552), .ZN(n11578) );
  NAND2_X1 U14224 ( .A1(n15095), .A2(n15214), .ZN(n11577) );
  AOI22_X1 U14225 ( .A1(n12490), .A2(n11578), .B1(n11577), .B2(n12650), .ZN(
        n11580) );
  INV_X1 U14226 ( .A(n15549), .ZN(n15573) );
  AOI22_X1 U14227 ( .A1(n15584), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n15573), .ZN(n11579) );
  OAI211_X1 U14228 ( .C1(n6804), .C2(n15196), .A(n11580), .B(n11579), .ZN(
        P1_U3293) );
  XNOR2_X1 U14229 ( .A(n11581), .B(n11582), .ZN(n15846) );
  INV_X1 U14230 ( .A(n15846), .ZN(n11594) );
  XNOR2_X1 U14231 ( .A(n11583), .B(n11582), .ZN(n11586) );
  OAI22_X1 U14232 ( .A1(n11873), .A2(n14471), .B1(n13839), .B2(n14473), .ZN(
        n11584) );
  INV_X1 U14233 ( .A(n11584), .ZN(n11585) );
  OAI21_X1 U14234 ( .B1(n11586), .B2(n14461), .A(n11585), .ZN(n11587) );
  AOI21_X1 U14235 ( .B1(n15846), .B2(n15818), .A(n11587), .ZN(n15848) );
  MUX2_X1 U14236 ( .A(n11588), .B(n15848), .S(n14499), .Z(n11593) );
  AOI21_X1 U14237 ( .B1(n11738), .B2(n6607), .A(n14482), .ZN(n11589) );
  AND2_X1 U14238 ( .A1(n11589), .A2(n11989), .ZN(n15841) );
  INV_X1 U14239 ( .A(n11590), .ZN(n11872) );
  OAI22_X1 U14240 ( .A1(n14486), .A2(n8988), .B1(n14406), .B2(n11872), .ZN(
        n11591) );
  AOI21_X1 U14241 ( .B1(n15767), .B2(n15841), .A(n11591), .ZN(n11592) );
  OAI211_X1 U14242 ( .C1(n11594), .C2(n14488), .A(n11593), .B(n11592), .ZN(
        P2_U3257) );
  XNOR2_X1 U14243 ( .A(n11595), .B(n11596), .ZN(n11602) );
  NAND2_X1 U14244 ( .A1(n12548), .A2(n15388), .ZN(n15692) );
  NOR2_X1 U14245 ( .A1(n11647), .A2(n15692), .ZN(n11601) );
  AOI21_X1 U14246 ( .B1(n14806), .B2(n15667), .A(n11597), .ZN(n11599) );
  OR2_X1 U14247 ( .A1(n14808), .A2(n15377), .ZN(n11598) );
  OAI211_X1 U14248 ( .C1(n15495), .C2(n11614), .A(n11599), .B(n11598), .ZN(
        n11600) );
  AOI211_X1 U14249 ( .C1(n11602), .C2(n15491), .A(n11601), .B(n11600), .ZN(
        n11603) );
  INV_X1 U14250 ( .A(n11603), .ZN(P1_U3221) );
  INV_X1 U14251 ( .A(n11604), .ZN(n11607) );
  OAI222_X1 U14252 ( .A1(n12702), .A2(n11606), .B1(n11978), .B2(n11607), .C1(
        n11605), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI222_X1 U14253 ( .A1(n15433), .A2(n11608), .B1(n6554), .B2(n11607), .C1(
        P1_U3086), .C2(n12430), .ZN(P1_U3335) );
  XNOR2_X1 U14254 ( .A(n11609), .B(n12658), .ZN(n15695) );
  XNOR2_X1 U14255 ( .A(n11610), .B(n12658), .ZN(n11611) );
  AOI222_X1 U14256 ( .A1(n11611), .A2(n15568), .B1(n15667), .B2(n15665), .C1(
        n14821), .C2(n15668), .ZN(n15690) );
  MUX2_X1 U14257 ( .A(n11612), .B(n15690), .S(n15178), .Z(n11618) );
  INV_X1 U14258 ( .A(n11912), .ZN(n11613) );
  AOI211_X1 U14259 ( .C1(n12548), .C2(n15522), .A(n15574), .B(n11613), .ZN(
        n15691) );
  INV_X1 U14260 ( .A(n12548), .ZN(n11615) );
  OAI22_X1 U14261 ( .A1(n15552), .A2(n11615), .B1(n11614), .B2(n15549), .ZN(
        n11616) );
  AOI21_X1 U14262 ( .B1(n15691), .B2(n15582), .A(n11616), .ZN(n11617) );
  OAI211_X1 U14263 ( .C1(n15214), .C2(n15695), .A(n11618), .B(n11617), .ZN(
        P1_U3285) );
  NAND2_X1 U14264 ( .A1(n11630), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14265 ( .A1(n11620), .A2(n11619), .ZN(n11622) );
  XNOR2_X1 U14266 ( .A(n11622), .B(n11621), .ZN(n15498) );
  INV_X1 U14267 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15497) );
  NAND2_X1 U14268 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  INV_X1 U14269 ( .A(n11621), .ZN(n15502) );
  OR2_X1 U14270 ( .A1(n11622), .A2(n15502), .ZN(n11624) );
  XNOR2_X1 U14271 ( .A(n11627), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n11623) );
  AOI21_X1 U14272 ( .B1(n15496), .B2(n11624), .A(n11623), .ZN(n11643) );
  AND2_X1 U14273 ( .A1(n11624), .A2(n11623), .ZN(n11625) );
  NAND2_X1 U14274 ( .A1(n15496), .A2(n11625), .ZN(n14942) );
  NAND2_X1 U14275 ( .A1(n14942), .A2(n15505), .ZN(n11642) );
  INV_X1 U14276 ( .A(n11627), .ZN(n12108) );
  NAND2_X1 U14277 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14726)
         );
  OAI21_X1 U14278 ( .B1(n15509), .B2(n10012), .A(n14726), .ZN(n11640) );
  INV_X1 U14279 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11626) );
  XNOR2_X1 U14280 ( .A(n11627), .B(n11626), .ZN(n11638) );
  AND2_X1 U14281 ( .A1(n11630), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11628) );
  OR2_X1 U14282 ( .A1(n11630), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U14283 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  INV_X1 U14284 ( .A(n11633), .ZN(n11635) );
  XNOR2_X1 U14285 ( .A(n11633), .B(n15502), .ZN(n15500) );
  INV_X1 U14286 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U14287 ( .A1(n15500), .A2(n15499), .ZN(n11634) );
  OAI21_X1 U14288 ( .B1(n15502), .B2(n11635), .A(n11634), .ZN(n11637) );
  INV_X1 U14289 ( .A(n12110), .ZN(n11636) );
  AOI211_X1 U14290 ( .C1(n11638), .C2(n11637), .A(n14962), .B(n11636), .ZN(
        n11639) );
  AOI211_X1 U14291 ( .C1(n15501), .C2(n12108), .A(n11640), .B(n11639), .ZN(
        n11641) );
  OAI21_X1 U14292 ( .B1(n11643), .B2(n11642), .A(n11641), .ZN(P1_U3259) );
  XNOR2_X1 U14293 ( .A(n11644), .B(n11645), .ZN(n11841) );
  XNOR2_X1 U14294 ( .A(n11841), .B(n11646), .ZN(n11655) );
  NAND2_X1 U14295 ( .A1(n15388), .A2(n12530), .ZN(n15671) );
  NOR2_X1 U14296 ( .A1(n11647), .A2(n15671), .ZN(n11654) );
  AOI21_X1 U14297 ( .B1(n14806), .B2(n15666), .A(n11648), .ZN(n11651) );
  OR2_X1 U14298 ( .A1(n15495), .A2(n11649), .ZN(n11650) );
  OAI211_X1 U14299 ( .C1(n11652), .C2(n14808), .A(n11651), .B(n11650), .ZN(
        n11653) );
  AOI211_X1 U14300 ( .C1(n11655), .C2(n15491), .A(n11654), .B(n11653), .ZN(
        n11656) );
  INV_X1 U14301 ( .A(n11656), .ZN(P1_U3239) );
  NAND2_X4 U14302 ( .A1(n11662), .A2(n6613), .ZN(n12385) );
  NAND2_X1 U14303 ( .A1(n15866), .A2(n12407), .ZN(n11666) );
  OAI21_X1 U14304 ( .B1(n12385), .B2(n11668), .A(n11667), .ZN(n11669) );
  NAND2_X1 U14305 ( .A1(n11747), .A2(n6682), .ZN(n11716) );
  XNOR2_X1 U14306 ( .A(n11670), .B(n12385), .ZN(n11673) );
  INV_X1 U14307 ( .A(n11671), .ZN(n11672) );
  XNOR2_X1 U14308 ( .A(n11673), .B(n11671), .ZN(n11717) );
  INV_X1 U14309 ( .A(n11673), .ZN(n11674) );
  NAND2_X1 U14310 ( .A1(n11674), .A2(n11671), .ZN(n11675) );
  NAND2_X1 U14311 ( .A1(n11715), .A2(n11675), .ZN(n12980) );
  XNOR2_X1 U14312 ( .A(n12385), .B(n15913), .ZN(n11677) );
  XNOR2_X1 U14313 ( .A(n11677), .B(n13150), .ZN(n12979) );
  NAND2_X1 U14314 ( .A1(n11677), .A2(n13150), .ZN(n11678) );
  XNOR2_X1 U14315 ( .A(n12385), .B(n15918), .ZN(n11679) );
  XNOR2_X1 U14316 ( .A(n11679), .B(n11803), .ZN(n13059) );
  INV_X1 U14317 ( .A(n11679), .ZN(n11680) );
  NAND2_X1 U14318 ( .A1(n11680), .A2(n11803), .ZN(n11681) );
  XNOR2_X1 U14319 ( .A(n12385), .B(n11682), .ZN(n12179) );
  XNOR2_X1 U14320 ( .A(n12179), .B(n12180), .ZN(n12177) );
  XOR2_X1 U14321 ( .A(n12178), .B(n12177), .Z(n11712) );
  NAND2_X1 U14322 ( .A1(n11687), .A2(n15928), .ZN(n11684) );
  OAI22_X1 U14323 ( .A1(n11688), .A2(n11684), .B1(n11697), .B2(n11683), .ZN(
        n11686) );
  NAND2_X1 U14324 ( .A1(n11688), .A2(n11687), .ZN(n11693) );
  NAND2_X1 U14325 ( .A1(n11697), .A2(n11689), .ZN(n11691) );
  NAND4_X1 U14326 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11694) );
  NAND2_X1 U14327 ( .A1(n11694), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11696) );
  INV_X1 U14328 ( .A(n11698), .ZN(n12943) );
  NAND2_X1 U14329 ( .A1(n12943), .A2(n11697), .ZN(n11695) );
  NAND2_X1 U14330 ( .A1(n11696), .A2(n11695), .ZN(n11719) );
  OR2_X2 U14331 ( .A1(n11719), .A2(n12941), .ZN(n13133) );
  INV_X1 U14332 ( .A(n11701), .ZN(n11699) );
  INV_X1 U14333 ( .A(n11803), .ZN(n13149) );
  NAND2_X1 U14334 ( .A1(n13130), .A2(n13149), .ZN(n11709) );
  NOR2_X1 U14335 ( .A1(n11702), .A2(n15928), .ZN(n11703) );
  NAND2_X1 U14336 ( .A1(n11704), .A2(n11703), .ZN(n11705) );
  INV_X1 U14337 ( .A(n11706), .ZN(n11707) );
  AOI21_X1 U14338 ( .B1(n15870), .B2(n15923), .A(n11707), .ZN(n11708) );
  OAI211_X1 U14339 ( .C1(n15874), .C2(n12183), .A(n11709), .B(n11708), .ZN(
        n11710) );
  AOI21_X1 U14340 ( .B1(n11808), .B2(n13133), .A(n11710), .ZN(n11711) );
  OAI21_X1 U14341 ( .B1(n11712), .B2(n15867), .A(n11711), .ZN(P3_U3167) );
  NAND2_X1 U14342 ( .A1(n13119), .A2(P3_U3897), .ZN(n11713) );
  OAI21_X1 U14343 ( .B1(P3_U3897), .B2(n11714), .A(n11713), .ZN(P3_U3516) );
  OAI21_X1 U14344 ( .B1(n11717), .B2(n11716), .A(n11715), .ZN(n11724) );
  NOR2_X1 U14345 ( .A1(n11719), .A2(n11718), .ZN(n15878) );
  INV_X1 U14346 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11722) );
  INV_X1 U14347 ( .A(n15874), .ZN(n13111) );
  AOI22_X1 U14348 ( .A1(n13111), .A2(n13150), .B1(n12809), .B2(n15870), .ZN(
        n11721) );
  NAND2_X1 U14349 ( .A1(n13130), .A2(n15866), .ZN(n11720) );
  OAI211_X1 U14350 ( .C1(n15878), .C2(n11722), .A(n11721), .B(n11720), .ZN(
        n11723) );
  AOI21_X1 U14351 ( .B1(n11724), .B2(n13128), .A(n11723), .ZN(n11725) );
  INV_X1 U14352 ( .A(n11725), .ZN(P3_U3177) );
  XOR2_X1 U14353 ( .A(n11726), .B(n11733), .Z(n15838) );
  NAND2_X1 U14354 ( .A1(n11727), .A2(n11728), .ZN(n11732) );
  INV_X1 U14355 ( .A(n11728), .ZN(n11729) );
  NOR3_X1 U14356 ( .A1(n11730), .A2(n11729), .A3(n11733), .ZN(n11731) );
  AOI211_X1 U14357 ( .C1(n11733), .C2(n11732), .A(n14461), .B(n11731), .ZN(
        n11736) );
  OAI22_X1 U14358 ( .A1(n13939), .A2(n14473), .B1(n11734), .B2(n14471), .ZN(
        n11735) );
  NOR2_X1 U14359 ( .A1(n11736), .A2(n11735), .ZN(n15837) );
  MUX2_X1 U14360 ( .A(n14116), .B(n15837), .S(n14499), .Z(n11744) );
  INV_X1 U14361 ( .A(n11737), .ZN(n11739) );
  AOI211_X1 U14362 ( .C1(n15834), .C2(n11739), .A(n14482), .B(n8989), .ZN(
        n15833) );
  OAI22_X1 U14363 ( .A1(n14486), .A2(n11741), .B1(n14406), .B2(n11740), .ZN(
        n11742) );
  AOI21_X1 U14364 ( .B1(n15833), .B2(n14457), .A(n11742), .ZN(n11743) );
  OAI211_X1 U14365 ( .C1(n14465), .C2(n15838), .A(n11744), .B(n11743), .ZN(
        P2_U3258) );
  INV_X1 U14366 ( .A(n12802), .ZN(n11745) );
  NAND3_X1 U14367 ( .A1(n12385), .A2(n11745), .A3(n12798), .ZN(n11746) );
  OAI211_X1 U14368 ( .C1(n11748), .C2(n12403), .A(n11747), .B(n11746), .ZN(
        n11752) );
  AOI22_X1 U14369 ( .A1(n13111), .A2(n11672), .B1(n12407), .B2(n15870), .ZN(
        n11750) );
  NAND2_X1 U14370 ( .A1(n13130), .A2(n11047), .ZN(n11749) );
  OAI211_X1 U14371 ( .C1(n15878), .C2(n12408), .A(n11750), .B(n11749), .ZN(
        n11751) );
  AOI21_X1 U14372 ( .B1(n11752), .B2(n13128), .A(n11751), .ZN(n11753) );
  INV_X1 U14373 ( .A(n11753), .ZN(P3_U3162) );
  INV_X1 U14374 ( .A(n11765), .ZN(n11928) );
  NAND2_X1 U14375 ( .A1(n11758), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n11924) );
  OAI21_X1 U14376 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11758), .A(n11924), 
        .ZN(n11759) );
  NAND2_X1 U14377 ( .A1(n11759), .A2(n15888), .ZN(n11769) );
  MUX2_X1 U14378 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13285), .Z(n11927) );
  XNOR2_X1 U14379 ( .A(n11927), .B(n11928), .ZN(n11762) );
  OAI21_X1 U14380 ( .B1(n11763), .B2(n11762), .A(n11933), .ZN(n11767) );
  NAND2_X1 U14381 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13088)
         );
  NAND2_X1 U14382 ( .A1(n15865), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11764) );
  OAI211_X1 U14383 ( .C1(n13317), .C2(n11765), .A(n13088), .B(n11764), .ZN(
        n11766) );
  AOI21_X1 U14384 ( .B1(n11767), .B2(n13154), .A(n11766), .ZN(n11768) );
  OAI211_X1 U14385 ( .C1(n11770), .C2(n13237), .A(n11769), .B(n11768), .ZN(
        P3_U3193) );
  INV_X1 U14386 ( .A(n11771), .ZN(n11773) );
  OAI222_X1 U14387 ( .A1(n14659), .A2(n11774), .B1(n11978), .B2(n11773), .C1(
        n11772), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U14388 ( .A(n11775), .B(n12804), .ZN(n15907) );
  NAND2_X1 U14389 ( .A1(n12936), .A2(n12755), .ZN(n12081) );
  INV_X1 U14390 ( .A(n12081), .ZN(n11776) );
  NAND2_X1 U14391 ( .A1(n12809), .A2(n15936), .ZN(n15908) );
  NOR2_X1 U14392 ( .A1(n15908), .A2(n12936), .ZN(n11781) );
  OAI21_X1 U14393 ( .B1(n11777), .B2(n12804), .A(n11793), .ZN(n11778) );
  NAND2_X1 U14394 ( .A1(n11778), .A2(n13562), .ZN(n11780) );
  AOI22_X1 U14395 ( .A1(n13567), .A2(n15866), .B1(n13150), .B2(n13566), .ZN(
        n11779) );
  OAI211_X1 U14396 ( .C1(n15907), .C2(n13433), .A(n11780), .B(n11779), .ZN(
        n15909) );
  AOI211_X1 U14397 ( .C1(n13579), .C2(P3_REG3_REG_2__SCAN_IN), .A(n11781), .B(
        n15909), .ZN(n11782) );
  MUX2_X1 U14398 ( .A(n11783), .B(n11782), .S(n13585), .Z(n11784) );
  OAI21_X1 U14399 ( .B1(n15907), .B2(n13436), .A(n11784), .ZN(P3_U3231) );
  OR2_X1 U14400 ( .A1(n11785), .A2(n11790), .ZN(n11786) );
  NAND2_X1 U14401 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  INV_X1 U14402 ( .A(n11788), .ZN(n15914) );
  INV_X1 U14403 ( .A(n13433), .ZN(n13413) );
  NAND2_X1 U14404 ( .A1(n11788), .A2(n13413), .ZN(n11798) );
  NAND2_X1 U14405 ( .A1(n11793), .A2(n11789), .ZN(n11791) );
  NAND2_X1 U14406 ( .A1(n11791), .A2(n11790), .ZN(n11794) );
  NAND2_X1 U14407 ( .A1(n11793), .A2(n11792), .ZN(n11830) );
  NAND3_X1 U14408 ( .A1(n11794), .A2(n13562), .A3(n11830), .ZN(n11797) );
  OAI22_X1 U14409 ( .A1(n11671), .A2(n13509), .B1(n11803), .B2(n13511), .ZN(
        n11795) );
  INV_X1 U14410 ( .A(n11795), .ZN(n11796) );
  NAND3_X1 U14411 ( .A1(n11798), .A2(n11797), .A3(n11796), .ZN(n15915) );
  MUX2_X1 U14412 ( .A(n15915), .B(P3_REG2_REG_3__SCAN_IN), .S(n13580), .Z(
        n11799) );
  INV_X1 U14413 ( .A(n11799), .ZN(n11801) );
  AOI22_X1 U14414 ( .A1(n13557), .A2(n12985), .B1(n13579), .B2(n9082), .ZN(
        n11800) );
  OAI211_X1 U14415 ( .C1(n15914), .C2(n13436), .A(n11801), .B(n11800), .ZN(
        P3_U3230) );
  XNOR2_X1 U14416 ( .A(n11802), .B(n12821), .ZN(n15924) );
  INV_X1 U14417 ( .A(n15924), .ZN(n11811) );
  OAI22_X1 U14418 ( .A1(n11803), .A2(n13509), .B1(n12183), .B2(n13511), .ZN(
        n11807) );
  NAND2_X1 U14419 ( .A1(n11804), .A2(n12821), .ZN(n11805) );
  AOI21_X1 U14420 ( .B1(n11819), .B2(n11805), .A(n13507), .ZN(n11806) );
  AOI211_X1 U14421 ( .C1(n15924), .C2(n13413), .A(n11807), .B(n11806), .ZN(
        n15926) );
  MUX2_X1 U14422 ( .A(n7341), .B(n15926), .S(n13585), .Z(n11810) );
  AOI22_X1 U14423 ( .A1(n13557), .A2(n15923), .B1(n13579), .B2(n11808), .ZN(
        n11809) );
  OAI211_X1 U14424 ( .C1(n11811), .C2(n13436), .A(n11810), .B(n11809), .ZN(
        P3_U3228) );
  OR2_X1 U14425 ( .A1(n11812), .A2(n12765), .ZN(n11813) );
  NAND2_X1 U14426 ( .A1(n11814), .A2(n11813), .ZN(n11820) );
  INV_X1 U14427 ( .A(n11820), .ZN(n15931) );
  INV_X1 U14428 ( .A(n11815), .ZN(n11816) );
  NAND2_X1 U14429 ( .A1(n11819), .A2(n11816), .ZN(n11950) );
  NAND2_X1 U14430 ( .A1(n11950), .A2(n13562), .ZN(n11824) );
  AOI21_X1 U14431 ( .B1(n11819), .B2(n11818), .A(n11817), .ZN(n11823) );
  NAND2_X1 U14432 ( .A1(n11820), .A2(n13413), .ZN(n11822) );
  INV_X1 U14433 ( .A(n12180), .ZN(n13148) );
  AOI22_X1 U14434 ( .A1(n13148), .A2(n13567), .B1(n13566), .B2(n13147), .ZN(
        n11821) );
  OAI211_X1 U14435 ( .C1(n11824), .C2(n11823), .A(n11822), .B(n11821), .ZN(
        n15932) );
  MUX2_X1 U14436 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15932), .S(n13585), .Z(
        n11825) );
  INV_X1 U14437 ( .A(n11825), .ZN(n11827) );
  AOI22_X1 U14438 ( .A1(n13557), .A2(n13109), .B1(n13579), .B2(n13112), .ZN(
        n11826) );
  OAI211_X1 U14439 ( .C1(n15931), .C2(n13436), .A(n11827), .B(n11826), .ZN(
        P3_U3227) );
  XNOR2_X1 U14440 ( .A(n11828), .B(n12815), .ZN(n11832) );
  INV_X1 U14441 ( .A(n11832), .ZN(n15919) );
  NAND2_X1 U14442 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  XNOR2_X1 U14443 ( .A(n11831), .B(n12762), .ZN(n11835) );
  NAND2_X1 U14444 ( .A1(n11832), .A2(n13413), .ZN(n11834) );
  AOI22_X1 U14445 ( .A1(n13148), .A2(n13566), .B1(n13567), .B2(n13150), .ZN(
        n11833) );
  OAI211_X1 U14446 ( .C1(n11835), .C2(n13507), .A(n11834), .B(n11833), .ZN(
        n15920) );
  MUX2_X1 U14447 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15920), .S(n13585), .Z(
        n11836) );
  INV_X1 U14448 ( .A(n11836), .ZN(n11838) );
  AOI22_X1 U14449 ( .A1(n13557), .A2(n13062), .B1(n13579), .B2(n13063), .ZN(
        n11837) );
  OAI211_X1 U14450 ( .C1(n15919), .C2(n13436), .A(n11838), .B(n11837), .ZN(
        P3_U3229) );
  AOI22_X1 U14451 ( .A1(n11841), .A2(n11840), .B1(n11644), .B2(n11839), .ZN(
        n11845) );
  XNOR2_X1 U14452 ( .A(n11843), .B(n11842), .ZN(n11844) );
  XNOR2_X1 U14453 ( .A(n11845), .B(n11844), .ZN(n11850) );
  NOR2_X1 U14454 ( .A1(n14809), .A2(n15683), .ZN(n11848) );
  NAND2_X1 U14455 ( .A1(n14806), .A2(n15531), .ZN(n11846) );
  NAND2_X1 U14456 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14899) );
  OAI211_X1 U14457 ( .C1(n14808), .C2(n15385), .A(n11846), .B(n14899), .ZN(
        n11847) );
  AOI211_X1 U14458 ( .C1(n14813), .C2(n15518), .A(n11848), .B(n11847), .ZN(
        n11849) );
  OAI21_X1 U14459 ( .B1(n11850), .B2(n14815), .A(n11849), .ZN(P1_U3213) );
  INV_X1 U14460 ( .A(SI_23_), .ZN(n11855) );
  NAND2_X1 U14461 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  OAI211_X1 U14462 ( .C1(n11855), .C2(n11854), .A(n11853), .B(n12945), .ZN(
        P3_U3272) );
  INV_X1 U14463 ( .A(n11858), .ZN(n11860) );
  NAND2_X1 U14464 ( .A1(n11860), .A2(n11859), .ZN(n11861) );
  XNOR2_X1 U14465 ( .A(n6607), .B(n13799), .ZN(n11863) );
  NAND2_X1 U14466 ( .A1(n13862), .A2(n14035), .ZN(n11864) );
  NAND2_X1 U14467 ( .A1(n11863), .A2(n11864), .ZN(n13732) );
  INV_X1 U14468 ( .A(n11863), .ZN(n11866) );
  INV_X1 U14469 ( .A(n11864), .ZN(n11865) );
  NAND2_X1 U14470 ( .A1(n11866), .A2(n11865), .ZN(n11867) );
  NAND2_X1 U14471 ( .A1(n13732), .A2(n11867), .ZN(n11870) );
  INV_X1 U14472 ( .A(n11870), .ZN(n11868) );
  INV_X1 U14473 ( .A(n13733), .ZN(n11869) );
  AOI21_X1 U14474 ( .B1(n11871), .B2(n11870), .A(n11869), .ZN(n11878) );
  NAND2_X1 U14475 ( .A1(n6531), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n14125) );
  OAI21_X1 U14476 ( .B1(n13950), .B2(n13839), .A(n14125), .ZN(n11875) );
  OAI22_X1 U14477 ( .A1(n13978), .A2(n11873), .B1(n13990), .B2(n11872), .ZN(
        n11874) );
  AOI211_X1 U14478 ( .C1(n6607), .C2(n14000), .A(n11875), .B(n11874), .ZN(
        n11877) );
  OAI21_X1 U14479 ( .B1(n11878), .B2(n14002), .A(n11877), .ZN(P2_U3193) );
  INV_X1 U14480 ( .A(n11879), .ZN(n11882) );
  OAI222_X1 U14481 ( .A1(n12702), .A2(n11881), .B1(n11978), .B2(n11882), .C1(
        n11880), .C2(n6531), .ZN(P2_U3306) );
  OAI222_X1 U14482 ( .A1(n15433), .A2(n11883), .B1(n6554), .B2(n11882), .C1(
        P1_U3086), .C2(n12646), .ZN(P1_U3334) );
  XNOR2_X1 U14483 ( .A(n11884), .B(n11885), .ZN(n15652) );
  XNOR2_X1 U14484 ( .A(n11886), .B(n11885), .ZN(n15656) );
  AOI21_X1 U14485 ( .B1(n15555), .B2(n12520), .A(n15574), .ZN(n11887) );
  NAND2_X1 U14486 ( .A1(n11887), .A2(n6850), .ZN(n15650) );
  NOR2_X1 U14487 ( .A1(n15185), .A2(n15650), .ZN(n11892) );
  INV_X1 U14488 ( .A(n15196), .ZN(n15158) );
  AOI22_X1 U14489 ( .A1(n15192), .A2(n15647), .B1(n15158), .B2(n15666), .ZN(
        n11890) );
  AOI22_X1 U14490 ( .A1(n15584), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n11888), 
        .B2(n15573), .ZN(n11889) );
  OAI211_X1 U14491 ( .C1(n12519), .C2(n15552), .A(n11890), .B(n11889), .ZN(
        n11891) );
  AOI211_X1 U14492 ( .C1(n15656), .C2(n15581), .A(n11892), .B(n11891), .ZN(
        n11893) );
  OAI21_X1 U14493 ( .B1(n15652), .B2(n15095), .A(n11893), .ZN(P1_U3289) );
  INV_X1 U14494 ( .A(n15930), .ZN(n15937) );
  XNOR2_X1 U14495 ( .A(n11894), .B(n12769), .ZN(n11947) );
  INV_X1 U14496 ( .A(n11947), .ZN(n11901) );
  INV_X1 U14497 ( .A(n11895), .ZN(n11896) );
  OR2_X1 U14498 ( .A1(n11895), .A2(n12835), .ZN(n11997) );
  OAI21_X1 U14499 ( .B1(n11896), .B2(n12769), .A(n11997), .ZN(n11899) );
  OAI22_X1 U14500 ( .A1(n11897), .A2(n13509), .B1(n12251), .B2(n13511), .ZN(
        n11898) );
  AOI21_X1 U14501 ( .B1(n11899), .B2(n13562), .A(n11898), .ZN(n11900) );
  OAI21_X1 U14502 ( .B1(n11947), .B2(n13433), .A(n11900), .ZN(n11942) );
  AOI21_X1 U14503 ( .B1(n15937), .B2(n11901), .A(n11942), .ZN(n12035) );
  AOI22_X1 U14504 ( .A1(n13675), .A2(n13003), .B1(P3_REG0_REG_8__SCAN_IN), 
        .B2(n15941), .ZN(n11902) );
  OAI21_X1 U14505 ( .B1(n12035), .B2(n15941), .A(n11902), .ZN(P3_U3414) );
  INV_X1 U14506 ( .A(n11903), .ZN(n11977) );
  AOI22_X1 U14507 ( .A1(n11904), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n15422), .ZN(n11905) );
  OAI21_X1 U14508 ( .B1(n11977), .B2(n6554), .A(n11905), .ZN(P1_U3331) );
  INV_X1 U14509 ( .A(n11906), .ZN(n11907) );
  AOI21_X1 U14510 ( .B1(n12657), .B2(n11908), .A(n11907), .ZN(n15393) );
  OR2_X1 U14511 ( .A1(n11909), .A2(n10164), .ZN(n12051) );
  NAND2_X1 U14512 ( .A1(n11909), .A2(n10164), .ZN(n11910) );
  AOI21_X1 U14513 ( .B1(n12051), .B2(n11910), .A(n15651), .ZN(n15390) );
  MUX2_X1 U14514 ( .A(n15390), .B(P1_REG2_REG_9__SCAN_IN), .S(n15584), .Z(
        n11911) );
  INV_X1 U14515 ( .A(n11911), .ZN(n11917) );
  AOI211_X1 U14516 ( .C1(n15389), .C2(n11912), .A(n15574), .B(n12144), .ZN(
        n15386) );
  AOI22_X1 U14517 ( .A1(n15192), .A2(n15514), .B1(n15573), .B2(n12133), .ZN(
        n11914) );
  NAND2_X1 U14518 ( .A1(n15212), .A2(n15389), .ZN(n11913) );
  OAI211_X1 U14519 ( .C1(n15384), .C2(n15196), .A(n11914), .B(n11913), .ZN(
        n11915) );
  AOI21_X1 U14520 ( .B1(n15386), .B2(n15582), .A(n11915), .ZN(n11916) );
  OAI211_X1 U14521 ( .C1(n15214), .C2(n15393), .A(n11917), .B(n11916), .ZN(
        P1_U3284) );
  XNOR2_X1 U14522 ( .A(n11938), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n13162) );
  INV_X1 U14523 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11919) );
  XOR2_X1 U14524 ( .A(n13162), .B(n13163), .Z(n11941) );
  INV_X1 U14525 ( .A(n11920), .ZN(n11922) );
  INV_X1 U14526 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11921) );
  XNOR2_X1 U14527 ( .A(n11938), .B(n11921), .ZN(n11923) );
  AOI21_X2 U14528 ( .B1(n11924), .B2(n11922), .A(n11923), .ZN(n13165) );
  AND3_X1 U14529 ( .A1(n11924), .A2(n11923), .A3(n11922), .ZN(n11925) );
  OAI21_X1 U14530 ( .B1(n13165), .B2(n11925), .A(n15888), .ZN(n11940) );
  INV_X1 U14531 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14532 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13025)
         );
  OAI21_X1 U14533 ( .B1(n15898), .B2(n11926), .A(n13025), .ZN(n11937) );
  MUX2_X1 U14534 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13285), .Z(n13168) );
  XNOR2_X1 U14535 ( .A(n13168), .B(n11938), .ZN(n11931) );
  INV_X1 U14536 ( .A(n11927), .ZN(n11929) );
  NAND2_X1 U14537 ( .A1(n11929), .A2(n11928), .ZN(n11932) );
  AND2_X1 U14538 ( .A1(n11931), .A2(n11932), .ZN(n11930) );
  INV_X1 U14539 ( .A(n13173), .ZN(n11935) );
  AOI21_X1 U14540 ( .B1(n11933), .B2(n11932), .A(n11931), .ZN(n11934) );
  NOR3_X1 U14541 ( .A1(n11935), .A2(n11934), .A3(n15892), .ZN(n11936) );
  AOI211_X1 U14542 ( .C1(n15886), .C2(n11938), .A(n11937), .B(n11936), .ZN(
        n11939) );
  OAI211_X1 U14543 ( .C1(n11941), .C2(n13237), .A(n11940), .B(n11939), .ZN(
        P3_U3194) );
  INV_X1 U14544 ( .A(n11942), .ZN(n11943) );
  MUX2_X1 U14545 ( .A(n11944), .B(n11943), .S(n13585), .Z(n11946) );
  AOI22_X1 U14546 ( .A1(n13557), .A2(n13003), .B1(n13579), .B2(n13004), .ZN(
        n11945) );
  OAI211_X1 U14547 ( .C1(n11947), .C2(n13436), .A(n11946), .B(n11945), .ZN(
        P3_U3225) );
  XNOR2_X1 U14548 ( .A(n11948), .B(n12829), .ZN(n15938) );
  INV_X1 U14549 ( .A(n15938), .ZN(n11957) );
  NAND2_X1 U14550 ( .A1(n11950), .A2(n11949), .ZN(n11951) );
  XNOR2_X1 U14551 ( .A(n11951), .B(n7235), .ZN(n11953) );
  INV_X1 U14552 ( .A(n12193), .ZN(n13146) );
  AOI22_X1 U14553 ( .A1(n13566), .A2(n13146), .B1(n12952), .B2(n13567), .ZN(
        n11952) );
  OAI21_X1 U14554 ( .B1(n11953), .B2(n13507), .A(n11952), .ZN(n11954) );
  AOI21_X1 U14555 ( .B1(n15938), .B2(n13413), .A(n11954), .ZN(n15940) );
  MUX2_X1 U14556 ( .A(n7313), .B(n15940), .S(n13585), .Z(n11956) );
  AOI22_X1 U14557 ( .A1(n13557), .A2(n15935), .B1(n13579), .B2(n12953), .ZN(
        n11955) );
  OAI211_X1 U14558 ( .C1(n11957), .C2(n13436), .A(n11956), .B(n11955), .ZN(
        P3_U3226) );
  INV_X1 U14559 ( .A(n11958), .ZN(n11959) );
  AOI22_X1 U14560 ( .A1(n11960), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11964), 
        .B2(n11959), .ZN(n11963) );
  INV_X1 U14561 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11961) );
  MUX2_X1 U14562 ( .A(n11961), .B(P2_REG2_REG_16__SCAN_IN), .S(n14173), .Z(
        n11962) );
  AOI211_X1 U14563 ( .C1(n11963), .C2(n11962), .A(n14197), .B(n14169), .ZN(
        n11975) );
  NAND2_X1 U14564 ( .A1(n11965), .A2(n11964), .ZN(n11966) );
  NAND2_X1 U14565 ( .A1(n11967), .A2(n11966), .ZN(n11970) );
  XNOR2_X1 U14566 ( .A(n14173), .B(n11968), .ZN(n11969) );
  NAND2_X1 U14567 ( .A1(n11970), .A2(n11969), .ZN(n14175) );
  OAI211_X1 U14568 ( .C1(n11970), .C2(n11969), .A(n14175), .B(n15744), .ZN(
        n11973) );
  NOR2_X1 U14569 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13909), .ZN(n11971) );
  AOI21_X1 U14570 ( .B1(n15747), .B2(n14173), .A(n11971), .ZN(n11972) );
  OAI211_X1 U14571 ( .C1(n15753), .C2(n7505), .A(n11973), .B(n11972), .ZN(
        n11974) );
  OR2_X1 U14572 ( .A1(n11975), .A2(n11974), .ZN(P2_U3230) );
  OAI222_X1 U14573 ( .A1(n12702), .A2(n11979), .B1(n11978), .B2(n11977), .C1(
        P2_U3088), .C2(n11976), .ZN(P2_U3303) );
  OR2_X1 U14574 ( .A1(n11980), .A2(n11984), .ZN(n11981) );
  AND2_X1 U14575 ( .A1(n11982), .A2(n11981), .ZN(n11991) );
  OAI22_X1 U14576 ( .A1(n13939), .A2(n14471), .B1(n13977), .B2(n14473), .ZN(
        n11987) );
  OR2_X1 U14577 ( .A1(n11983), .A2(n11984), .ZN(n12016) );
  NAND2_X1 U14578 ( .A1(n11983), .A2(n11984), .ZN(n11985) );
  AOI21_X1 U14579 ( .B1(n12016), .B2(n11985), .A(n14461), .ZN(n11986) );
  AOI211_X1 U14580 ( .C1(n11991), .C2(n15818), .A(n11987), .B(n11986), .ZN(
        n14606) );
  AOI211_X1 U14581 ( .C1(n14604), .C2(n11989), .A(n14482), .B(n11988), .ZN(
        n14603) );
  INV_X1 U14582 ( .A(n14604), .ZN(n13944) );
  AOI22_X1 U14583 ( .A1(n14484), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n13937), 
        .B2(n15760), .ZN(n11990) );
  OAI21_X1 U14584 ( .B1(n14486), .B2(n13944), .A(n11990), .ZN(n11993) );
  INV_X1 U14585 ( .A(n11991), .ZN(n14607) );
  NOR2_X1 U14586 ( .A1(n14607), .A2(n14488), .ZN(n11992) );
  AOI211_X1 U14587 ( .C1(n14603), .C2(n15767), .A(n11993), .B(n11992), .ZN(
        n11994) );
  OAI21_X1 U14588 ( .B1(n14484), .B2(n14606), .A(n11994), .ZN(P2_U3256) );
  XNOR2_X1 U14589 ( .A(n11995), .B(n12850), .ZN(n12269) );
  NAND2_X1 U14590 ( .A1(n11997), .A2(n11996), .ZN(n12040) );
  INV_X1 U14591 ( .A(n12042), .ZN(n12839) );
  OR2_X1 U14592 ( .A1(n12040), .A2(n12839), .ZN(n12041) );
  NAND2_X1 U14593 ( .A1(n12041), .A2(n11998), .ZN(n11999) );
  XNOR2_X1 U14594 ( .A(n11999), .B(n12838), .ZN(n12000) );
  NAND2_X1 U14595 ( .A1(n12000), .A2(n13562), .ZN(n12002) );
  AOI22_X1 U14596 ( .A1(n13144), .A2(n13566), .B1(n13567), .B2(n13145), .ZN(
        n12001) );
  NAND2_X1 U14597 ( .A1(n12002), .A2(n12001), .ZN(n12266) );
  AOI21_X1 U14598 ( .B1(n12269), .B2(n15905), .A(n12266), .ZN(n12174) );
  INV_X1 U14599 ( .A(n12847), .ZN(n12003) );
  AOI22_X1 U14600 ( .A1(n13675), .A2(n12003), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15941), .ZN(n12004) );
  OAI21_X1 U14601 ( .B1(n12174), .B2(n15941), .A(n12004), .ZN(P3_U3420) );
  INV_X1 U14602 ( .A(n12005), .ZN(n12006) );
  AOI21_X1 U14603 ( .B1(n12014), .B2(n12007), .A(n12006), .ZN(n12170) );
  AOI211_X1 U14604 ( .C1(n13842), .C2(n7513), .A(n14482), .B(n14506), .ZN(
        n12164) );
  INV_X1 U14605 ( .A(n12008), .ZN(n13838) );
  OAI22_X1 U14606 ( .A1(n14486), .A2(n12009), .B1(n14406), .B2(n13838), .ZN(
        n12010) );
  AOI21_X1 U14607 ( .B1(n12164), .B2(n14457), .A(n12010), .ZN(n12024) );
  NAND2_X1 U14608 ( .A1(n12016), .A2(n12012), .ZN(n12011) );
  NAND2_X1 U14609 ( .A1(n12011), .A2(n12014), .ZN(n14468) );
  INV_X1 U14610 ( .A(n12012), .ZN(n12013) );
  NOR2_X1 U14611 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  NAND2_X1 U14612 ( .A1(n12016), .A2(n12015), .ZN(n12017) );
  NAND2_X1 U14613 ( .A1(n14468), .A2(n12017), .ZN(n12018) );
  NAND2_X1 U14614 ( .A1(n12018), .A2(n15757), .ZN(n12020) );
  AOI22_X1 U14615 ( .A1(n14034), .A2(n14496), .B1(n14494), .B2(n14033), .ZN(
        n12019) );
  NAND2_X1 U14616 ( .A1(n12020), .A2(n12019), .ZN(n12163) );
  INV_X1 U14617 ( .A(n12163), .ZN(n12022) );
  MUX2_X1 U14618 ( .A(n12022), .B(n12021), .S(n14484), .Z(n12023) );
  OAI211_X1 U14619 ( .C1(n12170), .C2(n14465), .A(n12024), .B(n12023), .ZN(
        P2_U3255) );
  INV_X1 U14620 ( .A(n12025), .ZN(n12122) );
  AOI22_X1 U14621 ( .A1(n12026), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n15422), .ZN(n12027) );
  OAI21_X1 U14622 ( .B1(n12122), .B2(n6554), .A(n12027), .ZN(P1_U3330) );
  NAND2_X1 U14623 ( .A1(n6542), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12031) );
  NAND2_X1 U14624 ( .A1(n9066), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U14625 ( .A1(n12028), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12029) );
  AND3_X1 U14626 ( .A1(n12031), .A2(n12030), .A3(n12029), .ZN(n12032) );
  NAND2_X1 U14627 ( .A1(n13142), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n12034) );
  OAI21_X1 U14628 ( .B1(n13333), .B2(n13142), .A(n12034), .ZN(P3_U3522) );
  MUX2_X1 U14629 ( .A(n12036), .B(n12035), .S(n15954), .Z(n12037) );
  OAI21_X1 U14630 ( .B1(n12038), .B2(n13660), .A(n12037), .ZN(P3_U3467) );
  XNOR2_X1 U14631 ( .A(n12039), .B(n12042), .ZN(n12079) );
  INV_X1 U14632 ( .A(n12079), .ZN(n12046) );
  AOI22_X1 U14633 ( .A1(n13146), .A2(n13567), .B1(n13566), .B2(n13087), .ZN(
        n12045) );
  INV_X1 U14634 ( .A(n12040), .ZN(n12043) );
  OAI211_X1 U14635 ( .C1(n12043), .C2(n12042), .A(n13562), .B(n12041), .ZN(
        n12044) );
  OAI211_X1 U14636 ( .C1(n12079), .C2(n13433), .A(n12045), .B(n12044), .ZN(
        n12074) );
  AOI21_X1 U14637 ( .B1(n15937), .B2(n12046), .A(n12074), .ZN(n12171) );
  AOI22_X1 U14638 ( .A1(n13675), .A2(n12192), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15941), .ZN(n12047) );
  OAI21_X1 U14639 ( .B1(n12171), .B2(n15941), .A(n12047), .ZN(P3_U3417) );
  XNOR2_X1 U14640 ( .A(n12049), .B(n12052), .ZN(n15374) );
  NAND2_X1 U14641 ( .A1(n12051), .A2(n12050), .ZN(n12150) );
  INV_X1 U14642 ( .A(n15378), .ZN(n12562) );
  INV_X1 U14643 ( .A(n12660), .ZN(n12149) );
  NOR2_X1 U14644 ( .A1(n12150), .A2(n12149), .ZN(n15376) );
  OAI21_X1 U14645 ( .B1(n15384), .B2(n12562), .A(n12662), .ZN(n12054) );
  NAND2_X1 U14646 ( .A1(n12053), .A2(n12052), .ZN(n12089) );
  OAI211_X1 U14647 ( .C1(n15376), .C2(n12054), .A(n15568), .B(n12089), .ZN(
        n12056) );
  AOI22_X1 U14648 ( .A1(n14820), .A2(n15665), .B1(n15668), .B2(n15353), .ZN(
        n12055) );
  NAND2_X1 U14649 ( .A1(n12056), .A2(n12055), .ZN(n15370) );
  OR2_X1 U14650 ( .A1(n12058), .A2(n12062), .ZN(n12059) );
  AND3_X1 U14651 ( .A1(n12057), .A2(n12059), .A3(n15540), .ZN(n15371) );
  NAND2_X1 U14652 ( .A1(n15371), .A2(n15582), .ZN(n12061) );
  AOI22_X1 U14653 ( .A1(n15584), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12232), 
        .B2(n15573), .ZN(n12060) );
  OAI211_X1 U14654 ( .C1(n12062), .C2(n15552), .A(n12061), .B(n12060), .ZN(
        n12063) );
  AOI21_X1 U14655 ( .B1(n15370), .B2(n15178), .A(n12063), .ZN(n12064) );
  OAI21_X1 U14656 ( .B1(n15214), .B2(n15374), .A(n12064), .ZN(P1_U3282) );
  NOR2_X1 U14657 ( .A1(n6757), .A2(n12065), .ZN(n12066) );
  XNOR2_X1 U14658 ( .A(n12067), .B(n12066), .ZN(n12073) );
  NAND2_X1 U14659 ( .A1(n14806), .A2(n14821), .ZN(n12069) );
  OAI211_X1 U14660 ( .C1(n14808), .C2(n12565), .A(n12069), .B(n12068), .ZN(
        n12071) );
  NOR2_X1 U14661 ( .A1(n15378), .A2(n14809), .ZN(n12070) );
  AOI211_X1 U14662 ( .C1(n14813), .C2(n12146), .A(n12071), .B(n12070), .ZN(
        n12072) );
  OAI21_X1 U14663 ( .B1(n12073), .B2(n14815), .A(n12072), .ZN(P1_U3217) );
  INV_X1 U14664 ( .A(n12074), .ZN(n12075) );
  MUX2_X1 U14665 ( .A(n12076), .B(n12075), .S(n13585), .Z(n12078) );
  AOI22_X1 U14666 ( .A1(n13557), .A2(n12192), .B1(n13579), .B2(n12209), .ZN(
        n12077) );
  OAI211_X1 U14667 ( .C1(n12079), .C2(n13436), .A(n12078), .B(n12077), .ZN(
        P3_U3224) );
  XNOR2_X1 U14668 ( .A(n12080), .B(n12854), .ZN(n12138) );
  INV_X1 U14669 ( .A(n12138), .ZN(n12087) );
  NAND2_X1 U14670 ( .A1(n13433), .A2(n12081), .ZN(n12082) );
  XNOR2_X1 U14671 ( .A(n12241), .B(n12854), .ZN(n12083) );
  OAI222_X1 U14672 ( .A1(n13509), .A2(n12207), .B1(n13511), .B2(n13090), .C1(
        n12083), .C2(n13507), .ZN(n12137) );
  AOI22_X1 U14673 ( .A1(n13580), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n13579), 
        .B2(n13092), .ZN(n12084) );
  OAI21_X1 U14674 ( .B1(n13095), .B2(n13582), .A(n12084), .ZN(n12085) );
  AOI21_X1 U14675 ( .B1(n12137), .B2(n13574), .A(n12085), .ZN(n12086) );
  OAI21_X1 U14676 ( .B1(n12087), .B2(n13588), .A(n12086), .ZN(P3_U3222) );
  AND2_X1 U14677 ( .A1(n12089), .A2(n12088), .ZN(n12092) );
  NAND2_X1 U14678 ( .A1(n12091), .A2(n12090), .ZN(n12224) );
  AOI211_X1 U14679 ( .C1(n10124), .C2(n12092), .A(n15651), .B(n12224), .ZN(
        n15366) );
  INV_X1 U14680 ( .A(n15366), .ZN(n12103) );
  NAND2_X1 U14681 ( .A1(n15158), .A2(n15363), .ZN(n12094) );
  AOI22_X1 U14682 ( .A1(n15584), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12294), 
        .B2(n15573), .ZN(n12093) );
  OAI211_X1 U14683 ( .C1(n12565), .C2(n15162), .A(n12094), .B(n12093), .ZN(
        n12097) );
  AOI21_X1 U14684 ( .B1(n12057), .B2(n12098), .A(n6601), .ZN(n12095) );
  NAND2_X1 U14685 ( .A1(n12095), .A2(n12218), .ZN(n15365) );
  NOR2_X1 U14686 ( .A1(n15365), .A2(n15185), .ZN(n12096) );
  AOI211_X1 U14687 ( .C1(n15212), .C2(n12098), .A(n12097), .B(n12096), .ZN(
        n12102) );
  OAI21_X1 U14688 ( .B1(n12100), .B2(n10124), .A(n12099), .ZN(n15368) );
  NAND2_X1 U14689 ( .A1(n15368), .A2(n15581), .ZN(n12101) );
  OAI211_X1 U14690 ( .C1(n12103), .C2(n15584), .A(n12102), .B(n12101), .ZN(
        P1_U3281) );
  NAND2_X1 U14691 ( .A1(n12108), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14941) );
  NAND2_X1 U14692 ( .A1(n14942), .A2(n14941), .ZN(n12106) );
  MUX2_X1 U14693 ( .A(n12104), .B(P1_REG2_REG_17__SCAN_IN), .S(n14939), .Z(
        n12105) );
  NAND2_X1 U14694 ( .A1(n12106), .A2(n12105), .ZN(n14944) );
  OR2_X1 U14695 ( .A1(n14939), .A2(n12104), .ZN(n12107) );
  NAND2_X1 U14696 ( .A1(n14944), .A2(n12107), .ZN(n14953) );
  XNOR2_X1 U14697 ( .A(n14953), .B(n12113), .ZN(n14951) );
  XNOR2_X1 U14698 ( .A(n14951), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n12120) );
  NAND2_X1 U14699 ( .A1(n12108), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U14700 ( .A1(n12110), .A2(n12109), .ZN(n14935) );
  XNOR2_X1 U14701 ( .A(n14939), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14934) );
  NAND2_X1 U14702 ( .A1(n14935), .A2(n14934), .ZN(n14933) );
  INV_X1 U14703 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12111) );
  OR2_X1 U14704 ( .A1(n14939), .A2(n12111), .ZN(n12112) );
  NAND2_X1 U14705 ( .A1(n14933), .A2(n12112), .ZN(n12114) );
  INV_X1 U14706 ( .A(n12113), .ZN(n14952) );
  NAND2_X1 U14707 ( .A1(n12114), .A2(n14952), .ZN(n14948) );
  OR2_X1 U14708 ( .A1(n12114), .A2(n14952), .ZN(n12115) );
  AND2_X1 U14709 ( .A1(n14948), .A2(n12115), .ZN(n12116) );
  NAND2_X1 U14710 ( .A1(n12116), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14949) );
  OAI211_X1 U14711 ( .C1(n12116), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14949), 
        .B(n15504), .ZN(n12119) );
  NAND2_X1 U14712 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14788)
         );
  OAI21_X1 U14713 ( .B1(n15509), .B2(n10360), .A(n14788), .ZN(n12117) );
  AOI21_X1 U14714 ( .B1(n14952), .B2(n15501), .A(n12117), .ZN(n12118) );
  OAI211_X1 U14715 ( .C1(n12120), .C2(n14960), .A(n12119), .B(n12118), .ZN(
        P1_U3261) );
  OAI222_X1 U14716 ( .A1(P2_U3088), .A2(n12123), .B1(n11978), .B2(n12122), 
        .C1(n12121), .C2(n14659), .ZN(P2_U3302) );
  INV_X1 U14717 ( .A(n15389), .ZN(n12136) );
  INV_X1 U14718 ( .A(n12126), .ZN(n12130) );
  AOI21_X1 U14719 ( .B1(n12126), .B2(n12125), .A(n12124), .ZN(n12127) );
  NOR2_X1 U14720 ( .A1(n12127), .A2(n14815), .ZN(n12128) );
  OAI21_X1 U14721 ( .B1(n12130), .B2(n12129), .A(n12128), .ZN(n12135) );
  NAND2_X1 U14722 ( .A1(n14806), .A2(n15514), .ZN(n12131) );
  NAND2_X1 U14723 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14917) );
  OAI211_X1 U14724 ( .C1(n14808), .C2(n15384), .A(n12131), .B(n14917), .ZN(
        n12132) );
  AOI21_X1 U14725 ( .B1(n12133), .B2(n14813), .A(n12132), .ZN(n12134) );
  OAI211_X1 U14726 ( .C1(n12136), .C2(n14809), .A(n12135), .B(n12134), .ZN(
        P1_U3231) );
  AOI21_X1 U14727 ( .B1(n12138), .B2(n15905), .A(n12137), .ZN(n12142) );
  INV_X1 U14728 ( .A(n13095), .ZN(n12140) );
  AOI22_X1 U14729 ( .A1(n12140), .A2(n13675), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n15941), .ZN(n12139) );
  OAI21_X1 U14730 ( .B1(n12142), .B2(n15941), .A(n12139), .ZN(P3_U3423) );
  AOI22_X1 U14731 ( .A1(n12140), .A2(n13601), .B1(P3_REG1_REG_11__SCAN_IN), 
        .B2(n15951), .ZN(n12141) );
  OAI21_X1 U14732 ( .B1(n12142), .B2(n15951), .A(n12141), .ZN(P3_U3470) );
  XNOR2_X1 U14733 ( .A(n12143), .B(n12660), .ZN(n15383) );
  XNOR2_X1 U14734 ( .A(n12144), .B(n15378), .ZN(n12145) );
  OAI22_X1 U14735 ( .A1(n12145), .A2(n6601), .B1(n12565), .B2(n15628), .ZN(
        n15380) );
  NAND2_X1 U14736 ( .A1(n15192), .A2(n14821), .ZN(n12148) );
  AOI22_X1 U14737 ( .A1(n15584), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n12146), 
        .B2(n15573), .ZN(n12147) );
  OAI211_X1 U14738 ( .C1(n15378), .C2(n15552), .A(n12148), .B(n12147), .ZN(
        n12152) );
  AND2_X1 U14739 ( .A1(n12150), .A2(n12149), .ZN(n15375) );
  NOR3_X1 U14740 ( .A1(n15376), .A2(n15375), .A3(n15095), .ZN(n12151) );
  AOI211_X1 U14741 ( .C1(n15582), .C2(n15380), .A(n12152), .B(n12151), .ZN(
        n12153) );
  OAI21_X1 U14742 ( .B1(n15214), .B2(n15383), .A(n12153), .ZN(P1_U3283) );
  INV_X1 U14743 ( .A(n13345), .ZN(n12154) );
  NAND2_X1 U14744 ( .A1(n12154), .A2(P3_U3897), .ZN(n12155) );
  OAI21_X1 U14745 ( .B1(P3_U3897), .B2(n12156), .A(n12155), .ZN(P3_U3520) );
  INV_X1 U14746 ( .A(n12157), .ZN(n12161) );
  OAI222_X1 U14747 ( .A1(P2_U3088), .A2(n12159), .B1(n11978), .B2(n12161), 
        .C1(n12158), .C2(n12702), .ZN(P2_U3301) );
  OAI222_X1 U14748 ( .A1(P1_U3086), .A2(n12162), .B1(n6554), .B2(n12161), .C1(
        n12160), .C2(n15433), .ZN(P1_U3329) );
  INV_X1 U14749 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n12165) );
  AOI211_X1 U14750 ( .C1(n15835), .C2(n13842), .A(n12164), .B(n12163), .ZN(
        n12167) );
  MUX2_X1 U14751 ( .A(n12165), .B(n12167), .S(n15864), .Z(n12166) );
  OAI21_X1 U14752 ( .B1(n12170), .B2(n14586), .A(n12166), .ZN(P2_U3509) );
  INV_X1 U14753 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12168) );
  MUX2_X1 U14754 ( .A(n12168), .B(n12167), .S(n15850), .Z(n12169) );
  OAI21_X1 U14755 ( .B1(n12170), .B2(n14649), .A(n12169), .ZN(P2_U3460) );
  INV_X1 U14756 ( .A(n12192), .ZN(n12212) );
  MUX2_X1 U14757 ( .A(n12172), .B(n12171), .S(n15954), .Z(n12173) );
  OAI21_X1 U14758 ( .B1(n13660), .B2(n12212), .A(n12173), .ZN(P3_U3468) );
  MUX2_X1 U14759 ( .A(n12175), .B(n12174), .S(n15954), .Z(n12176) );
  OAI21_X1 U14760 ( .B1(n13660), .B2(n12847), .A(n12176), .ZN(P3_U3469) );
  INV_X1 U14761 ( .A(n15870), .ZN(n13136) );
  INV_X1 U14762 ( .A(n12179), .ZN(n12181) );
  NAND2_X1 U14763 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  INV_X1 U14764 ( .A(n13104), .ZN(n12185) );
  XNOR2_X1 U14765 ( .A(n12385), .B(n13109), .ZN(n12186) );
  XNOR2_X1 U14766 ( .A(n12186), .B(n12183), .ZN(n13105) );
  INV_X1 U14767 ( .A(n13105), .ZN(n12184) );
  INV_X1 U14768 ( .A(n12186), .ZN(n12187) );
  NAND2_X1 U14769 ( .A1(n12187), .A2(n12952), .ZN(n12188) );
  NAND2_X1 U14770 ( .A1(n13106), .A2(n12188), .ZN(n12196) );
  NAND2_X1 U14771 ( .A1(n12196), .A2(n12949), .ZN(n12948) );
  INV_X1 U14772 ( .A(n12949), .ZN(n12189) );
  AND2_X1 U14773 ( .A1(n12189), .A2(n13147), .ZN(n12198) );
  INV_X1 U14774 ( .A(n12198), .ZN(n12190) );
  NAND2_X1 U14775 ( .A1(n12948), .A2(n12190), .ZN(n13000) );
  XNOR2_X1 U14776 ( .A(n12385), .B(n13003), .ZN(n12194) );
  XNOR2_X1 U14777 ( .A(n12194), .B(n13146), .ZN(n12999) );
  NAND2_X1 U14778 ( .A1(n13000), .A2(n12999), .ZN(n12998) );
  INV_X1 U14779 ( .A(n12194), .ZN(n12191) );
  NAND2_X1 U14780 ( .A1(n12191), .A2(n13146), .ZN(n12199) );
  XNOR2_X1 U14781 ( .A(n12385), .B(n12192), .ZN(n12252) );
  XNOR2_X1 U14782 ( .A(n12252), .B(n13145), .ZN(n12201) );
  AOI21_X1 U14783 ( .B1(n12998), .B2(n12199), .A(n12201), .ZN(n12205) );
  NAND2_X1 U14784 ( .A1(n12194), .A2(n12193), .ZN(n12197) );
  AND2_X1 U14785 ( .A1(n12949), .A2(n12197), .ZN(n12195) );
  NAND2_X1 U14786 ( .A1(n12196), .A2(n12195), .ZN(n12203) );
  NAND2_X1 U14787 ( .A1(n12198), .A2(n12197), .ZN(n12200) );
  AND3_X1 U14788 ( .A1(n12201), .A2(n12200), .A3(n12199), .ZN(n12202) );
  INV_X1 U14789 ( .A(n12254), .ZN(n12204) );
  OAI21_X1 U14790 ( .B1(n12205), .B2(n12204), .A(n13128), .ZN(n12211) );
  NAND2_X1 U14791 ( .A1(n13130), .A2(n13146), .ZN(n12206) );
  NAND2_X1 U14792 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15896) );
  OAI211_X1 U14793 ( .C1(n15874), .C2(n12207), .A(n12206), .B(n15896), .ZN(
        n12208) );
  AOI21_X1 U14794 ( .B1(n12209), .B2(n13133), .A(n12208), .ZN(n12210) );
  OAI211_X1 U14795 ( .C1(n13136), .C2(n12212), .A(n12211), .B(n12210), .ZN(
        P3_U3171) );
  INV_X1 U14796 ( .A(n12663), .ZN(n12225) );
  INV_X1 U14797 ( .A(n12213), .ZN(n12278) );
  NAND2_X1 U14798 ( .A1(n12213), .A2(n12663), .ZN(n15190) );
  INV_X1 U14799 ( .A(n15190), .ZN(n12214) );
  AOI21_X1 U14800 ( .B1(n12225), .B2(n12278), .A(n12214), .ZN(n15361) );
  NAND2_X1 U14801 ( .A1(n15158), .A2(n15354), .ZN(n12216) );
  AOI22_X1 U14802 ( .A1(n15584), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n14768), 
        .B2(n15573), .ZN(n12215) );
  OAI211_X1 U14803 ( .C1(n12217), .C2(n15162), .A(n12216), .B(n12215), .ZN(
        n12221) );
  AOI21_X1 U14804 ( .B1(n12218), .B2(n15352), .A(n15574), .ZN(n12219) );
  NAND2_X1 U14805 ( .A1(n12219), .A2(n15198), .ZN(n15356) );
  NOR2_X1 U14806 ( .A1(n15356), .A2(n15185), .ZN(n12220) );
  AOI211_X1 U14807 ( .C1(n15212), .C2(n15352), .A(n12221), .B(n12220), .ZN(
        n12228) );
  INV_X1 U14808 ( .A(n12222), .ZN(n12223) );
  NAND2_X1 U14809 ( .A1(n12226), .A2(n12225), .ZN(n15203) );
  OAI211_X1 U14810 ( .C1(n12226), .C2(n12225), .A(n15568), .B(n15203), .ZN(
        n15359) );
  OR2_X1 U14811 ( .A1(n15359), .A2(n15584), .ZN(n12227) );
  OAI211_X1 U14812 ( .C1(n15361), .C2(n15214), .A(n12228), .B(n12227), .ZN(
        P1_U3280) );
  XOR2_X1 U14813 ( .A(n12230), .B(n12229), .Z(n12237) );
  AOI21_X1 U14814 ( .B1(n14779), .B2(n15353), .A(n12231), .ZN(n12234) );
  NAND2_X1 U14815 ( .A1(n14813), .A2(n12232), .ZN(n12233) );
  OAI211_X1 U14816 ( .C1(n15384), .C2(n14798), .A(n12234), .B(n12233), .ZN(
        n12235) );
  AOI21_X1 U14817 ( .B1(n14769), .B2(n15372), .A(n12235), .ZN(n12236) );
  OAI21_X1 U14818 ( .B1(n12237), .B2(n14815), .A(n12236), .ZN(P1_U3236) );
  OAI21_X1 U14819 ( .B1(n12239), .B2(n12774), .A(n12238), .ZN(n13657) );
  INV_X1 U14820 ( .A(n13657), .ZN(n12250) );
  OR2_X1 U14821 ( .A1(n12241), .A2(n12240), .ZN(n12243) );
  NAND2_X1 U14822 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  AOI211_X1 U14823 ( .C1(n12774), .C2(n12244), .A(n13507), .B(n7642), .ZN(
        n12246) );
  OAI22_X1 U14824 ( .A1(n13085), .A2(n13509), .B1(n13027), .B2(n13511), .ZN(
        n12245) );
  OR2_X1 U14825 ( .A1(n12246), .A2(n12245), .ZN(n13656) );
  INV_X1 U14826 ( .A(n13030), .ZN(n13712) );
  AOI22_X1 U14827 ( .A1(n13580), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13579), 
        .B2(n13029), .ZN(n12247) );
  OAI21_X1 U14828 ( .B1(n13712), .B2(n13582), .A(n12247), .ZN(n12248) );
  AOI21_X1 U14829 ( .B1(n13656), .B2(n13574), .A(n12248), .ZN(n12249) );
  OAI21_X1 U14830 ( .B1(n12250), .B2(n13588), .A(n12249), .ZN(P3_U3221) );
  NAND2_X1 U14831 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  XNOR2_X1 U14832 ( .A(n12847), .B(n12385), .ZN(n12303) );
  XNOR2_X1 U14833 ( .A(n12303), .B(n13087), .ZN(n12256) );
  AOI21_X1 U14834 ( .B1(n12255), .B2(n12256), .A(n15867), .ZN(n12258) );
  INV_X1 U14835 ( .A(n12256), .ZN(n12257) );
  NAND2_X1 U14836 ( .A1(n12258), .A2(n12305), .ZN(n12263) );
  NAND2_X1 U14837 ( .A1(n13130), .A2(n13145), .ZN(n12260) );
  OAI211_X1 U14838 ( .C1(n15874), .C2(n13085), .A(n12260), .B(n12259), .ZN(
        n12261) );
  AOI21_X1 U14839 ( .B1(n12264), .B2(n13133), .A(n12261), .ZN(n12262) );
  OAI211_X1 U14840 ( .C1(n13136), .C2(n12847), .A(n12263), .B(n12262), .ZN(
        P3_U3157) );
  INV_X1 U14841 ( .A(n12264), .ZN(n12265) );
  OAI22_X1 U14842 ( .A1(n13582), .A2(n12847), .B1(n12265), .B2(n13553), .ZN(
        n12268) );
  MUX2_X1 U14843 ( .A(n12266), .B(P3_REG2_REG_10__SCAN_IN), .S(n13580), .Z(
        n12267) );
  AOI211_X1 U14844 ( .C1(n13551), .C2(n12269), .A(n12268), .B(n12267), .ZN(
        n12270) );
  INV_X1 U14845 ( .A(n12270), .ZN(P3_U3223) );
  INV_X1 U14846 ( .A(n12271), .ZN(n12272) );
  OAI222_X1 U14847 ( .A1(n9637), .A2(P3_U3151), .B1(n13731), .B2(n12273), .C1(
        n13729), .C2(n12272), .ZN(P3_U3271) );
  XNOR2_X1 U14848 ( .A(n12275), .B(n12274), .ZN(n15343) );
  OAI211_X1 U14849 ( .C1(n12278), .C2(n12277), .A(n12276), .B(n12664), .ZN(
        n12280) );
  NAND2_X1 U14850 ( .A1(n12280), .A2(n12279), .ZN(n15341) );
  OAI211_X1 U14851 ( .C1(n15201), .C2(n15339), .A(n15174), .B(n15540), .ZN(
        n15338) );
  NOR2_X1 U14852 ( .A1(n15178), .A2(n15497), .ZN(n12284) );
  NOR2_X1 U14853 ( .A1(n14766), .A2(n15630), .ZN(n12281) );
  AOI21_X1 U14854 ( .B1(n14819), .B2(n15668), .A(n12281), .ZN(n15337) );
  INV_X1 U14855 ( .A(n14812), .ZN(n12282) );
  OAI22_X1 U14856 ( .A1(n15584), .A2(n15337), .B1(n12282), .B2(n15549), .ZN(
        n12283) );
  AOI211_X1 U14857 ( .C1(n12585), .C2(n15212), .A(n12284), .B(n12283), .ZN(
        n12285) );
  OAI21_X1 U14858 ( .B1(n15338), .B2(n15185), .A(n12285), .ZN(n12286) );
  AOI21_X1 U14859 ( .B1(n15341), .B2(n15581), .A(n12286), .ZN(n12287) );
  OAI21_X1 U14860 ( .B1(n15343), .B2(n15095), .A(n12287), .ZN(P1_U3278) );
  OAI211_X1 U14861 ( .C1(n12290), .C2(n12289), .A(n12288), .B(n15491), .ZN(
        n12296) );
  AOI21_X1 U14862 ( .B1(n14779), .B2(n15363), .A(n12291), .ZN(n12292) );
  OAI21_X1 U14863 ( .B1(n12565), .B2(n14798), .A(n12292), .ZN(n12293) );
  AOI21_X1 U14864 ( .B1(n12294), .B2(n14813), .A(n12293), .ZN(n12295) );
  OAI211_X1 U14865 ( .C1(n6549), .C2(n14809), .A(n12296), .B(n12295), .ZN(
        P1_U3224) );
  INV_X1 U14866 ( .A(n12297), .ZN(n12298) );
  OAI222_X1 U14867 ( .A1(n12300), .A2(P3_U3151), .B1(n13731), .B2(n12299), 
        .C1(n13725), .C2(n12298), .ZN(P3_U3270) );
  INV_X1 U14868 ( .A(n12301), .ZN(n12400) );
  OAI222_X1 U14869 ( .A1(n15433), .A2(n12302), .B1(n6554), .B2(n12400), .C1(
        P1_U3086), .C2(n12696), .ZN(P1_U3328) );
  NAND2_X1 U14870 ( .A1(n12303), .A2(n13087), .ZN(n12304) );
  XNOR2_X1 U14871 ( .A(n13095), .B(n11664), .ZN(n13019) );
  XNOR2_X1 U14872 ( .A(n13030), .B(n11664), .ZN(n13022) );
  NAND2_X1 U14873 ( .A1(n13022), .A2(n13143), .ZN(n12308) );
  OAI21_X1 U14874 ( .B1(n13085), .B2(n13019), .A(n12308), .ZN(n12310) );
  AND2_X1 U14875 ( .A1(n13019), .A2(n13085), .ZN(n12307) );
  INV_X1 U14876 ( .A(n13022), .ZN(n12306) );
  AOI22_X1 U14877 ( .A1(n12308), .A2(n12307), .B1(n13090), .B2(n12306), .ZN(
        n12309) );
  XNOR2_X1 U14878 ( .A(n13583), .B(n11664), .ZN(n12343) );
  XNOR2_X1 U14879 ( .A(n12343), .B(n13027), .ZN(n12311) );
  XNOR2_X1 U14880 ( .A(n12345), .B(n12311), .ZN(n12317) );
  NAND2_X1 U14881 ( .A1(n13130), .A2(n13143), .ZN(n12312) );
  NAND2_X1 U14882 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13175)
         );
  OAI211_X1 U14883 ( .C1(n15874), .C2(n12313), .A(n12312), .B(n13175), .ZN(
        n12315) );
  NOR2_X1 U14884 ( .A1(n13583), .A2(n13136), .ZN(n12314) );
  AOI211_X1 U14885 ( .C1(n13578), .C2(n13133), .A(n12315), .B(n12314), .ZN(
        n12316) );
  OAI21_X1 U14886 ( .B1(n12317), .B2(n15867), .A(n12316), .ZN(P3_U3174) );
  INV_X1 U14887 ( .A(n12318), .ZN(n15429) );
  OAI222_X1 U14888 ( .A1(n11978), .A2(n15429), .B1(P2_U3088), .B2(n12319), 
        .C1(n12734), .C2(n12702), .ZN(P2_U3298) );
  INV_X1 U14889 ( .A(SI_26_), .ZN(n12322) );
  INV_X1 U14890 ( .A(n12320), .ZN(n12321) );
  OAI222_X1 U14891 ( .A1(n12323), .A2(P3_U3151), .B1(n13731), .B2(n12322), 
        .C1(n13729), .C2(n12321), .ZN(P3_U3269) );
  INV_X1 U14892 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12329) );
  XNOR2_X1 U14893 ( .A(n12324), .B(n9569), .ZN(n13577) );
  NOR2_X1 U14894 ( .A1(n7642), .A2(n12325), .ZN(n12326) );
  XNOR2_X1 U14895 ( .A(n12326), .B(n9569), .ZN(n12328) );
  AOI22_X1 U14896 ( .A1(n13566), .A2(n13545), .B1(n13143), .B2(n13567), .ZN(
        n12327) );
  OAI21_X1 U14897 ( .B1(n12328), .B2(n13507), .A(n12327), .ZN(n13586) );
  AOI21_X1 U14898 ( .B1(n13577), .B2(n15905), .A(n13586), .ZN(n12331) );
  MUX2_X1 U14899 ( .A(n12329), .B(n12331), .S(n15943), .Z(n12330) );
  OAI21_X1 U14900 ( .B1(n13711), .B2(n13583), .A(n12330), .ZN(P3_U3429) );
  INV_X1 U14901 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13164) );
  MUX2_X1 U14902 ( .A(n13164), .B(n12331), .S(n15954), .Z(n12332) );
  OAI21_X1 U14903 ( .B1(n13660), .B2(n13583), .A(n12332), .ZN(P3_U3472) );
  XOR2_X1 U14904 ( .A(n12334), .B(n12333), .Z(n12335) );
  XNOR2_X1 U14905 ( .A(n12336), .B(n12335), .ZN(n12342) );
  NOR2_X1 U14906 ( .A1(n14809), .A2(n15659), .ZN(n12340) );
  NAND2_X1 U14907 ( .A1(n14806), .A2(n15532), .ZN(n12337) );
  NAND2_X1 U14908 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n14883) );
  OAI211_X1 U14909 ( .C1(n14808), .C2(n12338), .A(n12337), .B(n14883), .ZN(
        n12339) );
  AOI211_X1 U14910 ( .C1(n14813), .C2(n15536), .A(n12340), .B(n12339), .ZN(
        n12341) );
  OAI21_X1 U14911 ( .B1(n12342), .B2(n14815), .A(n12341), .ZN(P1_U3227) );
  INV_X1 U14912 ( .A(n12343), .ZN(n12344) );
  XNOR2_X1 U14913 ( .A(n13707), .B(n11664), .ZN(n12346) );
  XNOR2_X1 U14914 ( .A(n12346), .B(n13545), .ZN(n12965) );
  INV_X1 U14915 ( .A(n12346), .ZN(n12347) );
  XNOR2_X1 U14916 ( .A(n13651), .B(n11664), .ZN(n12348) );
  XNOR2_X1 U14917 ( .A(n12348), .B(n13565), .ZN(n13127) );
  NAND2_X1 U14918 ( .A1(n13126), .A2(n13127), .ZN(n13125) );
  NAND2_X1 U14919 ( .A1(n12348), .A2(n12968), .ZN(n12349) );
  XNOR2_X1 U14920 ( .A(n13541), .B(n11664), .ZN(n12351) );
  XNOR2_X1 U14921 ( .A(n13546), .B(n12351), .ZN(n13041) );
  NAND2_X1 U14922 ( .A1(n12351), .A2(n13546), .ZN(n12352) );
  XNOR2_X1 U14923 ( .A(n13643), .B(n11664), .ZN(n12353) );
  XNOR2_X1 U14924 ( .A(n12353), .B(n13527), .ZN(n13050) );
  INV_X1 U14925 ( .A(n12353), .ZN(n12354) );
  NAND2_X1 U14926 ( .A1(n12354), .A2(n13527), .ZN(n12355) );
  XNOR2_X1 U14927 ( .A(n13492), .B(n11664), .ZN(n13096) );
  AND2_X1 U14928 ( .A1(n13096), .A2(n13141), .ZN(n12358) );
  INV_X1 U14929 ( .A(n13096), .ZN(n12357) );
  XNOR2_X1 U14930 ( .A(n12990), .B(n12385), .ZN(n12359) );
  XNOR2_X1 U14931 ( .A(n12359), .B(n13499), .ZN(n12992) );
  INV_X1 U14932 ( .A(n12359), .ZN(n12360) );
  NAND2_X1 U14933 ( .A1(n12360), .A2(n13499), .ZN(n12361) );
  XNOR2_X1 U14934 ( .A(n13628), .B(n12385), .ZN(n12362) );
  XNOR2_X1 U14935 ( .A(n12362), .B(n13013), .ZN(n13069) );
  INV_X1 U14936 ( .A(n12362), .ZN(n12363) );
  NAND2_X1 U14937 ( .A1(n12363), .A2(n13013), .ZN(n12364) );
  XNOR2_X1 U14938 ( .A(n13459), .B(n11664), .ZN(n12366) );
  XNOR2_X1 U14939 ( .A(n12366), .B(n13140), .ZN(n13012) );
  INV_X1 U14940 ( .A(n12366), .ZN(n12367) );
  NAND2_X1 U14941 ( .A1(n12367), .A2(n13474), .ZN(n12368) );
  XNOR2_X1 U14942 ( .A(n13610), .B(n12385), .ZN(n12418) );
  INV_X1 U14943 ( .A(n12418), .ZN(n12369) );
  AOI22_X1 U14944 ( .A1(n12369), .A2(n13428), .B1(n6534), .B2(n13139), .ZN(
        n12372) );
  XNOR2_X1 U14945 ( .A(n13080), .B(n11664), .ZN(n12413) );
  INV_X1 U14946 ( .A(n12413), .ZN(n12414) );
  AND2_X1 U14947 ( .A1(n12372), .A2(n12370), .ZN(n12371) );
  INV_X1 U14948 ( .A(n12372), .ZN(n12374) );
  NAND2_X1 U14949 ( .A1(n12414), .A2(n13458), .ZN(n12373) );
  NOR2_X1 U14950 ( .A1(n12374), .A2(n12373), .ZN(n12379) );
  OAI21_X1 U14951 ( .B1(n6534), .B2(n13139), .A(n13428), .ZN(n12376) );
  NOR3_X1 U14952 ( .A1(n6534), .A2(n13139), .A3(n13428), .ZN(n12375) );
  AOI21_X1 U14953 ( .B1(n12418), .B2(n12376), .A(n12375), .ZN(n12377) );
  INV_X1 U14954 ( .A(n12377), .ZN(n12378) );
  NAND2_X1 U14955 ( .A1(n12381), .A2(n12380), .ZN(n13034) );
  XNOR2_X1 U14956 ( .A(n13399), .B(n11664), .ZN(n12382) );
  XNOR2_X1 U14957 ( .A(n12382), .B(n13410), .ZN(n13035) );
  INV_X1 U14958 ( .A(n12382), .ZN(n12383) );
  XNOR2_X1 U14959 ( .A(n9594), .B(n11664), .ZN(n12384) );
  XNOR2_X1 U14960 ( .A(n12384), .B(n13385), .ZN(n13118) );
  XNOR2_X1 U14961 ( .A(n13674), .B(n12385), .ZN(n12386) );
  XNOR2_X1 U14962 ( .A(n12386), .B(n13343), .ZN(n12959) );
  XNOR2_X1 U14963 ( .A(n13338), .B(n11664), .ZN(n12387) );
  AOI22_X1 U14964 ( .A1(n13349), .A2(n13133), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12389) );
  NAND2_X1 U14965 ( .A1(n13343), .A2(n13110), .ZN(n12388) );
  OAI211_X1 U14966 ( .C1(n13345), .C2(n15874), .A(n12389), .B(n12388), .ZN(
        n12390) );
  AOI21_X1 U14967 ( .B1(n9525), .B2(n15870), .A(n12390), .ZN(n12391) );
  OAI21_X1 U14968 ( .B1(n12392), .B2(n15867), .A(n12391), .ZN(P3_U3160) );
  XNOR2_X1 U14969 ( .A(n12708), .B(n12395), .ZN(n12393) );
  NAND2_X1 U14970 ( .A1(n12393), .A2(n10957), .ZN(n14512) );
  NAND2_X1 U14971 ( .A1(n12394), .A2(n14015), .ZN(n14514) );
  NOR2_X1 U14972 ( .A1(n14484), .A2(n14514), .ZN(n12712) );
  INV_X1 U14973 ( .A(n12395), .ZN(n14513) );
  NOR2_X1 U14974 ( .A1(n14513), .A2(n14486), .ZN(n12396) );
  AOI211_X1 U14975 ( .C1(P2_REG2_REG_31__SCAN_IN), .C2(n14484), .A(n12712), 
        .B(n12396), .ZN(n12397) );
  OAI21_X1 U14976 ( .B1(n14507), .B2(n14512), .A(n12397), .ZN(P2_U3234) );
  OAI222_X1 U14977 ( .A1(n14659), .A2(n12401), .B1(n11978), .B2(n12400), .C1(
        n12399), .C2(P2_U3088), .ZN(P2_U3300) );
  XNOR2_X1 U14978 ( .A(n12798), .B(n12802), .ZN(n15900) );
  OAI21_X1 U14979 ( .B1(n12798), .B2(n12403), .A(n12402), .ZN(n12404) );
  NAND2_X1 U14980 ( .A1(n12404), .A2(n13562), .ZN(n12406) );
  AOI22_X1 U14981 ( .A1(n11672), .A2(n13566), .B1(n13567), .B2(n11047), .ZN(
        n12405) );
  NAND2_X1 U14982 ( .A1(n12406), .A2(n12405), .ZN(n15902) );
  NAND2_X1 U14983 ( .A1(n12407), .A2(n15936), .ZN(n15901) );
  OAI22_X1 U14984 ( .A1(n13553), .A2(n12408), .B1(n15901), .B2(n12936), .ZN(
        n12409) );
  NOR2_X1 U14985 ( .A1(n15902), .A2(n12409), .ZN(n12411) );
  MUX2_X1 U14986 ( .A(n12411), .B(n12410), .S(n13580), .Z(n12412) );
  OAI21_X1 U14987 ( .B1(n15900), .B2(n13588), .A(n12412), .ZN(P3_U3232) );
  AOI22_X1 U14988 ( .A1(n13139), .A2(n13110), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12420) );
  NAND2_X1 U14989 ( .A1(n13414), .A2(n13133), .ZN(n12419) );
  OAI211_X1 U14990 ( .C1(n13410), .C2(n15874), .A(n12420), .B(n12419), .ZN(
        n12421) );
  AOI21_X1 U14991 ( .B1(n13610), .B2(n15870), .A(n12421), .ZN(n12422) );
  OAI222_X1 U14992 ( .A1(n13725), .A2(n12425), .B1(n12424), .B2(P3_U3151), 
        .C1(n12423), .C2(n13731), .ZN(P3_U3267) );
  INV_X1 U14993 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14973) );
  NAND2_X1 U14994 ( .A1(n10216), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U14995 ( .A1(n8145), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12427) );
  OAI211_X1 U14996 ( .C1(n12429), .C2(n14973), .A(n12428), .B(n12427), .ZN(
        n14971) );
  OAI21_X1 U14997 ( .B1(n12430), .B2(n14971), .A(n14817), .ZN(n12444) );
  INV_X1 U14998 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U14999 ( .A1(n15419), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15000 ( .A1(n12431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n12432) );
  AND2_X1 U15001 ( .A1(n12433), .A2(n12432), .ZN(n12437) );
  INV_X1 U15002 ( .A(n12437), .ZN(n12441) );
  NAND2_X1 U15003 ( .A1(n12434), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n12435) );
  OAI211_X1 U15004 ( .C1(P1_IR_REG_20__SCAN_IN), .C2(P1_IR_REG_22__SCAN_IN), 
        .A(n12435), .B(P1_IR_REG_31__SCAN_IN), .ZN(n12436) );
  OAI22_X1 U15005 ( .A1(n12438), .A2(n12437), .B1(n7763), .B2(n12436), .ZN(
        n12439) );
  INV_X1 U15006 ( .A(n12439), .ZN(n12440) );
  NAND2_X4 U15007 ( .A1(n12443), .A2(n12442), .ZN(n12625) );
  INV_X1 U15008 ( .A(n14817), .ZN(n12447) );
  AOI22_X1 U15009 ( .A1(n14971), .A2(n12625), .B1(n12646), .B2(n12445), .ZN(
        n12446) );
  INV_X1 U15010 ( .A(n15241), .ZN(n14988) );
  MUX2_X1 U15011 ( .A(n15241), .B(n15237), .S(n12625), .Z(n12455) );
  MUX2_X1 U15012 ( .A(n15223), .B(n15244), .S(n12625), .Z(n12463) );
  MUX2_X1 U15013 ( .A(n15252), .B(n15224), .S(n12642), .Z(n12464) );
  INV_X1 U15014 ( .A(n12464), .ZN(n12452) );
  NAND2_X1 U15015 ( .A1(n12465), .A2(n12452), .ZN(n12456) );
  INV_X1 U15016 ( .A(n12453), .ZN(n12458) );
  NAND2_X1 U15017 ( .A1(n12455), .A2(n12454), .ZN(n12457) );
  OAI22_X1 U15018 ( .A1(n12467), .A2(n12456), .B1(n12458), .B2(n12457), .ZN(
        n12462) );
  NAND2_X1 U15019 ( .A1(n12458), .A2(n12457), .ZN(n12460) );
  AND2_X1 U15020 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  MUX2_X1 U15021 ( .A(n15016), .B(n15255), .S(n12619), .Z(n12472) );
  MUX2_X1 U15022 ( .A(n15242), .B(n15003), .S(n12625), .Z(n12473) );
  INV_X1 U15023 ( .A(n12473), .ZN(n12468) );
  INV_X1 U15024 ( .A(n12472), .ZN(n12474) );
  NAND2_X1 U15025 ( .A1(n12474), .A2(n12468), .ZN(n12475) );
  NAND2_X1 U15026 ( .A1(n12476), .A2(n12475), .ZN(n12482) );
  MUX2_X1 U15027 ( .A(n15028), .B(n15020), .S(n12625), .Z(n12483) );
  INV_X1 U15028 ( .A(n12483), .ZN(n12478) );
  MUX2_X1 U15029 ( .A(n15251), .B(n15261), .S(n12642), .Z(n12484) );
  INV_X1 U15030 ( .A(n12484), .ZN(n12477) );
  MUX2_X1 U15031 ( .A(n15015), .B(n15034), .S(n12625), .Z(n12631) );
  INV_X1 U15032 ( .A(n12631), .ZN(n12481) );
  MUX2_X1 U15033 ( .A(n15274), .B(n15267), .S(n12642), .Z(n12632) );
  INV_X1 U15034 ( .A(n12632), .ZN(n12480) );
  INV_X1 U15035 ( .A(n12482), .ZN(n12485) );
  NAND3_X1 U15036 ( .A1(n12485), .A2(n12478), .A3(n12477), .ZN(n12486) );
  MUX2_X1 U15037 ( .A(n14766), .B(n15346), .S(n12619), .Z(n12584) );
  NAND2_X1 U15038 ( .A1(n12490), .A2(n12491), .ZN(n12489) );
  NAND2_X1 U15039 ( .A1(n15567), .A2(n12489), .ZN(n12494) );
  NAND2_X1 U15040 ( .A1(n12499), .A2(n12496), .ZN(n12498) );
  NAND2_X1 U15041 ( .A1(n12498), .A2(n12497), .ZN(n12506) );
  INV_X1 U15042 ( .A(n12499), .ZN(n12500) );
  NAND2_X1 U15043 ( .A1(n12500), .A2(n6804), .ZN(n12505) );
  OAI211_X1 U15044 ( .C1(n12501), .C2(n15566), .A(n6593), .B(n12625), .ZN(
        n12503) );
  NAND3_X1 U15045 ( .A1(n12501), .A2(n15566), .A3(n12625), .ZN(n12502) );
  NAND3_X1 U15046 ( .A1(n12506), .A2(n12505), .A3(n12504), .ZN(n12513) );
  MUX2_X1 U15047 ( .A(n15486), .B(n12508), .S(n12625), .Z(n12512) );
  MUX2_X1 U15048 ( .A(n15486), .B(n12508), .S(n12507), .Z(n12509) );
  INV_X1 U15049 ( .A(n12509), .ZN(n12510) );
  AOI21_X1 U15050 ( .B1(n12513), .B2(n12512), .A(n12510), .ZN(n12518) );
  OAI21_X1 U15051 ( .B1(n12513), .B2(n12512), .A(n12511), .ZN(n12517) );
  MUX2_X1 U15052 ( .A(n12515), .B(n12514), .S(n12619), .Z(n12516) );
  OAI21_X1 U15053 ( .B1(n12518), .B2(n12517), .A(n12516), .ZN(n12523) );
  MUX2_X1 U15054 ( .A(n15487), .B(n12519), .S(n12625), .Z(n12522) );
  MUX2_X1 U15055 ( .A(n15532), .B(n12520), .S(n12619), .Z(n12521) );
  NAND2_X1 U15056 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  MUX2_X1 U15057 ( .A(n15666), .B(n12526), .S(n12619), .Z(n12528) );
  MUX2_X1 U15058 ( .A(n12526), .B(n15666), .S(n12619), .Z(n12527) );
  INV_X1 U15059 ( .A(n12528), .ZN(n12529) );
  MUX2_X1 U15060 ( .A(n12530), .B(n15531), .S(n12619), .Z(n12534) );
  NAND2_X1 U15061 ( .A1(n12533), .A2(n12534), .ZN(n12532) );
  MUX2_X1 U15062 ( .A(n15531), .B(n12530), .S(n12619), .Z(n12531) );
  NAND2_X1 U15063 ( .A1(n12532), .A2(n12531), .ZN(n12545) );
  INV_X1 U15064 ( .A(n12533), .ZN(n12536) );
  INV_X1 U15065 ( .A(n12534), .ZN(n12535) );
  NAND2_X1 U15066 ( .A1(n12536), .A2(n12535), .ZN(n12542) );
  NAND2_X1 U15067 ( .A1(n12545), .A2(n12542), .ZN(n12537) );
  MUX2_X1 U15068 ( .A(n15667), .B(n12538), .S(n12619), .Z(n12541) );
  NAND2_X1 U15069 ( .A1(n12537), .A2(n12541), .ZN(n12540) );
  MUX2_X1 U15070 ( .A(n15667), .B(n12538), .S(n12625), .Z(n12539) );
  NAND2_X1 U15071 ( .A1(n12540), .A2(n12539), .ZN(n12547) );
  INV_X1 U15072 ( .A(n12541), .ZN(n12543) );
  AND2_X1 U15073 ( .A1(n12543), .A2(n12542), .ZN(n12544) );
  NAND2_X1 U15074 ( .A1(n12545), .A2(n12544), .ZN(n12546) );
  NAND2_X1 U15075 ( .A1(n12547), .A2(n12546), .ZN(n12551) );
  MUX2_X1 U15076 ( .A(n15514), .B(n12548), .S(n12625), .Z(n12552) );
  NAND2_X1 U15077 ( .A1(n12551), .A2(n12552), .ZN(n12550) );
  MUX2_X1 U15078 ( .A(n15514), .B(n12548), .S(n12619), .Z(n12549) );
  NAND2_X1 U15079 ( .A1(n12550), .A2(n12549), .ZN(n12556) );
  INV_X1 U15080 ( .A(n12551), .ZN(n12554) );
  INV_X1 U15081 ( .A(n12552), .ZN(n12553) );
  NAND2_X1 U15082 ( .A1(n12554), .A2(n12553), .ZN(n12555) );
  MUX2_X1 U15083 ( .A(n14821), .B(n15389), .S(n12619), .Z(n12558) );
  MUX2_X1 U15084 ( .A(n14821), .B(n15389), .S(n12625), .Z(n12557) );
  MUX2_X1 U15085 ( .A(n15362), .B(n15372), .S(n12619), .Z(n12568) );
  NAND2_X1 U15086 ( .A1(n15362), .A2(n12642), .ZN(n12560) );
  NAND2_X1 U15087 ( .A1(n15372), .A2(n12625), .ZN(n12559) );
  NAND3_X1 U15088 ( .A1(n12568), .A2(n12560), .A3(n12559), .ZN(n12561) );
  AND2_X1 U15089 ( .A1(n12569), .A2(n12561), .ZN(n12572) );
  MUX2_X1 U15090 ( .A(n15384), .B(n15378), .S(n12625), .Z(n12574) );
  MUX2_X1 U15091 ( .A(n14820), .B(n12562), .S(n12619), .Z(n12573) );
  NAND2_X1 U15092 ( .A1(n12574), .A2(n12573), .ZN(n12563) );
  OAI21_X1 U15093 ( .B1(n6549), .B2(n15353), .A(n12580), .ZN(n12571) );
  NAND2_X1 U15094 ( .A1(n12565), .A2(n12642), .ZN(n12566) );
  OAI21_X1 U15095 ( .B1(n15372), .B2(n12642), .A(n12566), .ZN(n12567) );
  NOR2_X1 U15096 ( .A1(n12568), .A2(n12567), .ZN(n12570) );
  AOI22_X1 U15097 ( .A1(n12571), .A2(n12625), .B1(n12570), .B2(n12569), .ZN(
        n12577) );
  INV_X1 U15098 ( .A(n12572), .ZN(n12575) );
  AOI21_X1 U15099 ( .B1(n12579), .B2(n15202), .A(n7645), .ZN(n12582) );
  NOR2_X1 U15100 ( .A1(n12580), .A2(n12625), .ZN(n12581) );
  MUX2_X1 U15101 ( .A(n15211), .B(n15354), .S(n12619), .Z(n12583) );
  MUX2_X1 U15102 ( .A(n12585), .B(n15344), .S(n12619), .Z(n12587) );
  MUX2_X1 U15103 ( .A(n15344), .B(n12585), .S(n12619), .Z(n12590) );
  INV_X1 U15104 ( .A(n12586), .ZN(n12589) );
  INV_X1 U15105 ( .A(n12587), .ZN(n12588) );
  MUX2_X1 U15106 ( .A(n15321), .B(n15332), .S(n12642), .Z(n12596) );
  NOR2_X1 U15107 ( .A1(n12592), .A2(n15329), .ZN(n12598) );
  MUX2_X1 U15108 ( .A(n12597), .B(n12598), .S(n12619), .Z(n12593) );
  INV_X1 U15109 ( .A(n12593), .ZN(n12594) );
  MUX2_X1 U15110 ( .A(n14819), .B(n15183), .S(n12625), .Z(n12595) );
  MUX2_X1 U15111 ( .A(n12598), .B(n12597), .S(n12619), .Z(n12599) );
  INV_X1 U15112 ( .A(n12602), .ZN(n12605) );
  MUX2_X1 U15113 ( .A(n15322), .B(n15315), .S(n12619), .Z(n12601) );
  INV_X1 U15114 ( .A(n12601), .ZN(n12604) );
  XNOR2_X1 U15115 ( .A(n15131), .B(n15314), .ZN(n15120) );
  INV_X1 U15116 ( .A(n15315), .ZN(n15143) );
  MUX2_X1 U15117 ( .A(n15143), .B(n15305), .S(n12619), .Z(n12600) );
  AOI21_X1 U15118 ( .B1(n12602), .B2(n12601), .A(n12600), .ZN(n12603) );
  NOR2_X1 U15119 ( .A1(n15314), .A2(n12625), .ZN(n12607) );
  NOR2_X1 U15120 ( .A1(n15145), .A2(n12642), .ZN(n12606) );
  MUX2_X1 U15121 ( .A(n12607), .B(n12606), .S(n15131), .Z(n12608) );
  MUX2_X1 U15122 ( .A(n15306), .B(n10129), .S(n12619), .Z(n12610) );
  MUX2_X1 U15123 ( .A(n10129), .B(n15306), .S(n12619), .Z(n12611) );
  MUX2_X1 U15124 ( .A(n15091), .B(n14818), .S(n12619), .Z(n12615) );
  MUX2_X1 U15125 ( .A(n14818), .B(n15091), .S(n12619), .Z(n12612) );
  NAND2_X1 U15126 ( .A1(n12613), .A2(n12612), .ZN(n12618) );
  INV_X1 U15127 ( .A(n12615), .ZN(n12616) );
  AND2_X1 U15128 ( .A1(n12618), .A2(n12617), .ZN(n12622) );
  MUX2_X1 U15129 ( .A(n15089), .B(n15076), .S(n12619), .Z(n12621) );
  MUX2_X1 U15130 ( .A(n7418), .B(n15294), .S(n12619), .Z(n12620) );
  NAND2_X1 U15131 ( .A1(n12622), .A2(n12621), .ZN(n12623) );
  NAND2_X1 U15132 ( .A1(n12624), .A2(n12623), .ZN(n12628) );
  MUX2_X1 U15133 ( .A(n15062), .B(n15045), .S(n12642), .Z(n12627) );
  MUX2_X1 U15134 ( .A(n14688), .B(n14752), .S(n12642), .Z(n12630) );
  MUX2_X1 U15135 ( .A(n15057), .B(n15276), .S(n12625), .Z(n12629) );
  OAI22_X1 U15136 ( .A1(n12628), .A2(n12627), .B1(n12630), .B2(n12629), .ZN(
        n12637) );
  MUX2_X1 U15137 ( .A(n15273), .B(n15285), .S(n12642), .Z(n12626) );
  AOI21_X1 U15138 ( .B1(n12628), .B2(n12627), .A(n12626), .ZN(n12636) );
  AOI22_X1 U15139 ( .A1(n12632), .A2(n12631), .B1(n12630), .B2(n12629), .ZN(
        n12633) );
  OAI21_X1 U15140 ( .B1(n12637), .B2(n12636), .A(n12635), .ZN(n12638) );
  NAND2_X1 U15141 ( .A1(n6604), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15142 ( .A1(n14971), .A2(n12642), .ZN(n12684) );
  NOR2_X1 U15143 ( .A1(n14971), .A2(n12642), .ZN(n12685) );
  NAND2_X1 U15144 ( .A1(n15215), .A2(n12685), .ZN(n12647) );
  NAND2_X1 U15145 ( .A1(n12643), .A2(n11002), .ZN(n12644) );
  NAND2_X1 U15146 ( .A1(n12644), .A2(n15149), .ZN(n12678) );
  NAND2_X1 U15147 ( .A1(n12646), .A2(n12645), .ZN(n12675) );
  AND2_X1 U15148 ( .A1(n12678), .A2(n12675), .ZN(n12681) );
  OAI211_X1 U15149 ( .C1(n15215), .C2(n12684), .A(n12647), .B(n12681), .ZN(
        n12676) );
  XOR2_X1 U15150 ( .A(n14817), .B(n14968), .Z(n12672) );
  XNOR2_X1 U15151 ( .A(n15143), .B(n15322), .ZN(n15138) );
  NAND2_X1 U15152 ( .A1(n12649), .A2(n12648), .ZN(n15578) );
  NOR3_X1 U15153 ( .A1(n15546), .A2(n15578), .A3(n12650), .ZN(n12654) );
  NAND4_X1 U15154 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12656) );
  NOR3_X1 U15155 ( .A1(n12656), .A2(n15512), .A3(n12655), .ZN(n12659) );
  NAND4_X1 U15156 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12661) );
  XNOR2_X1 U15157 ( .A(n15211), .B(n15354), .ZN(n15204) );
  NAND4_X1 U15158 ( .A1(n12665), .A2(n15170), .A3(n12664), .A4(n15204), .ZN(
        n12666) );
  NAND4_X1 U15159 ( .A1(n15039), .A2(n12667), .A3(n15108), .A4(n15055), .ZN(
        n12668) );
  NOR4_X1 U15160 ( .A1(n12669), .A2(n12668), .A3(n15082), .A4(n15069), .ZN(
        n12670) );
  NAND4_X1 U15161 ( .A1(n14983), .A2(n12670), .A3(n15007), .A4(n15013), .ZN(
        n12671) );
  XOR2_X1 U15162 ( .A(n15207), .B(n12673), .Z(n12674) );
  OAI22_X1 U15163 ( .A1(n12680), .A2(n12676), .B1(n12675), .B2(n12674), .ZN(
        n12695) );
  INV_X1 U15164 ( .A(n12678), .ZN(n12689) );
  NOR2_X1 U15165 ( .A1(n12677), .A2(n12678), .ZN(n12679) );
  INV_X1 U15166 ( .A(n12681), .ZN(n12686) );
  INV_X1 U15167 ( .A(n14971), .ZN(n12682) );
  OAI21_X1 U15168 ( .B1(n12686), .B2(n12682), .A(n12684), .ZN(n12683) );
  OAI21_X1 U15169 ( .B1(n12689), .B2(n12684), .A(n12683), .ZN(n12691) );
  INV_X1 U15170 ( .A(n12685), .ZN(n12688) );
  OAI21_X1 U15171 ( .B1(n12686), .B2(n14971), .A(n12688), .ZN(n12687) );
  OAI21_X1 U15172 ( .B1(n12689), .B2(n12688), .A(n12687), .ZN(n12690) );
  MUX2_X1 U15173 ( .A(n12691), .B(n12690), .S(n15215), .Z(n12692) );
  NAND2_X1 U15174 ( .A1(n12693), .A2(n12692), .ZN(n12694) );
  NOR2_X1 U15175 ( .A1(n12696), .A2(P1_U3086), .ZN(n12697) );
  NAND3_X1 U15176 ( .A1(n12698), .A2(n15665), .A3(n12697), .ZN(n12699) );
  OAI211_X1 U15177 ( .C1(n6608), .C2(n12701), .A(n12699), .B(P1_B_REG_SCAN_IN), 
        .ZN(n12700) );
  INV_X1 U15178 ( .A(n12704), .ZN(n12706) );
  INV_X1 U15179 ( .A(n12708), .ZN(n12709) );
  NOR2_X1 U15180 ( .A1(n14515), .A2(n14486), .ZN(n12711) );
  AOI211_X1 U15181 ( .C1(n14484), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12712), 
        .B(n12711), .ZN(n12713) );
  OAI21_X1 U15182 ( .B1(n14518), .B2(n14507), .A(n12713), .ZN(P2_U3235) );
  INV_X1 U15183 ( .A(n12714), .ZN(n12715) );
  NAND2_X1 U15184 ( .A1(n12715), .A2(n13585), .ZN(n12719) );
  NOR2_X1 U15185 ( .A1(n12716), .A2(n13553), .ZN(n13334) );
  NOR2_X1 U15186 ( .A1(n10240), .A2(n13582), .ZN(n12717) );
  AOI211_X1 U15187 ( .C1(n13580), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13334), 
        .B(n12717), .ZN(n12718) );
  OAI211_X1 U15188 ( .C1(n12720), .C2(n13588), .A(n12719), .B(n12718), .ZN(
        P3_U3204) );
  NAND2_X1 U15189 ( .A1(n12731), .A2(n15850), .ZN(n12729) );
  OR2_X1 U15190 ( .A1(n15850), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U15191 ( .A1(n12729), .A2(n12728), .ZN(n12730) );
  OAI21_X1 U15192 ( .B1(n12733), .B2(n14649), .A(n12730), .ZN(P2_U3496) );
  OAI21_X1 U15193 ( .B1(n12733), .B2(n14586), .A(n12732), .ZN(P2_U3528) );
  INV_X1 U15194 ( .A(SI_30_), .ZN(n12743) );
  NAND2_X1 U15195 ( .A1(n12734), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12735) );
  NAND2_X1 U15196 ( .A1(n12736), .A2(n12735), .ZN(n12738) );
  NAND2_X1 U15197 ( .A1(n15427), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12737) );
  XNOR2_X1 U15198 ( .A(n12739), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12740) );
  XNOR2_X1 U15199 ( .A(n12748), .B(n12740), .ZN(n12744) );
  INV_X1 U15200 ( .A(n12744), .ZN(n12741) );
  OAI222_X1 U15201 ( .A1(n13731), .A2(n12743), .B1(n12742), .B2(P3_U3151), 
        .C1(n13725), .C2(n12741), .ZN(P3_U3265) );
  NAND2_X1 U15202 ( .A1(n12744), .A2(n9490), .ZN(n12746) );
  NAND2_X1 U15203 ( .A1(n12751), .A2(SI_30_), .ZN(n12745) );
  NOR2_X1 U15204 ( .A1(n13664), .A2(n12930), .ZN(n12785) );
  INV_X1 U15205 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15425) );
  AND2_X1 U15206 ( .A1(n15425), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12747) );
  XNOR2_X1 U15207 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12749) );
  XNOR2_X1 U15208 ( .A(n12750), .B(n12749), .ZN(n13715) );
  NAND2_X1 U15209 ( .A1(n13715), .A2(n9490), .ZN(n12753) );
  NAND2_X1 U15210 ( .A1(n12751), .A2(SI_31_), .ZN(n12752) );
  AOI21_X1 U15211 ( .B1(n12785), .B2(n13331), .A(n12935), .ZN(n12792) );
  NAND3_X1 U15212 ( .A1(n12792), .A2(n12755), .A3(n12754), .ZN(n12759) );
  NAND2_X1 U15213 ( .A1(n12755), .A2(n13316), .ZN(n12791) );
  NAND2_X1 U15214 ( .A1(n13664), .A2(n13333), .ZN(n12756) );
  MUX2_X1 U15215 ( .A(n12759), .B(n12791), .S(n12758), .Z(n12760) );
  INV_X1 U15216 ( .A(n13407), .ZN(n13403) );
  NAND2_X1 U15217 ( .A1(n12895), .A2(n12896), .ZN(n13442) );
  INV_X1 U15218 ( .A(n13564), .ZN(n12868) );
  NOR2_X1 U15219 ( .A1(n12763), .A2(n12762), .ZN(n12767) );
  NOR2_X1 U15220 ( .A1(n12798), .A2(n12764), .ZN(n12766) );
  NAND4_X1 U15221 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n15868), .ZN(
        n12768) );
  NOR2_X1 U15222 ( .A1(n12768), .A2(n12804), .ZN(n12771) );
  NOR2_X1 U15223 ( .A1(n7235), .A2(n12769), .ZN(n12770) );
  NAND4_X1 U15224 ( .A1(n12838), .A2(n12839), .A3(n12771), .A4(n12770), .ZN(
        n12772) );
  NOR2_X1 U15225 ( .A1(n12854), .A2(n12772), .ZN(n12773) );
  AND4_X1 U15226 ( .A1(n9569), .A2(n13549), .A3(n12774), .A4(n12773), .ZN(
        n12775) );
  NAND4_X1 U15227 ( .A1(n13517), .A2(n13535), .A3(n12868), .A4(n12775), .ZN(
        n12776) );
  NOR2_X1 U15228 ( .A1(n12881), .A2(n12776), .ZN(n12779) );
  NAND2_X1 U15229 ( .A1(n12778), .A2(n12777), .ZN(n13480) );
  NAND2_X1 U15230 ( .A1(n12779), .A2(n13480), .ZN(n12780) );
  NOR2_X1 U15231 ( .A1(n13442), .A2(n12780), .ZN(n12781) );
  NAND4_X1 U15232 ( .A1(n13420), .A2(n13456), .A3(n12781), .A4(n7248), .ZN(
        n12782) );
  NOR3_X1 U15233 ( .A1(n13391), .A2(n13403), .A3(n12782), .ZN(n12783) );
  NAND4_X1 U15234 ( .A1(n13340), .A2(n13372), .A3(n12783), .A4(n13365), .ZN(
        n12784) );
  NOR2_X1 U15235 ( .A1(n12914), .A2(n12784), .ZN(n12787) );
  INV_X1 U15236 ( .A(n12785), .ZN(n12786) );
  INV_X1 U15237 ( .A(n13391), .ZN(n12903) );
  AND2_X1 U15238 ( .A1(n12830), .A2(n12796), .ZN(n12824) );
  NOR2_X1 U15239 ( .A1(n12799), .A2(n12801), .ZN(n12797) );
  OAI33_X1 U15240 ( .A1(n12800), .A2(n12799), .A3(n12798), .B1(n11665), .B2(
        n12797), .B3(n9602), .ZN(n12807) );
  NAND2_X1 U15241 ( .A1(n12802), .A2(n12801), .ZN(n12806) );
  MUX2_X1 U15242 ( .A(n12803), .B(n11665), .S(n9602), .Z(n12805) );
  AOI211_X1 U15243 ( .C1(n12807), .C2(n12806), .A(n12805), .B(n12804), .ZN(
        n12817) );
  NAND2_X1 U15244 ( .A1(n12812), .A2(n12808), .ZN(n12811) );
  OAI21_X1 U15245 ( .B1(n11671), .B2(n12809), .A(n12813), .ZN(n12810) );
  MUX2_X1 U15246 ( .A(n12811), .B(n12810), .S(n9602), .Z(n12816) );
  MUX2_X1 U15247 ( .A(n12813), .B(n12812), .S(n9602), .Z(n12814) );
  OAI211_X1 U15248 ( .C1(n12817), .C2(n12816), .A(n12815), .B(n12814), .ZN(
        n12822) );
  MUX2_X1 U15249 ( .A(n12819), .B(n12818), .S(n9602), .Z(n12820) );
  NAND3_X1 U15250 ( .A1(n12822), .A2(n12821), .A3(n12820), .ZN(n12823) );
  OAI21_X1 U15251 ( .B1(n12824), .B2(n12926), .A(n12823), .ZN(n12828) );
  AOI21_X1 U15252 ( .B1(n12827), .B2(n12825), .A(n9602), .ZN(n12826) );
  OAI21_X1 U15253 ( .B1(n12830), .B2(n9602), .A(n12829), .ZN(n12836) );
  INV_X1 U15254 ( .A(n15935), .ZN(n12831) );
  NAND2_X1 U15255 ( .A1(n13147), .A2(n12831), .ZN(n12833) );
  MUX2_X1 U15256 ( .A(n12833), .B(n12832), .S(n9602), .Z(n12834) );
  OAI211_X1 U15257 ( .C1(n12837), .C2(n12836), .A(n12835), .B(n12834), .ZN(
        n12840) );
  NAND3_X1 U15258 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(n12849) );
  INV_X1 U15259 ( .A(n12849), .ZN(n12842) );
  NAND2_X1 U15260 ( .A1(n12842), .A2(n12841), .ZN(n12844) );
  OAI211_X1 U15261 ( .C1(n12845), .C2(n12850), .A(n12844), .B(n12843), .ZN(
        n12853) );
  INV_X1 U15262 ( .A(n12846), .ZN(n12848) );
  OAI222_X1 U15263 ( .A1(n12851), .A2(n12850), .B1(n12849), .B2(n12848), .C1(
        n13087), .C2(n12847), .ZN(n12852) );
  NOR2_X1 U15264 ( .A1(n12855), .A2(n12854), .ZN(n12864) );
  NAND2_X1 U15265 ( .A1(n12860), .A2(n12856), .ZN(n12859) );
  NAND2_X1 U15266 ( .A1(n12861), .A2(n12857), .ZN(n12858) );
  MUX2_X1 U15267 ( .A(n12859), .B(n12858), .S(n9602), .Z(n12863) );
  MUX2_X1 U15268 ( .A(n12861), .B(n12860), .S(n9602), .Z(n12862) );
  OAI211_X1 U15269 ( .C1(n12864), .C2(n12863), .A(n9569), .B(n12862), .ZN(
        n12869) );
  MUX2_X1 U15270 ( .A(n12866), .B(n12865), .S(n9602), .Z(n12867) );
  NAND3_X1 U15271 ( .A1(n12869), .A2(n12868), .A3(n12867), .ZN(n12872) );
  MUX2_X1 U15272 ( .A(n12870), .B(n13531), .S(n9602), .Z(n12871) );
  NAND2_X1 U15273 ( .A1(n12876), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U15274 ( .A1(n12877), .A2(n13533), .ZN(n12874) );
  MUX2_X1 U15275 ( .A(n12875), .B(n12874), .S(n9602), .Z(n12879) );
  MUX2_X1 U15276 ( .A(n12877), .B(n12876), .S(n9602), .Z(n12878) );
  OAI211_X1 U15277 ( .C1(n12881), .C2(n13489), .A(n12880), .B(n12885), .ZN(
        n12884) );
  INV_X1 U15278 ( .A(n12882), .ZN(n12883) );
  MUX2_X1 U15279 ( .A(n12884), .B(n12883), .S(n9602), .Z(n12888) );
  MUX2_X1 U15280 ( .A(n12886), .B(n12885), .S(n9602), .Z(n12887) );
  NAND2_X1 U15281 ( .A1(n13628), .A2(n13482), .ZN(n12890) );
  MUX2_X1 U15282 ( .A(n12890), .B(n12889), .S(n9602), .Z(n12891) );
  NAND3_X1 U15283 ( .A1(n12892), .A2(n13456), .A3(n12891), .ZN(n12894) );
  INV_X1 U15284 ( .A(n13442), .ZN(n13444) );
  MUX2_X1 U15285 ( .A(n13440), .B(n13439), .S(n9602), .Z(n12893) );
  NAND3_X1 U15286 ( .A1(n12894), .A2(n13444), .A3(n12893), .ZN(n12898) );
  MUX2_X1 U15287 ( .A(n12896), .B(n12895), .S(n9602), .Z(n12897) );
  NAND4_X1 U15288 ( .A1(n13407), .A2(n13447), .A3(n9602), .A4(n13614), .ZN(
        n12902) );
  AOI21_X1 U15289 ( .B1(n13404), .B2(n13383), .A(n12899), .ZN(n12900) );
  MUX2_X1 U15290 ( .A(n12900), .B(n13383), .S(n9602), .Z(n12901) );
  MUX2_X1 U15291 ( .A(n12905), .B(n12904), .S(n9602), .Z(n12906) );
  MUX2_X1 U15292 ( .A(n12908), .B(n12907), .S(n9602), .Z(n12909) );
  NAND2_X1 U15293 ( .A1(n13343), .A2(n12926), .ZN(n12910) );
  NAND2_X1 U15294 ( .A1(n12913), .A2(n13340), .ZN(n12924) );
  NAND2_X1 U15295 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  NAND2_X1 U15296 ( .A1(n12918), .A2(n12917), .ZN(n12919) );
  NAND2_X1 U15297 ( .A1(n12919), .A2(n9602), .ZN(n12922) );
  NAND3_X1 U15298 ( .A1(n12927), .A2(n12926), .A3(n12925), .ZN(n12934) );
  INV_X1 U15299 ( .A(n12929), .ZN(n12932) );
  INV_X1 U15300 ( .A(n12930), .ZN(n13137) );
  AOI21_X1 U15301 ( .B1(n12930), .B2(n12929), .A(n13664), .ZN(n12931) );
  AOI21_X1 U15302 ( .B1(n12932), .B2(n13137), .A(n12931), .ZN(n12933) );
  NAND2_X1 U15303 ( .A1(n12939), .A2(n12937), .ZN(n12938) );
  NAND3_X1 U15304 ( .A1(n12943), .A2(n12942), .A3(n13285), .ZN(n12944) );
  OAI211_X1 U15305 ( .C1(n12946), .C2(n12945), .A(n12944), .B(P3_B_REG_SCAN_IN), .ZN(n12947) );
  OAI211_X1 U15306 ( .C1(n12196), .C2(n12949), .A(n12948), .B(n13128), .ZN(
        n12957) );
  INV_X1 U15307 ( .A(n12950), .ZN(n12951) );
  AOI21_X1 U15308 ( .B1(n15870), .B2(n15935), .A(n12951), .ZN(n12956) );
  AOI22_X1 U15309 ( .A1(n13111), .A2(n13146), .B1(n13110), .B2(n12952), .ZN(
        n12955) );
  NAND2_X1 U15310 ( .A1(n13133), .A2(n12953), .ZN(n12954) );
  NAND4_X1 U15311 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        P3_U3153) );
  XOR2_X1 U15312 ( .A(n12959), .B(n12958), .Z(n12964) );
  AOI22_X1 U15313 ( .A1(n13361), .A2(n13133), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12961) );
  NAND2_X1 U15314 ( .A1(n13385), .A2(n13130), .ZN(n12960) );
  OAI211_X1 U15315 ( .C1(n13358), .C2(n15874), .A(n12961), .B(n12960), .ZN(
        n12962) );
  AOI21_X1 U15316 ( .B1(n13674), .B2(n15870), .A(n12962), .ZN(n12963) );
  OAI21_X1 U15317 ( .B1(n12964), .B2(n15867), .A(n12963), .ZN(P3_U3154) );
  XNOR2_X1 U15318 ( .A(n12966), .B(n12965), .ZN(n12972) );
  NAND2_X1 U15319 ( .A1(n13130), .A2(n13568), .ZN(n12967) );
  NAND2_X1 U15320 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13196)
         );
  OAI211_X1 U15321 ( .C1(n15874), .C2(n12968), .A(n12967), .B(n13196), .ZN(
        n12970) );
  NOR2_X1 U15322 ( .A1(n13707), .A2(n13136), .ZN(n12969) );
  AOI211_X1 U15323 ( .C1(n13571), .C2(n13133), .A(n12970), .B(n12969), .ZN(
        n12971) );
  OAI21_X1 U15324 ( .B1(n12972), .B2(n15867), .A(n12971), .ZN(P3_U3155) );
  AOI22_X1 U15325 ( .A1(n13427), .A2(n13110), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12974) );
  NAND2_X1 U15326 ( .A1(n13423), .A2(n13133), .ZN(n12973) );
  OAI211_X1 U15327 ( .C1(n12975), .C2(n15874), .A(n12974), .B(n12973), .ZN(
        n12976) );
  AOI21_X1 U15328 ( .B1(n13614), .B2(n15870), .A(n12976), .ZN(n12977) );
  OAI21_X1 U15329 ( .B1(n12978), .B2(n15867), .A(n12977), .ZN(P3_U3156) );
  AOI21_X1 U15330 ( .B1(n12980), .B2(n12979), .A(n15867), .ZN(n12982) );
  NAND2_X1 U15331 ( .A1(n12982), .A2(n12981), .ZN(n12989) );
  INV_X1 U15332 ( .A(n12983), .ZN(n12984) );
  AOI21_X1 U15333 ( .B1(n15870), .B2(n12985), .A(n12984), .ZN(n12988) );
  AOI22_X1 U15334 ( .A1(n13111), .A2(n13149), .B1(n13110), .B2(n11672), .ZN(
        n12987) );
  NAND2_X1 U15335 ( .A1(n13133), .A2(n9082), .ZN(n12986) );
  NAND4_X1 U15336 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        P3_U3158) );
  INV_X1 U15337 ( .A(n12990), .ZN(n13696) );
  OAI211_X1 U15338 ( .C1(n12993), .C2(n12992), .A(n12991), .B(n13128), .ZN(
        n12997) );
  NAND2_X1 U15339 ( .A1(n13130), .A2(n13141), .ZN(n12994) );
  NAND2_X1 U15340 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13315)
         );
  OAI211_X1 U15341 ( .C1(n13482), .C2(n15874), .A(n12994), .B(n13315), .ZN(
        n12995) );
  AOI21_X1 U15342 ( .B1(n13483), .B2(n13133), .A(n12995), .ZN(n12996) );
  OAI211_X1 U15343 ( .C1(n13696), .C2(n13136), .A(n12997), .B(n12996), .ZN(
        P3_U3159) );
  OAI211_X1 U15344 ( .C1(n13000), .C2(n12999), .A(n12998), .B(n13128), .ZN(
        n13008) );
  INV_X1 U15345 ( .A(n13001), .ZN(n13002) );
  AOI21_X1 U15346 ( .B1(n15870), .B2(n13003), .A(n13002), .ZN(n13007) );
  AOI22_X1 U15347 ( .A1(n13111), .A2(n13145), .B1(n13110), .B2(n13147), .ZN(
        n13006) );
  NAND2_X1 U15348 ( .A1(n13133), .A2(n13004), .ZN(n13005) );
  NAND4_X1 U15349 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        P3_U3161) );
  INV_X1 U15350 ( .A(n13009), .ZN(n13010) );
  AOI21_X1 U15351 ( .B1(n13012), .B2(n13011), .A(n13010), .ZN(n13018) );
  AOI22_X1 U15352 ( .A1(n13013), .A2(n13110), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13015) );
  NAND2_X1 U15353 ( .A1(n13460), .A2(n13133), .ZN(n13014) );
  OAI211_X1 U15354 ( .C1(n13458), .C2(n15874), .A(n13015), .B(n13014), .ZN(
        n13016) );
  AOI21_X1 U15355 ( .B1(n13459), .B2(n15870), .A(n13016), .ZN(n13017) );
  OAI21_X1 U15356 ( .B1(n13018), .B2(n15867), .A(n13017), .ZN(P3_U3163) );
  INV_X1 U15357 ( .A(n13019), .ZN(n13020) );
  XOR2_X1 U15358 ( .A(n13021), .B(n13019), .Z(n13084) );
  NOR2_X1 U15359 ( .A1(n13084), .A2(n13085), .ZN(n13083) );
  AOI21_X1 U15360 ( .B1(n13021), .B2(n13020), .A(n13083), .ZN(n13024) );
  XNOR2_X1 U15361 ( .A(n13022), .B(n13143), .ZN(n13023) );
  XNOR2_X1 U15362 ( .A(n13024), .B(n13023), .ZN(n13033) );
  NAND2_X1 U15363 ( .A1(n13130), .A2(n13144), .ZN(n13026) );
  OAI211_X1 U15364 ( .C1(n15874), .C2(n13027), .A(n13026), .B(n13025), .ZN(
        n13028) );
  AOI21_X1 U15365 ( .B1(n13029), .B2(n13133), .A(n13028), .ZN(n13032) );
  NAND2_X1 U15366 ( .A1(n13030), .A2(n15870), .ZN(n13031) );
  OAI211_X1 U15367 ( .C1(n13033), .C2(n15867), .A(n13032), .B(n13031), .ZN(
        P3_U3164) );
  XOR2_X1 U15368 ( .A(n13035), .B(n13034), .Z(n13040) );
  AOI22_X1 U15369 ( .A1(n13395), .A2(n13133), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13037) );
  NAND2_X1 U15370 ( .A1(n13428), .A2(n13130), .ZN(n13036) );
  OAI211_X1 U15371 ( .C1(n13357), .C2(n15874), .A(n13037), .B(n13036), .ZN(
        n13038) );
  AOI21_X1 U15372 ( .B1(n13399), .B2(n15870), .A(n13038), .ZN(n13039) );
  OAI21_X1 U15373 ( .B1(n13040), .B2(n15867), .A(n13039), .ZN(P3_U3165) );
  INV_X1 U15374 ( .A(n13541), .ZN(n13647) );
  AOI21_X1 U15375 ( .B1(n13042), .B2(n13041), .A(n15867), .ZN(n13044) );
  NAND2_X1 U15376 ( .A1(n13044), .A2(n13043), .ZN(n13049) );
  NAND2_X1 U15377 ( .A1(n13130), .A2(n13565), .ZN(n13045) );
  NAND2_X1 U15378 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13252)
         );
  OAI211_X1 U15379 ( .C1(n15874), .C2(n13046), .A(n13045), .B(n13252), .ZN(
        n13047) );
  AOI21_X1 U15380 ( .B1(n13537), .B2(n13133), .A(n13047), .ZN(n13048) );
  OAI211_X1 U15381 ( .C1(n13647), .C2(n13136), .A(n13049), .B(n13048), .ZN(
        P3_U3166) );
  XNOR2_X1 U15382 ( .A(n13051), .B(n13050), .ZN(n13056) );
  NAND2_X1 U15383 ( .A1(n13130), .A2(n13546), .ZN(n13052) );
  NAND2_X1 U15384 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13274)
         );
  OAI211_X1 U15385 ( .C1(n13512), .C2(n15874), .A(n13052), .B(n13274), .ZN(
        n13054) );
  NOR2_X1 U15386 ( .A1(n13643), .A2(n13136), .ZN(n13053) );
  AOI211_X1 U15387 ( .C1(n13519), .C2(n13133), .A(n13054), .B(n13053), .ZN(
        n13055) );
  OAI21_X1 U15388 ( .B1(n13056), .B2(n15867), .A(n13055), .ZN(P3_U3168) );
  OAI21_X1 U15389 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n13060) );
  NAND2_X1 U15390 ( .A1(n13060), .A2(n13128), .ZN(n13067) );
  AOI21_X1 U15391 ( .B1(n15870), .B2(n13062), .A(n13061), .ZN(n13066) );
  AOI22_X1 U15392 ( .A1(n13111), .A2(n13148), .B1(n13110), .B2(n13150), .ZN(
        n13065) );
  NAND2_X1 U15393 ( .A1(n13133), .A2(n13063), .ZN(n13064) );
  NAND4_X1 U15394 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        P3_U3170) );
  INV_X1 U15395 ( .A(n13628), .ZN(n13075) );
  OAI211_X1 U15396 ( .C1(n13070), .C2(n13069), .A(n13068), .B(n13128), .ZN(
        n13074) );
  AOI22_X1 U15397 ( .A1(n13499), .A2(n13110), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13071) );
  OAI21_X1 U15398 ( .B1(n13474), .B2(n15874), .A(n13071), .ZN(n13072) );
  AOI21_X1 U15399 ( .B1(n13466), .B2(n13133), .A(n13072), .ZN(n13073) );
  OAI211_X1 U15400 ( .C1(n13075), .C2(n13136), .A(n13074), .B(n13073), .ZN(
        P3_U3173) );
  XNOR2_X1 U15401 ( .A(n13076), .B(n13427), .ZN(n13082) );
  AOI22_X1 U15402 ( .A1(n13140), .A2(n13110), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13078) );
  NAND2_X1 U15403 ( .A1(n13448), .A2(n13133), .ZN(n13077) );
  OAI211_X1 U15404 ( .C1(n13447), .C2(n15874), .A(n13078), .B(n13077), .ZN(
        n13079) );
  AOI21_X1 U15405 ( .B1(n13080), .B2(n15870), .A(n13079), .ZN(n13081) );
  OAI21_X1 U15406 ( .B1(n13082), .B2(n15867), .A(n13081), .ZN(P3_U3175) );
  AOI211_X1 U15407 ( .C1(n13085), .C2(n13084), .A(n15867), .B(n13083), .ZN(
        n13086) );
  INV_X1 U15408 ( .A(n13086), .ZN(n13094) );
  NAND2_X1 U15409 ( .A1(n13130), .A2(n13087), .ZN(n13089) );
  OAI211_X1 U15410 ( .C1(n15874), .C2(n13090), .A(n13089), .B(n13088), .ZN(
        n13091) );
  AOI21_X1 U15411 ( .B1(n13092), .B2(n13133), .A(n13091), .ZN(n13093) );
  OAI211_X1 U15412 ( .C1(n13136), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        P3_U3176) );
  XNOR2_X1 U15413 ( .A(n13096), .B(n13512), .ZN(n13097) );
  XNOR2_X1 U15414 ( .A(n13098), .B(n13097), .ZN(n13103) );
  NAND2_X1 U15415 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13301)
         );
  NAND2_X1 U15416 ( .A1(n13130), .A2(n13527), .ZN(n13099) );
  OAI211_X1 U15417 ( .C1(n13473), .C2(n15874), .A(n13301), .B(n13099), .ZN(
        n13100) );
  AOI21_X1 U15418 ( .B1(n13502), .B2(n13133), .A(n13100), .ZN(n13102) );
  NAND2_X1 U15419 ( .A1(n13492), .A2(n15870), .ZN(n13101) );
  OAI211_X1 U15420 ( .C1(n13103), .C2(n15867), .A(n13102), .B(n13101), .ZN(
        P3_U3178) );
  AOI21_X1 U15421 ( .B1(n13104), .B2(n13105), .A(n15867), .ZN(n13107) );
  NAND2_X1 U15422 ( .A1(n13107), .A2(n13106), .ZN(n13116) );
  AOI21_X1 U15423 ( .B1(n15870), .B2(n13109), .A(n13108), .ZN(n13115) );
  AOI22_X1 U15424 ( .A1(n13111), .A2(n13147), .B1(n13110), .B2(n13148), .ZN(
        n13114) );
  NAND2_X1 U15425 ( .A1(n13133), .A2(n13112), .ZN(n13113) );
  NAND4_X1 U15426 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        P3_U3179) );
  XOR2_X1 U15427 ( .A(n13118), .B(n13117), .Z(n13124) );
  AOI22_X1 U15428 ( .A1(n13375), .A2(n13133), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13121) );
  NAND2_X1 U15429 ( .A1(n13119), .A2(n13130), .ZN(n13120) );
  OAI211_X1 U15430 ( .C1(n13370), .C2(n15874), .A(n13121), .B(n13120), .ZN(
        n13122) );
  AOI21_X1 U15431 ( .B1(n9594), .B2(n15870), .A(n13122), .ZN(n13123) );
  OAI21_X1 U15432 ( .B1(n13124), .B2(n15867), .A(n13123), .ZN(P3_U3180) );
  OAI21_X1 U15433 ( .B1(n13127), .B2(n13126), .A(n13125), .ZN(n13129) );
  NAND2_X1 U15434 ( .A1(n13129), .A2(n13128), .ZN(n13135) );
  NAND2_X1 U15435 ( .A1(n13130), .A2(n13545), .ZN(n13131) );
  NAND2_X1 U15436 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13229)
         );
  OAI211_X1 U15437 ( .C1(n15874), .C2(n13510), .A(n13131), .B(n13229), .ZN(
        n13132) );
  AOI21_X1 U15438 ( .B1(n13552), .B2(n13133), .A(n13132), .ZN(n13134) );
  OAI211_X1 U15439 ( .C1(n13136), .C2(n13651), .A(n13135), .B(n13134), .ZN(
        P3_U3181) );
  MUX2_X1 U15440 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13137), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15441 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13138), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15442 ( .A(n13343), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13142), .Z(
        P3_U3518) );
  MUX2_X1 U15443 ( .A(n13385), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13142), .Z(
        P3_U3517) );
  MUX2_X1 U15444 ( .A(n13428), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13142), .Z(
        P3_U3515) );
  MUX2_X1 U15445 ( .A(n13139), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13142), .Z(
        P3_U3514) );
  MUX2_X1 U15446 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13427), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15447 ( .A(n13140), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13142), .Z(
        P3_U3512) );
  MUX2_X1 U15448 ( .A(n13499), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13142), .Z(
        P3_U3510) );
  MUX2_X1 U15449 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13141), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15450 ( .A(n13527), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13142), .Z(
        P3_U3508) );
  MUX2_X1 U15451 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13546), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15452 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13565), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15453 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13545), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15454 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13143), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15455 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13144), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15456 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13145), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15457 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13146), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15458 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13147), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15459 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13148), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15460 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13149), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15461 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13150), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15462 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n11672), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15463 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15866), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15464 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n11047), .S(P3_U3897), .Z(
        P3_U3491) );
  MUX2_X1 U15465 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13285), .Z(n13151) );
  AOI22_X1 U15466 ( .A1(n15888), .A2(P3_REG2_REG_0__SCAN_IN), .B1(n13154), 
        .B2(n13151), .ZN(n13153) );
  MUX2_X1 U15467 ( .A(n13317), .B(n13153), .S(n13152), .Z(n13161) );
  AOI22_X1 U15468 ( .A1(n15865), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n13160) );
  OR3_X1 U15469 ( .A1(n15888), .A2(n15895), .A3(n13154), .ZN(n13156) );
  NAND2_X1 U15470 ( .A1(n13156), .A2(n13155), .ZN(n13159) );
  NAND2_X1 U15471 ( .A1(n15895), .A2(n13157), .ZN(n13158) );
  NAND4_X1 U15472 ( .A1(n13161), .A2(n13160), .A3(n13159), .A4(n13158), .ZN(
        P3_U3182) );
  XNOR2_X1 U15473 ( .A(n13183), .B(n13185), .ZN(n13186) );
  XNOR2_X1 U15474 ( .A(n13186), .B(n13164), .ZN(n13182) );
  INV_X1 U15475 ( .A(n13185), .ZN(n13199) );
  OAI21_X1 U15476 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13166), .A(n13193), 
        .ZN(n13180) );
  NAND2_X1 U15477 ( .A1(n13168), .A2(n13167), .ZN(n13170) );
  MUX2_X1 U15478 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13285), .Z(n13198) );
  XNOR2_X1 U15479 ( .A(n13198), .B(n13199), .ZN(n13171) );
  AOI21_X1 U15480 ( .B1(n13173), .B2(n13170), .A(n13171), .ZN(n13169) );
  INV_X1 U15481 ( .A(n13169), .ZN(n13174) );
  AND2_X1 U15482 ( .A1(n13171), .A2(n13170), .ZN(n13172) );
  AOI21_X1 U15483 ( .B1(n13174), .B2(n13204), .A(n15892), .ZN(n13179) );
  NAND2_X1 U15484 ( .A1(n15886), .A2(n13199), .ZN(n13176) );
  OAI211_X1 U15485 ( .C1(n13177), .C2(n15898), .A(n13176), .B(n13175), .ZN(
        n13178) );
  AOI211_X1 U15486 ( .C1(n13180), .C2(n15888), .A(n13179), .B(n13178), .ZN(
        n13181) );
  OAI21_X1 U15487 ( .B1(n13182), .B2(n13237), .A(n13181), .ZN(P3_U3195) );
  INV_X1 U15488 ( .A(n13183), .ZN(n13184) );
  AOI22_X1 U15489 ( .A1(n13186), .A2(P3_REG1_REG_13__SCAN_IN), .B1(n13185), 
        .B2(n13184), .ZN(n13215) );
  NAND2_X1 U15490 ( .A1(n13195), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13223) );
  OR2_X1 U15491 ( .A1(n13195), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13187) );
  AND2_X1 U15492 ( .A1(n13223), .A2(n13187), .ZN(n13213) );
  XNOR2_X1 U15493 ( .A(n13215), .B(n13213), .ZN(n13212) );
  INV_X1 U15494 ( .A(n13193), .ZN(n13189) );
  NAND2_X1 U15495 ( .A1(n13195), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13222) );
  OR2_X1 U15496 ( .A1(n13195), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U15497 ( .A1(n13222), .A2(n13188), .ZN(n13191) );
  INV_X1 U15498 ( .A(n13191), .ZN(n13201) );
  NOR3_X1 U15499 ( .A1(n13189), .A2(n13190), .A3(n13201), .ZN(n13194) );
  INV_X1 U15500 ( .A(n13190), .ZN(n13192) );
  AOI21_X1 U15501 ( .B1(n13193), .B2(n13192), .A(n13191), .ZN(n13217) );
  OAI21_X1 U15502 ( .B1(n13194), .B2(n13217), .A(n15888), .ZN(n13211) );
  INV_X1 U15503 ( .A(n13195), .ZN(n13209) );
  INV_X1 U15504 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13197) );
  OAI21_X1 U15505 ( .B1(n15898), .B2(n13197), .A(n13196), .ZN(n13208) );
  INV_X1 U15506 ( .A(n13198), .ZN(n13200) );
  NAND2_X1 U15507 ( .A1(n13200), .A2(n13199), .ZN(n13203) );
  MUX2_X1 U15508 ( .A(n13213), .B(n13201), .S(n6821), .Z(n13202) );
  INV_X1 U15509 ( .A(n13225), .ZN(n13206) );
  AOI21_X1 U15510 ( .B1(n13204), .B2(n13203), .A(n13202), .ZN(n13205) );
  NOR3_X1 U15511 ( .A1(n13206), .A2(n13205), .A3(n15892), .ZN(n13207) );
  AOI211_X1 U15512 ( .C1(n15886), .C2(n13209), .A(n13208), .B(n13207), .ZN(
        n13210) );
  OAI211_X1 U15513 ( .C1(n13212), .C2(n13237), .A(n13211), .B(n13210), .ZN(
        P3_U3196) );
  INV_X1 U15514 ( .A(n13213), .ZN(n13214) );
  XNOR2_X1 U15515 ( .A(n13239), .B(n13226), .ZN(n13242) );
  XNOR2_X1 U15516 ( .A(n13242), .B(P3_REG1_REG_15__SCAN_IN), .ZN(n13238) );
  INV_X1 U15517 ( .A(n13222), .ZN(n13216) );
  INV_X1 U15518 ( .A(n13219), .ZN(n13218) );
  INV_X1 U15519 ( .A(n13226), .ZN(n13247) );
  NAND2_X1 U15520 ( .A1(n13219), .A2(n13247), .ZN(n13220) );
  OAI21_X1 U15521 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n13221), .A(n13260), 
        .ZN(n13235) );
  MUX2_X1 U15522 ( .A(n13223), .B(n13222), .S(n6821), .Z(n13224) );
  NAND2_X1 U15523 ( .A1(n13225), .A2(n13224), .ZN(n13245) );
  XNOR2_X1 U15524 ( .A(n13245), .B(n13226), .ZN(n13228) );
  MUX2_X1 U15525 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13285), .Z(n13227) );
  AOI21_X1 U15526 ( .B1(n13228), .B2(n13227), .A(n13246), .ZN(n13233) );
  OAI21_X1 U15527 ( .B1(n15898), .B2(n13230), .A(n13229), .ZN(n13231) );
  AOI21_X1 U15528 ( .B1(n15886), .B2(n13247), .A(n13231), .ZN(n13232) );
  OAI21_X1 U15529 ( .B1(n13233), .B2(n15892), .A(n13232), .ZN(n13234) );
  AOI21_X1 U15530 ( .B1(n13235), .B2(n15888), .A(n13234), .ZN(n13236) );
  OAI21_X1 U15531 ( .B1(n13238), .B2(n13237), .A(n13236), .ZN(P3_U3197) );
  INV_X1 U15532 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13241) );
  INV_X1 U15533 ( .A(n13239), .ZN(n13240) );
  XNOR2_X1 U15534 ( .A(n13272), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U15535 ( .A1(n13243), .A2(n13244), .ZN(n13270) );
  OAI21_X1 U15536 ( .B1(n13244), .B2(n13243), .A(n13270), .ZN(n13264) );
  INV_X1 U15537 ( .A(n13245), .ZN(n13248) );
  INV_X1 U15538 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13271) );
  MUX2_X1 U15539 ( .A(n13539), .B(n13271), .S(n13285), .Z(n13249) );
  NOR2_X1 U15540 ( .A1(n13272), .A2(n13249), .ZN(n13276) );
  NAND2_X1 U15541 ( .A1(n13272), .A2(n13249), .ZN(n13275) );
  INV_X1 U15542 ( .A(n13275), .ZN(n13250) );
  NOR2_X1 U15543 ( .A1(n13276), .A2(n13250), .ZN(n13251) );
  XNOR2_X1 U15544 ( .A(n13277), .B(n13251), .ZN(n13256) );
  OAI21_X1 U15545 ( .B1(n15898), .B2(n13253), .A(n13252), .ZN(n13254) );
  AOI21_X1 U15546 ( .B1(n15886), .B2(n13272), .A(n13254), .ZN(n13255) );
  OAI21_X1 U15547 ( .B1(n13256), .B2(n15892), .A(n13255), .ZN(n13263) );
  XNOR2_X1 U15548 ( .A(n13272), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13257) );
  INV_X1 U15549 ( .A(n13257), .ZN(n13259) );
  NAND3_X1 U15550 ( .A1(n13260), .A2(n13259), .A3(n13258), .ZN(n13261) );
  AOI21_X1 U15551 ( .B1(n13266), .B2(n13261), .A(n13329), .ZN(n13262) );
  AOI211_X1 U15552 ( .C1(n15895), .C2(n13264), .A(n13263), .B(n13262), .ZN(
        n13265) );
  INV_X1 U15553 ( .A(n13265), .ZN(P3_U3198) );
  INV_X1 U15554 ( .A(n13292), .ZN(n13268) );
  AOI21_X1 U15555 ( .B1(n13521), .B2(n13269), .A(n13268), .ZN(n13284) );
  XOR2_X1 U15556 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13299), .Z(n13282) );
  NAND2_X1 U15557 ( .A1(n15865), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13273) );
  OAI211_X1 U15558 ( .C1(n13317), .C2(n13294), .A(n13274), .B(n13273), .ZN(
        n13281) );
  MUX2_X1 U15559 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13285), .Z(n13287) );
  XNOR2_X1 U15560 ( .A(n13287), .B(n13294), .ZN(n13279) );
  AOI211_X1 U15561 ( .C1(n13279), .C2(n13278), .A(n15892), .B(n13286), .ZN(
        n13280) );
  AOI211_X1 U15562 ( .C1(n15895), .C2(n13282), .A(n13281), .B(n13280), .ZN(
        n13283) );
  OAI21_X1 U15563 ( .B1(n13284), .B2(n13329), .A(n13283), .ZN(P3_U3199) );
  MUX2_X1 U15564 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13285), .Z(n13289) );
  XNOR2_X1 U15565 ( .A(n13324), .B(n13323), .ZN(n13288) );
  NOR2_X1 U15566 ( .A1(n13288), .A2(n13289), .ZN(n13322) );
  AOI21_X1 U15567 ( .B1(n13289), .B2(n13288), .A(n13322), .ZN(n13306) );
  NAND2_X1 U15568 ( .A1(n13311), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13307) );
  OAI21_X1 U15569 ( .B1(n13311), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13307), 
        .ZN(n13290) );
  AND3_X1 U15570 ( .A1(n13292), .A2(n13291), .A3(n13290), .ZN(n13293) );
  OAI21_X1 U15571 ( .B1(n13308), .B2(n13293), .A(n15888), .ZN(n13305) );
  INV_X1 U15572 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13298) );
  INV_X1 U15573 ( .A(n13294), .ZN(n13297) );
  XNOR2_X1 U15574 ( .A(n13323), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13312) );
  XNOR2_X1 U15575 ( .A(n13313), .B(n13312), .ZN(n13303) );
  NAND2_X1 U15576 ( .A1(n15865), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13300) );
  OAI211_X1 U15577 ( .C1(n13317), .C2(n13311), .A(n13301), .B(n13300), .ZN(
        n13302) );
  AOI21_X1 U15578 ( .B1(n15895), .B2(n13303), .A(n13302), .ZN(n13304) );
  OAI211_X1 U15579 ( .C1(n13306), .C2(n15892), .A(n13305), .B(n13304), .ZN(
        P3_U3200) );
  XNOR2_X1 U15580 ( .A(n13316), .B(n13309), .ZN(n13318) );
  XNOR2_X1 U15581 ( .A(n13310), .B(n13318), .ZN(n13330) );
  XNOR2_X1 U15582 ( .A(n13316), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U15583 ( .A1(n15865), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13314) );
  OAI211_X1 U15584 ( .C1(n13317), .C2(n13316), .A(n13315), .B(n13314), .ZN(
        n13326) );
  INV_X1 U15585 ( .A(n13318), .ZN(n13320) );
  MUX2_X1 U15586 ( .A(n13321), .B(n13320), .S(n6821), .Z(n13325) );
  OAI21_X1 U15587 ( .B1(n13330), .B2(n13329), .A(n13328), .ZN(P3_U3201) );
  NOR2_X1 U15588 ( .A1(n13333), .A2(n13332), .ZN(n13661) );
  AOI21_X1 U15589 ( .B1(n13661), .B2(n13574), .A(n13334), .ZN(n13337) );
  NAND2_X1 U15590 ( .A1(n13580), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13335) );
  OAI211_X1 U15591 ( .C1(n13663), .C2(n13582), .A(n13337), .B(n13335), .ZN(
        P3_U3202) );
  INV_X1 U15592 ( .A(n13664), .ZN(n13593) );
  NAND2_X1 U15593 ( .A1(n13580), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13336) );
  OAI211_X1 U15594 ( .C1(n13593), .C2(n13582), .A(n13337), .B(n13336), .ZN(
        P3_U3203) );
  XNOR2_X1 U15595 ( .A(n13339), .B(n13338), .ZN(n13594) );
  INV_X1 U15596 ( .A(n13594), .ZN(n13353) );
  NAND2_X1 U15597 ( .A1(n13341), .A2(n13340), .ZN(n13342) );
  NAND2_X1 U15598 ( .A1(n13343), .A2(n13567), .ZN(n13344) );
  OAI21_X1 U15599 ( .B1(n13345), .B2(n13511), .A(n13344), .ZN(n13346) );
  INV_X1 U15600 ( .A(n13346), .ZN(n13347) );
  INV_X1 U15601 ( .A(n9525), .ZN(n13671) );
  AOI22_X1 U15602 ( .A1(n13349), .A2(n13579), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n13580), .ZN(n13350) );
  OAI21_X1 U15603 ( .B1(n13671), .B2(n13582), .A(n13350), .ZN(n13351) );
  AOI21_X1 U15604 ( .B1(n13595), .B2(n13574), .A(n13351), .ZN(n13352) );
  OAI21_X1 U15605 ( .B1(n13353), .B2(n13588), .A(n13352), .ZN(P3_U3205) );
  NAND2_X1 U15606 ( .A1(n13354), .A2(n13365), .ZN(n13355) );
  NAND2_X1 U15607 ( .A1(n13356), .A2(n13355), .ZN(n13360) );
  OAI22_X1 U15608 ( .A1(n13358), .A2(n13511), .B1(n13357), .B2(n13509), .ZN(
        n13359) );
  INV_X1 U15609 ( .A(n13361), .ZN(n13363) );
  INV_X1 U15610 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13362) );
  OAI22_X1 U15611 ( .A1(n13363), .A2(n13553), .B1(n13362), .B2(n13574), .ZN(
        n13364) );
  AOI21_X1 U15612 ( .B1(n13674), .B2(n13557), .A(n13364), .ZN(n13368) );
  XNOR2_X1 U15613 ( .A(n13366), .B(n13365), .ZN(n13597) );
  NAND2_X1 U15614 ( .A1(n13597), .A2(n13551), .ZN(n13367) );
  OAI211_X1 U15615 ( .C1(n13599), .C2(n13580), .A(n13368), .B(n13367), .ZN(
        P3_U3206) );
  XNOR2_X1 U15616 ( .A(n13369), .B(n13372), .ZN(n13374) );
  OAI22_X1 U15617 ( .A1(n13370), .A2(n13511), .B1(n13410), .B2(n13509), .ZN(
        n13373) );
  INV_X1 U15618 ( .A(n13605), .ZN(n13378) );
  AOI22_X1 U15619 ( .A1(n13375), .A2(n13579), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n13580), .ZN(n13376) );
  OAI21_X1 U15620 ( .B1(n7093), .B2(n13582), .A(n13376), .ZN(n13377) );
  AOI21_X1 U15621 ( .B1(n13378), .B2(n13418), .A(n13377), .ZN(n13379) );
  OAI21_X1 U15622 ( .B1(n13604), .B2(n13580), .A(n13379), .ZN(P3_U3207) );
  NAND2_X1 U15623 ( .A1(n13380), .A2(n13420), .ZN(n13402) );
  NAND2_X1 U15624 ( .A1(n13402), .A2(n13382), .ZN(n13405) );
  NAND2_X1 U15625 ( .A1(n13405), .A2(n13383), .ZN(n13384) );
  XNOR2_X1 U15626 ( .A(n13384), .B(n13391), .ZN(n13607) );
  AOI22_X1 U15627 ( .A1(n13385), .A2(n13566), .B1(n13567), .B2(n13428), .ZN(
        n13394) );
  AND2_X1 U15628 ( .A1(n13409), .A2(n13387), .ZN(n13392) );
  INV_X1 U15629 ( .A(n13388), .ZN(n13389) );
  NAND2_X1 U15630 ( .A1(n13409), .A2(n13389), .ZN(n13390) );
  OAI211_X1 U15631 ( .C1(n13392), .C2(n13391), .A(n13390), .B(n13562), .ZN(
        n13393) );
  NAND2_X1 U15632 ( .A1(n13609), .A2(n13585), .ZN(n13401) );
  INV_X1 U15633 ( .A(n13395), .ZN(n13397) );
  OAI22_X1 U15634 ( .A1(n13397), .A2(n13553), .B1(n13396), .B2(n13574), .ZN(
        n13398) );
  AOI21_X1 U15635 ( .B1(n13399), .B2(n13557), .A(n13398), .ZN(n13400) );
  OAI211_X1 U15636 ( .C1(n13436), .C2(n13607), .A(n13401), .B(n13400), .ZN(
        P3_U3208) );
  OAI21_X1 U15637 ( .B1(n13421), .B2(n13404), .A(n13403), .ZN(n13406) );
  NAND2_X1 U15638 ( .A1(n13406), .A2(n13405), .ZN(n13611) );
  NAND2_X1 U15639 ( .A1(n13386), .A2(n13407), .ZN(n13408) );
  AOI21_X1 U15640 ( .B1(n13409), .B2(n13408), .A(n13507), .ZN(n13412) );
  OAI22_X1 U15641 ( .A1(n13410), .A2(n13511), .B1(n13447), .B2(n13509), .ZN(
        n13411) );
  AOI211_X1 U15642 ( .C1(n13611), .C2(n13413), .A(n13412), .B(n13411), .ZN(
        n13613) );
  INV_X1 U15643 ( .A(n13610), .ZN(n13416) );
  AOI22_X1 U15644 ( .A1(n13414), .A2(n13579), .B1(n13580), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13415) );
  OAI21_X1 U15645 ( .B1(n13416), .B2(n13582), .A(n13415), .ZN(n13417) );
  AOI21_X1 U15646 ( .B1(n13611), .B2(n13418), .A(n13417), .ZN(n13419) );
  OAI21_X1 U15647 ( .B1(n13613), .B2(n13580), .A(n13419), .ZN(P3_U3209) );
  INV_X1 U15648 ( .A(n13380), .ZN(n13422) );
  INV_X1 U15649 ( .A(n13420), .ZN(n13430) );
  INV_X1 U15650 ( .A(n13616), .ZN(n13437) );
  INV_X1 U15651 ( .A(n13423), .ZN(n13425) );
  OAI22_X1 U15652 ( .A1(n13425), .A2(n13553), .B1(n13585), .B2(n13424), .ZN(
        n13426) );
  AOI21_X1 U15653 ( .B1(n13614), .B2(n13557), .A(n13426), .ZN(n13435) );
  AOI22_X1 U15654 ( .A1(n13428), .A2(n13566), .B1(n13567), .B2(n13427), .ZN(
        n13432) );
  OAI211_X1 U15655 ( .C1(n6704), .C2(n13430), .A(n13562), .B(n13429), .ZN(
        n13431) );
  OAI211_X1 U15656 ( .C1(n13437), .C2(n13433), .A(n13432), .B(n13431), .ZN(
        n13615) );
  NAND2_X1 U15657 ( .A1(n13615), .A2(n13585), .ZN(n13434) );
  OAI211_X1 U15658 ( .C1(n13437), .C2(n13436), .A(n13435), .B(n13434), .ZN(
        P3_U3210) );
  NAND2_X1 U15659 ( .A1(n13438), .A2(n13439), .ZN(n13441) );
  NAND2_X1 U15660 ( .A1(n13441), .A2(n13440), .ZN(n13443) );
  XNOR2_X1 U15661 ( .A(n13443), .B(n13442), .ZN(n13620) );
  INV_X1 U15662 ( .A(n13620), .ZN(n13452) );
  XNOR2_X1 U15663 ( .A(n13445), .B(n13444), .ZN(n13446) );
  OAI222_X1 U15664 ( .A1(n13511), .A2(n13447), .B1(n13509), .B2(n13474), .C1(
        n13507), .C2(n13446), .ZN(n13619) );
  AOI22_X1 U15665 ( .A1(n13448), .A2(n13579), .B1(n13580), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U15666 ( .B1(n13687), .B2(n13582), .A(n13449), .ZN(n13450) );
  AOI21_X1 U15667 ( .B1(n13619), .B2(n13574), .A(n13450), .ZN(n13451) );
  OAI21_X1 U15668 ( .B1(n13452), .B2(n13588), .A(n13451), .ZN(P3_U3211) );
  XOR2_X1 U15669 ( .A(n13438), .B(n13456), .Z(n13624) );
  INV_X1 U15670 ( .A(n13624), .ZN(n13464) );
  INV_X1 U15671 ( .A(n13453), .ZN(n13454) );
  AOI21_X1 U15672 ( .B1(n13456), .B2(n13455), .A(n13454), .ZN(n13457) );
  OAI222_X1 U15673 ( .A1(n13511), .A2(n13458), .B1(n13509), .B2(n13482), .C1(
        n13507), .C2(n13457), .ZN(n13623) );
  INV_X1 U15674 ( .A(n13459), .ZN(n13691) );
  AOI22_X1 U15675 ( .A1(n13460), .A2(n13579), .B1(n13580), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n13461) );
  OAI21_X1 U15676 ( .B1(n13691), .B2(n13582), .A(n13461), .ZN(n13462) );
  AOI21_X1 U15677 ( .B1(n13623), .B2(n13574), .A(n13462), .ZN(n13463) );
  OAI21_X1 U15678 ( .B1(n13464), .B2(n13588), .A(n13463), .ZN(P3_U3212) );
  OAI21_X1 U15679 ( .B1(n6676), .B2(n7248), .A(n13465), .ZN(n13631) );
  INV_X1 U15680 ( .A(n13466), .ZN(n13468) );
  INV_X1 U15681 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13467) );
  OAI22_X1 U15682 ( .A1(n13468), .A2(n13553), .B1(n13585), .B2(n13467), .ZN(
        n13469) );
  AOI21_X1 U15683 ( .B1(n13628), .B2(n13557), .A(n13469), .ZN(n13476) );
  XNOR2_X1 U15684 ( .A(n13471), .B(n13470), .ZN(n13472) );
  OAI222_X1 U15685 ( .A1(n13511), .A2(n13474), .B1(n13509), .B2(n13473), .C1(
        n13507), .C2(n13472), .ZN(n13627) );
  NAND2_X1 U15686 ( .A1(n13627), .A2(n13585), .ZN(n13475) );
  OAI211_X1 U15687 ( .C1(n13631), .C2(n13588), .A(n13476), .B(n13475), .ZN(
        P3_U3213) );
  NAND2_X1 U15688 ( .A1(n6836), .A2(n13517), .ZN(n13516) );
  NAND3_X1 U15689 ( .A1(n13516), .A2(n13496), .A3(n13489), .ZN(n13488) );
  NAND2_X1 U15690 ( .A1(n13488), .A2(n13477), .ZN(n13478) );
  XOR2_X1 U15691 ( .A(n13480), .B(n13478), .Z(n13633) );
  INV_X1 U15692 ( .A(n13633), .ZN(n13487) );
  XOR2_X1 U15693 ( .A(n13480), .B(n13479), .Z(n13481) );
  OAI222_X1 U15694 ( .A1(n13511), .A2(n13482), .B1(n13509), .B2(n13512), .C1(
        n13481), .C2(n13507), .ZN(n13632) );
  AOI22_X1 U15695 ( .A1(n13580), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13579), 
        .B2(n13483), .ZN(n13484) );
  OAI21_X1 U15696 ( .B1(n13696), .B2(n13582), .A(n13484), .ZN(n13485) );
  AOI21_X1 U15697 ( .B1(n13632), .B2(n13574), .A(n13485), .ZN(n13486) );
  OAI21_X1 U15698 ( .B1(n13487), .B2(n13588), .A(n13486), .ZN(P3_U3214) );
  INV_X1 U15699 ( .A(n13488), .ZN(n13491) );
  AOI21_X1 U15700 ( .B1(n13516), .B2(n13489), .A(n13496), .ZN(n13490) );
  NOR2_X1 U15701 ( .A1(n13491), .A2(n13490), .ZN(n13637) );
  INV_X1 U15702 ( .A(n13492), .ZN(n13700) );
  INV_X1 U15703 ( .A(n13508), .ZN(n13494) );
  INV_X1 U15704 ( .A(n13517), .ZN(n13493) );
  NAND2_X1 U15705 ( .A1(n13494), .A2(n13493), .ZN(n13515) );
  NAND2_X1 U15706 ( .A1(n13515), .A2(n13495), .ZN(n13497) );
  XNOR2_X1 U15707 ( .A(n13497), .B(n13496), .ZN(n13498) );
  NAND2_X1 U15708 ( .A1(n13498), .A2(n13562), .ZN(n13501) );
  AOI22_X1 U15709 ( .A1(n13499), .A2(n13566), .B1(n13567), .B2(n13527), .ZN(
        n13500) );
  NAND2_X1 U15710 ( .A1(n13501), .A2(n13500), .ZN(n13636) );
  NAND2_X1 U15711 ( .A1(n13636), .A2(n13585), .ZN(n13504) );
  AOI22_X1 U15712 ( .A1(n13580), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13579), 
        .B2(n13502), .ZN(n13503) );
  OAI211_X1 U15713 ( .C1(n13700), .C2(n13582), .A(n13504), .B(n13503), .ZN(
        n13505) );
  AOI21_X1 U15714 ( .B1(n13637), .B2(n13551), .A(n13505), .ZN(n13506) );
  INV_X1 U15715 ( .A(n13506), .ZN(P3_U3215) );
  AOI21_X1 U15716 ( .B1(n13508), .B2(n13517), .A(n13507), .ZN(n13514) );
  OAI22_X1 U15717 ( .A1(n13512), .A2(n13511), .B1(n13510), .B2(n13509), .ZN(
        n13513) );
  AOI21_X1 U15718 ( .B1(n13515), .B2(n13514), .A(n13513), .ZN(n13641) );
  OAI21_X1 U15719 ( .B1(n6836), .B2(n13517), .A(n13516), .ZN(n13640) );
  NAND2_X1 U15720 ( .A1(n13640), .A2(n13551), .ZN(n13525) );
  INV_X1 U15721 ( .A(n13643), .ZN(n13523) );
  INV_X1 U15722 ( .A(n13519), .ZN(n13520) );
  OAI22_X1 U15723 ( .A1(n13574), .A2(n13521), .B1(n13520), .B2(n13553), .ZN(
        n13522) );
  AOI21_X1 U15724 ( .B1(n13523), .B2(n13557), .A(n13522), .ZN(n13524) );
  OAI211_X1 U15725 ( .C1(n13580), .C2(n13641), .A(n13525), .B(n13524), .ZN(
        P3_U3216) );
  XNOR2_X1 U15726 ( .A(n13526), .B(n13535), .ZN(n13528) );
  AOI222_X1 U15727 ( .A1(n13562), .A2(n13528), .B1(n13565), .B2(n13567), .C1(
        n13527), .C2(n13566), .ZN(n13645) );
  OR2_X1 U15728 ( .A1(n13529), .A2(n13530), .ZN(n13532) );
  NAND2_X1 U15729 ( .A1(n13532), .A2(n13531), .ZN(n13550) );
  NAND2_X1 U15730 ( .A1(n13550), .A2(n13549), .ZN(n13548) );
  NAND2_X1 U15731 ( .A1(n13548), .A2(n13533), .ZN(n13536) );
  OAI21_X1 U15732 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13644) );
  NAND2_X1 U15733 ( .A1(n13644), .A2(n13551), .ZN(n13543) );
  INV_X1 U15734 ( .A(n13537), .ZN(n13538) );
  OAI22_X1 U15735 ( .A1(n13585), .A2(n13539), .B1(n13538), .B2(n13553), .ZN(
        n13540) );
  AOI21_X1 U15736 ( .B1(n13541), .B2(n13557), .A(n13540), .ZN(n13542) );
  OAI211_X1 U15737 ( .C1(n13580), .C2(n13645), .A(n13543), .B(n13542), .ZN(
        P3_U3217) );
  XNOR2_X1 U15738 ( .A(n13544), .B(n13549), .ZN(n13547) );
  AOI222_X1 U15739 ( .A1(n13562), .A2(n13547), .B1(n13546), .B2(n13566), .C1(
        n13545), .C2(n13567), .ZN(n13649) );
  OAI21_X1 U15740 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n13648) );
  NAND2_X1 U15741 ( .A1(n13648), .A2(n13551), .ZN(n13560) );
  INV_X1 U15742 ( .A(n13651), .ZN(n13558) );
  INV_X1 U15743 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13555) );
  INV_X1 U15744 ( .A(n13552), .ZN(n13554) );
  OAI22_X1 U15745 ( .A1(n13585), .A2(n13555), .B1(n13554), .B2(n13553), .ZN(
        n13556) );
  AOI21_X1 U15746 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(n13559) );
  OAI211_X1 U15747 ( .C1(n13580), .C2(n13649), .A(n13560), .B(n13559), .ZN(
        P3_U3218) );
  XNOR2_X1 U15748 ( .A(n13529), .B(n13564), .ZN(n13653) );
  INV_X1 U15749 ( .A(n13653), .ZN(n13576) );
  OAI211_X1 U15750 ( .C1(n13561), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13570) );
  AOI22_X1 U15751 ( .A1(n13568), .A2(n13567), .B1(n13566), .B2(n13565), .ZN(
        n13569) );
  NAND2_X1 U15752 ( .A1(n13570), .A2(n13569), .ZN(n13652) );
  AOI22_X1 U15753 ( .A1(n13580), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13579), 
        .B2(n13571), .ZN(n13572) );
  OAI21_X1 U15754 ( .B1(n13707), .B2(n13582), .A(n13572), .ZN(n13573) );
  AOI21_X1 U15755 ( .B1(n13652), .B2(n13574), .A(n13573), .ZN(n13575) );
  OAI21_X1 U15756 ( .B1(n13576), .B2(n13588), .A(n13575), .ZN(P3_U3219) );
  INV_X1 U15757 ( .A(n13577), .ZN(n13589) );
  AOI22_X1 U15758 ( .A1(n13580), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n13579), 
        .B2(n13578), .ZN(n13581) );
  OAI21_X1 U15759 ( .B1(n13583), .B2(n13582), .A(n13581), .ZN(n13584) );
  AOI21_X1 U15760 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13587) );
  OAI21_X1 U15761 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(P3_U3220) );
  NAND2_X1 U15762 ( .A1(n15951), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U15763 ( .A1(n13661), .A2(n15954), .ZN(n13592) );
  OAI211_X1 U15764 ( .C1(n13663), .C2(n13660), .A(n13590), .B(n13592), .ZN(
        P3_U3490) );
  NAND2_X1 U15765 ( .A1(n15951), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13591) );
  OAI211_X1 U15766 ( .C1(n13593), .C2(n13660), .A(n13592), .B(n13591), .ZN(
        P3_U3489) );
  INV_X1 U15767 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U15768 ( .A1(n13597), .A2(n15905), .ZN(n13598) );
  NAND2_X1 U15769 ( .A1(n13599), .A2(n13598), .ZN(n13672) );
  MUX2_X1 U15770 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13672), .S(n15954), .Z(
        n13600) );
  AOI21_X1 U15771 ( .B1(n13601), .B2(n13674), .A(n13600), .ZN(n13602) );
  INV_X1 U15772 ( .A(n13602), .ZN(P3_U3486) );
  NAND2_X1 U15773 ( .A1(n9594), .A2(n15936), .ZN(n13603) );
  MUX2_X1 U15774 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13677), .S(n15954), .Z(
        P3_U3485) );
  OAI22_X1 U15775 ( .A1(n13607), .A2(n15930), .B1(n13606), .B2(n15928), .ZN(
        n13608) );
  MUX2_X1 U15776 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13678), .S(n15954), .Z(
        P3_U3484) );
  AOI22_X1 U15777 ( .A1(n13611), .A2(n15937), .B1(n15936), .B2(n13610), .ZN(
        n13612) );
  NAND2_X1 U15778 ( .A1(n13613), .A2(n13612), .ZN(n13679) );
  MUX2_X1 U15779 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13679), .S(n15954), .Z(
        P3_U3483) );
  INV_X1 U15780 ( .A(n13614), .ZN(n13683) );
  INV_X1 U15781 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13617) );
  AOI21_X1 U15782 ( .B1(n15937), .B2(n13616), .A(n13615), .ZN(n13680) );
  MUX2_X1 U15783 ( .A(n13617), .B(n13680), .S(n15954), .Z(n13618) );
  OAI21_X1 U15784 ( .B1(n13683), .B2(n13660), .A(n13618), .ZN(P3_U3482) );
  INV_X1 U15785 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13621) );
  AOI21_X1 U15786 ( .B1(n13620), .B2(n15905), .A(n13619), .ZN(n13684) );
  MUX2_X1 U15787 ( .A(n13621), .B(n13684), .S(n15954), .Z(n13622) );
  OAI21_X1 U15788 ( .B1(n13687), .B2(n13660), .A(n13622), .ZN(P3_U3481) );
  AOI21_X1 U15789 ( .B1(n15905), .B2(n13624), .A(n13623), .ZN(n13688) );
  MUX2_X1 U15790 ( .A(n13625), .B(n13688), .S(n15954), .Z(n13626) );
  OAI21_X1 U15791 ( .B1(n13691), .B2(n13660), .A(n13626), .ZN(P3_U3480) );
  AOI21_X1 U15792 ( .B1(n15936), .B2(n13628), .A(n13627), .ZN(n13629) );
  OAI21_X1 U15793 ( .B1(n13631), .B2(n13630), .A(n13629), .ZN(n13692) );
  MUX2_X1 U15794 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13692), .S(n15954), .Z(
        P3_U3479) );
  INV_X1 U15795 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13634) );
  AOI21_X1 U15796 ( .B1(n13633), .B2(n15905), .A(n13632), .ZN(n13693) );
  MUX2_X1 U15797 ( .A(n13634), .B(n13693), .S(n15954), .Z(n13635) );
  OAI21_X1 U15798 ( .B1(n13696), .B2(n13660), .A(n13635), .ZN(P3_U3478) );
  INV_X1 U15799 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13638) );
  AOI21_X1 U15800 ( .B1(n13637), .B2(n15905), .A(n13636), .ZN(n13697) );
  MUX2_X1 U15801 ( .A(n13638), .B(n13697), .S(n15954), .Z(n13639) );
  OAI21_X1 U15802 ( .B1(n13700), .B2(n13660), .A(n13639), .ZN(P3_U3477) );
  NAND2_X1 U15803 ( .A1(n13640), .A2(n15905), .ZN(n13642) );
  OAI211_X1 U15804 ( .C1(n13643), .C2(n15928), .A(n13642), .B(n13641), .ZN(
        n13701) );
  MUX2_X1 U15805 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13701), .S(n15954), .Z(
        P3_U3476) );
  NAND2_X1 U15806 ( .A1(n13644), .A2(n15905), .ZN(n13646) );
  OAI211_X1 U15807 ( .C1(n13647), .C2(n15928), .A(n13646), .B(n13645), .ZN(
        n13702) );
  MUX2_X1 U15808 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13702), .S(n15954), .Z(
        P3_U3475) );
  NAND2_X1 U15809 ( .A1(n13648), .A2(n15905), .ZN(n13650) );
  OAI211_X1 U15810 ( .C1(n13651), .C2(n15928), .A(n13650), .B(n13649), .ZN(
        n13703) );
  MUX2_X1 U15811 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13703), .S(n15954), .Z(
        P3_U3474) );
  INV_X1 U15812 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13654) );
  AOI21_X1 U15813 ( .B1(n13653), .B2(n15905), .A(n13652), .ZN(n13704) );
  MUX2_X1 U15814 ( .A(n13654), .B(n13704), .S(n15954), .Z(n13655) );
  OAI21_X1 U15815 ( .B1(n13660), .B2(n13707), .A(n13655), .ZN(P3_U3473) );
  INV_X1 U15816 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13658) );
  AOI21_X1 U15817 ( .B1(n15905), .B2(n13657), .A(n13656), .ZN(n13708) );
  MUX2_X1 U15818 ( .A(n13658), .B(n13708), .S(n15954), .Z(n13659) );
  OAI21_X1 U15819 ( .B1(n13712), .B2(n13660), .A(n13659), .ZN(P3_U3471) );
  NAND2_X1 U15820 ( .A1(n15941), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U15821 ( .A1(n13661), .A2(n15943), .ZN(n13665) );
  OAI211_X1 U15822 ( .C1(n13663), .C2(n13711), .A(n13662), .B(n13665), .ZN(
        P3_U3458) );
  NAND2_X1 U15823 ( .A1(n13664), .A2(n13675), .ZN(n13666) );
  OAI211_X1 U15824 ( .C1(n15943), .C2(n13667), .A(n13666), .B(n13665), .ZN(
        P3_U3457) );
  OAI21_X1 U15825 ( .B1(n13671), .B2(n13711), .A(n13670), .ZN(P3_U3455) );
  MUX2_X1 U15826 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13672), .S(n15943), .Z(
        n13673) );
  AOI21_X1 U15827 ( .B1(n13675), .B2(n13674), .A(n13673), .ZN(n13676) );
  INV_X1 U15828 ( .A(n13676), .ZN(P3_U3454) );
  MUX2_X1 U15829 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13677), .S(n15943), .Z(
        P3_U3453) );
  MUX2_X1 U15830 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13678), .S(n15943), .Z(
        P3_U3452) );
  MUX2_X1 U15831 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13679), .S(n15943), .Z(
        P3_U3451) );
  INV_X1 U15832 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13681) );
  MUX2_X1 U15833 ( .A(n13681), .B(n13680), .S(n15943), .Z(n13682) );
  OAI21_X1 U15834 ( .B1(n13683), .B2(n13711), .A(n13682), .ZN(P3_U3450) );
  INV_X1 U15835 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13685) );
  MUX2_X1 U15836 ( .A(n13685), .B(n13684), .S(n15943), .Z(n13686) );
  OAI21_X1 U15837 ( .B1(n13687), .B2(n13711), .A(n13686), .ZN(P3_U3449) );
  INV_X1 U15838 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13689) );
  MUX2_X1 U15839 ( .A(n13689), .B(n13688), .S(n15943), .Z(n13690) );
  OAI21_X1 U15840 ( .B1(n13691), .B2(n13711), .A(n13690), .ZN(P3_U3448) );
  MUX2_X1 U15841 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13692), .S(n15943), .Z(
        P3_U3447) );
  INV_X1 U15842 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13694) );
  MUX2_X1 U15843 ( .A(n13694), .B(n13693), .S(n15943), .Z(n13695) );
  OAI21_X1 U15844 ( .B1(n13696), .B2(n13711), .A(n13695), .ZN(P3_U3446) );
  MUX2_X1 U15845 ( .A(n13698), .B(n13697), .S(n15943), .Z(n13699) );
  OAI21_X1 U15846 ( .B1(n13700), .B2(n13711), .A(n13699), .ZN(P3_U3444) );
  MUX2_X1 U15847 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13701), .S(n15943), .Z(
        P3_U3441) );
  MUX2_X1 U15848 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13702), .S(n15943), .Z(
        P3_U3438) );
  MUX2_X1 U15849 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13703), .S(n15943), .Z(
        P3_U3435) );
  INV_X1 U15850 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13705) );
  MUX2_X1 U15851 ( .A(n13705), .B(n13704), .S(n15943), .Z(n13706) );
  OAI21_X1 U15852 ( .B1(n13711), .B2(n13707), .A(n13706), .ZN(P3_U3432) );
  INV_X1 U15853 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13709) );
  MUX2_X1 U15854 ( .A(n13709), .B(n13708), .S(n15943), .Z(n13710) );
  OAI21_X1 U15855 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(P3_U3426) );
  MUX2_X1 U15856 ( .A(P3_D_REG_0__SCAN_IN), .B(n13714), .S(n13713), .Z(
        P3_U3376) );
  INV_X1 U15857 ( .A(n13715), .ZN(n13720) );
  NOR4_X1 U15858 ( .A1(n6857), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n9019), .ZN(n13717) );
  AOI21_X1 U15859 ( .B1(SI_31_), .B2(n13718), .A(n13717), .ZN(n13719) );
  OAI21_X1 U15860 ( .B1(n13720), .B2(n13729), .A(n13719), .ZN(P3_U3264) );
  INV_X1 U15861 ( .A(n13721), .ZN(n13724) );
  OAI222_X1 U15862 ( .A1(n13725), .A2(n13724), .B1(n13723), .B2(P3_U3151), 
        .C1(n13722), .C2(n13731), .ZN(P3_U3266) );
  INV_X1 U15863 ( .A(SI_27_), .ZN(n13730) );
  INV_X1 U15864 ( .A(n13726), .ZN(n13728) );
  OAI222_X1 U15865 ( .A1(n13731), .A2(n13730), .B1(n13729), .B2(n13728), .C1(
        P3_U3151), .C2(n13285), .ZN(P3_U3268) );
  XNOR2_X1 U15866 ( .A(n14604), .B(n13799), .ZN(n13734) );
  OR2_X1 U15867 ( .A1(n13839), .A2(n13800), .ZN(n13735) );
  NAND2_X1 U15868 ( .A1(n13734), .A2(n13735), .ZN(n13739) );
  INV_X1 U15869 ( .A(n13734), .ZN(n13737) );
  INV_X1 U15870 ( .A(n13735), .ZN(n13736) );
  NAND2_X1 U15871 ( .A1(n13737), .A2(n13736), .ZN(n13738) );
  AND2_X1 U15872 ( .A1(n13739), .A2(n13738), .ZN(n13935) );
  NAND2_X1 U15873 ( .A1(n13934), .A2(n13935), .ZN(n13933) );
  XNOR2_X1 U15874 ( .A(n13842), .B(n13864), .ZN(n13741) );
  NOR2_X1 U15875 ( .A1(n13977), .A2(n13800), .ZN(n13740) );
  XNOR2_X1 U15876 ( .A(n13741), .B(n13740), .ZN(n13837) );
  XNOR2_X1 U15877 ( .A(n14598), .B(n13799), .ZN(n13742) );
  NAND2_X1 U15878 ( .A1(n13862), .A2(n14033), .ZN(n13743) );
  NAND2_X1 U15879 ( .A1(n13742), .A2(n13743), .ZN(n13747) );
  INV_X1 U15880 ( .A(n13742), .ZN(n13745) );
  INV_X1 U15881 ( .A(n13743), .ZN(n13744) );
  NAND2_X1 U15882 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  AND2_X1 U15883 ( .A1(n13747), .A2(n13746), .ZN(n13973) );
  XNOR2_X1 U15884 ( .A(n14593), .B(n13864), .ZN(n13748) );
  NOR2_X1 U15885 ( .A1(n13958), .A2(n13800), .ZN(n13749) );
  NAND2_X1 U15886 ( .A1(n13748), .A2(n13749), .ZN(n13881) );
  INV_X1 U15887 ( .A(n13748), .ZN(n13751) );
  INV_X1 U15888 ( .A(n13749), .ZN(n13750) );
  NAND2_X1 U15889 ( .A1(n13751), .A2(n13750), .ZN(n13882) );
  XNOR2_X1 U15890 ( .A(n14589), .B(n13864), .ZN(n13752) );
  AND2_X1 U15891 ( .A1(n13862), .A2(n14032), .ZN(n13753) );
  NAND2_X1 U15892 ( .A1(n13752), .A2(n13753), .ZN(n13814) );
  INV_X1 U15893 ( .A(n13752), .ZN(n13755) );
  INV_X1 U15894 ( .A(n13753), .ZN(n13754) );
  NAND2_X1 U15895 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  NAND2_X1 U15896 ( .A1(n13814), .A2(n13756), .ZN(n13955) );
  XNOR2_X1 U15897 ( .A(n14583), .B(n13864), .ZN(n13757) );
  NAND2_X1 U15898 ( .A1(n13862), .A2(n14031), .ZN(n13758) );
  XNOR2_X1 U15899 ( .A(n13757), .B(n13758), .ZN(n13815) );
  XNOR2_X1 U15900 ( .A(n14578), .B(n13799), .ZN(n13905) );
  NAND2_X1 U15901 ( .A1(n14030), .A2(n13862), .ZN(n13903) );
  INV_X1 U15902 ( .A(n13757), .ZN(n13759) );
  AND2_X1 U15903 ( .A1(n13759), .A2(n13758), .ZN(n13899) );
  AOI21_X1 U15904 ( .B1(n13905), .B2(n13903), .A(n13899), .ZN(n13760) );
  XNOR2_X1 U15905 ( .A(n14573), .B(n13799), .ZN(n13898) );
  NAND2_X1 U15906 ( .A1(n14029), .A2(n13862), .ZN(n13897) );
  NAND2_X1 U15907 ( .A1(n13898), .A2(n13897), .ZN(n13914) );
  AND2_X1 U15908 ( .A1(n13760), .A2(n13914), .ZN(n13766) );
  NAND2_X1 U15909 ( .A1(n14028), .A2(n13862), .ZN(n13768) );
  XNOR2_X1 U15910 ( .A(n13767), .B(n13768), .ZN(n13915) );
  OAI21_X1 U15911 ( .B1(n13905), .B2(n13903), .A(n13897), .ZN(n13763) );
  INV_X1 U15912 ( .A(n13898), .ZN(n13762) );
  NOR2_X1 U15913 ( .A1(n13897), .A2(n13903), .ZN(n13761) );
  INV_X1 U15914 ( .A(n13905), .ZN(n13902) );
  AOI22_X1 U15915 ( .A1(n13763), .A2(n13762), .B1(n13761), .B2(n13902), .ZN(
        n13764) );
  NAND2_X1 U15916 ( .A1(n13915), .A2(n13764), .ZN(n13765) );
  XNOR2_X1 U15917 ( .A(n14562), .B(n13864), .ZN(n13847) );
  NAND2_X1 U15918 ( .A1(n14027), .A2(n13862), .ZN(n13846) );
  INV_X1 U15919 ( .A(n13846), .ZN(n13771) );
  NAND2_X1 U15920 ( .A1(n13847), .A2(n13771), .ZN(n13848) );
  XNOR2_X1 U15921 ( .A(n14557), .B(n13864), .ZN(n13774) );
  NOR2_X1 U15922 ( .A1(n14337), .A2(n13800), .ZN(n13775) );
  NOR2_X1 U15923 ( .A1(n13774), .A2(n13775), .ZN(n13850) );
  INV_X1 U15924 ( .A(n13767), .ZN(n13769) );
  AND2_X1 U15925 ( .A1(n13769), .A2(n13768), .ZN(n13845) );
  NOR2_X1 U15926 ( .A1(n13845), .A2(n13846), .ZN(n13772) );
  INV_X1 U15927 ( .A(n13845), .ZN(n13770) );
  OAI22_X1 U15928 ( .A1(n13772), .A2(n13847), .B1(n13771), .B2(n13770), .ZN(
        n13773) );
  INV_X1 U15929 ( .A(n13774), .ZN(n13777) );
  INV_X1 U15930 ( .A(n13775), .ZN(n13776) );
  NOR2_X1 U15931 ( .A1(n13777), .A2(n13776), .ZN(n13849) );
  NOR2_X1 U15932 ( .A1(n14349), .A2(n13800), .ZN(n13779) );
  XNOR2_X1 U15933 ( .A(n14553), .B(n13864), .ZN(n13778) );
  NOR2_X1 U15934 ( .A1(n13778), .A2(n13779), .ZN(n13780) );
  AOI21_X1 U15935 ( .B1(n13779), .B2(n13778), .A(n13780), .ZN(n13947) );
  INV_X1 U15936 ( .A(n13780), .ZN(n13781) );
  NAND2_X1 U15937 ( .A1(n14024), .A2(n13862), .ZN(n13783) );
  XNOR2_X1 U15938 ( .A(n14548), .B(n13864), .ZN(n13782) );
  XOR2_X1 U15939 ( .A(n13783), .B(n13782), .Z(n13873) );
  INV_X1 U15940 ( .A(n13782), .ZN(n13784) );
  XNOR2_X1 U15941 ( .A(n14543), .B(n13864), .ZN(n13788) );
  INV_X1 U15942 ( .A(n13788), .ZN(n13785) );
  XNOR2_X1 U15943 ( .A(n13789), .B(n13785), .ZN(n13824) );
  XNOR2_X1 U15944 ( .A(n14538), .B(n13864), .ZN(n13827) );
  NOR2_X1 U15945 ( .A1(n14287), .A2(n13800), .ZN(n13964) );
  INV_X1 U15946 ( .A(n13786), .ZN(n13787) );
  NAND2_X1 U15947 ( .A1(n13824), .A2(n13787), .ZN(n13792) );
  NOR2_X1 U15948 ( .A1(n14268), .A2(n13800), .ZN(n13826) );
  NAND2_X1 U15949 ( .A1(n13827), .A2(n13826), .ZN(n13790) );
  XNOR2_X1 U15950 ( .A(n14532), .B(n13864), .ZN(n13794) );
  NAND2_X1 U15951 ( .A1(n14021), .A2(n13862), .ZN(n13793) );
  XNOR2_X1 U15952 ( .A(n13794), .B(n13793), .ZN(n13925) );
  INV_X1 U15953 ( .A(n13793), .ZN(n13795) );
  NAND2_X1 U15954 ( .A1(n14020), .A2(n13862), .ZN(n13797) );
  XNOR2_X1 U15955 ( .A(n14527), .B(n13864), .ZN(n13796) );
  XOR2_X1 U15956 ( .A(n13797), .B(n13796), .Z(n13890) );
  INV_X1 U15957 ( .A(n13796), .ZN(n13798) );
  XNOR2_X1 U15958 ( .A(n14519), .B(n13799), .ZN(n13803) );
  OR2_X1 U15959 ( .A1(n13801), .A2(n13800), .ZN(n13802) );
  NAND2_X1 U15960 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  OAI21_X1 U15961 ( .B1(n13803), .B2(n13802), .A(n13804), .ZN(n13995) );
  XNOR2_X1 U15962 ( .A(n14225), .B(n13864), .ZN(n13858) );
  NAND2_X1 U15963 ( .A1(n14018), .A2(n13862), .ZN(n13857) );
  XNOR2_X1 U15964 ( .A(n13861), .B(n13860), .ZN(n13812) );
  INV_X1 U15965 ( .A(n14224), .ZN(n13806) );
  OAI22_X1 U15966 ( .A1(n13806), .A2(n13990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13805), .ZN(n13809) );
  NOR2_X1 U15967 ( .A1(n13807), .A2(n14014), .ZN(n13808) );
  AOI211_X1 U15968 ( .C1(n13992), .C2(n13810), .A(n13809), .B(n13808), .ZN(
        n13811) );
  OAI21_X1 U15969 ( .B1(n13812), .B2(n14002), .A(n13811), .ZN(P2_U3186) );
  AND2_X1 U15970 ( .A1(n13813), .A2(n13814), .ZN(n13816) );
  OAI21_X1 U15971 ( .B1(n13816), .B2(n13815), .A(n6864), .ZN(n13817) );
  NAND2_X1 U15972 ( .A1(n13817), .A2(n14004), .ZN(n13823) );
  INV_X1 U15973 ( .A(n13992), .ZN(n14009) );
  NAND2_X1 U15974 ( .A1(n14030), .A2(n14494), .ZN(n13819) );
  NAND2_X1 U15975 ( .A1(n14032), .A2(n14496), .ZN(n13818) );
  AND2_X1 U15976 ( .A1(n13819), .A2(n13818), .ZN(n14439) );
  OAI22_X1 U15977 ( .A1(n14009), .A2(n14439), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13820), .ZN(n13821) );
  AOI21_X1 U15978 ( .B1(n14442), .B2(n14011), .A(n13821), .ZN(n13822) );
  OAI211_X1 U15979 ( .C1(n14445), .C2(n14014), .A(n13823), .B(n13822), .ZN(
        P2_U3187) );
  AOI21_X1 U15980 ( .B1(n13965), .B2(n13964), .A(n13825), .ZN(n13829) );
  XNOR2_X1 U15981 ( .A(n13827), .B(n13826), .ZN(n13828) );
  XNOR2_X1 U15982 ( .A(n13829), .B(n13828), .ZN(n13835) );
  OAI22_X1 U15983 ( .A1(n14286), .A2(n13950), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13830), .ZN(n13833) );
  INV_X1 U15984 ( .A(n14291), .ZN(n13831) );
  OAI22_X1 U15985 ( .A1(n13978), .A2(n14287), .B1(n13990), .B2(n13831), .ZN(
        n13832) );
  AOI211_X1 U15986 ( .C1(n14538), .C2(n14000), .A(n13833), .B(n13832), .ZN(
        n13834) );
  OAI21_X1 U15987 ( .B1(n13835), .B2(n14002), .A(n13834), .ZN(P2_U3188) );
  XNOR2_X1 U15988 ( .A(n13836), .B(n13837), .ZN(n13844) );
  NAND2_X1 U15989 ( .A1(n6531), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U15990 ( .B1(n13950), .B2(n14472), .A(n14142), .ZN(n13841) );
  OAI22_X1 U15991 ( .A1(n13978), .A2(n13839), .B1(n13990), .B2(n13838), .ZN(
        n13840) );
  AOI211_X1 U15992 ( .C1(n13842), .C2(n14000), .A(n13841), .B(n13840), .ZN(
        n13843) );
  OAI21_X1 U15993 ( .B1(n13844), .B2(n14002), .A(n13843), .ZN(P2_U3189) );
  NOR2_X1 U15994 ( .A1(n6672), .A2(n13845), .ZN(n13986) );
  XNOR2_X1 U15995 ( .A(n13847), .B(n13846), .ZN(n13985) );
  NAND2_X1 U15996 ( .A1(n13986), .A2(n13985), .ZN(n13984) );
  NAND2_X1 U15997 ( .A1(n13984), .A2(n13848), .ZN(n13852) );
  NOR2_X1 U15998 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  XNOR2_X1 U15999 ( .A(n13852), .B(n13851), .ZN(n13856) );
  NAND2_X1 U16000 ( .A1(n6531), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14211) );
  OAI21_X1 U16001 ( .B1(n13978), .B2(n14348), .A(n14211), .ZN(n13854) );
  OAI22_X1 U16002 ( .A1(n13950), .A2(n14349), .B1(n13990), .B2(n14358), .ZN(
        n13853) );
  AOI211_X1 U16003 ( .C1(n14557), .C2(n14000), .A(n13854), .B(n13853), .ZN(
        n13855) );
  OAI21_X1 U16004 ( .B1(n13856), .B2(n14002), .A(n13855), .ZN(P2_U3191) );
  INV_X1 U16005 ( .A(n13857), .ZN(n13859) );
  NAND2_X1 U16006 ( .A1(n14017), .A2(n13862), .ZN(n13863) );
  XOR2_X1 U16007 ( .A(n13864), .B(n13863), .Z(n13865) );
  OAI22_X1 U16008 ( .A1(n14213), .A2(n13990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13866), .ZN(n13869) );
  NOR2_X1 U16009 ( .A1(n13867), .A2(n14014), .ZN(n13868) );
  AOI211_X1 U16010 ( .C1(n13992), .C2(n13870), .A(n13869), .B(n13868), .ZN(
        n13871) );
  OAI21_X1 U16011 ( .B1(n13872), .B2(n14002), .A(n13871), .ZN(P2_U3192) );
  XNOR2_X1 U16012 ( .A(n13874), .B(n13873), .ZN(n13879) );
  AOI22_X1 U16013 ( .A1(n14023), .A2(n14494), .B1(n14496), .B2(n14025), .ZN(
        n14319) );
  OAI22_X1 U16014 ( .A1(n14319), .A2(n14009), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13875), .ZN(n13876) );
  AOI21_X1 U16015 ( .B1(n14323), .B2(n14011), .A(n13876), .ZN(n13878) );
  NAND2_X1 U16016 ( .A1(n14548), .A2(n14000), .ZN(n13877) );
  OAI211_X1 U16017 ( .C1(n13879), .C2(n14002), .A(n13878), .B(n13877), .ZN(
        P2_U3195) );
  NAND2_X1 U16018 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  XNOR2_X1 U16019 ( .A(n13880), .B(n13883), .ZN(n13889) );
  INV_X1 U16020 ( .A(n14483), .ZN(n13884) );
  OAI22_X1 U16021 ( .A1(n13950), .A2(n14474), .B1(n13990), .B2(n13884), .ZN(
        n13886) );
  NAND2_X1 U16022 ( .A1(n6531), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15751) );
  OAI21_X1 U16023 ( .B1(n13978), .B2(n14472), .A(n15751), .ZN(n13885) );
  NOR2_X1 U16024 ( .A1(n13886), .A2(n13885), .ZN(n13888) );
  NAND2_X1 U16025 ( .A1(n14593), .A2(n14000), .ZN(n13887) );
  OAI211_X1 U16026 ( .C1(n13889), .C2(n14002), .A(n13888), .B(n13887), .ZN(
        P2_U3196) );
  XNOR2_X1 U16027 ( .A(n13891), .B(n13890), .ZN(n13896) );
  AOI22_X1 U16028 ( .A1(n14019), .A2(n14494), .B1(n14496), .B2(n14021), .ZN(
        n14250) );
  INV_X1 U16029 ( .A(n14250), .ZN(n13892) );
  AOI22_X1 U16030 ( .A1(n13892), .A2(n13992), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(n6531), .ZN(n13893) );
  OAI21_X1 U16031 ( .B1(n14257), .B2(n13990), .A(n13893), .ZN(n13894) );
  AOI21_X1 U16032 ( .B1(n14527), .B2(n14000), .A(n13894), .ZN(n13895) );
  OAI21_X1 U16033 ( .B1(n13896), .B2(n14002), .A(n13895), .ZN(P2_U3197) );
  XNOR2_X1 U16034 ( .A(n13898), .B(n13897), .ZN(n13907) );
  INV_X1 U16035 ( .A(n13899), .ZN(n13900) );
  NAND2_X1 U16036 ( .A1(n6864), .A2(n13900), .ZN(n13904) );
  XNOR2_X1 U16037 ( .A(n13904), .B(n13902), .ZN(n14007) );
  INV_X1 U16038 ( .A(n13903), .ZN(n14006) );
  NAND2_X1 U16039 ( .A1(n14007), .A2(n14006), .ZN(n14005) );
  OAI21_X1 U16040 ( .B1(n13905), .B2(n13904), .A(n14005), .ZN(n13906) );
  NOR2_X1 U16041 ( .A1(n13906), .A2(n13907), .ZN(n13917) );
  AOI21_X1 U16042 ( .B1(n13907), .B2(n13906), .A(n13917), .ZN(n13913) );
  NOR2_X1 U16043 ( .A1(n13990), .A2(n14407), .ZN(n13911) );
  AND2_X1 U16044 ( .A1(n14030), .A2(n14496), .ZN(n13908) );
  AOI21_X1 U16045 ( .B1(n14028), .B2(n14494), .A(n13908), .ZN(n14412) );
  OAI22_X1 U16046 ( .A1(n14009), .A2(n14412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13909), .ZN(n13910) );
  AOI211_X1 U16047 ( .C1(n14573), .C2(n14000), .A(n13911), .B(n13910), .ZN(
        n13912) );
  OAI21_X1 U16048 ( .B1(n13913), .B2(n14002), .A(n13912), .ZN(P2_U3198) );
  INV_X1 U16049 ( .A(n13914), .ZN(n13916) );
  NOR3_X1 U16050 ( .A1(n13917), .A2(n13916), .A3(n13915), .ZN(n13918) );
  OAI21_X1 U16051 ( .B1(n13918), .B2(n6672), .A(n14004), .ZN(n13923) );
  INV_X1 U16052 ( .A(n14390), .ZN(n13921) );
  AND2_X1 U16053 ( .A1(n14029), .A2(n14496), .ZN(n13919) );
  AOI21_X1 U16054 ( .B1(n14027), .B2(n14494), .A(n13919), .ZN(n14385) );
  OAI22_X1 U16055 ( .A1(n14009), .A2(n14385), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14170), .ZN(n13920) );
  AOI21_X1 U16056 ( .B1(n13921), .B2(n14011), .A(n13920), .ZN(n13922) );
  OAI211_X1 U16057 ( .C1(n13924), .C2(n14014), .A(n13923), .B(n13922), .ZN(
        P2_U3200) );
  XNOR2_X1 U16058 ( .A(n13926), .B(n13925), .ZN(n13932) );
  OAI22_X1 U16059 ( .A1(n14267), .A2(n13950), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13927), .ZN(n13930) );
  INV_X1 U16060 ( .A(n14269), .ZN(n13928) );
  OAI22_X1 U16061 ( .A1(n14268), .A2(n13978), .B1(n13928), .B2(n13990), .ZN(
        n13929) );
  AOI211_X1 U16062 ( .C1(n14532), .C2(n14000), .A(n13930), .B(n13929), .ZN(
        n13931) );
  OAI21_X1 U16063 ( .B1(n13932), .B2(n14002), .A(n13931), .ZN(P2_U3201) );
  OAI21_X1 U16064 ( .B1(n13935), .B2(n13934), .A(n13933), .ZN(n13936) );
  NAND2_X1 U16065 ( .A1(n13936), .A2(n14004), .ZN(n13943) );
  NAND2_X1 U16066 ( .A1(n6531), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n15728) );
  INV_X1 U16067 ( .A(n15728), .ZN(n13941) );
  INV_X1 U16068 ( .A(n13937), .ZN(n13938) );
  OAI22_X1 U16069 ( .A1(n13978), .A2(n13939), .B1(n13990), .B2(n13938), .ZN(
        n13940) );
  AOI211_X1 U16070 ( .C1(n13981), .C2(n14497), .A(n13941), .B(n13940), .ZN(
        n13942) );
  OAI211_X1 U16071 ( .C1(n13944), .C2(n14014), .A(n13943), .B(n13942), .ZN(
        P2_U3203) );
  INV_X1 U16072 ( .A(n14553), .ZN(n14341) );
  OAI21_X1 U16073 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n13948) );
  NAND2_X1 U16074 ( .A1(n13948), .A2(n14004), .ZN(n13954) );
  NOR2_X1 U16075 ( .A1(n13978), .A2(n14337), .ZN(n13952) );
  OAI22_X1 U16076 ( .A1(n13950), .A2(n14336), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13949), .ZN(n13951) );
  AOI211_X1 U16077 ( .C1(n14011), .C2(n14339), .A(n13952), .B(n13951), .ZN(
        n13953) );
  OAI211_X1 U16078 ( .C1(n14341), .C2(n14014), .A(n13954), .B(n13953), .ZN(
        P2_U3205) );
  INV_X1 U16079 ( .A(n14589), .ZN(n14455) );
  AOI21_X1 U16080 ( .B1(n13956), .B2(n13955), .A(n14002), .ZN(n13957) );
  NAND2_X1 U16081 ( .A1(n13957), .A2(n13813), .ZN(n13963) );
  OR2_X1 U16082 ( .A1(n13958), .A2(n14471), .ZN(n13960) );
  NAND2_X1 U16083 ( .A1(n14031), .A2(n14494), .ZN(n13959) );
  AND2_X1 U16084 ( .A1(n13960), .A2(n13959), .ZN(n14460) );
  OAI22_X1 U16085 ( .A1(n14009), .A2(n14460), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14154), .ZN(n13961) );
  AOI21_X1 U16086 ( .B1(n14453), .B2(n14011), .A(n13961), .ZN(n13962) );
  OAI211_X1 U16087 ( .C1(n14455), .C2(n14014), .A(n13963), .B(n13962), .ZN(
        P2_U3206) );
  XNOR2_X1 U16088 ( .A(n13965), .B(n13964), .ZN(n13971) );
  OR2_X1 U16089 ( .A1(n14268), .A2(n14473), .ZN(n13967) );
  NAND2_X1 U16090 ( .A1(n14024), .A2(n14496), .ZN(n13966) );
  NAND2_X1 U16091 ( .A1(n13967), .A2(n13966), .ZN(n14301) );
  AOI22_X1 U16092 ( .A1(n14301), .A2(n13992), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(n6531), .ZN(n13968) );
  OAI21_X1 U16093 ( .B1(n14307), .B2(n13990), .A(n13968), .ZN(n13969) );
  AOI21_X1 U16094 ( .B1(n14543), .B2(n14000), .A(n13969), .ZN(n13970) );
  OAI21_X1 U16095 ( .B1(n13971), .B2(n14002), .A(n13970), .ZN(P2_U3207) );
  OAI21_X1 U16096 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13975) );
  NAND2_X1 U16097 ( .A1(n13975), .A2(n14004), .ZN(n13983) );
  INV_X1 U16098 ( .A(n14501), .ZN(n13976) );
  OAI22_X1 U16099 ( .A1(n13978), .A2(n13977), .B1(n13990), .B2(n13976), .ZN(
        n13979) );
  AOI211_X1 U16100 ( .C1(n13981), .C2(n14495), .A(n13980), .B(n13979), .ZN(
        n13982) );
  OAI211_X1 U16101 ( .C1(n14505), .C2(n14014), .A(n13983), .B(n13982), .ZN(
        P2_U3208) );
  OAI211_X1 U16102 ( .C1(n13986), .C2(n13985), .A(n13984), .B(n14004), .ZN(
        n13994) );
  OAI22_X1 U16103 ( .A1(n14337), .A2(n14473), .B1(n13987), .B2(n14471), .ZN(
        n14366) );
  NOR2_X1 U16104 ( .A1(n13988), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14184) );
  INV_X1 U16105 ( .A(n14369), .ZN(n13989) );
  NOR2_X1 U16106 ( .A1(n13990), .A2(n13989), .ZN(n13991) );
  AOI211_X1 U16107 ( .C1(n13992), .C2(n14366), .A(n14184), .B(n13991), .ZN(
        n13993) );
  OAI211_X1 U16108 ( .C1(n14371), .C2(n14014), .A(n13994), .B(n13993), .ZN(
        P2_U3210) );
  AOI21_X1 U16109 ( .B1(n13996), .B2(n13995), .A(n6699), .ZN(n14003) );
  AND2_X1 U16110 ( .A1(n14020), .A2(n14496), .ZN(n13997) );
  AOI21_X1 U16111 ( .B1(n14018), .B2(n14494), .A(n13997), .ZN(n14244) );
  AOI22_X1 U16112 ( .A1(n14238), .A2(n14011), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(n6531), .ZN(n13998) );
  OAI21_X1 U16113 ( .B1(n14244), .B2(n14009), .A(n13998), .ZN(n13999) );
  AOI21_X1 U16114 ( .B1(n14519), .B2(n14000), .A(n13999), .ZN(n14001) );
  OAI21_X1 U16115 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(P2_U3212) );
  OAI211_X1 U16116 ( .C1(n14007), .C2(n14006), .A(n14005), .B(n14004), .ZN(
        n14013) );
  AOI22_X1 U16117 ( .A1(n14029), .A2(n14494), .B1(n14496), .B2(n14031), .ZN(
        n14431) );
  OAI22_X1 U16118 ( .A1(n14009), .A2(n14431), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14008), .ZN(n14010) );
  AOI21_X1 U16119 ( .B1(n14423), .B2(n14011), .A(n14010), .ZN(n14012) );
  OAI211_X1 U16120 ( .C1(n14425), .C2(n14014), .A(n14013), .B(n14012), .ZN(
        P2_U3213) );
  MUX2_X1 U16121 ( .A(n14015), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14042), .Z(
        P2_U3562) );
  MUX2_X1 U16122 ( .A(n14016), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14042), .Z(
        P2_U3561) );
  MUX2_X1 U16123 ( .A(n14017), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14042), .Z(
        P2_U3559) );
  MUX2_X1 U16124 ( .A(n14018), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14042), .Z(
        P2_U3558) );
  MUX2_X1 U16125 ( .A(n14019), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14042), .Z(
        P2_U3557) );
  MUX2_X1 U16126 ( .A(n14020), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14042), .Z(
        P2_U3556) );
  MUX2_X1 U16127 ( .A(n14021), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14042), .Z(
        P2_U3555) );
  MUX2_X1 U16128 ( .A(n14022), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14042), .Z(
        P2_U3554) );
  MUX2_X1 U16129 ( .A(n14023), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14042), .Z(
        P2_U3553) );
  MUX2_X1 U16130 ( .A(n14024), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14042), .Z(
        P2_U3552) );
  MUX2_X1 U16131 ( .A(n14025), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14042), .Z(
        P2_U3551) );
  MUX2_X1 U16132 ( .A(n14026), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14042), .Z(
        P2_U3550) );
  MUX2_X1 U16133 ( .A(n14027), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14042), .Z(
        P2_U3549) );
  MUX2_X1 U16134 ( .A(n14028), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14042), .Z(
        P2_U3548) );
  MUX2_X1 U16135 ( .A(n14029), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14042), .Z(
        P2_U3547) );
  MUX2_X1 U16136 ( .A(n14030), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14042), .Z(
        P2_U3546) );
  MUX2_X1 U16137 ( .A(n14031), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14042), .Z(
        P2_U3545) );
  MUX2_X1 U16138 ( .A(n14032), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14042), .Z(
        P2_U3544) );
  MUX2_X1 U16139 ( .A(n14495), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14042), .Z(
        P2_U3543) );
  MUX2_X1 U16140 ( .A(n14033), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14042), .Z(
        P2_U3542) );
  MUX2_X1 U16141 ( .A(n14497), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14042), .Z(
        P2_U3541) );
  MUX2_X1 U16142 ( .A(n14034), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14042), .Z(
        P2_U3540) );
  MUX2_X1 U16143 ( .A(n14035), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14042), .Z(
        P2_U3539) );
  MUX2_X1 U16144 ( .A(n14036), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14042), .Z(
        P2_U3538) );
  MUX2_X1 U16145 ( .A(n14037), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14042), .Z(
        P2_U3537) );
  MUX2_X1 U16146 ( .A(n14038), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14042), .Z(
        P2_U3536) );
  MUX2_X1 U16147 ( .A(n14039), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14042), .Z(
        P2_U3535) );
  MUX2_X1 U16148 ( .A(n14040), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14042), .Z(
        P2_U3534) );
  MUX2_X1 U16149 ( .A(n14041), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14042), .Z(
        P2_U3533) );
  MUX2_X1 U16150 ( .A(n6596), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14042), .Z(
        P2_U3532) );
  MUX2_X1 U16151 ( .A(n9670), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14042), .Z(
        P2_U3531) );
  OAI211_X1 U16152 ( .C1(n14045), .C2(n14044), .A(n15744), .B(n14043), .ZN(
        n14053) );
  NOR2_X1 U16153 ( .A1(n15441), .A2(n15753), .ZN(n14046) );
  AOI21_X1 U16154 ( .B1(n6531), .B2(P2_REG3_REG_2__SCAN_IN), .A(n14046), .ZN(
        n14052) );
  OAI211_X1 U16155 ( .C1(n14048), .C2(n14047), .A(n15734), .B(n14060), .ZN(
        n14051) );
  NAND2_X1 U16156 ( .A1(n15747), .A2(n14049), .ZN(n14050) );
  NAND4_X1 U16157 ( .A1(n14053), .A2(n14052), .A3(n14051), .A4(n14050), .ZN(
        P2_U3216) );
  OAI211_X1 U16158 ( .C1(n14056), .C2(n14055), .A(n15744), .B(n14054), .ZN(
        n14066) );
  NOR2_X1 U16159 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11371), .ZN(n14057) );
  AOI21_X1 U16160 ( .B1(n15747), .B2(n14058), .A(n14057), .ZN(n14065) );
  NAND2_X1 U16161 ( .A1(n15715), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n14064) );
  MUX2_X1 U16162 ( .A(n11379), .B(P2_REG2_REG_3__SCAN_IN), .S(n14058), .Z(
        n14061) );
  NAND3_X1 U16163 ( .A1(n14061), .A2(n14060), .A3(n14059), .ZN(n14062) );
  NAND3_X1 U16164 ( .A1(n15734), .A2(n14076), .A3(n14062), .ZN(n14063) );
  NAND4_X1 U16165 ( .A1(n14066), .A2(n14065), .A3(n14064), .A4(n14063), .ZN(
        P2_U3217) );
  OAI211_X1 U16166 ( .C1(n14069), .C2(n14068), .A(n15744), .B(n14067), .ZN(
        n14081) );
  INV_X1 U16167 ( .A(n14070), .ZN(n14071) );
  AOI21_X1 U16168 ( .B1(n15747), .B2(n14072), .A(n14071), .ZN(n14080) );
  NAND2_X1 U16169 ( .A1(n15715), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14079) );
  MUX2_X1 U16170 ( .A(n14073), .B(P2_REG2_REG_4__SCAN_IN), .S(n14072), .Z(
        n14074) );
  NAND3_X1 U16171 ( .A1(n14076), .A2(n14075), .A3(n14074), .ZN(n14077) );
  NAND3_X1 U16172 ( .A1(n15734), .A2(n14090), .A3(n14077), .ZN(n14078) );
  NAND4_X1 U16173 ( .A1(n14081), .A2(n14080), .A3(n14079), .A4(n14078), .ZN(
        P2_U3218) );
  OAI211_X1 U16174 ( .C1(n14084), .C2(n14083), .A(n15744), .B(n14082), .ZN(
        n14096) );
  INV_X1 U16175 ( .A(n14085), .ZN(n14086) );
  AOI21_X1 U16176 ( .B1(n15747), .B2(n14087), .A(n14086), .ZN(n14095) );
  NAND2_X1 U16177 ( .A1(n15715), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n14094) );
  MUX2_X1 U16178 ( .A(n14088), .B(P2_REG2_REG_5__SCAN_IN), .S(n14087), .Z(
        n14091) );
  NAND3_X1 U16179 ( .A1(n14091), .A2(n14090), .A3(n14089), .ZN(n14092) );
  NAND3_X1 U16180 ( .A1(n15734), .A2(n14105), .A3(n14092), .ZN(n14093) );
  NAND4_X1 U16181 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        P2_U3219) );
  OAI211_X1 U16182 ( .C1(n14099), .C2(n14098), .A(n15744), .B(n14097), .ZN(
        n14110) );
  INV_X1 U16183 ( .A(n14100), .ZN(n14101) );
  AOI21_X1 U16184 ( .B1(n15747), .B2(n14102), .A(n14101), .ZN(n14109) );
  MUX2_X1 U16185 ( .A(n11557), .B(P2_REG2_REG_6__SCAN_IN), .S(n14102), .Z(
        n14103) );
  NAND3_X1 U16186 ( .A1(n14105), .A2(n14104), .A3(n14103), .ZN(n14106) );
  NAND3_X1 U16187 ( .A1(n15734), .A2(n14119), .A3(n14106), .ZN(n14108) );
  NAND2_X1 U16188 ( .A1(n15715), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14107) );
  NAND4_X1 U16189 ( .A1(n14110), .A2(n14109), .A3(n14108), .A4(n14107), .ZN(
        P2_U3220) );
  OAI211_X1 U16190 ( .C1(n14113), .C2(n14112), .A(n15744), .B(n14111), .ZN(
        n14124) );
  NOR2_X1 U16191 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8609), .ZN(n14114) );
  AOI21_X1 U16192 ( .B1(n15747), .B2(n14115), .A(n14114), .ZN(n14123) );
  MUX2_X1 U16193 ( .A(n14116), .B(P2_REG2_REG_7__SCAN_IN), .S(n14115), .Z(
        n14117) );
  NAND3_X1 U16194 ( .A1(n14119), .A2(n14118), .A3(n14117), .ZN(n14120) );
  NAND3_X1 U16195 ( .A1(n15734), .A2(n14132), .A3(n14120), .ZN(n14122) );
  NAND2_X1 U16196 ( .A1(n15715), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n14121) );
  NAND4_X1 U16197 ( .A1(n14124), .A2(n14123), .A3(n14122), .A4(n14121), .ZN(
        P2_U3221) );
  OAI21_X1 U16198 ( .B1(n14206), .B2(n14129), .A(n14125), .ZN(n14126) );
  AOI21_X1 U16199 ( .B1(n15715), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n14126), .ZN(
        n14137) );
  OAI211_X1 U16200 ( .C1(n14128), .C2(n14127), .A(n15744), .B(n15719), .ZN(
        n14136) );
  MUX2_X1 U16201 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11588), .S(n14129), .Z(
        n14130) );
  NAND3_X1 U16202 ( .A1(n14132), .A2(n14131), .A3(n14130), .ZN(n14133) );
  NAND3_X1 U16203 ( .A1(n15734), .A2(n14134), .A3(n14133), .ZN(n14135) );
  NAND3_X1 U16204 ( .A1(n14137), .A2(n14136), .A3(n14135), .ZN(P2_U3222) );
  AOI21_X1 U16205 ( .B1(n14139), .B2(n14138), .A(n14207), .ZN(n14141) );
  NAND2_X1 U16206 ( .A1(n14141), .A2(n14140), .ZN(n14150) );
  OAI21_X1 U16207 ( .B1(n14206), .B2(n14143), .A(n14142), .ZN(n14144) );
  AOI21_X1 U16208 ( .B1(n15715), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n14144), 
        .ZN(n14149) );
  OAI211_X1 U16209 ( .C1(n14147), .C2(n14146), .A(n15734), .B(n14145), .ZN(
        n14148) );
  NAND3_X1 U16210 ( .A1(n14150), .A2(n14149), .A3(n14148), .ZN(P2_U3224) );
  OAI211_X1 U16211 ( .C1(n14153), .C2(n14152), .A(n14151), .B(n15734), .ZN(
        n14164) );
  NOR2_X1 U16212 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14154), .ZN(n14157) );
  NOR2_X1 U16213 ( .A1(n14206), .A2(n14155), .ZN(n14156) );
  AOI211_X1 U16214 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n15715), .A(n14157), 
        .B(n14156), .ZN(n14163) );
  AOI21_X1 U16215 ( .B1(n14159), .B2(n14158), .A(n14207), .ZN(n14161) );
  NAND2_X1 U16216 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  NAND3_X1 U16217 ( .A1(n14164), .A2(n14163), .A3(n14162), .ZN(P2_U3227) );
  INV_X1 U16218 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14183) );
  MUX2_X1 U16219 ( .A(n14183), .B(P2_REG2_REG_17__SCAN_IN), .S(n14186), .Z(
        n14166) );
  NAND2_X1 U16220 ( .A1(n14166), .A2(n7041), .ZN(n14168) );
  MUX2_X1 U16221 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14183), .S(n14186), .Z(
        n14167) );
  OAI211_X1 U16222 ( .C1(n14169), .C2(n14168), .A(n14181), .B(n15734), .ZN(
        n14180) );
  NOR2_X1 U16223 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14170), .ZN(n14172) );
  NOR2_X1 U16224 ( .A1(n14206), .A2(n14182), .ZN(n14171) );
  AOI211_X1 U16225 ( .C1(n15715), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n14172), 
        .B(n14171), .ZN(n14179) );
  NAND2_X1 U16226 ( .A1(n14173), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n14174) );
  NAND2_X1 U16227 ( .A1(n14175), .A2(n14174), .ZN(n14177) );
  INV_X1 U16228 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14569) );
  XNOR2_X1 U16229 ( .A(n14186), .B(n14569), .ZN(n14176) );
  NAND2_X1 U16230 ( .A1(n14177), .A2(n14176), .ZN(n14188) );
  OAI211_X1 U16231 ( .C1(n14177), .C2(n14176), .A(n14188), .B(n15744), .ZN(
        n14178) );
  NAND3_X1 U16232 ( .A1(n14180), .A2(n14179), .A3(n14178), .ZN(P2_U3231) );
  NOR2_X1 U16233 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n6644), .ZN(n14200) );
  AOI21_X1 U16234 ( .B1(n6644), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14200), .ZN(
        n14198) );
  INV_X1 U16235 ( .A(n14184), .ZN(n14185) );
  OAI21_X1 U16236 ( .B1(n14206), .B2(n7042), .A(n14185), .ZN(n14195) );
  INV_X1 U16237 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14193) );
  NAND2_X1 U16238 ( .A1(n14186), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U16239 ( .A1(n14188), .A2(n14187), .ZN(n14190) );
  AND2_X1 U16240 ( .A1(n14190), .A2(n14189), .ZN(n14202) );
  NOR2_X1 U16241 ( .A1(n14190), .A2(n14189), .ZN(n14191) );
  OR2_X1 U16242 ( .A1(n14202), .A2(n14191), .ZN(n14192) );
  NOR2_X1 U16243 ( .A1(n14192), .A2(n14193), .ZN(n14203) );
  AOI211_X1 U16244 ( .C1(n14193), .C2(n14192), .A(n14207), .B(n14203), .ZN(
        n14194) );
  AOI211_X1 U16245 ( .C1(n15715), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14195), 
        .B(n14194), .ZN(n14196) );
  OAI21_X1 U16246 ( .B1(n14198), .B2(n14197), .A(n14196), .ZN(P2_U3232) );
  NOR2_X1 U16247 ( .A1(n14200), .A2(n14199), .ZN(n14201) );
  XOR2_X1 U16248 ( .A(n14201), .B(P2_REG2_REG_19__SCAN_IN), .Z(n14210) );
  NOR2_X1 U16249 ( .A1(n14203), .A2(n14202), .ZN(n14205) );
  XOR2_X1 U16250 ( .A(n14205), .B(n14204), .Z(n14209) );
  OAI21_X1 U16251 ( .B1(n14209), .B2(n14207), .A(n14206), .ZN(n14208) );
  INV_X1 U16252 ( .A(n14212), .ZN(n14217) );
  OAI22_X1 U16253 ( .A1(n14215), .A2(n14214), .B1(n14213), .B2(n14406), .ZN(
        n14216) );
  OAI21_X1 U16254 ( .B1(n14217), .B2(n14216), .A(n14499), .ZN(n14220) );
  AOI22_X1 U16255 ( .A1(n14218), .A2(n15759), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14484), .ZN(n14219) );
  OAI211_X1 U16256 ( .C1(n14221), .C2(n14465), .A(n14220), .B(n14219), .ZN(
        P2_U3237) );
  NAND3_X1 U16257 ( .A1(n14223), .A2(n14222), .A3(n15768), .ZN(n14231) );
  AOI22_X1 U16258 ( .A1(n14224), .A2(n15760), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14484), .ZN(n14227) );
  NAND2_X1 U16259 ( .A1(n14225), .A2(n15759), .ZN(n14226) );
  OAI211_X1 U16260 ( .C1(n14228), .C2(n14507), .A(n14227), .B(n14226), .ZN(
        n14229) );
  INV_X1 U16261 ( .A(n14229), .ZN(n14230) );
  OAI211_X1 U16262 ( .C1(n14232), .C2(n14484), .A(n14231), .B(n14230), .ZN(
        P2_U3238) );
  OAI21_X1 U16263 ( .B1(n14234), .B2(n14241), .A(n14233), .ZN(n14613) );
  INV_X1 U16264 ( .A(n14613), .ZN(n14248) );
  OAI21_X1 U16265 ( .B1(n14235), .B2(n8844), .A(n10957), .ZN(n14237) );
  NOR2_X1 U16266 ( .A1(n14237), .A2(n14236), .ZN(n14520) );
  AOI22_X1 U16267 ( .A1(n14238), .A2(n15760), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14484), .ZN(n14239) );
  OAI21_X1 U16268 ( .B1(n8844), .B2(n14486), .A(n14239), .ZN(n14240) );
  AOI21_X1 U16269 ( .B1(n14520), .B2(n15767), .A(n14240), .ZN(n14247) );
  XNOR2_X1 U16270 ( .A(n14242), .B(n14241), .ZN(n14243) );
  NAND2_X1 U16271 ( .A1(n14243), .A2(n15757), .ZN(n14245) );
  NAND2_X1 U16272 ( .A1(n14522), .A2(n14499), .ZN(n14246) );
  OAI211_X1 U16273 ( .C1(n14248), .C2(n14465), .A(n14247), .B(n14246), .ZN(
        P2_U3239) );
  XOR2_X1 U16274 ( .A(n14254), .B(n14249), .Z(n14251) );
  INV_X1 U16275 ( .A(n14525), .ZN(n14264) );
  AOI21_X1 U16276 ( .B1(n14252), .B2(n14254), .A(n14253), .ZN(n14524) );
  INV_X1 U16277 ( .A(n14527), .ZN(n14261) );
  NAND2_X1 U16278 ( .A1(n14270), .A2(n14527), .ZN(n14255) );
  NAND2_X1 U16279 ( .A1(n14255), .A2(n10957), .ZN(n14256) );
  NOR2_X1 U16280 ( .A1(n14235), .A2(n14256), .ZN(n14526) );
  NAND2_X1 U16281 ( .A1(n14526), .A2(n15767), .ZN(n14260) );
  INV_X1 U16282 ( .A(n14257), .ZN(n14258) );
  AOI22_X1 U16283 ( .A1(n14258), .A2(n15760), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14484), .ZN(n14259) );
  OAI211_X1 U16284 ( .C1(n14261), .C2(n14486), .A(n14260), .B(n14259), .ZN(
        n14262) );
  AOI21_X1 U16285 ( .B1(n14524), .B2(n15768), .A(n14262), .ZN(n14263) );
  OAI21_X1 U16286 ( .B1(n14484), .B2(n14264), .A(n14263), .ZN(P2_U3240) );
  XOR2_X1 U16287 ( .A(n14273), .B(n14265), .Z(n14266) );
  OAI222_X1 U16288 ( .A1(n14471), .A2(n14268), .B1(n14473), .B2(n14267), .C1(
        n14266), .C2(n14461), .ZN(n14530) );
  AOI21_X1 U16289 ( .B1(n14269), .B2(n15760), .A(n14530), .ZN(n14280) );
  AOI211_X1 U16290 ( .C1(n14532), .C2(n14281), .A(n14482), .B(n8990), .ZN(
        n14531) );
  INV_X1 U16291 ( .A(n14532), .ZN(n14272) );
  OAI22_X1 U16292 ( .A1(n14272), .A2(n14486), .B1(n14499), .B2(n14271), .ZN(
        n14278) );
  AND2_X1 U16293 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  OR2_X1 U16294 ( .A1(n14276), .A2(n14275), .ZN(n14621) );
  NOR2_X1 U16295 ( .A1(n14621), .A2(n14465), .ZN(n14277) );
  AOI211_X1 U16296 ( .C1(n14531), .C2(n14457), .A(n14278), .B(n14277), .ZN(
        n14279) );
  OAI21_X1 U16297 ( .B1(n14280), .B2(n14484), .A(n14279), .ZN(P2_U3241) );
  INV_X1 U16298 ( .A(n14305), .ZN(n14283) );
  INV_X1 U16299 ( .A(n14281), .ZN(n14282) );
  AOI211_X1 U16300 ( .C1(n14538), .C2(n14283), .A(n14482), .B(n14282), .ZN(
        n14537) );
  AOI21_X1 U16301 ( .B1(n14289), .B2(n14284), .A(n6700), .ZN(n14285) );
  OAI222_X1 U16302 ( .A1(n14471), .A2(n14287), .B1(n14473), .B2(n14286), .C1(
        n14285), .C2(n14461), .ZN(n14536) );
  AOI21_X1 U16303 ( .B1(n14537), .B2(n6547), .A(n14536), .ZN(n14296) );
  OAI21_X1 U16304 ( .B1(n14290), .B2(n14289), .A(n14288), .ZN(n14535) );
  AOI22_X1 U16305 ( .A1(n14484), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14291), 
        .B2(n15760), .ZN(n14292) );
  OAI21_X1 U16306 ( .B1(n14293), .B2(n14486), .A(n14292), .ZN(n14294) );
  AOI21_X1 U16307 ( .B1(n14535), .B2(n15768), .A(n14294), .ZN(n14295) );
  OAI21_X1 U16308 ( .B1(n14296), .B2(n14484), .A(n14295), .ZN(P2_U3242) );
  OAI21_X1 U16309 ( .B1(n14298), .B2(n14299), .A(n14297), .ZN(n14629) );
  XNOR2_X1 U16310 ( .A(n14300), .B(n14299), .ZN(n14303) );
  INV_X1 U16311 ( .A(n14301), .ZN(n14302) );
  OAI21_X1 U16312 ( .B1(n14303), .B2(n14461), .A(n14302), .ZN(n14541) );
  NAND2_X1 U16313 ( .A1(n14541), .A2(n14499), .ZN(n14313) );
  INV_X1 U16314 ( .A(n14304), .ZN(n14306) );
  AOI211_X1 U16315 ( .C1(n14543), .C2(n14306), .A(n14482), .B(n14305), .ZN(
        n14542) );
  INV_X1 U16316 ( .A(n14307), .ZN(n14308) );
  AOI22_X1 U16317 ( .A1(n14484), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14308), 
        .B2(n15760), .ZN(n14309) );
  OAI21_X1 U16318 ( .B1(n14310), .B2(n14486), .A(n14309), .ZN(n14311) );
  AOI21_X1 U16319 ( .B1(n14542), .B2(n14457), .A(n14311), .ZN(n14312) );
  OAI211_X1 U16320 ( .C1(n14465), .C2(n14629), .A(n14313), .B(n14312), .ZN(
        P2_U3243) );
  AOI21_X1 U16321 ( .B1(n14316), .B2(n14315), .A(n14314), .ZN(n14633) );
  XNOR2_X1 U16322 ( .A(n14317), .B(n14318), .ZN(n14320) );
  OAI21_X1 U16323 ( .B1(n14320), .B2(n14461), .A(n14319), .ZN(n14546) );
  NAND2_X1 U16324 ( .A1(n14546), .A2(n14499), .ZN(n14327) );
  NAND2_X1 U16325 ( .A1(n6610), .A2(n14548), .ZN(n14321) );
  NAND2_X1 U16326 ( .A1(n14321), .A2(n10957), .ZN(n14322) );
  NOR2_X1 U16327 ( .A1(n14304), .A2(n14322), .ZN(n14547) );
  AOI22_X1 U16328 ( .A1(n14484), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14323), 
        .B2(n15760), .ZN(n14324) );
  OAI21_X1 U16329 ( .B1(n7509), .B2(n14486), .A(n14324), .ZN(n14325) );
  AOI21_X1 U16330 ( .B1(n14547), .B2(n14457), .A(n14325), .ZN(n14326) );
  OAI211_X1 U16331 ( .C1(n14465), .C2(n14633), .A(n14327), .B(n14326), .ZN(
        P2_U3244) );
  OR2_X1 U16332 ( .A1(n14328), .A2(n14334), .ZN(n14329) );
  NAND2_X1 U16333 ( .A1(n14330), .A2(n14329), .ZN(n14637) );
  INV_X1 U16334 ( .A(n14331), .ZN(n14332) );
  AOI21_X1 U16335 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n14335) );
  OAI222_X1 U16336 ( .A1(n14471), .A2(n14337), .B1(n14473), .B2(n14336), .C1(
        n14335), .C2(n14461), .ZN(n14551) );
  NAND2_X1 U16337 ( .A1(n14551), .A2(n14499), .ZN(n14344) );
  AOI211_X1 U16338 ( .C1(n14553), .C2(n14338), .A(n14482), .B(n6786), .ZN(
        n14552) );
  AOI22_X1 U16339 ( .A1(n14484), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14339), 
        .B2(n15760), .ZN(n14340) );
  OAI21_X1 U16340 ( .B1(n14341), .B2(n14486), .A(n14340), .ZN(n14342) );
  AOI21_X1 U16341 ( .B1(n14552), .B2(n15767), .A(n14342), .ZN(n14343) );
  OAI211_X1 U16342 ( .C1(n14465), .C2(n14637), .A(n14344), .B(n14343), .ZN(
        P2_U3245) );
  NAND2_X1 U16343 ( .A1(n14346), .A2(n14345), .ZN(n14347) );
  XNOR2_X1 U16344 ( .A(n14347), .B(n14351), .ZN(n14355) );
  OAI22_X1 U16345 ( .A1(n14349), .A2(n14473), .B1(n14348), .B2(n14471), .ZN(
        n14354) );
  OAI21_X1 U16346 ( .B1(n14352), .B2(n14351), .A(n14350), .ZN(n14560) );
  NOR2_X1 U16347 ( .A1(n14560), .A2(n8920), .ZN(n14353) );
  AOI211_X1 U16348 ( .C1(n14355), .C2(n15757), .A(n14354), .B(n14353), .ZN(
        n14559) );
  INV_X1 U16349 ( .A(n14368), .ZN(n14357) );
  INV_X1 U16350 ( .A(n14338), .ZN(n14356) );
  AOI211_X1 U16351 ( .C1(n14557), .C2(n14357), .A(n14482), .B(n14356), .ZN(
        n14556) );
  INV_X1 U16352 ( .A(n14358), .ZN(n14359) );
  AOI22_X1 U16353 ( .A1(n14484), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14359), 
        .B2(n15760), .ZN(n14360) );
  OAI21_X1 U16354 ( .B1(n14361), .B2(n14486), .A(n14360), .ZN(n14363) );
  NOR2_X1 U16355 ( .A1(n14560), .A2(n14488), .ZN(n14362) );
  AOI211_X1 U16356 ( .C1(n14556), .C2(n15767), .A(n14363), .B(n14362), .ZN(
        n14364) );
  OAI21_X1 U16357 ( .B1(n14559), .B2(n14484), .A(n14364), .ZN(P2_U3246) );
  XNOR2_X1 U16358 ( .A(n14365), .B(n14376), .ZN(n14367) );
  AOI21_X1 U16359 ( .B1(n14367), .B2(n15757), .A(n14366), .ZN(n14564) );
  AOI211_X1 U16360 ( .C1(n14562), .C2(n14394), .A(n14482), .B(n14368), .ZN(
        n14561) );
  AOI22_X1 U16361 ( .A1(n14484), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14369), 
        .B2(n15760), .ZN(n14370) );
  OAI21_X1 U16362 ( .B1(n14371), .B2(n14486), .A(n14370), .ZN(n14379) );
  INV_X1 U16363 ( .A(n14373), .ZN(n14388) );
  NAND2_X1 U16364 ( .A1(n14372), .A2(n14388), .ZN(n14387) );
  INV_X1 U16365 ( .A(n14374), .ZN(n14375) );
  NAND2_X1 U16366 ( .A1(n14387), .A2(n14375), .ZN(n14377) );
  XNOR2_X1 U16367 ( .A(n14377), .B(n14376), .ZN(n14565) );
  NOR2_X1 U16368 ( .A1(n14565), .A2(n14465), .ZN(n14378) );
  AOI211_X1 U16369 ( .C1(n14561), .C2(n14457), .A(n14379), .B(n14378), .ZN(
        n14380) );
  OAI21_X1 U16370 ( .B1(n14484), .B2(n14564), .A(n14380), .ZN(P2_U3247) );
  NAND3_X1 U16371 ( .A1(n14381), .A2(n14388), .A3(n14382), .ZN(n14383) );
  NAND3_X1 U16372 ( .A1(n14384), .A2(n15757), .A3(n14383), .ZN(n14386) );
  NAND2_X1 U16373 ( .A1(n14386), .A2(n14385), .ZN(n14566) );
  OAI21_X1 U16374 ( .B1(n14372), .B2(n14388), .A(n14387), .ZN(n14643) );
  NAND2_X1 U16375 ( .A1(n14484), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14389) );
  OAI21_X1 U16376 ( .B1(n14406), .B2(n14390), .A(n14389), .ZN(n14391) );
  AOI21_X1 U16377 ( .B1(n14568), .B2(n15759), .A(n14391), .ZN(n14396) );
  AOI21_X1 U16378 ( .B1(n14405), .B2(n14568), .A(n14482), .ZN(n14393) );
  AND2_X1 U16379 ( .A1(n14394), .A2(n14393), .ZN(n14567) );
  NAND2_X1 U16380 ( .A1(n14567), .A2(n14457), .ZN(n14395) );
  OAI211_X1 U16381 ( .C1(n14643), .C2(n14465), .A(n14396), .B(n14395), .ZN(
        n14397) );
  AOI21_X1 U16382 ( .B1(n14499), .B2(n14566), .A(n14397), .ZN(n14398) );
  INV_X1 U16383 ( .A(n14398), .ZN(P2_U3248) );
  INV_X1 U16384 ( .A(n14400), .ZN(n14402) );
  AOI21_X1 U16385 ( .B1(n14399), .B2(n14402), .A(n14401), .ZN(n14417) );
  NAND2_X1 U16386 ( .A1(n14417), .A2(n14430), .ZN(n14416) );
  NAND2_X1 U16387 ( .A1(n14416), .A2(n14403), .ZN(n14404) );
  XNOR2_X1 U16388 ( .A(n14404), .B(n14410), .ZN(n14575) );
  AOI211_X1 U16389 ( .C1(n14573), .C2(n14420), .A(n14482), .B(n14392), .ZN(
        n14572) );
  NOR2_X1 U16390 ( .A1(n7518), .A2(n14486), .ZN(n14409) );
  OAI22_X1 U16391 ( .A1(n14499), .A2(n11961), .B1(n14407), .B2(n14406), .ZN(
        n14408) );
  AOI211_X1 U16392 ( .C1(n14572), .C2(n15767), .A(n14409), .B(n14408), .ZN(
        n14415) );
  OAI211_X1 U16393 ( .C1(n14411), .C2(n14410), .A(n14381), .B(n15757), .ZN(
        n14413) );
  NAND2_X1 U16394 ( .A1(n14413), .A2(n14412), .ZN(n14571) );
  NAND2_X1 U16395 ( .A1(n14571), .A2(n14499), .ZN(n14414) );
  OAI211_X1 U16396 ( .C1(n14575), .C2(n14465), .A(n14415), .B(n14414), .ZN(
        P2_U3249) );
  OAI21_X1 U16397 ( .B1(n14417), .B2(n14430), .A(n14416), .ZN(n14418) );
  INV_X1 U16398 ( .A(n14418), .ZN(n14580) );
  INV_X1 U16399 ( .A(n14419), .ZN(n14422) );
  INV_X1 U16400 ( .A(n14420), .ZN(n14421) );
  AOI211_X1 U16401 ( .C1(n14578), .C2(n14422), .A(n14482), .B(n14421), .ZN(
        n14577) );
  AOI22_X1 U16402 ( .A1(n14484), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14423), 
        .B2(n15760), .ZN(n14424) );
  OAI21_X1 U16403 ( .B1(n14425), .B2(n14486), .A(n14424), .ZN(n14426) );
  AOI21_X1 U16404 ( .B1(n14577), .B2(n15767), .A(n14426), .ZN(n14434) );
  INV_X1 U16405 ( .A(n14428), .ZN(n14429) );
  AOI21_X1 U16406 ( .B1(n14430), .B2(n14427), .A(n14429), .ZN(n14432) );
  OAI21_X1 U16407 ( .B1(n14432), .B2(n14461), .A(n14431), .ZN(n14576) );
  NAND2_X1 U16408 ( .A1(n14576), .A2(n14499), .ZN(n14433) );
  OAI211_X1 U16409 ( .C1(n14580), .C2(n14465), .A(n14434), .B(n14433), .ZN(
        P2_U3250) );
  INV_X1 U16410 ( .A(n14399), .ZN(n14449) );
  NAND2_X1 U16411 ( .A1(n14449), .A2(n14459), .ZN(n14448) );
  NAND2_X1 U16412 ( .A1(n14448), .A2(n14435), .ZN(n14436) );
  XOR2_X1 U16413 ( .A(n14438), .B(n14436), .Z(n14650) );
  XNOR2_X1 U16414 ( .A(n14437), .B(n14438), .ZN(n14440) );
  OAI21_X1 U16415 ( .B1(n14440), .B2(n14461), .A(n14439), .ZN(n14581) );
  INV_X1 U16416 ( .A(n14452), .ZN(n14441) );
  AOI211_X1 U16417 ( .C1(n14583), .C2(n14441), .A(n14482), .B(n14419), .ZN(
        n14582) );
  NAND2_X1 U16418 ( .A1(n14582), .A2(n15767), .ZN(n14444) );
  AOI22_X1 U16419 ( .A1(n14484), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14442), 
        .B2(n15760), .ZN(n14443) );
  OAI211_X1 U16420 ( .C1(n14445), .C2(n14486), .A(n14444), .B(n14443), .ZN(
        n14446) );
  AOI21_X1 U16421 ( .B1(n14499), .B2(n14581), .A(n14446), .ZN(n14447) );
  OAI21_X1 U16422 ( .B1(n14650), .B2(n14465), .A(n14447), .ZN(P2_U3251) );
  OAI21_X1 U16423 ( .B1(n14449), .B2(n14459), .A(n14448), .ZN(n14651) );
  INV_X1 U16424 ( .A(n14651), .ZN(n14466) );
  NAND2_X1 U16425 ( .A1(n14481), .A2(n14589), .ZN(n14450) );
  NAND2_X1 U16426 ( .A1(n14450), .A2(n10957), .ZN(n14451) );
  NOR2_X1 U16427 ( .A1(n14452), .A2(n14451), .ZN(n14588) );
  AOI22_X1 U16428 ( .A1(n14484), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14453), 
        .B2(n15760), .ZN(n14454) );
  OAI21_X1 U16429 ( .B1(n14455), .B2(n14486), .A(n14454), .ZN(n14456) );
  AOI21_X1 U16430 ( .B1(n14588), .B2(n14457), .A(n14456), .ZN(n14464) );
  XOR2_X1 U16431 ( .A(n14458), .B(n14459), .Z(n14462) );
  OAI21_X1 U16432 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n14587) );
  NAND2_X1 U16433 ( .A1(n14587), .A2(n14499), .ZN(n14463) );
  OAI211_X1 U16434 ( .C1(n14466), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        P2_U3252) );
  NAND2_X1 U16435 ( .A1(n14468), .A2(n14467), .ZN(n14493) );
  NAND2_X1 U16436 ( .A1(n14493), .A2(n14503), .ZN(n14492) );
  NAND2_X1 U16437 ( .A1(n14492), .A2(n14469), .ZN(n14470) );
  XOR2_X1 U16438 ( .A(n14470), .B(n14475), .Z(n14479) );
  OAI22_X1 U16439 ( .A1(n14474), .A2(n14473), .B1(n14472), .B2(n14471), .ZN(
        n14478) );
  XNOR2_X1 U16440 ( .A(n14476), .B(n14475), .ZN(n14596) );
  NOR2_X1 U16441 ( .A1(n14596), .A2(n8920), .ZN(n14477) );
  AOI211_X1 U16442 ( .C1(n15757), .C2(n14479), .A(n14478), .B(n14477), .ZN(
        n14595) );
  AOI211_X1 U16443 ( .C1(n14593), .C2(n14480), .A(n14482), .B(n7516), .ZN(
        n14592) );
  INV_X1 U16444 ( .A(n14593), .ZN(n14487) );
  AOI22_X1 U16445 ( .A1(n14484), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n14483), 
        .B2(n15760), .ZN(n14485) );
  OAI21_X1 U16446 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14490) );
  NOR2_X1 U16447 ( .A1(n14596), .A2(n14488), .ZN(n14489) );
  AOI211_X1 U16448 ( .C1(n14592), .C2(n14457), .A(n14490), .B(n14489), .ZN(
        n14491) );
  OAI21_X1 U16449 ( .B1(n14595), .B2(n14484), .A(n14491), .ZN(P2_U3253) );
  OAI21_X1 U16450 ( .B1(n14493), .B2(n14503), .A(n14492), .ZN(n14498) );
  AOI222_X1 U16451 ( .A1(n14498), .A2(n15757), .B1(n14497), .B2(n14496), .C1(
        n14495), .C2(n14494), .ZN(n14602) );
  MUX2_X1 U16452 ( .A(n14500), .B(n14602), .S(n14499), .Z(n14511) );
  AOI22_X1 U16453 ( .A1(n15759), .A2(n14598), .B1(n15760), .B2(n14501), .ZN(
        n14510) );
  NAND2_X1 U16454 ( .A1(n14504), .A2(n14503), .ZN(n14597) );
  NAND3_X1 U16455 ( .A1(n14502), .A2(n14597), .A3(n15768), .ZN(n14509) );
  OAI211_X1 U16456 ( .C1(n14506), .C2(n14505), .A(n10957), .B(n14480), .ZN(
        n14599) );
  OR2_X1 U16457 ( .A1(n14599), .A2(n14507), .ZN(n14508) );
  NAND4_X1 U16458 ( .A1(n14511), .A2(n14510), .A3(n14509), .A4(n14508), .ZN(
        P2_U3254) );
  OAI211_X1 U16459 ( .C1(n14513), .C2(n15843), .A(n14512), .B(n14514), .ZN(
        n14608) );
  MUX2_X1 U16460 ( .A(n14608), .B(P2_REG1_REG_31__SCAN_IN), .S(n8995), .Z(
        P2_U3530) );
  INV_X1 U16461 ( .A(n14516), .ZN(n14517) );
  MUX2_X1 U16462 ( .A(n14609), .B(P2_REG1_REG_30__SCAN_IN), .S(n8995), .Z(
        P2_U3529) );
  INV_X1 U16463 ( .A(n14586), .ZN(n14590) );
  AND2_X1 U16464 ( .A1(n14519), .A2(n15835), .ZN(n14521) );
  MUX2_X1 U16465 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14611), .S(n15864), .Z(
        n14523) );
  INV_X1 U16466 ( .A(n14524), .ZN(n14617) );
  INV_X1 U16467 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14528) );
  MUX2_X1 U16468 ( .A(n14528), .B(n14614), .S(n15864), .Z(n14529) );
  OAI21_X1 U16469 ( .B1(n14586), .B2(n14617), .A(n14529), .ZN(P2_U3524) );
  INV_X1 U16470 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14533) );
  AOI211_X1 U16471 ( .C1(n15835), .C2(n14532), .A(n14531), .B(n14530), .ZN(
        n14618) );
  MUX2_X1 U16472 ( .A(n14533), .B(n14618), .S(n15864), .Z(n14534) );
  OAI21_X1 U16473 ( .B1(n14586), .B2(n14621), .A(n14534), .ZN(P2_U3523) );
  INV_X1 U16474 ( .A(n14535), .ZN(n14625) );
  INV_X1 U16475 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14539) );
  MUX2_X1 U16476 ( .A(n14539), .B(n14622), .S(n15864), .Z(n14540) );
  OAI21_X1 U16477 ( .B1(n14625), .B2(n14586), .A(n14540), .ZN(P2_U3522) );
  AOI211_X1 U16478 ( .C1(n15835), .C2(n14543), .A(n14542), .B(n14541), .ZN(
        n14626) );
  MUX2_X1 U16479 ( .A(n14544), .B(n14626), .S(n15864), .Z(n14545) );
  OAI21_X1 U16480 ( .B1(n14586), .B2(n14629), .A(n14545), .ZN(P2_U3521) );
  AOI211_X1 U16481 ( .C1(n15835), .C2(n14548), .A(n14547), .B(n14546), .ZN(
        n14630) );
  MUX2_X1 U16482 ( .A(n14549), .B(n14630), .S(n15864), .Z(n14550) );
  OAI21_X1 U16483 ( .B1(n14633), .B2(n14586), .A(n14550), .ZN(P2_U3520) );
  INV_X1 U16484 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14554) );
  AOI211_X1 U16485 ( .C1(n15835), .C2(n14553), .A(n14552), .B(n14551), .ZN(
        n14634) );
  MUX2_X1 U16486 ( .A(n14554), .B(n14634), .S(n15864), .Z(n14555) );
  OAI21_X1 U16487 ( .B1(n14586), .B2(n14637), .A(n14555), .ZN(P2_U3519) );
  AOI21_X1 U16488 ( .B1(n15835), .B2(n14557), .A(n14556), .ZN(n14558) );
  OAI211_X1 U16489 ( .C1(n15808), .C2(n14560), .A(n14559), .B(n14558), .ZN(
        n14638) );
  MUX2_X1 U16490 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14638), .S(n15864), .Z(
        P2_U3518) );
  AOI21_X1 U16491 ( .B1(n15835), .B2(n14562), .A(n14561), .ZN(n14563) );
  OAI211_X1 U16492 ( .C1(n10269), .C2(n14565), .A(n14564), .B(n14563), .ZN(
        n14639) );
  MUX2_X1 U16493 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14639), .S(n15864), .Z(
        P2_U3517) );
  AOI211_X1 U16494 ( .C1(n15835), .C2(n14568), .A(n14567), .B(n14566), .ZN(
        n14640) );
  MUX2_X1 U16495 ( .A(n14569), .B(n14640), .S(n15864), .Z(n14570) );
  OAI21_X1 U16496 ( .B1(n14586), .B2(n14643), .A(n14570), .ZN(P2_U3516) );
  AOI211_X1 U16497 ( .C1(n15835), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14574) );
  OAI21_X1 U16498 ( .B1(n10269), .B2(n14575), .A(n14574), .ZN(n14644) );
  MUX2_X1 U16499 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14644), .S(n15864), .Z(
        P2_U3515) );
  AOI211_X1 U16500 ( .C1(n15835), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        n14579) );
  OAI21_X1 U16501 ( .B1(n10269), .B2(n14580), .A(n14579), .ZN(n14645) );
  MUX2_X1 U16502 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14645), .S(n15864), .Z(
        P2_U3514) );
  AOI211_X1 U16503 ( .C1(n15835), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14646) );
  MUX2_X1 U16504 ( .A(n14584), .B(n14646), .S(n15864), .Z(n14585) );
  OAI21_X1 U16505 ( .B1(n14650), .B2(n14586), .A(n14585), .ZN(P2_U3513) );
  AOI211_X1 U16506 ( .C1(n15835), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14653) );
  AOI22_X1 U16507 ( .A1(n14651), .A2(n14590), .B1(P2_REG1_REG_13__SCAN_IN), 
        .B2(n8995), .ZN(n14591) );
  OAI21_X1 U16508 ( .B1(n14653), .B2(n8995), .A(n14591), .ZN(P2_U3512) );
  AOI21_X1 U16509 ( .B1(n15835), .B2(n14593), .A(n14592), .ZN(n14594) );
  OAI211_X1 U16510 ( .C1(n14596), .C2(n15808), .A(n14595), .B(n14594), .ZN(
        n14654) );
  MUX2_X1 U16511 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14654), .S(n15864), .Z(
        P2_U3511) );
  NAND3_X1 U16512 ( .A1(n14502), .A2(n15797), .A3(n14597), .ZN(n14601) );
  NAND2_X1 U16513 ( .A1(n14598), .A2(n15835), .ZN(n14600) );
  NAND4_X1 U16514 ( .A1(n14602), .A2(n14601), .A3(n14600), .A4(n14599), .ZN(
        n14655) );
  MUX2_X1 U16515 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14655), .S(n15864), .Z(
        P2_U3510) );
  AOI21_X1 U16516 ( .B1(n15835), .B2(n14604), .A(n14603), .ZN(n14605) );
  OAI211_X1 U16517 ( .C1(n15808), .C2(n14607), .A(n14606), .B(n14605), .ZN(
        n14656) );
  MUX2_X1 U16518 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14656), .S(n15864), .Z(
        P2_U3508) );
  MUX2_X1 U16519 ( .A(n14608), .B(P2_REG0_REG_31__SCAN_IN), .S(n9003), .Z(
        P2_U3498) );
  MUX2_X1 U16520 ( .A(n14609), .B(P2_REG0_REG_30__SCAN_IN), .S(n9003), .Z(
        P2_U3497) );
  MUX2_X1 U16521 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14610), .S(n15850), .Z(
        P2_U3494) );
  MUX2_X1 U16522 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14611), .S(n15850), .Z(
        n14612) );
  INV_X1 U16523 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14615) );
  MUX2_X1 U16524 ( .A(n14615), .B(n14614), .S(n15850), .Z(n14616) );
  OAI21_X1 U16525 ( .B1(n14617), .B2(n14649), .A(n14616), .ZN(P2_U3492) );
  INV_X1 U16526 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14619) );
  MUX2_X1 U16527 ( .A(n14619), .B(n14618), .S(n15850), .Z(n14620) );
  OAI21_X1 U16528 ( .B1(n14621), .B2(n14649), .A(n14620), .ZN(P2_U3491) );
  INV_X1 U16529 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14623) );
  MUX2_X1 U16530 ( .A(n14623), .B(n14622), .S(n15850), .Z(n14624) );
  OAI21_X1 U16531 ( .B1(n14625), .B2(n14649), .A(n14624), .ZN(P2_U3490) );
  INV_X1 U16532 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14627) );
  MUX2_X1 U16533 ( .A(n14627), .B(n14626), .S(n15850), .Z(n14628) );
  OAI21_X1 U16534 ( .B1(n14629), .B2(n14649), .A(n14628), .ZN(P2_U3489) );
  INV_X1 U16535 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14631) );
  MUX2_X1 U16536 ( .A(n14631), .B(n14630), .S(n15850), .Z(n14632) );
  OAI21_X1 U16537 ( .B1(n14633), .B2(n14649), .A(n14632), .ZN(P2_U3488) );
  INV_X1 U16538 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14635) );
  MUX2_X1 U16539 ( .A(n14635), .B(n14634), .S(n15850), .Z(n14636) );
  OAI21_X1 U16540 ( .B1(n14637), .B2(n14649), .A(n14636), .ZN(P2_U3487) );
  MUX2_X1 U16541 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14638), .S(n15850), .Z(
        P2_U3486) );
  MUX2_X1 U16542 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14639), .S(n15850), .Z(
        P2_U3484) );
  INV_X1 U16543 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14641) );
  MUX2_X1 U16544 ( .A(n14641), .B(n14640), .S(n15850), .Z(n14642) );
  OAI21_X1 U16545 ( .B1(n14643), .B2(n14649), .A(n14642), .ZN(P2_U3481) );
  MUX2_X1 U16546 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14644), .S(n15850), .Z(
        P2_U3478) );
  MUX2_X1 U16547 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14645), .S(n15850), .Z(
        P2_U3475) );
  INV_X1 U16548 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14647) );
  MUX2_X1 U16549 ( .A(n14647), .B(n14646), .S(n15850), .Z(n14648) );
  OAI21_X1 U16550 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(P2_U3472) );
  AOI22_X1 U16551 ( .A1(n14651), .A2(n9001), .B1(P2_REG0_REG_13__SCAN_IN), 
        .B2(n9003), .ZN(n14652) );
  OAI21_X1 U16552 ( .B1(n14653), .B2(n9003), .A(n14652), .ZN(P2_U3469) );
  MUX2_X1 U16553 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14654), .S(n15850), .Z(
        P2_U3466) );
  MUX2_X1 U16554 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14655), .S(n15850), .Z(
        P2_U3463) );
  MUX2_X1 U16555 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14656), .S(n15850), .Z(
        P2_U3457) );
  INV_X1 U16556 ( .A(n14657), .ZN(n15424) );
  NAND3_X1 U16557 ( .A1(n14658), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14661) );
  OAI22_X1 U16558 ( .A1(n8514), .A2(n14661), .B1(n14660), .B2(n14659), .ZN(
        n14662) );
  INV_X1 U16559 ( .A(n14662), .ZN(n14663) );
  OAI21_X1 U16560 ( .B1(n15424), .B2(n11978), .A(n14663), .ZN(P2_U3296) );
  INV_X1 U16561 ( .A(n14664), .ZN(n15431) );
  AOI21_X1 U16562 ( .B1(n14666), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14665), 
        .ZN(n14667) );
  OAI21_X1 U16563 ( .B1(n15431), .B2(n11978), .A(n14667), .ZN(P2_U3299) );
  MUX2_X1 U16564 ( .A(n14668), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16565 ( .A(n14669), .B(n6658), .Z(n14676) );
  AOI21_X1 U16566 ( .B1(n14779), .B2(n15344), .A(n14670), .ZN(n14672) );
  NAND2_X1 U16567 ( .A1(n14813), .A2(n15193), .ZN(n14671) );
  OAI211_X1 U16568 ( .C1(n14673), .C2(n14798), .A(n14672), .B(n14671), .ZN(
        n14674) );
  AOI21_X1 U16569 ( .B1(n15211), .B2(n14769), .A(n14674), .ZN(n14675) );
  OAI21_X1 U16570 ( .B1(n14676), .B2(n14815), .A(n14675), .ZN(P1_U3215) );
  XNOR2_X1 U16571 ( .A(n14678), .B(n14681), .ZN(n14701) );
  NAND2_X1 U16572 ( .A1(n14677), .A2(n14701), .ZN(n14774) );
  XNOR2_X1 U16573 ( .A(n14680), .B(n14679), .ZN(n14776) );
  NAND2_X1 U16574 ( .A1(n14682), .A2(n14681), .ZN(n14773) );
  AND2_X1 U16575 ( .A1(n14683), .A2(n14742), .ZN(n14684) );
  AOI21_X1 U16576 ( .B1(n14775), .B2(n14685), .A(n14684), .ZN(n14686) );
  OAI21_X1 U16577 ( .B1(n14745), .B2(n14686), .A(n15491), .ZN(n14692) );
  NOR2_X1 U16578 ( .A1(n15058), .A2(n15495), .ZN(n14690) );
  OAI22_X1 U16579 ( .A1(n14688), .A2(n14808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14687), .ZN(n14689) );
  AOI211_X1 U16580 ( .C1(n14806), .C2(n15294), .A(n14690), .B(n14689), .ZN(
        n14691) );
  OAI211_X1 U16581 ( .C1(n15285), .C2(n14809), .A(n14692), .B(n14691), .ZN(
        P1_U3216) );
  AND2_X1 U16582 ( .A1(n14784), .A2(n14693), .ZN(n14696) );
  OAI211_X1 U16583 ( .C1(n14696), .C2(n14695), .A(n15491), .B(n14694), .ZN(
        n14700) );
  NOR2_X1 U16584 ( .A1(n15495), .A2(n15125), .ZN(n14698) );
  NAND2_X1 U16585 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14966)
         );
  OAI21_X1 U16586 ( .B1(n14808), .B2(n15129), .A(n14966), .ZN(n14697) );
  AOI211_X1 U16587 ( .C1(n14806), .C2(n15305), .A(n14698), .B(n14697), .ZN(
        n14699) );
  OAI211_X1 U16588 ( .C1(n15309), .C2(n14809), .A(n14700), .B(n14699), .ZN(
        P1_U3219) );
  OAI21_X1 U16589 ( .B1(n14677), .B2(n14701), .A(n14774), .ZN(n14702) );
  NAND2_X1 U16590 ( .A1(n14702), .A2(n15491), .ZN(n14707) );
  NOR2_X1 U16591 ( .A1(n15085), .A2(n15495), .ZN(n14705) );
  OAI22_X1 U16592 ( .A1(n15089), .A2(n14808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14703), .ZN(n14704) );
  AOI211_X1 U16593 ( .C1(n14806), .C2(n15306), .A(n14705), .B(n14704), .ZN(
        n14706) );
  OAI211_X1 U16594 ( .C1(n7436), .C2(n14809), .A(n14707), .B(n14706), .ZN(
        P1_U3223) );
  INV_X1 U16595 ( .A(n14708), .ZN(n14746) );
  INV_X1 U16596 ( .A(n14709), .ZN(n14711) );
  NOR3_X1 U16597 ( .A1(n14746), .A2(n14711), .A3(n14710), .ZN(n14714) );
  INV_X1 U16598 ( .A(n14712), .ZN(n14713) );
  OAI21_X1 U16599 ( .B1(n14714), .B2(n14713), .A(n15491), .ZN(n14718) );
  AOI22_X1 U16600 ( .A1(n15057), .A2(n14806), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14715) );
  OAI21_X1 U16601 ( .B1(n15029), .B2(n15495), .A(n14715), .ZN(n14716) );
  AOI21_X1 U16602 ( .B1(n14779), .B2(n15028), .A(n14716), .ZN(n14717) );
  OAI211_X1 U16603 ( .C1(n15267), .C2(n14809), .A(n14718), .B(n14717), .ZN(
        P1_U3225) );
  XNOR2_X1 U16604 ( .A(n14720), .B(n14721), .ZN(n14805) );
  INV_X1 U16605 ( .A(n14719), .ZN(n14804) );
  NOR2_X1 U16606 ( .A1(n14805), .A2(n14804), .ZN(n14803) );
  AOI21_X1 U16607 ( .B1(n14721), .B2(n14720), .A(n14803), .ZN(n14725) );
  XNOR2_X1 U16608 ( .A(n14723), .B(n14722), .ZN(n14724) );
  XNOR2_X1 U16609 ( .A(n14725), .B(n14724), .ZN(n14731) );
  OAI21_X1 U16610 ( .B1(n14808), .B2(n15181), .A(n14726), .ZN(n14727) );
  AOI21_X1 U16611 ( .B1(n14806), .B2(n15344), .A(n14727), .ZN(n14728) );
  OAI21_X1 U16612 ( .B1(n15176), .B2(n15495), .A(n14728), .ZN(n14729) );
  AOI21_X1 U16613 ( .B1(n15183), .B2(n14769), .A(n14729), .ZN(n14730) );
  OAI21_X1 U16614 ( .B1(n14731), .B2(n14815), .A(n14730), .ZN(P1_U3226) );
  XNOR2_X1 U16615 ( .A(n14734), .B(n14733), .ZN(n14735) );
  XNOR2_X1 U16616 ( .A(n14732), .B(n14735), .ZN(n14741) );
  NOR2_X1 U16617 ( .A1(n14736), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14937) );
  AOI21_X1 U16618 ( .B1(n14779), .B2(n15305), .A(n14937), .ZN(n14738) );
  NAND2_X1 U16619 ( .A1(n14813), .A2(n15159), .ZN(n14737) );
  OAI211_X1 U16620 ( .C1(n15321), .C2(n14798), .A(n14738), .B(n14737), .ZN(
        n14739) );
  AOI21_X1 U16621 ( .B1(n15325), .B2(n14769), .A(n14739), .ZN(n14740) );
  OAI21_X1 U16622 ( .B1(n14741), .B2(n14815), .A(n14740), .ZN(P1_U3228) );
  INV_X1 U16623 ( .A(n14742), .ZN(n14744) );
  NOR3_X1 U16624 ( .A1(n14745), .A2(n14744), .A3(n14743), .ZN(n14747) );
  AOI22_X1 U16625 ( .A1(n15015), .A2(n14779), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14748) );
  OAI21_X1 U16626 ( .B1(n15273), .B2(n14798), .A(n14748), .ZN(n14749) );
  AOI21_X1 U16627 ( .B1(n15044), .B2(n14813), .A(n14749), .ZN(n14750) );
  OAI211_X1 U16628 ( .C1(n14752), .C2(n14809), .A(n14751), .B(n14750), .ZN(
        P1_U3229) );
  XNOR2_X1 U16629 ( .A(n14754), .B(n14753), .ZN(n14760) );
  OAI22_X1 U16630 ( .A1(n15098), .A2(n14808), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14755), .ZN(n14756) );
  AOI21_X1 U16631 ( .B1(n14806), .B2(n15145), .A(n14756), .ZN(n14757) );
  OAI21_X1 U16632 ( .B1(n15104), .B2(n15495), .A(n14757), .ZN(n14758) );
  AOI21_X1 U16633 ( .B1(n10129), .B2(n14769), .A(n14758), .ZN(n14759) );
  OAI21_X1 U16634 ( .B1(n14760), .B2(n14815), .A(n14759), .ZN(P1_U3233) );
  AOI21_X1 U16635 ( .B1(n14763), .B2(n14762), .A(n14761), .ZN(n14772) );
  NAND2_X1 U16636 ( .A1(n14806), .A2(n15353), .ZN(n14765) );
  OAI211_X1 U16637 ( .C1(n14808), .C2(n14766), .A(n14765), .B(n14764), .ZN(
        n14767) );
  AOI21_X1 U16638 ( .B1(n14768), .B2(n14813), .A(n14767), .ZN(n14771) );
  NAND2_X1 U16639 ( .A1(n15352), .A2(n14769), .ZN(n14770) );
  OAI211_X1 U16640 ( .C1(n14772), .C2(n14815), .A(n14771), .B(n14770), .ZN(
        P1_U3234) );
  AND2_X1 U16641 ( .A1(n14774), .A2(n14773), .ZN(n14777) );
  OAI211_X1 U16642 ( .C1(n14777), .C2(n14776), .A(n15491), .B(n14775), .ZN(
        n14783) );
  INV_X1 U16643 ( .A(n14778), .ZN(n15074) );
  AOI22_X1 U16644 ( .A1(n15045), .A2(n14779), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14780) );
  OAI21_X1 U16645 ( .B1(n15098), .B2(n14798), .A(n14780), .ZN(n14781) );
  AOI21_X1 U16646 ( .B1(n15074), .B2(n14813), .A(n14781), .ZN(n14782) );
  OAI211_X1 U16647 ( .C1(n14809), .C2(n15076), .A(n14783), .B(n14782), .ZN(
        P1_U3235) );
  OAI21_X1 U16648 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(n14787) );
  NAND2_X1 U16649 ( .A1(n14787), .A2(n15491), .ZN(n14792) );
  NAND2_X1 U16650 ( .A1(n14806), .A2(n15329), .ZN(n14789) );
  OAI211_X1 U16651 ( .C1(n14808), .C2(n15314), .A(n14789), .B(n14788), .ZN(
        n14790) );
  AOI21_X1 U16652 ( .B1(n15144), .B2(n14813), .A(n14790), .ZN(n14791) );
  OAI211_X1 U16653 ( .C1(n15315), .C2(n14809), .A(n14792), .B(n14791), .ZN(
        P1_U3238) );
  OAI21_X1 U16654 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14796) );
  NAND2_X1 U16655 ( .A1(n14796), .A2(n15491), .ZN(n14802) );
  OAI22_X1 U16656 ( .A1(n15274), .A2(n14798), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14797), .ZN(n14800) );
  NOR2_X1 U16657 ( .A1(n15242), .A2(n14808), .ZN(n14799) );
  AOI211_X1 U16658 ( .C1(n14813), .C2(n15017), .A(n14800), .B(n14799), .ZN(
        n14801) );
  OAI211_X1 U16659 ( .C1(n15261), .C2(n14809), .A(n14802), .B(n14801), .ZN(
        P1_U3240) );
  AOI21_X1 U16660 ( .B1(n14805), .B2(n14804), .A(n14803), .ZN(n14816) );
  NAND2_X1 U16661 ( .A1(n14806), .A2(n15354), .ZN(n14807) );
  NAND2_X1 U16662 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15507)
         );
  OAI211_X1 U16663 ( .C1(n14808), .C2(n15321), .A(n14807), .B(n15507), .ZN(
        n14811) );
  NOR2_X1 U16664 ( .A1(n15339), .A2(n14809), .ZN(n14810) );
  AOI211_X1 U16665 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  OAI21_X1 U16666 ( .B1(n14816), .B2(n14815), .A(n14814), .ZN(P1_U3241) );
  MUX2_X1 U16667 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14971), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16668 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14817), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16669 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14988), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16670 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15223), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16671 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15016), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16672 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15028), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16673 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15015), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16674 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15057), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16675 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15045), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16676 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15294), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16677 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14818), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16678 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15306), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16679 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15145), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16680 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15305), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16681 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15329), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16682 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14819), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16683 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15344), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16684 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15354), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16685 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15363), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16686 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15353), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16687 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15362), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16688 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14820), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16689 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14821), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16690 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15514), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16691 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15667), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16692 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15531), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16693 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15666), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16694 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15532), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16695 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15647), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16696 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15562), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16697 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15566), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16698 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15567), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16699 ( .A1(n15509), .A2(n14823), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14822), .ZN(n14824) );
  AOI21_X1 U16700 ( .B1(n14825), .B2(n15501), .A(n14824), .ZN(n14831) );
  NAND2_X1 U16701 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14833) );
  OAI211_X1 U16702 ( .C1(n10714), .C2(n14826), .A(n15505), .B(n14847), .ZN(
        n14830) );
  OAI211_X1 U16703 ( .C1(n14828), .C2(n14827), .A(n15504), .B(n14841), .ZN(
        n14829) );
  NAND3_X1 U16704 ( .A1(n14831), .A2(n14830), .A3(n14829), .ZN(P1_U3244) );
  MUX2_X1 U16705 ( .A(n14834), .B(n14833), .S(n14832), .Z(n14837) );
  NAND2_X1 U16706 ( .A1(n14835), .A2(n7559), .ZN(n14836) );
  OAI211_X1 U16707 ( .C1(n14837), .C2(n15430), .A(P1_U4016), .B(n14836), .ZN(
        n14882) );
  OAI22_X1 U16708 ( .A1(n15509), .A2(n10013), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14838), .ZN(n14839) );
  AOI21_X1 U16709 ( .B1(n14844), .B2(n15501), .A(n14839), .ZN(n14852) );
  MUX2_X1 U16710 ( .A(n10685), .B(P1_REG1_REG_2__SCAN_IN), .S(n14844), .Z(
        n14842) );
  NAND3_X1 U16711 ( .A1(n14842), .A2(n14841), .A3(n14840), .ZN(n14843) );
  NAND3_X1 U16712 ( .A1(n15504), .A2(n14861), .A3(n14843), .ZN(n14851) );
  MUX2_X1 U16713 ( .A(n14845), .B(P1_REG2_REG_2__SCAN_IN), .S(n14844), .Z(
        n14848) );
  NAND3_X1 U16714 ( .A1(n14848), .A2(n14847), .A3(n14846), .ZN(n14849) );
  NAND3_X1 U16715 ( .A1(n15505), .A2(n14856), .A3(n14849), .ZN(n14850) );
  NAND4_X1 U16716 ( .A1(n14882), .A2(n14852), .A3(n14851), .A4(n14850), .ZN(
        P1_U3245) );
  AND2_X1 U16717 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15482) );
  NOR2_X1 U16718 ( .A1(n14957), .A2(n14859), .ZN(n14854) );
  AOI211_X1 U16719 ( .C1(n14938), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n15482), .B(
        n14854), .ZN(n14866) );
  MUX2_X1 U16720 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10717), .S(n14859), .Z(
        n14857) );
  NAND3_X1 U16721 ( .A1(n14857), .A2(n14856), .A3(n14855), .ZN(n14858) );
  NAND3_X1 U16722 ( .A1(n15505), .A2(n14871), .A3(n14858), .ZN(n14865) );
  MUX2_X1 U16723 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n15703), .S(n14859), .Z(
        n14862) );
  NAND3_X1 U16724 ( .A1(n14862), .A2(n14861), .A3(n14860), .ZN(n14863) );
  NAND3_X1 U16725 ( .A1(n15504), .A2(n14876), .A3(n14863), .ZN(n14864) );
  NAND3_X1 U16726 ( .A1(n14866), .A2(n14865), .A3(n14864), .ZN(P1_U3246) );
  NOR2_X1 U16727 ( .A1(n14957), .A2(n14873), .ZN(n14867) );
  AOI211_X1 U16728 ( .C1(n14938), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n14868), .B(
        n14867), .ZN(n14881) );
  MUX2_X1 U16729 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10720), .S(n14873), .Z(
        n14869) );
  NAND3_X1 U16730 ( .A1(n14871), .A2(n14870), .A3(n14869), .ZN(n14872) );
  NAND3_X1 U16731 ( .A1(n15505), .A2(n14889), .A3(n14872), .ZN(n14880) );
  MUX2_X1 U16732 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10691), .S(n14873), .Z(
        n14874) );
  NAND3_X1 U16733 ( .A1(n14876), .A2(n14875), .A3(n14874), .ZN(n14877) );
  NAND3_X1 U16734 ( .A1(n15504), .A2(n14878), .A3(n14877), .ZN(n14879) );
  NAND4_X1 U16735 ( .A1(n14882), .A2(n14881), .A3(n14880), .A4(n14879), .ZN(
        P1_U3247) );
  OAI21_X1 U16736 ( .B1(n15509), .B2(n10045), .A(n14883), .ZN(n14884) );
  AOI21_X1 U16737 ( .B1(n14885), .B2(n15501), .A(n14884), .ZN(n14898) );
  MUX2_X1 U16738 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10723), .S(n14886), .Z(
        n14887) );
  NAND3_X1 U16739 ( .A1(n14889), .A2(n14888), .A3(n14887), .ZN(n14890) );
  NAND3_X1 U16740 ( .A1(n15505), .A2(n14891), .A3(n14890), .ZN(n14897) );
  OAI21_X1 U16741 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(n14895) );
  NAND2_X1 U16742 ( .A1(n15504), .A2(n14895), .ZN(n14896) );
  NAND3_X1 U16743 ( .A1(n14898), .A2(n14897), .A3(n14896), .ZN(P1_U3248) );
  INV_X1 U16744 ( .A(n14908), .ZN(n14902) );
  OAI21_X1 U16745 ( .B1(n15509), .B2(n14900), .A(n14899), .ZN(n14901) );
  AOI21_X1 U16746 ( .B1(n14902), .B2(n15501), .A(n14901), .ZN(n14916) );
  MUX2_X1 U16747 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10730), .S(n14908), .Z(
        n14903) );
  NAND3_X1 U16748 ( .A1(n14905), .A2(n14904), .A3(n14903), .ZN(n14906) );
  NAND3_X1 U16749 ( .A1(n15505), .A2(n14907), .A3(n14906), .ZN(n14915) );
  MUX2_X1 U16750 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10696), .S(n14908), .Z(
        n14909) );
  NAND3_X1 U16751 ( .A1(n14911), .A2(n14910), .A3(n14909), .ZN(n14912) );
  NAND3_X1 U16752 ( .A1(n15504), .A2(n14913), .A3(n14912), .ZN(n14914) );
  NAND3_X1 U16753 ( .A1(n14916), .A2(n14915), .A3(n14914), .ZN(P1_U3250) );
  INV_X1 U16754 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14918) );
  OAI21_X1 U16755 ( .B1(n15509), .B2(n14918), .A(n14917), .ZN(n14919) );
  AOI21_X1 U16756 ( .B1(n14924), .B2(n15501), .A(n14919), .ZN(n14932) );
  OAI21_X1 U16757 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n14923) );
  NAND2_X1 U16758 ( .A1(n15504), .A2(n14923), .ZN(n14931) );
  MUX2_X1 U16759 ( .A(n10733), .B(P1_REG2_REG_9__SCAN_IN), .S(n14924), .Z(
        n14925) );
  NAND3_X1 U16760 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14928) );
  NAND3_X1 U16761 ( .A1(n15505), .A2(n14929), .A3(n14928), .ZN(n14930) );
  NAND3_X1 U16762 ( .A1(n14932), .A2(n14931), .A3(n14930), .ZN(P1_U3252) );
  OAI211_X1 U16763 ( .C1(n14935), .C2(n14934), .A(n14933), .B(n15504), .ZN(
        n14947) );
  NOR2_X1 U16764 ( .A1(n14957), .A2(n14939), .ZN(n14936) );
  AOI211_X1 U16765 ( .C1(n14938), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n14937), 
        .B(n14936), .ZN(n14946) );
  MUX2_X1 U16766 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n12104), .S(n14939), .Z(
        n14940) );
  NAND3_X1 U16767 ( .A1(n14942), .A2(n14941), .A3(n14940), .ZN(n14943) );
  NAND3_X1 U16768 ( .A1(n14944), .A2(n15505), .A3(n14943), .ZN(n14945) );
  NAND3_X1 U16769 ( .A1(n14947), .A2(n14946), .A3(n14945), .ZN(P1_U3260) );
  NAND2_X1 U16770 ( .A1(n14949), .A2(n14948), .ZN(n14950) );
  XNOR2_X1 U16771 ( .A(n14950), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14963) );
  NAND2_X1 U16772 ( .A1(n14963), .A2(n15504), .ZN(n14959) );
  NAND2_X1 U16773 ( .A1(n14951), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14955) );
  NAND2_X1 U16774 ( .A1(n14953), .A2(n14952), .ZN(n14954) );
  NAND2_X1 U16775 ( .A1(n14955), .A2(n14954), .ZN(n14956) );
  XNOR2_X1 U16776 ( .A(n14956), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U16777 ( .A1(n14961), .A2(n15505), .ZN(n14958) );
  NAND3_X1 U16778 ( .A1(n14959), .A2(n14958), .A3(n14957), .ZN(n14965) );
  OAI22_X1 U16779 ( .A1(n14963), .A2(n14962), .B1(n14961), .B2(n14960), .ZN(
        n14964) );
  NOR2_X2 U16780 ( .A1(n14976), .A2(n14968), .ZN(n14969) );
  XNOR2_X1 U16781 ( .A(n14969), .B(n15215), .ZN(n14970) );
  NAND2_X1 U16782 ( .A1(n14970), .A2(n15540), .ZN(n15216) );
  NAND2_X1 U16783 ( .A1(n14972), .A2(n14971), .ZN(n15218) );
  NOR2_X1 U16784 ( .A1(n15584), .A2(n15218), .ZN(n14979) );
  NOR2_X1 U16785 ( .A1(n15178), .A2(n14973), .ZN(n14974) );
  AOI211_X1 U16786 ( .C1(n15215), .C2(n15212), .A(n14979), .B(n14974), .ZN(
        n14975) );
  OAI21_X1 U16787 ( .B1(n15216), .B2(n15185), .A(n14975), .ZN(P1_U3263) );
  XNOR2_X1 U16788 ( .A(n14976), .B(n15220), .ZN(n14977) );
  NAND2_X1 U16789 ( .A1(n14977), .A2(n15540), .ZN(n15219) );
  NOR2_X1 U16790 ( .A1(n15220), .A2(n15552), .ZN(n14978) );
  AOI211_X1 U16791 ( .C1(n15584), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14979), 
        .B(n14978), .ZN(n14980) );
  OAI21_X1 U16792 ( .B1(n15185), .B2(n15219), .A(n14980), .ZN(P1_U3264) );
  XNOR2_X1 U16793 ( .A(n15232), .B(n14983), .ZN(n15240) );
  INV_X1 U16794 ( .A(n15240), .ZN(n14994) );
  OAI211_X1 U16795 ( .C1(n14998), .C2(n15224), .A(n15540), .B(n14984), .ZN(
        n15246) );
  NOR2_X1 U16796 ( .A1(n15246), .A2(n15185), .ZN(n14992) );
  INV_X1 U16797 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14985) );
  OAI22_X1 U16798 ( .A1(n14986), .A2(n15549), .B1(n14985), .B2(n15178), .ZN(
        n14987) );
  AOI21_X1 U16799 ( .B1(n14988), .B2(n15158), .A(n14987), .ZN(n14990) );
  NAND2_X1 U16800 ( .A1(n15016), .A2(n15192), .ZN(n14989) );
  OAI211_X1 U16801 ( .C1(n15224), .C2(n15552), .A(n14990), .B(n14989), .ZN(
        n14991) );
  AOI211_X1 U16802 ( .C1(n15248), .C2(n15581), .A(n14992), .B(n14991), .ZN(
        n14993) );
  OAI21_X1 U16803 ( .B1(n14994), .B2(n15095), .A(n14993), .ZN(P1_U3265) );
  OAI21_X1 U16804 ( .B1(n6680), .B2(n15007), .A(n14995), .ZN(n14996) );
  NAND2_X1 U16805 ( .A1(n14996), .A2(n15568), .ZN(n15257) );
  INV_X1 U16806 ( .A(n14997), .ZN(n15014) );
  AOI211_X1 U16807 ( .C1(n15255), .C2(n15014), .A(n15574), .B(n14998), .ZN(
        n15253) );
  AOI22_X1 U16808 ( .A1(n14999), .A2(n15573), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15584), .ZN(n15000) );
  OAI21_X1 U16809 ( .B1(n15252), .B2(n15196), .A(n15000), .ZN(n15001) );
  AOI21_X1 U16810 ( .B1(n15192), .B2(n15028), .A(n15001), .ZN(n15002) );
  OAI21_X1 U16811 ( .B1(n15003), .B2(n15552), .A(n15002), .ZN(n15008) );
  INV_X1 U16812 ( .A(n15004), .ZN(n15005) );
  OAI21_X1 U16813 ( .B1(n15257), .B2(n15584), .A(n15009), .ZN(P1_U3266) );
  XNOR2_X1 U16814 ( .A(n15011), .B(n15010), .ZN(n15265) );
  XNOR2_X1 U16815 ( .A(n15012), .B(n15013), .ZN(n15263) );
  OAI211_X1 U16816 ( .C1(n15261), .C2(n6646), .A(n15014), .B(n15540), .ZN(
        n15260) );
  AOI22_X1 U16817 ( .A1(n15016), .A2(n15668), .B1(n15665), .B2(n15015), .ZN(
        n15259) );
  AOI22_X1 U16818 ( .A1(n15017), .A2(n15573), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15584), .ZN(n15018) );
  OAI21_X1 U16819 ( .B1(n15259), .B2(n15584), .A(n15018), .ZN(n15019) );
  AOI21_X1 U16820 ( .B1(n15020), .B2(n15212), .A(n15019), .ZN(n15021) );
  OAI21_X1 U16821 ( .B1(n15260), .B2(n15185), .A(n15021), .ZN(n15022) );
  AOI21_X1 U16822 ( .B1(n15263), .B2(n15581), .A(n15022), .ZN(n15023) );
  OAI21_X1 U16823 ( .B1(n15265), .B2(n15095), .A(n15023), .ZN(P1_U3267) );
  NAND2_X1 U16824 ( .A1(n15038), .A2(n15024), .ZN(n15025) );
  XNOR2_X1 U16825 ( .A(n15025), .B(n15026), .ZN(n15272) );
  XNOR2_X1 U16826 ( .A(n15027), .B(n15026), .ZN(n15270) );
  INV_X1 U16827 ( .A(n15270), .ZN(n15032) );
  AOI211_X1 U16828 ( .C1(n15034), .C2(n15042), .A(n15574), .B(n6646), .ZN(
        n15269) );
  AOI22_X1 U16829 ( .A1(n15028), .A2(n15668), .B1(n15665), .B2(n15057), .ZN(
        n15266) );
  OAI21_X1 U16830 ( .B1(n15029), .B2(n15549), .A(n15266), .ZN(n15030) );
  AOI21_X1 U16831 ( .B1(n15269), .B2(n15207), .A(n15030), .ZN(n15031) );
  OAI21_X1 U16832 ( .B1(n15032), .B2(n15095), .A(n15031), .ZN(n15033) );
  NAND2_X1 U16833 ( .A1(n15033), .A2(n15178), .ZN(n15036) );
  AOI22_X1 U16834 ( .A1(n15034), .A2(n15212), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15584), .ZN(n15035) );
  OAI211_X1 U16835 ( .C1(n15272), .C2(n15214), .A(n15036), .B(n15035), .ZN(
        P1_U3268) );
  XNOR2_X1 U16836 ( .A(n15037), .B(n15039), .ZN(n15281) );
  INV_X1 U16837 ( .A(n15281), .ZN(n15052) );
  AOI21_X1 U16838 ( .B1(n15041), .B2(n15276), .A(n6601), .ZN(n15043) );
  NAND2_X1 U16839 ( .A1(n15043), .A2(n15042), .ZN(n15277) );
  AOI22_X1 U16840 ( .A1(n15044), .A2(n15573), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15584), .ZN(n15047) );
  NAND2_X1 U16841 ( .A1(n15192), .A2(n15045), .ZN(n15046) );
  OAI211_X1 U16842 ( .C1(n15274), .C2(n15196), .A(n15047), .B(n15046), .ZN(
        n15048) );
  AOI21_X1 U16843 ( .B1(n15276), .B2(n15212), .A(n15048), .ZN(n15049) );
  OAI21_X1 U16844 ( .B1(n15277), .B2(n15185), .A(n15049), .ZN(n15050) );
  AOI21_X1 U16845 ( .B1(n6896), .B2(n15581), .A(n15050), .ZN(n15051) );
  OAI21_X1 U16846 ( .B1(n15052), .B2(n15095), .A(n15051), .ZN(P1_U3269) );
  XNOR2_X1 U16847 ( .A(n15053), .B(n15055), .ZN(n15289) );
  OAI21_X1 U16848 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15287) );
  INV_X1 U16849 ( .A(n15095), .ZN(n15187) );
  OAI211_X1 U16850 ( .C1(n15073), .C2(n15285), .A(n15041), .B(n15540), .ZN(
        n15284) );
  AOI22_X1 U16851 ( .A1(n15057), .A2(n15668), .B1(n15665), .B2(n15294), .ZN(
        n15283) );
  NOR2_X1 U16852 ( .A1(n15283), .A2(n15584), .ZN(n15061) );
  OAI22_X1 U16853 ( .A1(n15178), .A2(n15059), .B1(n15058), .B2(n15549), .ZN(
        n15060) );
  AOI211_X1 U16854 ( .C1(n15062), .C2(n15212), .A(n15061), .B(n15060), .ZN(
        n15063) );
  OAI21_X1 U16855 ( .B1(n15284), .B2(n15185), .A(n15063), .ZN(n15064) );
  AOI21_X1 U16856 ( .B1(n15287), .B2(n15187), .A(n15064), .ZN(n15065) );
  OAI21_X1 U16857 ( .B1(n15214), .B2(n15289), .A(n15065), .ZN(P1_U3270) );
  NAND2_X1 U16858 ( .A1(n15066), .A2(n15082), .ZN(n15081) );
  NAND2_X1 U16859 ( .A1(n15081), .A2(n15067), .ZN(n15068) );
  XOR2_X1 U16860 ( .A(n15069), .B(n15068), .Z(n15293) );
  OAI222_X1 U16861 ( .A1(n15630), .A2(n15098), .B1(n15628), .B2(n15273), .C1(
        n15070), .C2(n15651), .ZN(n15290) );
  NAND2_X1 U16862 ( .A1(n15290), .A2(n15178), .ZN(n15079) );
  NAND2_X1 U16863 ( .A1(n15083), .A2(n7418), .ZN(n15071) );
  NAND2_X1 U16864 ( .A1(n15071), .A2(n15540), .ZN(n15072) );
  NOR2_X1 U16865 ( .A1(n15073), .A2(n15072), .ZN(n15291) );
  AOI22_X1 U16866 ( .A1(P1_REG2_REG_22__SCAN_IN), .A2(n15584), .B1(n15074), 
        .B2(n15573), .ZN(n15075) );
  OAI21_X1 U16867 ( .B1(n15076), .B2(n15552), .A(n15075), .ZN(n15077) );
  AOI21_X1 U16868 ( .B1(n15291), .B2(n15582), .A(n15077), .ZN(n15078) );
  OAI211_X1 U16869 ( .C1(n15293), .C2(n15214), .A(n15079), .B(n15078), .ZN(
        P1_U3271) );
  XNOR2_X1 U16870 ( .A(n15080), .B(n15082), .ZN(n15300) );
  OAI21_X1 U16871 ( .B1(n15066), .B2(n15082), .A(n15081), .ZN(n15298) );
  NAND2_X1 U16872 ( .A1(n15084), .A2(n15083), .ZN(n15296) );
  OR2_X1 U16873 ( .A1(n15162), .A2(n15129), .ZN(n15088) );
  NOR2_X1 U16874 ( .A1(n15085), .A2(n15549), .ZN(n15086) );
  AOI21_X1 U16875 ( .B1(n15584), .B2(P1_REG2_REG_21__SCAN_IN), .A(n15086), 
        .ZN(n15087) );
  OAI211_X1 U16876 ( .C1(n15089), .C2(n15196), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U16877 ( .B1(n15091), .B2(n15212), .A(n15090), .ZN(n15092) );
  OAI21_X1 U16878 ( .B1(n15296), .B2(n15185), .A(n15092), .ZN(n15093) );
  AOI21_X1 U16879 ( .B1(n15298), .B2(n15581), .A(n15093), .ZN(n15094) );
  OAI21_X1 U16880 ( .B1(n15300), .B2(n15095), .A(n15094), .ZN(P1_U3272) );
  OAI21_X1 U16881 ( .B1(n15139), .B2(n15138), .A(n15096), .ZN(n15119) );
  OR2_X1 U16882 ( .A1(n15119), .A2(n15120), .ZN(n15121) );
  OAI21_X1 U16883 ( .B1(n15309), .B2(n15145), .A(n15121), .ZN(n15097) );
  AOI21_X1 U16884 ( .B1(n15097), .B2(n10188), .A(n15651), .ZN(n15101) );
  OAI22_X1 U16885 ( .A1(n15098), .A2(n15628), .B1(n15314), .B2(n15630), .ZN(
        n15099) );
  AOI21_X1 U16886 ( .B1(n15101), .B2(n15100), .A(n15099), .ZN(n15303) );
  AOI211_X1 U16887 ( .C1(n10129), .C2(n15102), .A(n15574), .B(n15103), .ZN(
        n15301) );
  INV_X1 U16888 ( .A(n10129), .ZN(n15107) );
  INV_X1 U16889 ( .A(n15104), .ZN(n15105) );
  AOI22_X1 U16890 ( .A1(n15584), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n15105), 
        .B2(n15573), .ZN(n15106) );
  OAI21_X1 U16891 ( .B1(n15107), .B2(n15552), .A(n15106), .ZN(n15113) );
  NAND2_X1 U16892 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  NAND2_X1 U16893 ( .A1(n15111), .A2(n15110), .ZN(n15304) );
  NOR2_X1 U16894 ( .A1(n15304), .A2(n15214), .ZN(n15112) );
  AOI211_X1 U16895 ( .C1(n15301), .C2(n15582), .A(n15113), .B(n15112), .ZN(
        n15114) );
  OAI21_X1 U16896 ( .B1(n15303), .B2(n15584), .A(n15114), .ZN(P1_U3273) );
  INV_X1 U16897 ( .A(n15136), .ZN(n15117) );
  AOI22_X1 U16898 ( .A1(n15117), .A2(n15116), .B1(n15322), .B2(n15315), .ZN(
        n15118) );
  XNOR2_X1 U16899 ( .A(n15118), .B(n15120), .ZN(n15313) );
  INV_X1 U16900 ( .A(n15119), .ZN(n15123) );
  INV_X1 U16901 ( .A(n15120), .ZN(n15122) );
  OAI21_X1 U16902 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15311) );
  OAI211_X1 U16903 ( .C1(n15124), .C2(n15309), .A(n15540), .B(n15102), .ZN(
        n15308) );
  NAND2_X1 U16904 ( .A1(n15192), .A2(n15305), .ZN(n15128) );
  INV_X1 U16905 ( .A(n15125), .ZN(n15126) );
  AOI22_X1 U16906 ( .A1(n15584), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n15126), 
        .B2(n15573), .ZN(n15127) );
  OAI211_X1 U16907 ( .C1(n15129), .C2(n15196), .A(n15128), .B(n15127), .ZN(
        n15130) );
  AOI21_X1 U16908 ( .B1(n15131), .B2(n15212), .A(n15130), .ZN(n15132) );
  OAI21_X1 U16909 ( .B1(n15308), .B2(n15185), .A(n15132), .ZN(n15133) );
  AOI21_X1 U16910 ( .B1(n15311), .B2(n15187), .A(n15133), .ZN(n15134) );
  OAI21_X1 U16911 ( .B1(n15214), .B2(n15313), .A(n15134), .ZN(P1_U3274) );
  INV_X1 U16912 ( .A(n15138), .ZN(n15135) );
  XNOR2_X1 U16913 ( .A(n15136), .B(n15135), .ZN(n15148) );
  INV_X1 U16914 ( .A(n15137), .ZN(n15678) );
  XOR2_X1 U16915 ( .A(n15139), .B(n15138), .Z(n15140) );
  AOI222_X1 U16916 ( .A1(n15148), .A2(n15678), .B1(n15568), .B2(n15140), .C1(
        n15329), .C2(n15665), .ZN(n15319) );
  INV_X1 U16917 ( .A(n15141), .ZN(n15142) );
  AOI211_X1 U16918 ( .C1(n15143), .C2(n15142), .A(n6601), .B(n15124), .ZN(
        n15317) );
  AOI22_X1 U16919 ( .A1(n15584), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15144), 
        .B2(n15573), .ZN(n15147) );
  NAND2_X1 U16920 ( .A1(n15158), .A2(n15145), .ZN(n15146) );
  OAI211_X1 U16921 ( .C1(n15315), .C2(n15552), .A(n15147), .B(n15146), .ZN(
        n15151) );
  INV_X1 U16922 ( .A(n15148), .ZN(n15320) );
  OR2_X1 U16923 ( .A1(n15584), .A2(n15149), .ZN(n15521) );
  NOR2_X1 U16924 ( .A1(n15320), .A2(n15521), .ZN(n15150) );
  AOI211_X1 U16925 ( .C1(n15317), .C2(n15582), .A(n15151), .B(n15150), .ZN(
        n15152) );
  OAI21_X1 U16926 ( .B1(n15319), .B2(n15584), .A(n15152), .ZN(P1_U3275) );
  XNOR2_X1 U16927 ( .A(n15153), .B(n15156), .ZN(n15328) );
  AOI211_X1 U16928 ( .C1(n15156), .C2(n15155), .A(n15651), .B(n15154), .ZN(
        n15157) );
  INV_X1 U16929 ( .A(n15157), .ZN(n15327) );
  NAND2_X1 U16930 ( .A1(n15158), .A2(n15305), .ZN(n15161) );
  AOI22_X1 U16931 ( .A1(n15584), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15159), 
        .B2(n15573), .ZN(n15160) );
  OAI211_X1 U16932 ( .C1(n15321), .C2(n15162), .A(n15161), .B(n15160), .ZN(
        n15163) );
  AOI21_X1 U16933 ( .B1(n15325), .B2(n15212), .A(n15163), .ZN(n15167) );
  NAND2_X1 U16934 ( .A1(n7638), .A2(n15325), .ZN(n15164) );
  NAND2_X1 U16935 ( .A1(n15164), .A2(n15540), .ZN(n15165) );
  NOR2_X1 U16936 ( .A1(n15141), .A2(n15165), .ZN(n15323) );
  NAND2_X1 U16937 ( .A1(n15323), .A2(n15582), .ZN(n15166) );
  OAI211_X1 U16938 ( .C1(n15327), .C2(n15584), .A(n15167), .B(n15166), .ZN(
        n15168) );
  INV_X1 U16939 ( .A(n15168), .ZN(n15169) );
  OAI21_X1 U16940 ( .B1(n15214), .B2(n15328), .A(n15169), .ZN(P1_U3276) );
  XNOR2_X1 U16941 ( .A(n15171), .B(n15170), .ZN(n15336) );
  XNOR2_X1 U16942 ( .A(n15172), .B(n15173), .ZN(n15334) );
  INV_X1 U16943 ( .A(n15174), .ZN(n15175) );
  OAI211_X1 U16944 ( .C1(n15175), .C2(n15332), .A(n15540), .B(n7638), .ZN(
        n15331) );
  INV_X1 U16945 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15177) );
  OAI22_X1 U16946 ( .A1(n15178), .A2(n15177), .B1(n15176), .B2(n15549), .ZN(
        n15179) );
  AOI21_X1 U16947 ( .B1(n15192), .B2(n15344), .A(n15179), .ZN(n15180) );
  OAI21_X1 U16948 ( .B1(n15181), .B2(n15196), .A(n15180), .ZN(n15182) );
  AOI21_X1 U16949 ( .B1(n15183), .B2(n15212), .A(n15182), .ZN(n15184) );
  OAI21_X1 U16950 ( .B1(n15331), .B2(n15185), .A(n15184), .ZN(n15186) );
  AOI21_X1 U16951 ( .B1(n15334), .B2(n15187), .A(n15186), .ZN(n15188) );
  OAI21_X1 U16952 ( .B1(n15214), .B2(n15336), .A(n15188), .ZN(P1_U3277) );
  NAND2_X1 U16953 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  XNOR2_X1 U16954 ( .A(n15191), .B(n15204), .ZN(n15351) );
  NAND2_X1 U16955 ( .A1(n15192), .A2(n15363), .ZN(n15195) );
  AOI22_X1 U16956 ( .A1(n15584), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15193), 
        .B2(n15573), .ZN(n15194) );
  OAI211_X1 U16957 ( .C1(n15197), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        n15210) );
  NAND2_X1 U16958 ( .A1(n15198), .A2(n15211), .ZN(n15199) );
  NAND2_X1 U16959 ( .A1(n15199), .A2(n15540), .ZN(n15200) );
  NOR2_X1 U16960 ( .A1(n15201), .A2(n15200), .ZN(n15348) );
  NAND2_X1 U16961 ( .A1(n15203), .A2(n15202), .ZN(n15205) );
  XNOR2_X1 U16962 ( .A(n15205), .B(n15204), .ZN(n15206) );
  NOR2_X1 U16963 ( .A1(n15206), .A2(n15651), .ZN(n15349) );
  AOI21_X1 U16964 ( .B1(n15348), .B2(n15207), .A(n15349), .ZN(n15208) );
  NOR2_X1 U16965 ( .A1(n15208), .A2(n15584), .ZN(n15209) );
  AOI211_X1 U16966 ( .C1(n15212), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15213) );
  OAI21_X1 U16967 ( .B1(n15214), .B2(n15351), .A(n15213), .ZN(P1_U3279) );
  INV_X1 U16968 ( .A(n15215), .ZN(n15217) );
  MUX2_X1 U16969 ( .A(n15396), .B(P1_REG1_REG_31__SCAN_IN), .S(n15711), .Z(
        P1_U3559) );
  MUX2_X1 U16970 ( .A(n15397), .B(P1_REG1_REG_30__SCAN_IN), .S(n15711), .Z(
        P1_U3558) );
  INV_X1 U16971 ( .A(n15227), .ZN(n15221) );
  NAND2_X1 U16972 ( .A1(n15222), .A2(n15221), .ZN(n15231) );
  NAND2_X1 U16973 ( .A1(n15224), .A2(n15223), .ZN(n15225) );
  NOR2_X1 U16974 ( .A1(n15228), .A2(n15225), .ZN(n15226) );
  AOI211_X1 U16975 ( .C1(n15228), .C2(n15227), .A(n15651), .B(n15226), .ZN(
        n15229) );
  OAI211_X1 U16976 ( .C1(n15232), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        n15238) );
  OAI21_X1 U16977 ( .B1(n15252), .B2(n15630), .A(n15233), .ZN(n15234) );
  INV_X1 U16978 ( .A(n15234), .ZN(n15236) );
  OAI211_X1 U16979 ( .C1(n15694), .C2(n15239), .A(n15238), .B(n6693), .ZN(
        n15398) );
  MUX2_X1 U16980 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15398), .S(n15714), .Z(
        P1_U3557) );
  NAND2_X1 U16981 ( .A1(n15240), .A2(n15568), .ZN(n15250) );
  INV_X1 U16982 ( .A(n15694), .ZN(n15655) );
  OAI22_X1 U16983 ( .A1(n15242), .A2(n15630), .B1(n15241), .B2(n15628), .ZN(
        n15243) );
  AOI21_X1 U16984 ( .B1(n15244), .B2(n15388), .A(n15243), .ZN(n15245) );
  NAND2_X1 U16985 ( .A1(n15246), .A2(n15245), .ZN(n15247) );
  NAND2_X1 U16986 ( .A1(n15250), .A2(n15249), .ZN(n15399) );
  MUX2_X1 U16987 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15399), .S(n15714), .Z(
        P1_U3556) );
  OAI22_X1 U16988 ( .A1(n15252), .A2(n15628), .B1(n15251), .B2(n15630), .ZN(
        n15254) );
  AOI211_X1 U16989 ( .C1(n15255), .C2(n15388), .A(n15254), .B(n15253), .ZN(
        n15256) );
  OAI211_X1 U16990 ( .C1(n15694), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15400) );
  MUX2_X1 U16991 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15400), .S(n15714), .Z(
        P1_U3555) );
  OAI211_X1 U16992 ( .C1(n15261), .C2(n15682), .A(n15260), .B(n15259), .ZN(
        n15262) );
  AOI21_X1 U16993 ( .B1(n15263), .B2(n15655), .A(n15262), .ZN(n15264) );
  OAI21_X1 U16994 ( .B1(n15265), .B2(n15651), .A(n15264), .ZN(n15401) );
  MUX2_X1 U16995 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15401), .S(n15714), .Z(
        P1_U3554) );
  OAI21_X1 U16996 ( .B1(n15267), .B2(n15682), .A(n15266), .ZN(n15268) );
  AOI211_X1 U16997 ( .C1(n15270), .C2(n15568), .A(n15269), .B(n15268), .ZN(
        n15271) );
  OAI21_X1 U16998 ( .B1(n15694), .B2(n15272), .A(n15271), .ZN(n15402) );
  MUX2_X1 U16999 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15402), .S(n15714), .Z(
        P1_U3553) );
  OAI22_X1 U17000 ( .A1(n15274), .A2(n15628), .B1(n15273), .B2(n15630), .ZN(
        n15275) );
  AOI21_X1 U17001 ( .B1(n15276), .B2(n15388), .A(n15275), .ZN(n15278) );
  OAI211_X1 U17002 ( .C1(n15279), .C2(n15694), .A(n15278), .B(n15277), .ZN(
        n15280) );
  INV_X1 U17003 ( .A(n15282), .ZN(n15403) );
  MUX2_X1 U17004 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15403), .S(n15714), .Z(
        P1_U3552) );
  OAI211_X1 U17005 ( .C1(n15285), .C2(n15682), .A(n15284), .B(n15283), .ZN(
        n15286) );
  AOI21_X1 U17006 ( .B1(n15287), .B2(n15568), .A(n15286), .ZN(n15288) );
  OAI21_X1 U17007 ( .B1(n15694), .B2(n15289), .A(n15288), .ZN(n15404) );
  MUX2_X1 U17008 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15404), .S(n15714), .Z(
        P1_U3551) );
  AOI211_X1 U17009 ( .C1(n7418), .C2(n15388), .A(n15291), .B(n15290), .ZN(
        n15292) );
  MUX2_X1 U17010 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15405), .S(n15714), .Z(
        P1_U3550) );
  AOI22_X1 U17011 ( .A1(n15294), .A2(n15668), .B1(n15665), .B2(n15306), .ZN(
        n15295) );
  OAI211_X1 U17012 ( .C1(n7436), .C2(n15682), .A(n15296), .B(n15295), .ZN(
        n15297) );
  AOI21_X1 U17013 ( .B1(n15298), .B2(n15655), .A(n15297), .ZN(n15299) );
  OAI21_X1 U17014 ( .B1(n15300), .B2(n15651), .A(n15299), .ZN(n15406) );
  MUX2_X1 U17015 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15406), .S(n15714), .Z(
        P1_U3549) );
  AOI21_X1 U17016 ( .B1(n10129), .B2(n15388), .A(n15301), .ZN(n15302) );
  OAI211_X1 U17017 ( .C1(n15694), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15407) );
  MUX2_X1 U17018 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15407), .S(n15714), .Z(
        P1_U3548) );
  AOI22_X1 U17019 ( .A1(n15668), .A2(n15306), .B1(n15305), .B2(n15665), .ZN(
        n15307) );
  OAI211_X1 U17020 ( .C1(n15309), .C2(n15682), .A(n15308), .B(n15307), .ZN(
        n15310) );
  AOI21_X1 U17021 ( .B1(n15311), .B2(n15568), .A(n15310), .ZN(n15312) );
  OAI21_X1 U17022 ( .B1(n15694), .B2(n15313), .A(n15312), .ZN(n15408) );
  MUX2_X1 U17023 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15408), .S(n15714), .Z(
        P1_U3547) );
  OAI22_X1 U17024 ( .A1(n15315), .A2(n15682), .B1(n15314), .B2(n15628), .ZN(
        n15316) );
  NOR2_X1 U17025 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  OAI211_X1 U17026 ( .C1(n15320), .C2(n15674), .A(n15319), .B(n15318), .ZN(
        n15409) );
  MUX2_X1 U17027 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15409), .S(n15714), .Z(
        P1_U3546) );
  OAI22_X1 U17028 ( .A1(n15322), .A2(n15628), .B1(n15321), .B2(n15630), .ZN(
        n15324) );
  AOI211_X1 U17029 ( .C1(n15325), .C2(n15388), .A(n15324), .B(n15323), .ZN(
        n15326) );
  OAI211_X1 U17030 ( .C1(n15694), .C2(n15328), .A(n15327), .B(n15326), .ZN(
        n15410) );
  MUX2_X1 U17031 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15410), .S(n15714), .Z(
        P1_U3545) );
  AOI22_X1 U17032 ( .A1(n15329), .A2(n15668), .B1(n15665), .B2(n15344), .ZN(
        n15330) );
  OAI211_X1 U17033 ( .C1(n15332), .C2(n15682), .A(n15331), .B(n15330), .ZN(
        n15333) );
  AOI21_X1 U17034 ( .B1(n15334), .B2(n15568), .A(n15333), .ZN(n15335) );
  OAI21_X1 U17035 ( .B1(n15694), .B2(n15336), .A(n15335), .ZN(n15411) );
  MUX2_X1 U17036 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15411), .S(n15714), .Z(
        P1_U3544) );
  OAI211_X1 U17037 ( .C1(n15339), .C2(n15682), .A(n15338), .B(n15337), .ZN(
        n15340) );
  AOI21_X1 U17038 ( .B1(n15341), .B2(n15655), .A(n15340), .ZN(n15342) );
  OAI21_X1 U17039 ( .B1(n15343), .B2(n15651), .A(n15342), .ZN(n15412) );
  MUX2_X1 U17040 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15412), .S(n15714), .Z(
        P1_U3543) );
  AOI22_X1 U17041 ( .A1(n15363), .A2(n15665), .B1(n15668), .B2(n15344), .ZN(
        n15345) );
  OAI21_X1 U17042 ( .B1(n15346), .B2(n15682), .A(n15345), .ZN(n15347) );
  NOR3_X1 U17043 ( .A1(n15349), .A2(n15348), .A3(n15347), .ZN(n15350) );
  OAI21_X1 U17044 ( .B1(n15694), .B2(n15351), .A(n15350), .ZN(n15413) );
  MUX2_X1 U17045 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15413), .S(n15714), .Z(
        P1_U3542) );
  INV_X1 U17046 ( .A(n15352), .ZN(n15357) );
  AOI22_X1 U17047 ( .A1(n15354), .A2(n15668), .B1(n15665), .B2(n15353), .ZN(
        n15355) );
  OAI211_X1 U17048 ( .C1(n15357), .C2(n15682), .A(n15356), .B(n15355), .ZN(
        n15358) );
  INV_X1 U17049 ( .A(n15358), .ZN(n15360) );
  OAI211_X1 U17050 ( .C1(n15361), .C2(n15694), .A(n15360), .B(n15359), .ZN(
        n15414) );
  MUX2_X1 U17051 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15414), .S(n15714), .Z(
        P1_U3541) );
  AOI22_X1 U17052 ( .A1(n15363), .A2(n15668), .B1(n15665), .B2(n15362), .ZN(
        n15364) );
  OAI211_X1 U17053 ( .C1(n6549), .C2(n15682), .A(n15365), .B(n15364), .ZN(
        n15367) );
  AOI211_X1 U17054 ( .C1(n15655), .C2(n15368), .A(n15367), .B(n15366), .ZN(
        n15369) );
  INV_X1 U17055 ( .A(n15369), .ZN(n15415) );
  MUX2_X1 U17056 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15415), .S(n15714), .Z(
        P1_U3540) );
  AOI211_X1 U17057 ( .C1(n15372), .C2(n15388), .A(n15371), .B(n15370), .ZN(
        n15373) );
  OAI21_X1 U17058 ( .B1(n15694), .B2(n15374), .A(n15373), .ZN(n15416) );
  MUX2_X1 U17059 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15416), .S(n15714), .Z(
        P1_U3539) );
  NOR3_X1 U17060 ( .A1(n15376), .A2(n15375), .A3(n15651), .ZN(n15381) );
  OAI22_X1 U17061 ( .A1(n15378), .A2(n15682), .B1(n15377), .B2(n15630), .ZN(
        n15379) );
  NOR3_X1 U17062 ( .A1(n15381), .A2(n15380), .A3(n15379), .ZN(n15382) );
  OAI21_X1 U17063 ( .B1(n15694), .B2(n15383), .A(n15382), .ZN(n15417) );
  MUX2_X1 U17064 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15417), .S(n15714), .Z(
        P1_U3538) );
  OAI22_X1 U17065 ( .A1(n15385), .A2(n15630), .B1(n15384), .B2(n15628), .ZN(
        n15387) );
  AOI211_X1 U17066 ( .C1(n15389), .C2(n15388), .A(n15387), .B(n15386), .ZN(
        n15392) );
  INV_X1 U17067 ( .A(n15390), .ZN(n15391) );
  OAI211_X1 U17068 ( .C1(n15393), .C2(n15694), .A(n15392), .B(n15391), .ZN(
        n15418) );
  MUX2_X1 U17069 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15418), .S(n15714), .Z(
        P1_U3537) );
  AND2_X2 U17070 ( .A1(n15395), .A2(n15394), .ZN(n15700) );
  MUX2_X1 U17071 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15398), .S(n15700), .Z(
        P1_U3525) );
  MUX2_X1 U17072 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15399), .S(n15700), .Z(
        P1_U3524) );
  MUX2_X1 U17073 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15400), .S(n15700), .Z(
        P1_U3523) );
  MUX2_X1 U17074 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15401), .S(n15700), .Z(
        P1_U3522) );
  MUX2_X1 U17075 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15402), .S(n15700), .Z(
        P1_U3521) );
  MUX2_X1 U17076 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15403), .S(n15700), .Z(
        P1_U3520) );
  MUX2_X1 U17077 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15404), .S(n15700), .Z(
        P1_U3519) );
  MUX2_X1 U17078 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15406), .S(n15700), .Z(
        P1_U3517) );
  MUX2_X1 U17079 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15407), .S(n15700), .Z(
        P1_U3516) );
  MUX2_X1 U17080 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15408), .S(n15700), .Z(
        P1_U3515) );
  MUX2_X1 U17081 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15409), .S(n15700), .Z(
        P1_U3513) );
  MUX2_X1 U17082 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15410), .S(n15700), .Z(
        P1_U3510) );
  MUX2_X1 U17083 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15411), .S(n15700), .Z(
        P1_U3507) );
  MUX2_X1 U17084 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15412), .S(n15700), .Z(
        P1_U3504) );
  MUX2_X1 U17085 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15413), .S(n15700), .Z(
        P1_U3501) );
  MUX2_X1 U17086 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15414), .S(n15700), .Z(
        P1_U3498) );
  MUX2_X1 U17087 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15415), .S(n15700), .Z(
        P1_U3495) );
  MUX2_X1 U17088 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15416), .S(n15700), .Z(
        P1_U3492) );
  MUX2_X1 U17089 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15417), .S(n15700), .Z(
        P1_U3489) );
  MUX2_X1 U17090 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n15418), .S(n15700), .Z(
        P1_U3486) );
  NOR4_X1 U17091 ( .A1(n15420), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15419), .A4(
        P1_U3086), .ZN(n15421) );
  AOI21_X1 U17092 ( .B1(n15422), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15421), 
        .ZN(n15423) );
  OAI21_X1 U17093 ( .B1(n15424), .B2(n6554), .A(n15423), .ZN(P1_U3324) );
  OAI222_X1 U17094 ( .A1(n6554), .A2(n12426), .B1(P1_U3086), .B2(n15426), .C1(
        n15425), .C2(n15433), .ZN(P1_U3325) );
  OAI222_X1 U17095 ( .A1(n6554), .A2(n15429), .B1(P1_U3086), .B2(n15428), .C1(
        n15427), .C2(n15433), .ZN(P1_U3326) );
  OAI222_X1 U17096 ( .A1(n15433), .A2(n15432), .B1(n6554), .B2(n15431), .C1(
        P1_U3086), .C2(n15430), .ZN(P1_U3327) );
  MUX2_X1 U17097 ( .A(n6608), .B(n15434), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U17098 ( .A(n15435), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U17099 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15436) );
  OAI21_X1 U17100 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15436), 
        .ZN(U28) );
  AOI21_X1 U17101 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15437) );
  OAI21_X1 U17102 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15437), 
        .ZN(U29) );
  OAI21_X1 U17103 ( .B1(n15440), .B2(n15439), .A(n15438), .ZN(n15442) );
  XOR2_X1 U17104 ( .A(n15442), .B(n15441), .Z(SUB_1596_U61) );
  AOI21_X1 U17105 ( .B1(n15445), .B2(n15444), .A(n15443), .ZN(SUB_1596_U57) );
  AOI21_X1 U17106 ( .B1(n15448), .B2(n15447), .A(n15446), .ZN(n15449) );
  XOR2_X1 U17107 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15449), .Z(SUB_1596_U55) );
  AOI21_X1 U17108 ( .B1(n15730), .B2(n15450), .A(n15451), .ZN(SUB_1596_U54) );
  OAI21_X1 U17109 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n15455) );
  XNOR2_X1 U17110 ( .A(n15455), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  AOI21_X1 U17111 ( .B1(n15457), .B2(n15456), .A(n6742), .ZN(SUB_1596_U63) );
  OAI21_X1 U17112 ( .B1(n15460), .B2(n15459), .A(n15458), .ZN(SUB_1596_U69) );
  AOI21_X1 U17113 ( .B1(n15463), .B2(n15462), .A(n15461), .ZN(n15464) );
  XNOR2_X1 U17114 ( .A(n7497), .B(n15464), .ZN(SUB_1596_U68) );
  OAI21_X1 U17115 ( .B1(n15467), .B2(n15466), .A(n15465), .ZN(n15468) );
  XNOR2_X1 U17116 ( .A(n15468), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U17117 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n15472) );
  XNOR2_X1 U17118 ( .A(n15472), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U17119 ( .A1(n15477), .A2(n15476), .B1(n15477), .B2(n15475), .C1(
        n15474), .C2(n15473), .ZN(SUB_1596_U65) );
  OAI21_X1 U17120 ( .B1(n15480), .B2(n15479), .A(n15478), .ZN(n15481) );
  XNOR2_X1 U17121 ( .A(n15481), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NOR2_X1 U17122 ( .A1(n15682), .A2(n10156), .ZN(n15641) );
  AOI21_X1 U17123 ( .B1(n15483), .B2(n15641), .A(n15482), .ZN(n15494) );
  XOR2_X1 U17124 ( .A(n15484), .B(n15485), .Z(n15492) );
  OR2_X1 U17125 ( .A1(n15486), .A2(n15630), .ZN(n15489) );
  OR2_X1 U17126 ( .A1(n15487), .A2(n15628), .ZN(n15488) );
  NAND2_X1 U17127 ( .A1(n15489), .A2(n15488), .ZN(n15640) );
  AOI22_X1 U17128 ( .A1(n15492), .A2(n15491), .B1(n15490), .B2(n15640), .ZN(
        n15493) );
  OAI211_X1 U17129 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n15495), .A(n15494), .B(
        n15493), .ZN(P1_U3218) );
  OAI21_X1 U17130 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15506) );
  XNOR2_X1 U17131 ( .A(n15500), .B(n15499), .ZN(n15503) );
  AOI222_X1 U17132 ( .A1(n15506), .A2(n15505), .B1(n15504), .B2(n15503), .C1(
        n15502), .C2(n15501), .ZN(n15508) );
  OAI211_X1 U17133 ( .C1(n15510), .C2(n15509), .A(n15508), .B(n15507), .ZN(
        P1_U3258) );
  XNOR2_X1 U17134 ( .A(n15511), .B(n15512), .ZN(n15687) );
  XNOR2_X1 U17135 ( .A(n15513), .B(n15512), .ZN(n15516) );
  AOI22_X1 U17136 ( .A1(n15668), .A2(n15514), .B1(n15531), .B2(n15665), .ZN(
        n15515) );
  OAI21_X1 U17137 ( .B1(n15516), .B2(n15651), .A(n15515), .ZN(n15517) );
  AOI21_X1 U17138 ( .B1(n15678), .B2(n15687), .A(n15517), .ZN(n15684) );
  AOI22_X1 U17139 ( .A1(n15584), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n15518), 
        .B2(n15573), .ZN(n15519) );
  OAI21_X1 U17140 ( .B1(n15552), .B2(n15683), .A(n15519), .ZN(n15520) );
  INV_X1 U17141 ( .A(n15520), .ZN(n15526) );
  INV_X1 U17142 ( .A(n15521), .ZN(n15558) );
  OAI211_X1 U17143 ( .C1(n15523), .C2(n15683), .A(n15540), .B(n15522), .ZN(
        n15681) );
  INV_X1 U17144 ( .A(n15681), .ZN(n15524) );
  AOI22_X1 U17145 ( .A1(n15687), .A2(n15558), .B1(n15582), .B2(n15524), .ZN(
        n15525) );
  OAI211_X1 U17146 ( .C1(n15584), .C2(n15684), .A(n15526), .B(n15525), .ZN(
        P1_U3286) );
  XNOR2_X1 U17147 ( .A(n15528), .B(n15529), .ZN(n15663) );
  XNOR2_X1 U17148 ( .A(n15530), .B(n15529), .ZN(n15534) );
  AOI22_X1 U17149 ( .A1(n15532), .A2(n15665), .B1(n15668), .B2(n15531), .ZN(
        n15533) );
  OAI21_X1 U17150 ( .B1(n15534), .B2(n15651), .A(n15533), .ZN(n15535) );
  AOI21_X1 U17151 ( .B1(n15678), .B2(n15663), .A(n15535), .ZN(n15660) );
  AOI22_X1 U17152 ( .A1(n15584), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15536), 
        .B2(n15573), .ZN(n15537) );
  OAI21_X1 U17153 ( .B1(n15552), .B2(n15659), .A(n15537), .ZN(n15538) );
  INV_X1 U17154 ( .A(n15538), .ZN(n15544) );
  INV_X1 U17155 ( .A(n6753), .ZN(n15541) );
  OAI211_X1 U17156 ( .C1(n15659), .C2(n7442), .A(n15541), .B(n15540), .ZN(
        n15658) );
  INV_X1 U17157 ( .A(n15658), .ZN(n15542) );
  AOI22_X1 U17158 ( .A1(n15663), .A2(n15558), .B1(n15582), .B2(n15542), .ZN(
        n15543) );
  OAI211_X1 U17159 ( .C1(n15584), .C2(n15660), .A(n15544), .B(n15543), .ZN(
        P1_U3288) );
  XNOR2_X1 U17160 ( .A(n15545), .B(n15546), .ZN(n15645) );
  XNOR2_X1 U17161 ( .A(n15547), .B(n15546), .ZN(n15548) );
  NOR2_X1 U17162 ( .A1(n15548), .A2(n15651), .ZN(n15643) );
  AOI211_X1 U17163 ( .C1(n15678), .C2(n15645), .A(n15640), .B(n15643), .ZN(
        n15561) );
  NOR2_X1 U17164 ( .A1(n15549), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15550) );
  AOI21_X1 U17165 ( .B1(n15584), .B2(P1_REG2_REG_3__SCAN_IN), .A(n15550), .ZN(
        n15551) );
  OAI21_X1 U17166 ( .B1(n15552), .B2(n10156), .A(n15551), .ZN(n15553) );
  INV_X1 U17167 ( .A(n15553), .ZN(n15560) );
  INV_X1 U17168 ( .A(n15554), .ZN(n15556) );
  AOI211_X1 U17169 ( .C1(n15557), .C2(n15556), .A(n15574), .B(n10211), .ZN(
        n15642) );
  AOI22_X1 U17170 ( .A1(n15558), .A2(n15645), .B1(n15642), .B2(n15582), .ZN(
        n15559) );
  OAI211_X1 U17171 ( .C1(n15584), .C2(n15561), .A(n15560), .B(n15559), .ZN(
        P1_U3290) );
  NAND2_X1 U17172 ( .A1(n15562), .A2(n15668), .ZN(n15620) );
  OAI21_X1 U17173 ( .B1(n6593), .B2(n15563), .A(n15620), .ZN(n15572) );
  OAI21_X1 U17174 ( .B1(n15578), .B2(n15564), .A(n15568), .ZN(n15571) );
  OAI21_X1 U17175 ( .B1(n6593), .B2(n12492), .A(n15565), .ZN(n15575) );
  XNOR2_X1 U17176 ( .A(n15575), .B(n15566), .ZN(n15569) );
  AOI21_X1 U17177 ( .B1(n15569), .B2(n15568), .A(n15567), .ZN(n15570) );
  AOI21_X1 U17178 ( .B1(n15630), .B2(n15571), .A(n15570), .ZN(n15623) );
  AOI211_X1 U17179 ( .C1(n15573), .C2(P1_REG3_REG_1__SCAN_IN), .A(n15572), .B(
        n15623), .ZN(n15585) );
  NOR2_X1 U17180 ( .A1(n15575), .A2(n6601), .ZN(n15619) );
  INV_X1 U17181 ( .A(n15576), .ZN(n15580) );
  OAI22_X1 U17182 ( .A1(n15580), .A2(n15579), .B1(n15578), .B2(n15577), .ZN(
        n15625) );
  AOI222_X1 U17183 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n15584), .B1(n15582), 
        .B2(n15619), .C1(n15625), .C2(n15581), .ZN(n15583) );
  OAI21_X1 U17184 ( .B1(n15585), .B2(n15584), .A(n15583), .ZN(P1_U3292) );
  NOR2_X1 U17185 ( .A1(n15616), .A2(n15586), .ZN(P1_U3294) );
  INV_X1 U17186 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15587) );
  NOR2_X1 U17187 ( .A1(n15616), .A2(n15587), .ZN(P1_U3295) );
  INV_X1 U17188 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15588) );
  NOR2_X1 U17189 ( .A1(n15616), .A2(n15588), .ZN(P1_U3296) );
  INV_X1 U17190 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15589) );
  NOR2_X1 U17191 ( .A1(n15616), .A2(n15589), .ZN(P1_U3297) );
  INV_X1 U17192 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15590) );
  NOR2_X1 U17193 ( .A1(n15616), .A2(n15590), .ZN(P1_U3298) );
  INV_X1 U17194 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15591) );
  NOR2_X1 U17195 ( .A1(n15616), .A2(n15591), .ZN(P1_U3299) );
  INV_X1 U17196 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15592) );
  NOR2_X1 U17197 ( .A1(n15616), .A2(n15592), .ZN(P1_U3300) );
  NOR2_X1 U17198 ( .A1(n15616), .A2(n15593), .ZN(P1_U3301) );
  NOR2_X1 U17199 ( .A1(n15616), .A2(n15594), .ZN(P1_U3302) );
  NOR2_X1 U17200 ( .A1(n15616), .A2(n15595), .ZN(P1_U3303) );
  INV_X1 U17201 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15596) );
  NOR2_X1 U17202 ( .A1(n15616), .A2(n15596), .ZN(P1_U3304) );
  INV_X1 U17203 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15597) );
  NOR2_X1 U17204 ( .A1(n15616), .A2(n15597), .ZN(P1_U3305) );
  INV_X1 U17205 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15598) );
  NOR2_X1 U17206 ( .A1(n15616), .A2(n15598), .ZN(P1_U3306) );
  INV_X1 U17207 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15599) );
  NOR2_X1 U17208 ( .A1(n15616), .A2(n15599), .ZN(P1_U3307) );
  INV_X1 U17209 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15600) );
  NOR2_X1 U17210 ( .A1(n15616), .A2(n15600), .ZN(P1_U3308) );
  INV_X1 U17211 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15601) );
  NOR2_X1 U17212 ( .A1(n15616), .A2(n15601), .ZN(P1_U3309) );
  NOR2_X1 U17213 ( .A1(n15616), .A2(n15602), .ZN(P1_U3310) );
  NOR2_X1 U17214 ( .A1(n15616), .A2(n15603), .ZN(P1_U3311) );
  INV_X1 U17215 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15604) );
  NOR2_X1 U17216 ( .A1(n15616), .A2(n15604), .ZN(P1_U3312) );
  NOR2_X1 U17217 ( .A1(n15616), .A2(n15605), .ZN(P1_U3313) );
  INV_X1 U17218 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15606) );
  NOR2_X1 U17219 ( .A1(n15616), .A2(n15606), .ZN(P1_U3314) );
  INV_X1 U17220 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15607) );
  NOR2_X1 U17221 ( .A1(n15616), .A2(n15607), .ZN(P1_U3315) );
  INV_X1 U17222 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15608) );
  NOR2_X1 U17223 ( .A1(n15616), .A2(n15608), .ZN(P1_U3316) );
  INV_X1 U17224 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15609) );
  NOR2_X1 U17225 ( .A1(n15616), .A2(n15609), .ZN(P1_U3317) );
  INV_X1 U17226 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15610) );
  NOR2_X1 U17227 ( .A1(n15616), .A2(n15610), .ZN(P1_U3318) );
  INV_X1 U17228 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15611) );
  NOR2_X1 U17229 ( .A1(n15616), .A2(n15611), .ZN(P1_U3319) );
  INV_X1 U17230 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15612) );
  NOR2_X1 U17231 ( .A1(n15616), .A2(n15612), .ZN(P1_U3320) );
  INV_X1 U17232 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15613) );
  NOR2_X1 U17233 ( .A1(n15616), .A2(n15613), .ZN(P1_U3321) );
  INV_X1 U17234 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15614) );
  NOR2_X1 U17235 ( .A1(n15616), .A2(n15614), .ZN(P1_U3322) );
  INV_X1 U17236 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15615) );
  NOR2_X1 U17237 ( .A1(n15616), .A2(n15615), .ZN(P1_U3323) );
  INV_X1 U17238 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U17239 ( .A1(n15700), .A2(n15618), .B1(n15617), .B2(n15698), .ZN(
        P1_U3459) );
  INV_X1 U17240 ( .A(n15619), .ZN(n15621) );
  OAI211_X1 U17241 ( .C1(n6593), .C2(n15682), .A(n15621), .B(n15620), .ZN(
        n15624) );
  AOI211_X1 U17242 ( .C1(n15655), .C2(n15625), .A(n15624), .B(n15623), .ZN(
        n15701) );
  INV_X1 U17243 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U17244 ( .A1(n15700), .A2(n15701), .B1(n15626), .B2(n15698), .ZN(
        P1_U3462) );
  INV_X1 U17245 ( .A(n15636), .ZN(n15638) );
  INV_X1 U17246 ( .A(n15627), .ZN(n15632) );
  OAI22_X1 U17247 ( .A1(n6804), .A2(n15630), .B1(n15629), .B2(n15628), .ZN(
        n15631) );
  NOR4_X1 U17248 ( .A1(n15634), .A2(n15633), .A3(n15632), .A4(n15631), .ZN(
        n15635) );
  OAI21_X1 U17249 ( .B1(n15674), .B2(n15636), .A(n15635), .ZN(n15637) );
  AOI21_X1 U17250 ( .B1(n15678), .B2(n15638), .A(n15637), .ZN(n15702) );
  INV_X1 U17251 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15639) );
  AOI22_X1 U17252 ( .A1(n15700), .A2(n15702), .B1(n15639), .B2(n15698), .ZN(
        P1_U3465) );
  OR4_X1 U17253 ( .A1(n15643), .A2(n15642), .A3(n15641), .A4(n15640), .ZN(
        n15644) );
  AOI21_X1 U17254 ( .B1(n15655), .B2(n15645), .A(n15644), .ZN(n15704) );
  INV_X1 U17255 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U17256 ( .A1(n15700), .A2(n15704), .B1(n15646), .B2(n15698), .ZN(
        P1_U3468) );
  AOI22_X1 U17257 ( .A1(n15647), .A2(n15665), .B1(n15668), .B2(n15666), .ZN(
        n15649) );
  NAND3_X1 U17258 ( .A1(n15650), .A2(n15649), .A3(n15648), .ZN(n15654) );
  NOR2_X1 U17259 ( .A1(n15652), .A2(n15651), .ZN(n15653) );
  AOI211_X1 U17260 ( .C1(n15656), .C2(n15655), .A(n15654), .B(n15653), .ZN(
        n15705) );
  INV_X1 U17261 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U17262 ( .A1(n15700), .A2(n15705), .B1(n15657), .B2(n15698), .ZN(
        P1_U3471) );
  INV_X1 U17263 ( .A(n15674), .ZN(n15688) );
  OAI21_X1 U17264 ( .B1(n15659), .B2(n15682), .A(n15658), .ZN(n15662) );
  INV_X1 U17265 ( .A(n15660), .ZN(n15661) );
  AOI211_X1 U17266 ( .C1(n15688), .C2(n15663), .A(n15662), .B(n15661), .ZN(
        n15707) );
  INV_X1 U17267 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U17268 ( .A1(n15700), .A2(n15707), .B1(n15664), .B2(n15698), .ZN(
        P1_U3474) );
  INV_X1 U17269 ( .A(n15675), .ZN(n15679) );
  AOI22_X1 U17270 ( .A1(n15668), .A2(n15667), .B1(n15666), .B2(n15665), .ZN(
        n15672) );
  INV_X1 U17271 ( .A(n15669), .ZN(n15670) );
  NAND4_X1 U17272 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15677) );
  NOR2_X1 U17273 ( .A1(n15675), .A2(n15674), .ZN(n15676) );
  AOI211_X1 U17274 ( .C1(n15679), .C2(n15678), .A(n15677), .B(n15676), .ZN(
        n15709) );
  INV_X1 U17275 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U17276 ( .A1(n15700), .A2(n15709), .B1(n15680), .B2(n15698), .ZN(
        P1_U3477) );
  OAI21_X1 U17277 ( .B1(n15683), .B2(n15682), .A(n15681), .ZN(n15686) );
  INV_X1 U17278 ( .A(n15684), .ZN(n15685) );
  AOI211_X1 U17279 ( .C1(n15688), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n15710) );
  INV_X1 U17280 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15689) );
  AOI22_X1 U17281 ( .A1(n15700), .A2(n15710), .B1(n15689), .B2(n15698), .ZN(
        P1_U3480) );
  INV_X1 U17282 ( .A(n15690), .ZN(n15697) );
  INV_X1 U17283 ( .A(n15691), .ZN(n15693) );
  OAI211_X1 U17284 ( .C1(n15695), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        n15696) );
  NOR2_X1 U17285 ( .A1(n15697), .A2(n15696), .ZN(n15713) );
  INV_X1 U17286 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15699) );
  AOI22_X1 U17287 ( .A1(n15700), .A2(n15713), .B1(n15699), .B2(n15698), .ZN(
        P1_U3483) );
  AOI22_X1 U17288 ( .A1(n15714), .A2(n15701), .B1(n10686), .B2(n15711), .ZN(
        P1_U3529) );
  AOI22_X1 U17289 ( .A1(n15714), .A2(n15702), .B1(n10685), .B2(n15711), .ZN(
        P1_U3530) );
  AOI22_X1 U17290 ( .A1(n15714), .A2(n15704), .B1(n15703), .B2(n15711), .ZN(
        P1_U3531) );
  AOI22_X1 U17291 ( .A1(n15714), .A2(n15705), .B1(n10691), .B2(n15711), .ZN(
        P1_U3532) );
  AOI22_X1 U17292 ( .A1(n15714), .A2(n15707), .B1(n15706), .B2(n15711), .ZN(
        P1_U3533) );
  AOI22_X1 U17293 ( .A1(n15714), .A2(n15709), .B1(n15708), .B2(n15711), .ZN(
        P1_U3534) );
  AOI22_X1 U17294 ( .A1(n15714), .A2(n15710), .B1(n10696), .B2(n15711), .ZN(
        P1_U3535) );
  AOI22_X1 U17295 ( .A1(n15714), .A2(n15713), .B1(n15712), .B2(n15711), .ZN(
        P1_U3536) );
  NOR2_X1 U17296 ( .A1(n15715), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U17297 ( .B1(n15717), .B2(n6770), .A(n15716), .ZN(n15727) );
  INV_X1 U17298 ( .A(n15718), .ZN(n15726) );
  INV_X1 U17299 ( .A(n15719), .ZN(n15722) );
  OAI21_X1 U17300 ( .B1(n15722), .B2(n15721), .A(n15720), .ZN(n15724) );
  NAND2_X1 U17301 ( .A1(n15724), .A2(n15723), .ZN(n15725) );
  AOI222_X1 U17302 ( .A1(n15727), .A2(n15734), .B1(n15726), .B2(n15747), .C1(
        n15725), .C2(n15744), .ZN(n15729) );
  OAI211_X1 U17303 ( .C1(n15730), .C2(n15753), .A(n15729), .B(n15728), .ZN(
        P2_U3223) );
  AND3_X1 U17304 ( .A1(n15733), .A2(n15732), .A3(n15731), .ZN(n15735) );
  OAI21_X1 U17305 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15750) );
  NAND2_X1 U17306 ( .A1(n15738), .A2(n15737), .ZN(n15741) );
  INV_X1 U17307 ( .A(n15739), .ZN(n15740) );
  NAND2_X1 U17308 ( .A1(n15741), .A2(n15740), .ZN(n15743) );
  NAND2_X1 U17309 ( .A1(n15743), .A2(n15742), .ZN(n15745) );
  NAND2_X1 U17310 ( .A1(n15745), .A2(n15744), .ZN(n15749) );
  NAND2_X1 U17311 ( .A1(n15747), .A2(n15746), .ZN(n15748) );
  AND3_X1 U17312 ( .A1(n15750), .A2(n15749), .A3(n15748), .ZN(n15752) );
  OAI211_X1 U17313 ( .C1(n7497), .C2(n15753), .A(n15752), .B(n15751), .ZN(
        P2_U3226) );
  XNOR2_X1 U17314 ( .A(n15754), .B(n15755), .ZN(n15758) );
  AOI21_X1 U17315 ( .B1(n15758), .B2(n15757), .A(n15756), .ZN(n15794) );
  AOI222_X1 U17316 ( .A1(P2_REG2_REG_2__SCAN_IN), .A2(n14484), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n15760), .C1(n15764), .C2(n15759), .ZN(
        n15770) );
  XNOR2_X1 U17317 ( .A(n15762), .B(n15761), .ZN(n15798) );
  NAND2_X1 U17318 ( .A1(n15764), .A2(n15763), .ZN(n15765) );
  NAND2_X1 U17319 ( .A1(n15765), .A2(n10957), .ZN(n15766) );
  NOR2_X1 U17320 ( .A1(n11369), .A2(n15766), .ZN(n15791) );
  AOI22_X1 U17321 ( .A1(n15768), .A2(n15798), .B1(n15791), .B2(n15767), .ZN(
        n15769) );
  OAI211_X1 U17322 ( .C1(n14484), .C2(n15794), .A(n15770), .B(n15769), .ZN(
        P2_U3263) );
  INV_X1 U17323 ( .A(n15781), .ZN(n15783) );
  NOR2_X1 U17324 ( .A1(n15783), .A2(n15771), .ZN(n15777) );
  AND2_X1 U17325 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15778), .ZN(P2_U3266) );
  AND2_X1 U17326 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15778), .ZN(P2_U3267) );
  AND2_X1 U17327 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15778), .ZN(P2_U3268) );
  NOR2_X1 U17328 ( .A1(n15777), .A2(n15772), .ZN(P2_U3269) );
  NOR2_X1 U17329 ( .A1(n15777), .A2(n15773), .ZN(P2_U3270) );
  AND2_X1 U17330 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15778), .ZN(P2_U3271) );
  AND2_X1 U17331 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15778), .ZN(P2_U3272) );
  AND2_X1 U17332 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15778), .ZN(P2_U3273) );
  AND2_X1 U17333 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15778), .ZN(P2_U3274) );
  AND2_X1 U17334 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15778), .ZN(P2_U3275) );
  AND2_X1 U17335 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15778), .ZN(P2_U3276) );
  NOR2_X1 U17336 ( .A1(n15777), .A2(n15774), .ZN(P2_U3277) );
  AND2_X1 U17337 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15778), .ZN(P2_U3278) );
  AND2_X1 U17338 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15778), .ZN(P2_U3279) );
  AND2_X1 U17339 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15778), .ZN(P2_U3280) );
  AND2_X1 U17340 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15778), .ZN(P2_U3281) );
  AND2_X1 U17341 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15778), .ZN(P2_U3282) );
  NOR2_X1 U17342 ( .A1(n15777), .A2(n15775), .ZN(P2_U3283) );
  AND2_X1 U17343 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15778), .ZN(P2_U3284) );
  AND2_X1 U17344 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15778), .ZN(P2_U3285) );
  AND2_X1 U17345 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15778), .ZN(P2_U3286) );
  AND2_X1 U17346 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15778), .ZN(P2_U3287) );
  AND2_X1 U17347 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15778), .ZN(P2_U3288) );
  AND2_X1 U17348 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15778), .ZN(P2_U3289) );
  AND2_X1 U17349 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15778), .ZN(P2_U3290) );
  AND2_X1 U17350 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15778), .ZN(P2_U3291) );
  AND2_X1 U17351 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15778), .ZN(P2_U3292) );
  AND2_X1 U17352 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15778), .ZN(P2_U3293) );
  NOR2_X1 U17353 ( .A1(n15777), .A2(n15776), .ZN(P2_U3294) );
  AND2_X1 U17354 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15778), .ZN(P2_U3295) );
  AOI22_X1 U17355 ( .A1(n15781), .A2(n15780), .B1(n15779), .B2(n15783), .ZN(
        P2_U3416) );
  AOI21_X1 U17356 ( .B1(n15784), .B2(n15783), .A(n15782), .ZN(P2_U3417) );
  INV_X1 U17357 ( .A(n15785), .ZN(n15789) );
  OAI21_X1 U17358 ( .B1(n15843), .B2(n8535), .A(n15786), .ZN(n15788) );
  AOI211_X1 U17359 ( .C1(n15789), .C2(n15797), .A(n15788), .B(n15787), .ZN(
        n15852) );
  INV_X1 U17360 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U17361 ( .A1(n15850), .A2(n15852), .B1(n15790), .B2(n9003), .ZN(
        P2_U3433) );
  INV_X1 U17362 ( .A(n15791), .ZN(n15792) );
  OAI21_X1 U17363 ( .B1(n15793), .B2(n15843), .A(n15792), .ZN(n15796) );
  INV_X1 U17364 ( .A(n15794), .ZN(n15795) );
  AOI211_X1 U17365 ( .C1(n15798), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15854) );
  AOI22_X1 U17366 ( .A1(n15850), .A2(n15854), .B1(n15799), .B2(n9003), .ZN(
        P2_U3436) );
  INV_X1 U17367 ( .A(n15800), .ZN(n15801) );
  AOI21_X1 U17368 ( .B1(n8920), .B2(n15808), .A(n15801), .ZN(n15806) );
  OAI211_X1 U17369 ( .C1(n15804), .C2(n15843), .A(n15803), .B(n15802), .ZN(
        n15805) );
  NOR2_X1 U17370 ( .A1(n15806), .A2(n15805), .ZN(n15855) );
  INV_X1 U17371 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U17372 ( .A1(n15850), .A2(n15855), .B1(n15807), .B2(n9003), .ZN(
        P2_U3439) );
  INV_X1 U17373 ( .A(n15808), .ZN(n15845) );
  INV_X1 U17374 ( .A(n15809), .ZN(n15814) );
  OAI21_X1 U17375 ( .B1(n15811), .B2(n15843), .A(n15810), .ZN(n15813) );
  AOI211_X1 U17376 ( .C1(n15845), .C2(n15814), .A(n15813), .B(n15812), .ZN(
        n15857) );
  AOI22_X1 U17377 ( .A1(n15850), .A2(n15857), .B1(n15815), .B2(n9003), .ZN(
        P2_U3442) );
  INV_X1 U17378 ( .A(n15816), .ZN(n15817) );
  OAI21_X1 U17379 ( .B1(n15818), .B2(n15845), .A(n15817), .ZN(n15824) );
  AND2_X1 U17380 ( .A1(n15835), .A2(n15819), .ZN(n15820) );
  NOR2_X1 U17381 ( .A1(n15821), .A2(n15820), .ZN(n15822) );
  AND3_X1 U17382 ( .A1(n15824), .A2(n15823), .A3(n15822), .ZN(n15858) );
  INV_X1 U17383 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U17384 ( .A1(n15850), .A2(n15858), .B1(n15825), .B2(n9003), .ZN(
        P2_U3445) );
  AOI21_X1 U17385 ( .B1(n15835), .B2(n15827), .A(n15826), .ZN(n15828) );
  OAI211_X1 U17386 ( .C1(n10269), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        n15831) );
  INV_X1 U17387 ( .A(n15831), .ZN(n15860) );
  INV_X1 U17388 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15832) );
  AOI22_X1 U17389 ( .A1(n15850), .A2(n15860), .B1(n15832), .B2(n9003), .ZN(
        P2_U3448) );
  AOI21_X1 U17390 ( .B1(n15835), .B2(n15834), .A(n15833), .ZN(n15836) );
  OAI211_X1 U17391 ( .C1(n10269), .C2(n15838), .A(n15837), .B(n15836), .ZN(
        n15839) );
  INV_X1 U17392 ( .A(n15839), .ZN(n15862) );
  INV_X1 U17393 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15840) );
  AOI22_X1 U17394 ( .A1(n15850), .A2(n15862), .B1(n15840), .B2(n9003), .ZN(
        P2_U3451) );
  INV_X1 U17395 ( .A(n15841), .ZN(n15842) );
  OAI21_X1 U17396 ( .B1(n8988), .B2(n15843), .A(n15842), .ZN(n15844) );
  AOI21_X1 U17397 ( .B1(n15846), .B2(n15845), .A(n15844), .ZN(n15847) );
  AND2_X1 U17398 ( .A1(n15848), .A2(n15847), .ZN(n15863) );
  AOI22_X1 U17399 ( .A1(n15850), .A2(n15863), .B1(n15849), .B2(n9003), .ZN(
        P2_U3454) );
  INV_X1 U17400 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n15851) );
  AOI22_X1 U17401 ( .A1(n15864), .A2(n15852), .B1(n15851), .B2(n8995), .ZN(
        P2_U3500) );
  AOI22_X1 U17402 ( .A1(n15864), .A2(n15854), .B1(n15853), .B2(n8995), .ZN(
        P2_U3501) );
  AOI22_X1 U17403 ( .A1(n15864), .A2(n15855), .B1(n10897), .B2(n8995), .ZN(
        P2_U3502) );
  AOI22_X1 U17404 ( .A1(n15864), .A2(n15857), .B1(n15856), .B2(n8995), .ZN(
        P2_U3503) );
  AOI22_X1 U17405 ( .A1(n15864), .A2(n15858), .B1(n10900), .B2(n8995), .ZN(
        P2_U3504) );
  AOI22_X1 U17406 ( .A1(n15864), .A2(n15860), .B1(n15859), .B2(n8995), .ZN(
        P2_U3505) );
  AOI22_X1 U17407 ( .A1(n15864), .A2(n15862), .B1(n15861), .B2(n8995), .ZN(
        P2_U3506) );
  AOI22_X1 U17408 ( .A1(n15864), .A2(n15863), .B1(n10904), .B2(n8995), .ZN(
        P2_U3507) );
  NOR2_X1 U17409 ( .A1(P3_U3897), .A2(n15865), .ZN(P3_U3150) );
  INV_X1 U17410 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15877) );
  INV_X1 U17411 ( .A(n15866), .ZN(n15873) );
  OR2_X1 U17412 ( .A1(n15868), .A2(n15867), .ZN(n15872) );
  NAND2_X1 U17413 ( .A1(n15870), .A2(n15869), .ZN(n15871) );
  OAI211_X1 U17414 ( .C1(n15874), .C2(n15873), .A(n15872), .B(n15871), .ZN(
        n15875) );
  INV_X1 U17415 ( .A(n15875), .ZN(n15876) );
  OAI21_X1 U17416 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(P3_U3172) );
  XNOR2_X1 U17417 ( .A(n15879), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n15894) );
  INV_X1 U17418 ( .A(n15880), .ZN(n15882) );
  NAND2_X1 U17419 ( .A1(n15882), .A2(n15881), .ZN(n15883) );
  XNOR2_X1 U17420 ( .A(n15884), .B(n15883), .ZN(n15891) );
  OAI21_X1 U17421 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15885), .A(n11462), .ZN(
        n15889) );
  AOI22_X1 U17422 ( .A1(n15889), .A2(n15888), .B1(n15887), .B2(n15886), .ZN(
        n15890) );
  OAI21_X1 U17423 ( .B1(n15892), .B2(n15891), .A(n15890), .ZN(n15893) );
  AOI21_X1 U17424 ( .B1(n15895), .B2(n15894), .A(n15893), .ZN(n15897) );
  OAI211_X1 U17425 ( .C1(n15899), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        P3_U3191) );
  INV_X1 U17426 ( .A(n15900), .ZN(n15904) );
  INV_X1 U17427 ( .A(n15901), .ZN(n15903) );
  AOI211_X1 U17428 ( .C1(n15905), .C2(n15904), .A(n15903), .B(n15902), .ZN(
        n15944) );
  INV_X1 U17429 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15906) );
  AOI22_X1 U17430 ( .A1(n15943), .A2(n15944), .B1(n15906), .B2(n15941), .ZN(
        P3_U3393) );
  INV_X1 U17431 ( .A(n15907), .ZN(n15911) );
  INV_X1 U17432 ( .A(n15908), .ZN(n15910) );
  AOI211_X1 U17433 ( .C1(n15911), .C2(n15937), .A(n15910), .B(n15909), .ZN(
        n15945) );
  AOI22_X1 U17434 ( .A1(n15943), .A2(n15945), .B1(n15912), .B2(n15941), .ZN(
        P3_U3396) );
  OAI22_X1 U17435 ( .A1(n15914), .A2(n15930), .B1(n15928), .B2(n15913), .ZN(
        n15916) );
  NOR2_X1 U17436 ( .A1(n15916), .A2(n15915), .ZN(n15947) );
  INV_X1 U17437 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U17438 ( .A1(n15943), .A2(n15947), .B1(n15917), .B2(n15941), .ZN(
        P3_U3399) );
  OAI22_X1 U17439 ( .A1(n15919), .A2(n15930), .B1(n15928), .B2(n15918), .ZN(
        n15921) );
  NOR2_X1 U17440 ( .A1(n15921), .A2(n15920), .ZN(n15948) );
  INV_X1 U17441 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U17442 ( .A1(n15943), .A2(n15948), .B1(n15922), .B2(n15941), .ZN(
        P3_U3402) );
  AOI22_X1 U17443 ( .A1(n15924), .A2(n15937), .B1(n15936), .B2(n15923), .ZN(
        n15925) );
  AND2_X1 U17444 ( .A1(n15926), .A2(n15925), .ZN(n15949) );
  INV_X1 U17445 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15927) );
  AOI22_X1 U17446 ( .A1(n15943), .A2(n15949), .B1(n15927), .B2(n15941), .ZN(
        P3_U3405) );
  OAI22_X1 U17447 ( .A1(n15931), .A2(n15930), .B1(n15929), .B2(n15928), .ZN(
        n15933) );
  NOR2_X1 U17448 ( .A1(n15933), .A2(n15932), .ZN(n15950) );
  INV_X1 U17449 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15934) );
  AOI22_X1 U17450 ( .A1(n15943), .A2(n15950), .B1(n15934), .B2(n15941), .ZN(
        P3_U3408) );
  AOI22_X1 U17451 ( .A1(n15938), .A2(n15937), .B1(n15936), .B2(n15935), .ZN(
        n15939) );
  AND2_X1 U17452 ( .A1(n15940), .A2(n15939), .ZN(n15953) );
  INV_X1 U17453 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15942) );
  AOI22_X1 U17454 ( .A1(n15943), .A2(n15953), .B1(n15942), .B2(n15941), .ZN(
        P3_U3411) );
  AOI22_X1 U17455 ( .A1(n15954), .A2(n15944), .B1(n11187), .B2(n15951), .ZN(
        P3_U3460) );
  AOI22_X1 U17456 ( .A1(n15954), .A2(n15945), .B1(n9023), .B2(n15951), .ZN(
        P3_U3461) );
  INV_X1 U17457 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15946) );
  AOI22_X1 U17458 ( .A1(n15954), .A2(n15947), .B1(n15946), .B2(n15951), .ZN(
        P3_U3462) );
  AOI22_X1 U17459 ( .A1(n15954), .A2(n15948), .B1(n11080), .B2(n15951), .ZN(
        P3_U3463) );
  AOI22_X1 U17460 ( .A1(n15954), .A2(n15949), .B1(n7067), .B2(n15951), .ZN(
        P3_U3464) );
  AOI22_X1 U17461 ( .A1(n15954), .A2(n15950), .B1(n11251), .B2(n15951), .ZN(
        P3_U3465) );
  INV_X1 U17462 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15952) );
  AOI22_X1 U17463 ( .A1(n15954), .A2(n15953), .B1(n15952), .B2(n15951), .ZN(
        P3_U3466) );
  AOI21_X1 U17464 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(SUB_1596_U59) );
  OAI21_X1 U17465 ( .B1(n15960), .B2(n15959), .A(n15958), .ZN(SUB_1596_U58) );
  XOR2_X1 U17466 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15961), .Z(SUB_1596_U53) );
  OAI21_X1 U17467 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(SUB_1596_U56) );
  OAI21_X1 U17468 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(n15968) );
  XNOR2_X1 U17469 ( .A(n15968), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17470 ( .B1(n15971), .B2(n15970), .A(n15969), .ZN(SUB_1596_U5) );
  INV_X1 U10190 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8029) );
  INV_X1 U10191 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7968) );
  BUF_X2 U7667 ( .A(n8542), .Z(n7309) );
  AND2_X1 U11547 ( .A1(n9024), .A2(n12742), .ZN(n9345) );
  CLKBUF_X3 U7355 ( .A(n7794), .Z(n6537) );
  NAND2_X1 U7832 ( .A1(n15124), .A2(n15309), .ZN(n15102) );
  CLKBUF_X1 U7305 ( .A(n9815), .Z(n6600) );
  CLKBUF_X1 U7311 ( .A(n12619), .Z(n12642) );
  INV_X1 U7327 ( .A(n11301), .ZN(n11335) );
  CLKBUF_X1 U7343 ( .A(n7931), .Z(n8450) );
  CLKBUF_X1 U7354 ( .A(n7976), .Z(n8145) );
  BUF_X1 U7369 ( .A(n15622), .Z(n6593) );
  CLKBUF_X1 U7399 ( .A(n9556), .Z(n12804) );
  CLKBUF_X1 U7406 ( .A(n13319), .Z(n6821) );
  CLKBUF_X1 U7635 ( .A(n11876), .Z(n6607) );
  CLKBUF_X1 U7639 ( .A(n7767), .Z(n6608) );
  AND2_X1 U7802 ( .A1(n7832), .A2(n10567), .ZN(n15975) );
endmodule

