

module b14_C_SARLock_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828;

  CLKBUF_X1 U2396 ( .A(n4507), .Z(n2153) );
  OAI21_X1 U2397 ( .B1(n2812), .B2(n2811), .A(n4716), .ZN(n4507) );
  NOR4_X1 U2398 ( .A1(n3595), .A2(n3594), .A3(n3983), .A4(n3593), .ZN(n3596)
         );
  OR2_X1 U2399 ( .A1(n2636), .A2(n3414), .ZN(n2644) );
  INV_X2 U2400 ( .A(n3335), .ZN(n3386) );
  INV_X2 U2401 ( .A(n4712), .ZN(n4700) );
  NAND2_X1 U2402 ( .A1(n2687), .A2(n2720), .ZN(n2930) );
  XNOR2_X2 U2403 ( .A(n2680), .B(n2679), .ZN(n2687) );
  XNOR2_X2 U2404 ( .A(n2414), .B(IR_REG_2__SCAN_IN), .ZN(n4489) );
  NOR2_X2 U2405 ( .A1(n2521), .A2(n3163), .ZN(n2541) );
  XNOR2_X2 U2406 ( .A(n2725), .B(n2724), .ZN(n2744) );
  NAND2_X2 U2407 ( .A1(n2748), .A2(IR_REG_31__SCAN_IN), .ZN(n2725) );
  AND2_X4 U2408 ( .A1(n2385), .A2(n2384), .ZN(n2407) );
  XNOR2_X2 U2409 ( .A(n2379), .B(IR_REG_29__SCAN_IN), .ZN(n2385) );
  INV_X1 U2410 ( .A(n2838), .ZN(n2832) );
  CLKBUF_X2 U2411 ( .A(n2405), .Z(n3290) );
  INV_X1 U2412 ( .A(IR_REG_3__SCAN_IN), .ZN(n4369) );
  AND2_X1 U2413 ( .A1(n2240), .A2(n2239), .ZN(n3875) );
  OAI21_X1 U2414 ( .B1(n3214), .B2(n2550), .A(n2549), .ZN(n3264) );
  NAND2_X1 U2415 ( .A1(n2995), .A2(n2994), .ZN(n3037) );
  INV_X1 U2416 ( .A(n2691), .ZN(n2154) );
  INV_X1 U2417 ( .A(n2418), .ZN(n4676) );
  INV_X1 U2418 ( .A(n2841), .ZN(n2831) );
  NOR2_X1 U2419 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  AND4_X1 U2420 ( .A1(n2477), .A2(n2476), .A3(n2475), .A4(n2474), .ZN(n3090)
         );
  NAND2_X1 U2421 ( .A1(n2678), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  BUF_X4 U2422 ( .A(n2415), .Z(n3526) );
  NAND2_X1 U2423 ( .A1(n2610), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  OR2_X1 U2424 ( .A1(n2591), .A2(n2361), .ZN(n2165) );
  AND2_X1 U2425 ( .A1(n4321), .A2(n2579), .ZN(n2366) );
  AND2_X1 U2426 ( .A1(n2372), .A2(n2353), .ZN(n2352) );
  XNOR2_X1 U2427 ( .A(n2295), .B(IR_REG_1__SCAN_IN), .ZN(n4490) );
  AND4_X1 U2428 ( .A1(n2246), .A2(n2245), .A3(n2244), .A4(n2243), .ZN(n2370)
         );
  INV_X1 U2429 ( .A(IR_REG_13__SCAN_IN), .ZN(n2353) );
  NOR2_X1 U2430 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2246)
         );
  NOR2_X1 U2431 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2245)
         );
  NOR2_X1 U2432 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2244)
         );
  NOR2_X1 U2433 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2726)
         );
  INV_X1 U2434 ( .A(IR_REG_20__SCAN_IN), .ZN(n2679) );
  NOR2_X1 U2435 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2369)
         );
  NOR2_X1 U2436 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2243)
         );
  OAI21_X1 U2437 ( .B1(n3421), .B2(n3420), .A(n3327), .ZN(n3477) );
  NAND2_X4 U2438 ( .A1(n2798), .A2(n2797), .ZN(n2838) );
  INV_X4 U2439 ( .A(n2838), .ZN(n2839) );
  NAND3_X4 U2440 ( .A1(n2747), .A2(n2746), .A3(n2765), .ZN(n2798) );
  XNOR2_X2 U2441 ( .A(n2728), .B(IR_REG_25__SCAN_IN), .ZN(n2745) );
  NOR2_X1 U2442 ( .A1(n3694), .A2(n2946), .ZN(n2262) );
  AND2_X1 U2443 ( .A1(n2930), .A2(n2828), .ZN(n3335) );
  NAND2_X1 U2444 ( .A1(n2290), .A2(n2289), .ZN(n2671) );
  NAND2_X1 U2445 ( .A1(n3835), .A2(n3850), .ZN(n2289) );
  NAND2_X1 U2446 ( .A1(n2661), .A2(n2291), .ZN(n2290) );
  NAND2_X1 U2447 ( .A1(n3864), .A2(n3844), .ZN(n2291) );
  INV_X1 U2448 ( .A(n2569), .ZN(n2373) );
  INV_X1 U2449 ( .A(n4512), .ZN(n2333) );
  INV_X1 U2450 ( .A(n2215), .ZN(n2212) );
  NOR2_X1 U2451 ( .A1(n2436), .A2(n2251), .ZN(n2250) );
  INV_X1 U2452 ( .A(n2420), .ZN(n2251) );
  NAND2_X1 U2453 ( .A1(n2418), .A2(n4055), .ZN(n3616) );
  NAND2_X1 U2454 ( .A1(n4680), .A2(n4681), .ZN(n4683) );
  INV_X1 U2455 ( .A(IR_REG_25__SCAN_IN), .ZN(n4286) );
  AND2_X1 U2456 ( .A1(n4318), .A2(n2363), .ZN(n2362) );
  INV_X1 U2457 ( .A(IR_REG_17__SCAN_IN), .ZN(n2363) );
  INV_X1 U2458 ( .A(n2357), .ZN(n2356) );
  AOI21_X1 U2459 ( .B1(n2357), .B2(n2355), .A(n2180), .ZN(n2354) );
  AOI21_X1 U2460 ( .B1(n3201), .B2(n3202), .A(n2179), .ZN(n2357) );
  XNOR2_X1 U2461 ( .A(n2835), .B(n3386), .ZN(n2855) );
  OAI211_X1 U2462 ( .C1(n2391), .C2(IR_REG_28__SCAN_IN), .A(n2393), .B(n2392), 
        .ZN(n2415) );
  NAND2_X1 U2463 ( .A1(n2798), .A2(n4730), .ZN(n2796) );
  NAND2_X1 U2464 ( .A1(n4588), .A2(n4589), .ZN(n4587) );
  XNOR2_X1 U2465 ( .A(n3771), .B(n2292), .ZN(n4600) );
  NOR2_X1 U2466 ( .A1(n3845), .A2(n3831), .ZN(n2670) );
  NOR2_X1 U2467 ( .A1(n3847), .A2(n3869), .ZN(n2660) );
  AND2_X1 U2468 ( .A1(n2510), .A2(n2173), .ZN(n2271) );
  NOR2_X1 U2469 ( .A1(n2262), .A2(n2468), .ZN(n2259) );
  NAND2_X1 U2470 ( .A1(n2682), .A2(n2611), .ZN(n2678) );
  INV_X1 U2471 ( .A(IR_REG_19__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U2472 ( .A1(n3554), .A2(n2714), .ZN(n4702) );
  OR2_X1 U2473 ( .A1(n2757), .A2(n3392), .ZN(n3280) );
  NAND2_X1 U2474 ( .A1(n2374), .A2(n2362), .ZN(n2361) );
  NOR3_X1 U2475 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .A3(
        IR_REG_20__SCAN_IN), .ZN(n2374) );
  INV_X1 U2476 ( .A(n2273), .ZN(n2272) );
  OR2_X1 U2477 ( .A1(n2730), .A2(n2276), .ZN(n2275) );
  NOR2_X1 U2478 ( .A1(n4648), .A2(n4647), .ZN(n4649) );
  NAND2_X1 U2479 ( .A1(n3309), .A2(n2333), .ZN(n2332) );
  AOI21_X1 U2480 ( .B1(n2345), .B2(n2348), .A(n3448), .ZN(n2344) );
  NAND2_X1 U2481 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  OR2_X1 U2482 ( .A1(n4549), .A2(n2470), .ZN(n3736) );
  NAND2_X1 U2483 ( .A1(n3735), .A2(n4546), .ZN(n3737) );
  NOR2_X1 U2484 ( .A1(n3918), .A2(n2642), .ZN(n2241) );
  AND2_X1 U2485 ( .A1(n3899), .A2(n2710), .ZN(n3918) );
  INV_X1 U2486 ( .A(n3637), .ZN(n2235) );
  INV_X1 U2487 ( .A(n3636), .ZN(n2234) );
  NOR2_X1 U2488 ( .A1(n2213), .A2(n3004), .ZN(n2210) );
  NOR2_X1 U2489 ( .A1(n2693), .A2(n2216), .ZN(n2215) );
  INV_X1 U2490 ( .A(n3622), .ZN(n2216) );
  NAND2_X1 U2491 ( .A1(n4020), .A2(n3300), .ZN(n2320) );
  NAND2_X1 U2492 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2688) );
  INV_X1 U2493 ( .A(IR_REG_9__SCAN_IN), .ZN(n4313) );
  INV_X1 U2494 ( .A(IR_REG_7__SCAN_IN), .ZN(n2502) );
  INV_X1 U2495 ( .A(n3507), .ZN(n2338) );
  AND2_X1 U2496 ( .A1(n2339), .A2(n2338), .ZN(n2337) );
  NAND2_X1 U2497 ( .A1(n3104), .A2(n3103), .ZN(n2351) );
  NOR2_X1 U2498 ( .A1(n2604), .A2(n4420), .ZN(n2615) );
  NOR2_X1 U2499 ( .A1(n3497), .A2(n3498), .ZN(n3319) );
  NAND2_X1 U2500 ( .A1(n3042), .A2(n3041), .ZN(n2328) );
  AND2_X1 U2501 ( .A1(n3359), .A2(n3360), .ZN(n2350) );
  NAND2_X1 U2502 ( .A1(n2615), .A2(REG3_REG_20__SCAN_IN), .ZN(n2635) );
  AND2_X1 U2503 ( .A1(n3160), .A2(n3159), .ZN(n3197) );
  XNOR2_X1 U2504 ( .A(n2844), .B(n3335), .ZN(n2849) );
  AOI21_X1 U2505 ( .B1(n2344), .B2(n2341), .A(n2340), .ZN(n2339) );
  INV_X1 U2506 ( .A(n3449), .ZN(n2340) );
  INV_X1 U2507 ( .A(n2345), .ZN(n2341) );
  INV_X1 U2508 ( .A(n2344), .ZN(n2342) );
  AND2_X1 U2509 ( .A1(n3303), .A2(n3302), .ZN(n4512) );
  OR2_X1 U2510 ( .A1(n2421), .A2(n3511), .ZN(n2388) );
  OR2_X1 U2511 ( .A1(n2421), .A2(n3452), .ZN(n2657) );
  NAND2_X1 U2512 ( .A1(n3721), .A2(n3722), .ZN(n3720) );
  INV_X1 U2513 ( .A(n4488), .ZN(n2434) );
  XNOR2_X1 U2514 ( .A(n3729), .B(n3756), .ZN(n2884) );
  NAND2_X1 U2515 ( .A1(n2884), .A2(REG1_REG_4__SCAN_IN), .ZN(n3731) );
  NOR2_X1 U2516 ( .A1(n4527), .A2(n3732), .ZN(n3733) );
  AND2_X1 U2517 ( .A1(n3753), .A2(REG1_REG_5__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U2518 ( .A1(n4587), .A2(n2183), .ZN(n3743) );
  NAND2_X1 U2519 ( .A1(n4590), .A2(n2177), .ZN(n3771) );
  OAI21_X1 U2520 ( .B1(n4612), .B2(n4608), .A(n2294), .ZN(n3775) );
  OR2_X1 U2521 ( .A1(n3774), .A2(REG2_REG_13__SCAN_IN), .ZN(n2294) );
  NAND2_X1 U2522 ( .A1(n2188), .A2(n3791), .ZN(n3786) );
  INV_X1 U2523 ( .A(n2189), .ZN(n2188) );
  AND2_X1 U2524 ( .A1(n3531), .A2(n3660), .ZN(n3829) );
  AOI21_X1 U2525 ( .B1(n3875), .B2(n2652), .A(n2651), .ZN(n3857) );
  AND2_X1 U2526 ( .A1(n3906), .A2(n3888), .ZN(n2651) );
  AOI21_X1 U2527 ( .B1(n3950), .B2(n3564), .A(n3566), .ZN(n3934) );
  NOR2_X1 U2528 ( .A1(n4000), .A2(n2285), .ZN(n2284) );
  INV_X1 U2529 ( .A(n2593), .ZN(n2285) );
  INV_X1 U2530 ( .A(n2283), .ZN(n2282) );
  OAI21_X1 U2531 ( .B1(n4000), .B2(n2288), .A(n2158), .ZN(n2283) );
  AND2_X1 U2532 ( .A1(n3972), .A2(n3973), .ZN(n4000) );
  INV_X1 U2533 ( .A(n4033), .ZN(n4026) );
  NAND2_X1 U2534 ( .A1(n2552), .A2(REG3_REG_14__SCAN_IN), .ZN(n2563) );
  AOI21_X1 U2535 ( .B1(n2266), .B2(n2269), .A(n2178), .ZN(n2263) );
  AOI21_X1 U2536 ( .B1(n2271), .B2(n2156), .A(n2170), .ZN(n2270) );
  AOI21_X1 U2537 ( .B1(n2259), .B2(n2459), .A(n2163), .ZN(n2257) );
  INV_X1 U2538 ( .A(n4051), .ZN(n2247) );
  OR2_X1 U2539 ( .A1(n3831), .A2(n3844), .ZN(n2309) );
  AND2_X1 U2540 ( .A1(n4684), .A2(n4805), .ZN(n4778) );
  AND2_X1 U2541 ( .A1(n2755), .A2(n2923), .ZN(n2760) );
  AND2_X1 U2542 ( .A1(n4710), .A2(n2721), .ZN(n4803) );
  INV_X1 U2543 ( .A(n2796), .ZN(n2810) );
  NOR2_X1 U2544 ( .A1(n2312), .A2(n2361), .ZN(n2311) );
  AND2_X1 U2545 ( .A1(n2364), .A2(n2412), .ZN(n2418) );
  AND3_X1 U2546 ( .A1(n2410), .A2(n2409), .A3(n2408), .ZN(n2364) );
  OAI21_X1 U2547 ( .B1(n3526), .B2(n2434), .A(n2433), .ZN(n3620) );
  NAND2_X1 U2548 ( .A1(n3526), .A2(DATAI_3_), .ZN(n2433) );
  MUX2_X1 U2549 ( .A(n4490), .B(DATAI_1_), .S(n2415), .Z(n4690) );
  NAND2_X1 U2550 ( .A1(n2938), .A2(n2937), .ZN(n2943) );
  INV_X1 U2551 ( .A(n4519), .ZN(n3517) );
  NAND4_X1 U2552 ( .A1(n2428), .A2(n2427), .A3(n2426), .A4(n2425), .ZN(n4046)
         );
  NAND2_X1 U2553 ( .A1(n2785), .A2(REG1_REG_3__SCAN_IN), .ZN(n2883) );
  NOR2_X1 U2554 ( .A1(n4539), .A2(n2461), .ZN(n4538) );
  NAND2_X1 U2555 ( .A1(n4591), .A2(n4592), .ZN(n4590) );
  XNOR2_X1 U2556 ( .A(n3743), .B(n2292), .ZN(n4605) );
  NAND2_X1 U2557 ( .A1(n3786), .A2(n2187), .ZN(n3748) );
  NAND2_X1 U2558 ( .A1(n2189), .A2(n4485), .ZN(n2187) );
  NOR2_X1 U2559 ( .A1(n4649), .A2(n2186), .ZN(n3803) );
  AND2_X1 U2560 ( .A1(n3702), .A2(n3698), .ZN(n4646) );
  AOI21_X1 U2561 ( .B1(n3796), .B2(n2299), .A(n2298), .ZN(n2297) );
  OR2_X1 U2562 ( .A1(n3796), .A2(n3808), .ZN(n2301) );
  AOI21_X1 U2563 ( .B1(n3278), .B2(n3277), .A(n3276), .ZN(n3279) );
  AND2_X1 U2564 ( .A1(n3832), .A2(n3392), .ZN(n3276) );
  NAND2_X1 U2565 ( .A1(n2198), .A2(n3293), .ZN(n4070) );
  NAND2_X1 U2566 ( .A1(n3285), .A2(n4702), .ZN(n2198) );
  OAI21_X1 U2567 ( .B1(n3404), .B2(n4678), .A(n3291), .ZN(n3292) );
  NAND2_X1 U2568 ( .A1(n2678), .A2(n2613), .ZN(n3811) );
  INV_X1 U2569 ( .A(n2682), .ZN(n2612) );
  NOR2_X1 U2570 ( .A1(n2315), .A2(n2361), .ZN(n2314) );
  NAND2_X1 U2571 ( .A1(n2164), .A2(n2366), .ZN(n2315) );
  INV_X1 U2572 ( .A(n3799), .ZN(n3807) );
  NOR2_X1 U2573 ( .A1(n2175), .A2(n2256), .ZN(n2255) );
  INV_X1 U2574 ( .A(n3243), .ZN(n2359) );
  INV_X1 U2575 ( .A(n3201), .ZN(n2355) );
  INV_X1 U2576 ( .A(n3241), .ZN(n2358) );
  XNOR2_X1 U2577 ( .A(n2829), .B(n3386), .ZN(n2894) );
  INV_X1 U2578 ( .A(n3808), .ZN(n2300) );
  NAND2_X1 U2579 ( .A1(n3548), .A2(n2205), .ZN(n2204) );
  INV_X1 U2580 ( .A(n3656), .ZN(n2205) );
  INV_X1 U2581 ( .A(n3662), .ZN(n2206) );
  OR2_X1 U2582 ( .A1(n3877), .A2(n2204), .ZN(n2202) );
  AND2_X1 U2583 ( .A1(n3542), .A2(n3541), .ZN(n3652) );
  NAND2_X1 U2584 ( .A1(n2219), .A2(n2217), .ZN(n3953) );
  NOR2_X1 U2585 ( .A1(n3648), .A2(n2218), .ZN(n2217) );
  INV_X1 U2586 ( .A(n2221), .ZN(n2218) );
  NOR2_X1 U2587 ( .A1(n4361), .A2(n2572), .ZN(n2573) );
  AOI21_X1 U2588 ( .B1(n2224), .B2(n2223), .A(n2222), .ZN(n2221) );
  INV_X1 U2589 ( .A(n3537), .ZN(n2223) );
  NAND2_X1 U2590 ( .A1(n2220), .A2(n2224), .ZN(n2219) );
  INV_X1 U2591 ( .A(n3228), .ZN(n2220) );
  AND2_X1 U2592 ( .A1(n3604), .A2(n3537), .ZN(n3571) );
  AND2_X1 U2593 ( .A1(n3598), .A2(n2182), .ZN(n2232) );
  AOI21_X1 U2594 ( .B1(n3606), .B2(n2232), .A(n2231), .ZN(n2230) );
  INV_X1 U2595 ( .A(n3603), .ZN(n2231) );
  AOI21_X1 U2596 ( .B1(n2268), .B2(n2270), .A(n2267), .ZN(n2266) );
  INV_X1 U2597 ( .A(n4659), .ZN(n2267) );
  INV_X1 U2598 ( .A(n2271), .ZN(n2268) );
  INV_X1 U2599 ( .A(n2270), .ZN(n2269) );
  AND2_X1 U2600 ( .A1(n3095), .A2(n3067), .ZN(n2323) );
  OR2_X1 U2601 ( .A1(n3863), .A2(n3881), .ZN(n2310) );
  NAND2_X1 U2602 ( .A1(n3096), .A2(n2322), .ZN(n3143) );
  AND2_X1 U2603 ( .A1(n2157), .A2(n3156), .ZN(n2322) );
  INV_X1 U2604 ( .A(n3088), .ZN(n3095) );
  NAND2_X1 U2605 ( .A1(n2690), .A2(n3615), .ZN(n4681) );
  INV_X1 U2606 ( .A(IR_REG_16__SCAN_IN), .ZN(n4321) );
  NAND2_X1 U2607 ( .A1(IR_REG_30__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2276) );
  OAI22_X1 U2608 ( .A1(n2367), .A2(n2276), .B1(IR_REG_31__SCAN_IN), .B2(
        IR_REG_30__SCAN_IN), .ZN(n2273) );
  AND2_X1 U2609 ( .A1(n2366), .A2(n4326), .ZN(n2313) );
  INV_X1 U2610 ( .A(IR_REG_23__SCAN_IN), .ZN(n4319) );
  INV_X1 U2611 ( .A(n2362), .ZN(n2360) );
  INV_X1 U2612 ( .A(IR_REG_14__SCAN_IN), .ZN(n2372) );
  INV_X1 U2613 ( .A(n2423), .ZN(n2406) );
  AOI21_X1 U2614 ( .B1(n2347), .B2(n3468), .A(n2346), .ZN(n2345) );
  NOR2_X1 U2615 ( .A1(n3359), .A2(n3360), .ZN(n2346) );
  INV_X1 U2616 ( .A(n2350), .ZN(n2347) );
  NOR2_X1 U2617 ( .A1(n3468), .A2(n2349), .ZN(n2348) );
  INV_X1 U2618 ( .A(n3359), .ZN(n2349) );
  INV_X1 U2619 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4361) );
  INV_X1 U2620 ( .A(n2331), .ZN(n2330) );
  AOI21_X1 U2621 ( .B1(n2161), .B2(n2331), .A(n3310), .ZN(n2329) );
  AND2_X1 U2622 ( .A1(n4497), .A2(n2332), .ZN(n2331) );
  NOR2_X1 U2623 ( .A1(n3073), .A2(n2327), .ZN(n2326) );
  INV_X1 U2624 ( .A(n3046), .ZN(n2327) );
  OR2_X1 U2625 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  OR2_X1 U2626 ( .A1(n2635), .A2(n2382), .ZN(n2636) );
  NAND2_X1 U2627 ( .A1(n3437), .A2(n3436), .ZN(n3341) );
  AND2_X1 U2628 ( .A1(n2721), .A2(n2751), .ZN(n4707) );
  NAND2_X1 U2629 ( .A1(n3299), .A2(n2160), .ZN(n4509) );
  AOI21_X1 U2630 ( .B1(n3299), .B2(n3298), .A(n3309), .ZN(n4511) );
  NAND2_X1 U2631 ( .A1(n3708), .A2(n3709), .ZN(n3707) );
  NAND2_X1 U2632 ( .A1(n3720), .A2(n2784), .ZN(n2881) );
  NAND2_X1 U2633 ( .A1(n4532), .A2(n2168), .ZN(n3759) );
  XNOR2_X1 U2634 ( .A(n3738), .B(n4746), .ZN(n4558) );
  NAND2_X1 U2635 ( .A1(n4578), .A2(n3742), .ZN(n4588) );
  NAND2_X1 U2636 ( .A1(n4616), .A2(n2184), .ZN(n3745) );
  NAND2_X1 U2637 ( .A1(n4634), .A2(n3747), .ZN(n2189) );
  AND2_X1 U2638 ( .A1(n2300), .A2(n2303), .ZN(n2298) );
  NOR2_X1 U2639 ( .A1(n2303), .A2(n2300), .ZN(n2299) );
  AND4_X1 U2640 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n3514)
         );
  AND2_X1 U2641 ( .A1(n3526), .A2(DATAI_28_), .ZN(n3392) );
  AND2_X1 U2642 ( .A1(n3532), .A2(n3523), .ZN(n3572) );
  NAND2_X1 U2643 ( .A1(n2201), .A2(n2199), .ZN(n3282) );
  AOI21_X1 U2644 ( .B1(n2162), .B2(n2204), .A(n2200), .ZN(n2199) );
  NAND2_X1 U2645 ( .A1(n3877), .A2(n2162), .ZN(n2201) );
  INV_X1 U2646 ( .A(n3531), .ZN(n2200) );
  NOR2_X1 U2647 ( .A1(n2662), .A2(n4394), .ZN(n2672) );
  NAND2_X1 U2648 ( .A1(n2202), .A2(n2162), .ZN(n3828) );
  AND2_X1 U2649 ( .A1(n3575), .A2(n3574), .ZN(n3842) );
  INV_X1 U2650 ( .A(n2643), .ZN(n2239) );
  NAND2_X1 U2651 ( .A1(n2242), .A2(n2241), .ZN(n2240) );
  AND2_X1 U2652 ( .A1(n3526), .A2(DATAI_24_), .ZN(n3881) );
  AND2_X1 U2653 ( .A1(n3526), .A2(DATAI_23_), .ZN(n3903) );
  AND4_X1 U2654 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(n3906)
         );
  AND2_X1 U2655 ( .A1(n3526), .A2(DATAI_21_), .ZN(n3937) );
  OR2_X1 U2656 ( .A1(n2280), .A2(n2614), .ZN(n2279) );
  AND2_X1 U2657 ( .A1(n2282), .A2(n2166), .ZN(n2280) );
  NAND2_X1 U2658 ( .A1(n2594), .A2(REG3_REG_18__SCAN_IN), .ZN(n2604) );
  AND2_X1 U2659 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2573), .ZN(n2594) );
  NAND2_X1 U2660 ( .A1(n2219), .A2(n2221), .ZN(n4009) );
  NAND2_X1 U2661 ( .A1(n3261), .A2(n3605), .ZN(n3228) );
  OAI21_X1 U2662 ( .B1(n3138), .B2(n2229), .A(n2227), .ZN(n3261) );
  INV_X1 U2663 ( .A(n2230), .ZN(n2229) );
  AOI21_X1 U2664 ( .B1(n2228), .B2(n2230), .A(n2701), .ZN(n2227) );
  INV_X1 U2665 ( .A(n2232), .ZN(n2228) );
  NAND2_X1 U2666 ( .A1(n2226), .A2(n2230), .ZN(n3539) );
  NAND2_X1 U2667 ( .A1(n3138), .A2(n2232), .ZN(n2226) );
  OAI22_X1 U2668 ( .A1(n3142), .A2(n2540), .B1(n4658), .B2(n3185), .ZN(n3214)
         );
  AND2_X1 U2669 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2381) );
  OAI21_X1 U2670 ( .B1(n3138), .B2(n3606), .A(n3598), .ZN(n3215) );
  INV_X1 U2671 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U2672 ( .A1(n3096), .A2(n2157), .ZN(n4666) );
  OR2_X1 U2673 ( .A1(n2512), .A2(n4215), .ZN(n2521) );
  OAI21_X1 U2674 ( .B1(n3066), .B2(n2156), .A(n2510), .ZN(n3119) );
  INV_X1 U2675 ( .A(n2237), .ZN(n2236) );
  AOI21_X1 U2676 ( .B1(n2237), .B2(n2235), .A(n2234), .ZN(n2233) );
  AND2_X1 U2677 ( .A1(n3631), .A2(n2238), .ZN(n2237) );
  INV_X1 U2678 ( .A(n3082), .ZN(n3067) );
  NAND2_X1 U2679 ( .A1(n3096), .A2(n2323), .ZN(n3128) );
  NOR2_X1 U2680 ( .A1(n2472), .A2(n2471), .ZN(n2482) );
  NOR2_X1 U2681 ( .A1(n2995), .A2(n3029), .ZN(n3096) );
  OAI21_X1 U2682 ( .B1(n2978), .B2(n2209), .A(n2207), .ZN(n2989) );
  AND2_X1 U2683 ( .A1(n3634), .A2(n2208), .ZN(n2207) );
  INV_X1 U2684 ( .A(n2946), .ZN(n3010) );
  NAND2_X1 U2685 ( .A1(n2214), .A2(n3627), .ZN(n3005) );
  NAND2_X1 U2686 ( .A1(n2978), .A2(n2215), .ZN(n2214) );
  AND2_X1 U2687 ( .A1(n2984), .A2(n2915), .ZN(n3011) );
  NAND2_X1 U2688 ( .A1(n2154), .A2(n2250), .ZN(n2248) );
  NAND2_X1 U2689 ( .A1(n4051), .A2(n2250), .ZN(n2249) );
  INV_X1 U2690 ( .A(n2907), .ZN(n2915) );
  NAND2_X1 U2691 ( .A1(n2978), .A2(n3622), .ZN(n2912) );
  NOR2_X1 U2692 ( .A1(n4762), .A2(n3620), .ZN(n2984) );
  OR2_X1 U2693 ( .A1(n4681), .A2(n3613), .ZN(n4671) );
  NAND2_X1 U2694 ( .A1(n4480), .A2(n2791), .ZN(n4678) );
  AND2_X1 U2695 ( .A1(n2772), .A2(n2743), .ZN(n2924) );
  INV_X1 U2696 ( .A(n2840), .ZN(n4706) );
  INV_X1 U2697 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4420) );
  NOR2_X1 U2698 ( .A1(n3907), .A2(n2310), .ZN(n3867) );
  NOR2_X1 U2699 ( .A1(n3907), .A2(n3881), .ZN(n3886) );
  OR2_X1 U2700 ( .A1(n4092), .A2(n3903), .ZN(n3907) );
  OR2_X1 U2701 ( .A1(n3943), .A2(n3929), .ZN(n4092) );
  NAND2_X1 U2702 ( .A1(n3960), .A2(n3944), .ZN(n3943) );
  AND2_X1 U2703 ( .A1(n3984), .A2(n3962), .ZN(n3960) );
  NAND2_X1 U2704 ( .A1(n2319), .A2(n2318), .ZN(n2317) );
  NOR2_X1 U2705 ( .A1(n4495), .A2(n3994), .ZN(n2318) );
  INV_X1 U2706 ( .A(n2320), .ZN(n2319) );
  NOR2_X1 U2707 ( .A1(n4001), .A2(n3424), .ZN(n3984) );
  AOI21_X1 U2708 ( .B1(n4018), .B2(n2593), .A(n2286), .ZN(n3999) );
  INV_X1 U2709 ( .A(n3464), .ZN(n4020) );
  NOR3_X1 U2710 ( .A1(n4122), .A2(n4495), .A3(n4508), .ZN(n4034) );
  NOR2_X1 U2711 ( .A1(n4122), .A2(n4508), .ZN(n4037) );
  INV_X1 U2712 ( .A(n3216), .ZN(n3221) );
  NAND2_X1 U2713 ( .A1(n3222), .A2(n3221), .ZN(n3269) );
  NOR2_X1 U2714 ( .A1(n3143), .A2(n3172), .ZN(n3222) );
  AND2_X1 U2715 ( .A1(n3096), .A2(n3095), .ZN(n4787) );
  INV_X1 U2716 ( .A(n4778), .ZN(n4797) );
  NAND2_X1 U2717 ( .A1(n3011), .A2(n3010), .ZN(n3009) );
  NAND2_X1 U2718 ( .A1(n2307), .A2(n2306), .ZN(n2995) );
  INV_X1 U2719 ( .A(n3009), .ZN(n2307) );
  NAND2_X1 U2720 ( .A1(n2260), .A2(n2261), .ZN(n2998) );
  INV_X1 U2721 ( .A(n2262), .ZN(n2261) );
  OR2_X1 U2722 ( .A1(n3003), .A2(n2459), .ZN(n2260) );
  INV_X1 U2723 ( .A(IR_REG_22__SCAN_IN), .ZN(n2375) );
  INV_X1 U2724 ( .A(IR_REG_26__SCAN_IN), .ZN(n4326) );
  INV_X1 U2725 ( .A(IR_REG_28__SCAN_IN), .ZN(n4328) );
  INV_X1 U2726 ( .A(IR_REG_29__SCAN_IN), .ZN(n4327) );
  INV_X1 U2727 ( .A(IR_REG_27__SCAN_IN), .ZN(n4320) );
  XNOR2_X1 U2728 ( .A(n2689), .B(IR_REG_28__SCAN_IN), .ZN(n2875) );
  INV_X1 U2729 ( .A(IR_REG_15__SCAN_IN), .ZN(n2579) );
  OR2_X1 U2730 ( .A1(n2528), .A2(IR_REG_10__SCAN_IN), .ZN(n2529) );
  NOR2_X1 U2731 ( .A1(n2505), .A2(n2504), .ZN(n2507) );
  AND2_X1 U2732 ( .A1(n2336), .A2(n3506), .ZN(n2335) );
  INV_X1 U2733 ( .A(n3687), .ZN(n3263) );
  AND4_X1 U2734 ( .A1(n2527), .A2(n2526), .A3(n2525), .A4(n2524), .ZN(n3158)
         );
  INV_X1 U2735 ( .A(n3986), .ZN(n3424) );
  XNOR2_X1 U2736 ( .A(n2849), .B(n2850), .ZN(n3429) );
  INV_X1 U2737 ( .A(n3937), .ZN(n3944) );
  INV_X1 U2738 ( .A(n3172), .ZN(n3185) );
  INV_X1 U2739 ( .A(n2343), .ZN(n3447) );
  OAI21_X1 U2740 ( .B1(n3410), .B2(n2348), .A(n2345), .ZN(n2343) );
  AND4_X1 U2741 ( .A1(n2568), .A2(n2567), .A3(n2566), .A4(n2565), .ZN(n4492)
         );
  AND4_X1 U2742 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n2944)
         );
  AOI21_X1 U2743 ( .B1(n3410), .B2(n3360), .A(n3359), .ZN(n3467) );
  INV_X1 U2744 ( .A(n2897), .ZN(n2325) );
  INV_X1 U2745 ( .A(n3691), .ZN(n3080) );
  NAND2_X1 U2746 ( .A1(n3526), .A2(DATAI_20_), .ZN(n3962) );
  OAI21_X1 U2747 ( .B1(n3526), .B2(n2417), .A(n2416), .ZN(n4055) );
  INV_X1 U2748 ( .A(n3995), .ZN(n3502) );
  AND4_X1 U2749 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n4491)
         );
  OAI21_X1 U2750 ( .B1(n3410), .B2(n2342), .A(n2339), .ZN(n3510) );
  AND4_X1 U2751 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n4502)
         );
  AND4_X1 U2752 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n4505)
         );
  INV_X1 U2753 ( .A(n3431), .ZN(n4503) );
  INV_X1 U2754 ( .A(n3519), .ZN(n4514) );
  NAND2_X1 U2755 ( .A1(n2825), .A2(STATE_REG_SCAN_IN), .ZN(n4519) );
  INV_X1 U2756 ( .A(n3514), .ZN(n3845) );
  NAND4_X1 U2757 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .ZN(n3864)
         );
  NAND4_X1 U2758 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n3882)
         );
  AND4_X1 U2759 ( .A1(n2624), .A2(n2623), .A3(n2622), .A4(n2621), .ZN(n3956)
         );
  INV_X1 U2760 ( .A(n4011), .ZN(n3979) );
  INV_X1 U2761 ( .A(n3158), .ZN(n3689) );
  INV_X1 U2762 ( .A(n2944), .ZN(n3695) );
  INV_X1 U2763 ( .A(U4043), .ZN(n3696) );
  NAND4_X1 U2764 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n3697)
         );
  OR2_X1 U2765 ( .A1(n2405), .A2(n2397), .ZN(n2402) );
  AND2_X1 U2766 ( .A1(n2780), .A2(n2779), .ZN(n3702) );
  XNOR2_X1 U2767 ( .A(n2881), .B(n2434), .ZN(n2785) );
  NAND2_X1 U2768 ( .A1(n3755), .A2(n2305), .ZN(n4533) );
  NAND2_X1 U2769 ( .A1(n4533), .A2(n4534), .ZN(n4532) );
  AND2_X1 U2770 ( .A1(n3731), .A2(n3730), .ZN(n4529) );
  XNOR2_X1 U2771 ( .A(n3759), .B(n2304), .ZN(n4543) );
  NOR2_X1 U2772 ( .A1(n4538), .A2(n3734), .ZN(n4549) );
  NAND2_X1 U2773 ( .A1(n4580), .A2(n3769), .ZN(n4591) );
  NAND2_X1 U2774 ( .A1(n4604), .A2(n3744), .ZN(n4617) );
  NAND2_X1 U2775 ( .A1(n4617), .A2(n4618), .ZN(n4616) );
  NAND2_X1 U2776 ( .A1(n4599), .A2(n3773), .ZN(n4612) );
  XNOR2_X1 U2777 ( .A(n3745), .B(n2293), .ZN(n4626) );
  XNOR2_X1 U2778 ( .A(n3775), .B(n2293), .ZN(n4622) );
  NOR2_X1 U2779 ( .A1(n4622), .A2(n3271), .ZN(n4621) );
  NOR2_X1 U2780 ( .A1(n3788), .A2(n3787), .ZN(n4648) );
  AND2_X1 U2781 ( .A1(n2781), .A2(n2780), .ZN(n4645) );
  INV_X1 U2782 ( .A(n3802), .ZN(n2192) );
  INV_X1 U2783 ( .A(n2671), .ZN(n3824) );
  NAND2_X1 U2784 ( .A1(n4018), .A2(n2284), .ZN(n2281) );
  OR2_X1 U2785 ( .A1(n3269), .A2(n3268), .ZN(n4122) );
  NAND2_X1 U2786 ( .A1(n2265), .A2(n2270), .ZN(n4660) );
  NAND2_X1 U2787 ( .A1(n3066), .A2(n2271), .ZN(n2265) );
  NAND2_X1 U2788 ( .A1(n2258), .A2(n2257), .ZN(n2953) );
  OR2_X1 U2789 ( .A1(n4700), .A2(n2931), .ZN(n4693) );
  NAND2_X1 U2790 ( .A1(n4050), .A2(n2420), .ZN(n2977) );
  OR2_X1 U2791 ( .A1(n4692), .A2(n4055), .ZN(n4762) );
  NAND2_X1 U2792 ( .A1(n2810), .A2(n2809), .ZN(n4716) );
  INV_X1 U2793 ( .A(n4828), .ZN(n4826) );
  OAI21_X1 U2794 ( .B1(n4072), .B2(n4778), .A(n2197), .ZN(n2196) );
  NAND2_X1 U2795 ( .A1(n4071), .A2(n4811), .ZN(n2197) );
  AND2_X1 U2796 ( .A1(n2744), .A2(n3399), .ZN(n2774) );
  NAND2_X1 U2797 ( .A1(n2773), .A2(n2810), .ZN(n4729) );
  INV_X1 U2798 ( .A(n2875), .ZN(n4480) );
  XNOR2_X1 U2799 ( .A(n2732), .B(IR_REG_26__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U2800 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2732) );
  AND2_X1 U2801 ( .A1(n2777), .A2(STATE_REG_SCAN_IN), .ZN(n4730) );
  XNOR2_X1 U2802 ( .A(n2685), .B(IR_REG_22__SCAN_IN), .ZN(n4482) );
  INV_X1 U2803 ( .A(IR_REG_21__SCAN_IN), .ZN(n2683) );
  INV_X1 U2804 ( .A(n3811), .ZN(n4484) );
  AND3_X1 U2805 ( .A1(n2371), .A2(n2370), .A3(n2353), .ZN(n2558) );
  AND2_X1 U2806 ( .A1(n2443), .A2(n2432), .ZN(n4488) );
  NAND2_X1 U2807 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2295)
         );
  NAND2_X1 U2808 ( .A1(n2191), .A2(n4646), .ZN(n2190) );
  XNOR2_X1 U2809 ( .A(n3803), .B(n2192), .ZN(n2191) );
  AOI21_X1 U2810 ( .B1(n2302), .B2(n4610), .A(n3812), .ZN(n3813) );
  OR2_X1 U2811 ( .A1(n3819), .A2(n4130), .ZN(n2762) );
  OR2_X1 U2812 ( .A1(n3819), .A2(n4478), .ZN(n2758) );
  OR3_X1 U2813 ( .A1(n3907), .A2(n2310), .A3(n3844), .ZN(n2155) );
  NOR2_X1 U2814 ( .A1(n3690), .A2(n3082), .ZN(n2156) );
  AND2_X1 U2815 ( .A1(n2373), .A2(n2314), .ZN(n2730) );
  AND2_X1 U2816 ( .A1(n2323), .A2(n3129), .ZN(n2157) );
  OR2_X1 U2817 ( .A1(n3979), .A2(n3994), .ZN(n2158) );
  AND2_X1 U2818 ( .A1(n3114), .A2(n3108), .ZN(n2159) );
  AND2_X1 U2819 ( .A1(n3298), .A2(n3309), .ZN(n2160) );
  NOR2_X1 U2820 ( .A1(n2160), .A2(n2181), .ZN(n2161) );
  INV_X1 U2821 ( .A(n3844), .ZN(n3850) );
  AND2_X1 U2822 ( .A1(n3526), .A2(DATAI_26_), .ZN(n3844) );
  NAND2_X1 U2823 ( .A1(n2247), .A2(n2691), .ZN(n4050) );
  AND2_X1 U2824 ( .A1(n2206), .A2(n3829), .ZN(n2162) );
  AND2_X1 U2825 ( .A1(n3693), .A2(n2993), .ZN(n2163) );
  NOR2_X1 U2826 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2413)
         );
  INV_X1 U2827 ( .A(n2371), .ZN(n2457) );
  INV_X1 U2828 ( .A(n2661), .ZN(n3838) );
  AND3_X1 U2829 ( .A1(n2726), .A2(n2375), .A3(n4286), .ZN(n2164) );
  NAND2_X1 U2830 ( .A1(n2376), .A2(IR_REG_31__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U2831 ( .A1(n4706), .A2(n4690), .ZN(n2690) );
  NAND2_X1 U2832 ( .A1(n3502), .A2(n3986), .ZN(n2166) );
  AND2_X1 U2833 ( .A1(n3410), .A2(n2350), .ZN(n2167) );
  OR2_X1 U2834 ( .A1(n4751), .A2(n3758), .ZN(n2168) );
  NOR2_X1 U2835 ( .A1(n3801), .A2(n3800), .ZN(n2169) );
  AND2_X1 U2836 ( .A1(n3164), .A2(n3129), .ZN(n2170) );
  INV_X1 U2837 ( .A(n2203), .ZN(n3858) );
  INV_X1 U2838 ( .A(n2288), .ZN(n2286) );
  NAND2_X1 U2839 ( .A1(n4491), .A2(n4020), .ZN(n2288) );
  INV_X1 U2840 ( .A(IR_REG_30__SCAN_IN), .ZN(n2277) );
  AND2_X1 U2841 ( .A1(n2367), .A2(n2277), .ZN(n2171) );
  AND2_X1 U2842 ( .A1(n2284), .A2(n2287), .ZN(n2172) );
  NAND2_X1 U2843 ( .A1(n4656), .A2(n3121), .ZN(n2173) );
  AND2_X1 U2844 ( .A1(n2202), .A2(n2206), .ZN(n2174) );
  INV_X1 U2845 ( .A(n2614), .ZN(n2287) );
  AND2_X1 U2846 ( .A1(n2695), .A2(n3637), .ZN(n2175) );
  NAND2_X1 U2847 ( .A1(n3690), .A2(n3067), .ZN(n2176) );
  INV_X1 U2848 ( .A(n3760), .ZN(n2304) );
  NOR3_X1 U2849 ( .A1(n3907), .A2(n2310), .A3(n2309), .ZN(n2308) );
  INV_X1 U2850 ( .A(n2993), .ZN(n2306) );
  OAI21_X1 U2851 ( .B1(n3232), .B2(n2571), .A(n2570), .ZN(n4032) );
  NAND2_X1 U2852 ( .A1(n2281), .A2(n2282), .ZN(n3982) );
  INV_X1 U2853 ( .A(n3634), .ZN(n2211) );
  NOR2_X1 U2854 ( .A1(n2591), .A2(IR_REG_17__SCAN_IN), .ZN(n2600) );
  AOI21_X1 U2855 ( .B1(n3934), .B2(n2626), .A(n2625), .ZN(n3915) );
  INV_X1 U2856 ( .A(n3915), .ZN(n2242) );
  NAND2_X1 U2857 ( .A1(n2351), .A2(n3108), .ZN(n3112) );
  NAND2_X1 U2858 ( .A1(n2373), .A2(n2366), .ZN(n2591) );
  OR2_X1 U2859 ( .A1(n4595), .A2(n3770), .ZN(n2177) );
  AND2_X1 U2860 ( .A1(n3158), .A2(n3156), .ZN(n2178) );
  AND2_X1 U2861 ( .A1(n4033), .A2(n2225), .ZN(n2224) );
  XNOR2_X1 U2862 ( .A(n3206), .B(n3335), .ZN(n3243) );
  AND2_X1 U2863 ( .A1(n2359), .A2(n3241), .ZN(n2179) );
  INV_X1 U2864 ( .A(n2701), .ZN(n3592) );
  AND2_X1 U2865 ( .A1(n3243), .A2(n2358), .ZN(n2180) );
  AND2_X1 U2866 ( .A1(n3298), .A2(n2333), .ZN(n2181) );
  INV_X1 U2867 ( .A(n3772), .ZN(n2292) );
  NAND2_X1 U2868 ( .A1(n3687), .A2(n3221), .ZN(n2182) );
  NAND2_X1 U2869 ( .A1(n2328), .A2(n3046), .ZN(n3072) );
  NAND2_X1 U2870 ( .A1(n2264), .A2(n2263), .ZN(n3142) );
  INV_X1 U2871 ( .A(n3647), .ZN(n2222) );
  NAND2_X1 U2872 ( .A1(n2898), .A2(n2324), .ZN(n2938) );
  NAND2_X1 U2873 ( .A1(n2898), .A2(n2897), .ZN(n2902) );
  NAND2_X1 U2874 ( .A1(n2371), .A2(n2370), .ZN(n2547) );
  OR2_X1 U2875 ( .A1(n4595), .A2(n2523), .ZN(n2183) );
  NOR2_X1 U2876 ( .A1(n4122), .A2(n2317), .ZN(n2321) );
  INV_X1 U2877 ( .A(n2316), .ZN(n4019) );
  NOR3_X1 U2878 ( .A1(n4122), .A2(n2320), .A3(n4495), .ZN(n2316) );
  INV_X1 U2879 ( .A(n4736), .ZN(n2293) );
  OR2_X1 U2880 ( .A1(n4739), .A2(n4271), .ZN(n2184) );
  AND2_X1 U2881 ( .A1(n3526), .A2(DATAI_25_), .ZN(n3863) );
  INV_X1 U2882 ( .A(n3831), .ZN(n3403) );
  AND2_X1 U2883 ( .A1(n3526), .A2(DATAI_27_), .ZN(n3831) );
  NAND2_X1 U2884 ( .A1(n2730), .A2(n2367), .ZN(n2185) );
  AND2_X1 U2885 ( .A1(n4652), .A2(n4274), .ZN(n2186) );
  NOR2_X2 U2886 ( .A1(n4003), .A2(n4798), .ZN(n4696) );
  NOR2_X2 U2887 ( .A1(n3748), .A2(REG1_REG_16__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U2888 ( .A1(n2169), .A2(n2190), .ZN(U3258) );
  NAND2_X1 U2889 ( .A1(n4549), .A2(n2470), .ZN(n3735) );
  XNOR2_X1 U2890 ( .A(n3733), .B(n2304), .ZN(n4539) );
  NAND2_X2 U2891 ( .A1(n2193), .A2(n2380), .ZN(n2423) );
  NAND3_X1 U2892 ( .A1(n2380), .A2(n2193), .A3(REG1_REG_1__SCAN_IN), .ZN(n2194) );
  NAND2_X2 U2893 ( .A1(n2384), .A2(n2193), .ZN(n2421) );
  NAND3_X1 U2894 ( .A1(n2384), .A2(n2193), .A3(REG3_REG_1__SCAN_IN), .ZN(n2195) );
  INV_X1 U2895 ( .A(n2385), .ZN(n2193) );
  NAND4_X1 U2896 ( .A1(n2395), .A2(n2195), .A3(n2396), .A4(n2194), .ZN(n2840)
         );
  OR2_X2 U2897 ( .A1(n4070), .A2(n2196), .ZN(n4134) );
  OR2_X1 U2898 ( .A1(n3877), .A2(n3656), .ZN(n2203) );
  INV_X1 U2899 ( .A(n3627), .ZN(n2213) );
  NAND2_X1 U2900 ( .A1(n2210), .A2(n2212), .ZN(n2208) );
  INV_X1 U2901 ( .A(n2210), .ZN(n2209) );
  OAI21_X1 U2902 ( .B1(n3228), .B2(n3233), .A(n3537), .ZN(n4027) );
  NAND2_X1 U2903 ( .A1(n3233), .A2(n3537), .ZN(n2225) );
  OAI21_X1 U2904 ( .B1(n2949), .B2(n2236), .A(n2233), .ZN(n3062) );
  OAI21_X1 U2905 ( .B1(n2949), .B2(n2696), .A(n3637), .ZN(n3087) );
  NAND2_X1 U2906 ( .A1(n2696), .A2(n3637), .ZN(n2238) );
  AOI21_X1 U2907 ( .B1(n3936), .B2(n3654), .A(n3544), .ZN(n3877) );
  OAI21_X1 U2908 ( .B1(n3953), .B2(n3649), .A(n2708), .ZN(n2709) );
  NAND2_X1 U2909 ( .A1(n2692), .A2(n2154), .ZN(n4045) );
  AOI21_X1 U2910 ( .B1(n3282), .B2(n3523), .A(n3281), .ZN(n3283) );
  NAND2_X1 U2911 ( .A1(n2700), .A2(n3609), .ZN(n3138) );
  INV_X1 U2912 ( .A(n2709), .ZN(n3936) );
  NAND2_X1 U2913 ( .A1(n2979), .A2(n3584), .ZN(n2978) );
  NAND2_X1 U2914 ( .A1(n2698), .A2(n3632), .ZN(n3120) );
  NAND2_X1 U2915 ( .A1(n2694), .A2(n3628), .ZN(n2949) );
  NAND2_X1 U2916 ( .A1(n2313), .A2(n2164), .ZN(n2312) );
  NAND2_X1 U2917 ( .A1(n2373), .A2(n2311), .ZN(n2376) );
  INV_X1 U2918 ( .A(n2380), .ZN(n2384) );
  NAND2_X1 U2919 ( .A1(n2730), .A2(n2171), .ZN(n2274) );
  NAND3_X1 U2920 ( .A1(n2370), .A2(n2371), .A3(n2352), .ZN(n2569) );
  AND3_X2 U2921 ( .A1(n2413), .A2(n4369), .A3(n2369), .ZN(n2371) );
  NAND3_X1 U2922 ( .A1(n2249), .A2(n2435), .A3(n2248), .ZN(n2918) );
  NAND2_X1 U2923 ( .A1(n3003), .A2(n2255), .ZN(n2254) );
  NAND2_X1 U2924 ( .A1(n3003), .A2(n2259), .ZN(n2258) );
  NAND2_X1 U2925 ( .A1(n2254), .A2(n2252), .ZN(n3086) );
  INV_X1 U2926 ( .A(n2253), .ZN(n2252) );
  OAI21_X1 U2927 ( .B1(n2175), .B2(n2257), .A(n2480), .ZN(n2253) );
  INV_X1 U2928 ( .A(n2259), .ZN(n2256) );
  NAND2_X1 U2929 ( .A1(n3066), .A2(n2266), .ZN(n2264) );
  NAND3_X1 U2930 ( .A1(n2275), .A2(n2274), .A3(n2272), .ZN(n2380) );
  NAND2_X1 U2931 ( .A1(n4018), .A2(n2172), .ZN(n2278) );
  NAND2_X1 U2932 ( .A1(n2278), .A2(n2279), .ZN(n3950) );
  MUX2_X1 U2933 ( .A(REG2_REG_1__SCAN_IN), .B(n2775), .S(n4490), .Z(n3708) );
  NOR2_X1 U2934 ( .A1(n3795), .A2(n3796), .ZN(n3806) );
  NAND2_X1 U2935 ( .A1(n3795), .A2(n2299), .ZN(n2296) );
  OAI211_X1 U2936 ( .C1(n3795), .C2(n2301), .A(n2297), .B(n2296), .ZN(n2302)
         );
  AND2_X1 U2937 ( .A1(n3807), .A2(REG2_REG_18__SCAN_IN), .ZN(n2303) );
  OR2_X1 U2938 ( .A1(n3757), .A2(n3756), .ZN(n2305) );
  INV_X1 U2939 ( .A(n2308), .ZN(n2757) );
  INV_X1 U2940 ( .A(n2321), .ZN(n4001) );
  NOR2_X1 U2941 ( .A1(n2903), .A2(n2325), .ZN(n2324) );
  XNOR2_X1 U2942 ( .A(n2936), .B(n2935), .ZN(n2903) );
  NAND2_X1 U2943 ( .A1(n2328), .A2(n2326), .ZN(n3075) );
  OAI21_X1 U2944 ( .B1(n3299), .B2(n2330), .A(n2329), .ZN(n3457) );
  NAND2_X1 U2945 ( .A1(n3410), .A2(n2337), .ZN(n2334) );
  NAND2_X1 U2946 ( .A1(n2334), .A2(n2335), .ZN(n3401) );
  NAND3_X1 U2947 ( .A1(n2339), .A2(n2342), .A3(n2338), .ZN(n2336) );
  NAND2_X1 U2948 ( .A1(n2351), .A2(n2159), .ZN(n3155) );
  OAI21_X1 U2949 ( .B1(n3203), .B2(n2356), .A(n2354), .ZN(n3253) );
  OAI21_X1 U2950 ( .B1(n3203), .B2(n3202), .A(n3201), .ZN(n3242) );
  NOR2_X1 U2951 ( .A1(n2591), .A2(n2360), .ZN(n2602) );
  OR2_X1 U2952 ( .A1(n2405), .A2(n2404), .ZN(n2410) );
  OR2_X1 U2953 ( .A1(n2421), .A2(n2398), .ZN(n2400) );
  OAI21_X2 U2954 ( .B1(n3086), .B2(n2492), .A(n2491), .ZN(n3066) );
  OAI21_X2 U2955 ( .B1(n2671), .B2(n2670), .A(n2669), .ZN(n3278) );
  NAND2_X1 U2956 ( .A1(n2391), .A2(IR_REG_27__SCAN_IN), .ZN(n2392) );
  AOI22_X2 U2957 ( .A1(n4032), .A2(n4026), .B1(n4495), .B2(n4013), .ZN(n4018)
         );
  NAND2_X2 U2958 ( .A1(n3488), .A2(n3352), .ZN(n3410) );
  NAND2_X2 U2959 ( .A1(n3489), .A2(n3490), .ZN(n3488) );
  OAI21_X1 U2960 ( .B1(n4706), .B2(n3384), .A(n2845), .ZN(n2850) );
  INV_X4 U2961 ( .A(n3384), .ZN(n2830) );
  NAND2_X4 U2962 ( .A1(n2841), .A2(n4798), .ZN(n3384) );
  AND2_X1 U2963 ( .A1(n3340), .A2(n3339), .ZN(n2365) );
  INV_X1 U2964 ( .A(n4489), .ZN(n2417) );
  AND4_X1 U2965 ( .A1(n4326), .A2(n4328), .A3(n4320), .A4(n4327), .ZN(n2367)
         );
  OR2_X1 U2966 ( .A1(n3882), .A2(n3863), .ZN(n2368) );
  INV_X1 U2967 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2494) );
  INV_X1 U2968 ( .A(n4546), .ZN(n4748) );
  NAND2_X2 U2969 ( .A1(n2929), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U2970 ( .A1(n3618), .A2(n3616), .ZN(n2691) );
  NAND2_X1 U2971 ( .A1(n3620), .A2(n2841), .ZN(n2826) );
  NAND2_X1 U2972 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  NAND2_X1 U2973 ( .A1(n2697), .A2(n2176), .ZN(n2698) );
  INV_X1 U2974 ( .A(IR_REG_18__SCAN_IN), .ZN(n4318) );
  INV_X1 U2975 ( .A(n3113), .ZN(n3114) );
  NAND2_X1 U2976 ( .A1(n4690), .A2(n2841), .ZN(n2842) );
  NOR2_X1 U2977 ( .A1(n2644), .A2(n3471), .ZN(n2653) );
  OR2_X1 U2978 ( .A1(n3123), .A2(n3067), .ZN(n2510) );
  AND2_X1 U2979 ( .A1(n3697), .A2(n4689), .ZN(n4680) );
  OR2_X1 U2980 ( .A1(n2655), .A2(n3512), .ZN(n2662) );
  NAND2_X1 U2981 ( .A1(n2385), .A2(n2380), .ZN(n2405) );
  OR2_X1 U2982 ( .A1(n3514), .A2(n3403), .ZN(n2669) );
  AND2_X1 U2983 ( .A1(n3424), .A2(n3995), .ZN(n2614) );
  OR2_X1 U2984 ( .A1(n4502), .A2(n4495), .ZN(n3647) );
  INV_X1 U2985 ( .A(n4705), .ZN(n4675) );
  AND2_X1 U2986 ( .A1(n3526), .A2(DATAI_22_), .ZN(n3929) );
  AND2_X1 U2987 ( .A1(n4482), .A2(n2720), .ZN(n2791) );
  INV_X1 U2988 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2471) );
  AND2_X1 U2989 ( .A1(n3411), .A2(n3412), .ZN(n3352) );
  INV_X1 U2990 ( .A(n3690), .ZN(n3123) );
  AND2_X1 U2991 ( .A1(n3338), .A2(n3337), .ZN(n3436) );
  INV_X1 U2992 ( .A(n3882), .ZN(n3847) );
  INV_X1 U2993 ( .A(n3432), .ZN(n4504) );
  INV_X1 U2994 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4215) );
  INV_X1 U2995 ( .A(n3292), .ZN(n3293) );
  INV_X1 U2996 ( .A(n3864), .ZN(n3835) );
  INV_X1 U2997 ( .A(n3922), .ZN(n3885) );
  AND2_X1 U2998 ( .A1(n3647), .A2(n3651), .ZN(n4033) );
  INV_X1 U2999 ( .A(n3571), .ZN(n3233) );
  INV_X1 U3000 ( .A(n4696), .ZN(n4040) );
  INV_X1 U3001 ( .A(n3521), .ZN(n3528) );
  INV_X1 U3002 ( .A(n4702), .ZN(n4015) );
  AND2_X1 U3003 ( .A1(n2733), .A2(n2765), .ZN(n2772) );
  NAND2_X1 U3004 ( .A1(n2482), .A2(REG3_REG_8__SCAN_IN), .ZN(n2495) );
  OR2_X1 U3005 ( .A1(n2495), .A2(n2494), .ZN(n2512) );
  AND2_X1 U3006 ( .A1(n2541), .A2(n2381), .ZN(n2552) );
  AND3_X1 U3007 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2462) );
  OR2_X1 U3008 ( .A1(n2563), .A2(n2562), .ZN(n2572) );
  AND4_X1 U3009 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n3404)
         );
  AND4_X1 U3010 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n3442)
         );
  AND4_X1 U3011 ( .A1(n2599), .A2(n2598), .A3(n2597), .A4(n2596), .ZN(n4011)
         );
  NAND2_X1 U3012 ( .A1(n4626), .A2(REG1_REG_14__SCAN_IN), .ZN(n4625) );
  AND2_X1 U3013 ( .A1(n3702), .A2(n3675), .ZN(n4610) );
  INV_X1 U3014 ( .A(n3967), .ZN(n4042) );
  INV_X1 U3015 ( .A(n4678), .ZN(n4655) );
  AOI21_X1 U3016 ( .B1(n2772), .B2(n4362), .A(n2774), .ZN(n2790) );
  INV_X1 U3017 ( .A(n3863), .ZN(n3869) );
  INV_X1 U3018 ( .A(n3881), .ZN(n3888) );
  INV_X1 U3019 ( .A(n4803), .ZN(n4805) );
  INV_X1 U3020 ( .A(n4798), .ZN(n4811) );
  INV_X1 U3021 ( .A(n2765), .ZN(n3399) );
  INV_X1 U3022 ( .A(IR_REG_31__SCAN_IN), .ZN(n2767) );
  AND2_X1 U3023 ( .A1(n2489), .A2(n2479), .ZN(n4546) );
  INV_X1 U3024 ( .A(n4730), .ZN(n2806) );
  OR3_X1 U3025 ( .A1(n2812), .A2(n2796), .A3(n2795), .ZN(n3519) );
  INV_X1 U3026 ( .A(n3404), .ZN(n3832) );
  INV_X1 U3027 ( .A(n3442), .ZN(n3938) );
  INV_X1 U3028 ( .A(n4492), .ZN(n3685) );
  INV_X1 U3029 ( .A(n4610), .ZN(n4639) );
  NAND2_X1 U3030 ( .A1(n3702), .A2(n2875), .ZN(n4653) );
  AND2_X1 U3031 ( .A1(n4693), .A2(n2954), .ZN(n3967) );
  NAND2_X1 U3032 ( .A1(n4828), .A2(n4811), .ZN(n4130) );
  AND2_X2 U3033 ( .A1(n2760), .A2(n2790), .ZN(n4828) );
  NAND2_X1 U3034 ( .A1(n4813), .A2(n4811), .ZN(n4478) );
  NAND2_X1 U3035 ( .A1(n2760), .A2(n2928), .ZN(n4812) );
  INV_X1 U3036 ( .A(n4729), .ZN(n4728) );
  NOR2_X1 U3037 ( .A1(n2509), .A2(n2508), .ZN(n4486) );
  NAND2_X1 U3038 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .ZN(n2377) );
  AND2_X1 U3039 ( .A1(n2688), .A2(n2377), .ZN(n2378) );
  NAND2_X1 U3040 ( .A1(n2391), .A2(n2378), .ZN(n2379) );
  NAND2_X1 U3041 ( .A1(n2407), .A2(REG2_REG_26__SCAN_IN), .ZN(n2390) );
  INV_X1 U3042 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4137) );
  OR2_X1 U3043 ( .A1(n3290), .A2(n4137), .ZN(n2389) );
  NAND2_X1 U3044 ( .A1(n2462), .A2(REG3_REG_6__SCAN_IN), .ZN(n2472) );
  INV_X1 U3045 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U3046 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2382) );
  INV_X1 U3047 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3414) );
  INV_X1 U3048 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U3049 ( .A1(n2653), .A2(REG3_REG_25__SCAN_IN), .ZN(n2655) );
  INV_X1 U3050 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U3051 ( .A1(n2655), .A2(n3512), .ZN(n2383) );
  NAND2_X1 U3052 ( .A1(n2662), .A2(n2383), .ZN(n3511) );
  INV_X1 U3053 ( .A(REG1_REG_26__SCAN_IN), .ZN(n2386) );
  OR2_X1 U3054 ( .A1(n2423), .A2(n2386), .ZN(n2387) );
  NAND2_X1 U3055 ( .A1(n4320), .A2(IR_REG_28__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3056 ( .A1(n2407), .A2(REG2_REG_1__SCAN_IN), .ZN(n2396) );
  INV_X1 U3057 ( .A(n2405), .ZN(n2394) );
  NAND2_X1 U3058 ( .A1(n2394), .A2(REG0_REG_1__SCAN_IN), .ZN(n2395) );
  INV_X1 U3059 ( .A(n4690), .ZN(n2756) );
  NAND2_X1 U3060 ( .A1(n2756), .A2(n2840), .ZN(n3615) );
  INV_X1 U3061 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U3062 ( .A1(n2407), .A2(REG2_REG_0__SCAN_IN), .ZN(n2401) );
  INV_X1 U3063 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2398) );
  INV_X1 U3064 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2800) );
  OR2_X1 U3065 ( .A1(n2423), .A2(n2800), .ZN(n2399) );
  MUX2_X1 U3066 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2415), .Z(n4689) );
  NAND2_X1 U3067 ( .A1(n2840), .A2(n4690), .ZN(n2403) );
  NAND2_X1 U3068 ( .A1(n4683), .A2(n2403), .ZN(n4051) );
  INV_X1 U3069 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3070 ( .A1(n2406), .A2(REG1_REG_2__SCAN_IN), .ZN(n2409) );
  NAND2_X1 U3071 ( .A1(n2407), .A2(REG2_REG_2__SCAN_IN), .ZN(n2408) );
  INV_X1 U3072 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3073 ( .A1(n2421), .A2(n2411), .ZN(n2412) );
  OR2_X1 U3074 ( .A1(n2413), .A2(n2767), .ZN(n2414) );
  NAND2_X1 U3075 ( .A1(n2415), .A2(DATAI_2_), .ZN(n2416) );
  INV_X1 U3076 ( .A(n4055), .ZN(n2419) );
  NAND2_X1 U3077 ( .A1(n4676), .A2(n2419), .ZN(n3618) );
  NAND2_X1 U3078 ( .A1(n2418), .A2(n2419), .ZN(n2420) );
  NAND2_X1 U3079 ( .A1(n2407), .A2(REG2_REG_3__SCAN_IN), .ZN(n2428) );
  OR2_X1 U3080 ( .A1(n2421), .A2(REG3_REG_3__SCAN_IN), .ZN(n2427) );
  INV_X1 U3081 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2422) );
  OR2_X1 U3082 ( .A1(n2423), .A2(n2422), .ZN(n2426) );
  INV_X1 U3083 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2424) );
  OR2_X1 U3084 ( .A1(n2405), .A2(n2424), .ZN(n2425) );
  INV_X1 U3085 ( .A(IR_REG_2__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3086 ( .A1(n2413), .A2(n2429), .ZN(n2430) );
  NAND2_X1 U3087 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3088 ( .A1(n2431), .A2(n4369), .ZN(n2443) );
  OR2_X1 U3089 ( .A1(n2431), .A2(n4369), .ZN(n2432) );
  NOR2_X1 U3090 ( .A1(n4046), .A2(n3620), .ZN(n2436) );
  NAND2_X1 U3091 ( .A1(n4046), .A2(n3620), .ZN(n2435) );
  NAND2_X1 U3092 ( .A1(n2407), .A2(REG2_REG_4__SCAN_IN), .ZN(n2442) );
  INV_X1 U3093 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2437) );
  OR2_X1 U3094 ( .A1(n2405), .A2(n2437), .ZN(n2441) );
  INV_X1 U3095 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3096 ( .A1(n2423), .A2(n2438), .ZN(n2440) );
  XNOR2_X1 U3097 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n2911) );
  OR2_X1 U3098 ( .A1(n2421), .A2(n2911), .ZN(n2439) );
  NAND2_X1 U3099 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2444) );
  XNOR2_X1 U3100 ( .A(n2444), .B(IR_REG_4__SCAN_IN), .ZN(n4487) );
  MUX2_X1 U3101 ( .A(n4487), .B(DATAI_4_), .S(n3526), .Z(n2907) );
  NAND2_X1 U3102 ( .A1(n2944), .A2(n2907), .ZN(n3623) );
  NAND2_X1 U3103 ( .A1(n3695), .A2(n2915), .ZN(n3627) );
  NAND2_X1 U3104 ( .A1(n3623), .A2(n3627), .ZN(n3589) );
  NAND2_X1 U3105 ( .A1(n2918), .A2(n3589), .ZN(n2446) );
  NAND2_X1 U3106 ( .A1(n3695), .A2(n2907), .ZN(n2445) );
  NAND2_X1 U3107 ( .A1(n2446), .A2(n2445), .ZN(n3003) );
  NAND2_X1 U3108 ( .A1(n2407), .A2(REG2_REG_5__SCAN_IN), .ZN(n2456) );
  INV_X1 U3109 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3110 ( .A1(n3290), .A2(n2447), .ZN(n2455) );
  INV_X1 U3111 ( .A(n2462), .ZN(n2451) );
  INV_X1 U3112 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U3113 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2448) );
  NAND2_X1 U3114 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  NAND2_X1 U3115 ( .A1(n2451), .A2(n2450), .ZN(n3012) );
  OR2_X1 U3116 ( .A1(n2421), .A2(n3012), .ZN(n2454) );
  INV_X1 U3117 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2452) );
  OR2_X1 U3118 ( .A1(n2423), .A2(n2452), .ZN(n2453) );
  NAND4_X1 U3119 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n3694)
         );
  NAND2_X1 U3120 ( .A1(n2457), .A2(IR_REG_31__SCAN_IN), .ZN(n2458) );
  XNOR2_X1 U3121 ( .A(n2458), .B(IR_REG_5__SCAN_IN), .ZN(n3753) );
  MUX2_X1 U3122 ( .A(n3753), .B(DATAI_5_), .S(n3526), .Z(n2946) );
  AND2_X1 U3123 ( .A1(n3694), .A2(n2946), .ZN(n2459) );
  NAND2_X1 U3124 ( .A1(n2407), .A2(REG2_REG_6__SCAN_IN), .ZN(n2466) );
  INV_X1 U3125 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2460) );
  OR2_X1 U3126 ( .A1(n3290), .A2(n2460), .ZN(n2465) );
  INV_X1 U3127 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2461) );
  OR2_X1 U3128 ( .A1(n2423), .A2(n2461), .ZN(n2464) );
  OAI21_X1 U3129 ( .B1(n2462), .B2(REG3_REG_6__SCAN_IN), .A(n2472), .ZN(n2996)
         );
  OR2_X1 U3130 ( .A1(n2421), .A2(n2996), .ZN(n2463) );
  NAND4_X1 U3131 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), .ZN(n3693)
         );
  OR2_X1 U3132 ( .A1(n2457), .A2(IR_REG_5__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U3133 ( .A1(n2505), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3134 ( .A(n2467), .B(IR_REG_6__SCAN_IN), .ZN(n3760) );
  MUX2_X1 U3135 ( .A(n3760), .B(DATAI_6_), .S(n3526), .Z(n2993) );
  NOR2_X1 U3136 ( .A1(n3693), .A2(n2993), .ZN(n2468) );
  NAND2_X1 U3137 ( .A1(n2407), .A2(REG2_REG_7__SCAN_IN), .ZN(n2477) );
  INV_X1 U3138 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3139 ( .A1(n3290), .A2(n2469), .ZN(n2476) );
  INV_X1 U3140 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2470) );
  OR2_X1 U3141 ( .A1(n2423), .A2(n2470), .ZN(n2475) );
  AND2_X1 U3142 ( .A1(n2472), .A2(n2471), .ZN(n2473) );
  OR2_X1 U3143 ( .A1(n2473), .A2(n2482), .ZN(n3032) );
  OR2_X1 U3144 ( .A1(n2421), .A2(n3032), .ZN(n2474) );
  OAI21_X1 U3145 ( .B1(n2505), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2478) );
  NAND2_X1 U3146 ( .A1(n2478), .A2(n2502), .ZN(n2489) );
  OR2_X1 U3147 ( .A1(n2478), .A2(n2502), .ZN(n2479) );
  MUX2_X1 U31480 ( .A(n4546), .B(DATAI_7_), .S(n3526), .Z(n3029) );
  NAND2_X1 U31490 ( .A1(n3090), .A2(n3029), .ZN(n2695) );
  INV_X1 U3150 ( .A(n3090), .ZN(n3692) );
  INV_X1 U3151 ( .A(n3029), .ZN(n3022) );
  NAND2_X1 U3152 ( .A1(n3692), .A2(n3022), .ZN(n3637) );
  NAND2_X1 U3153 ( .A1(n3692), .A2(n3029), .ZN(n2480) );
  NAND2_X1 U3154 ( .A1(n2407), .A2(REG2_REG_8__SCAN_IN), .ZN(n2488) );
  INV_X1 U3155 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2481) );
  OR2_X1 U3156 ( .A1(n3290), .A2(n2481), .ZN(n2487) );
  OR2_X1 U3157 ( .A1(n2482), .A2(REG3_REG_8__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3158 ( .A1(n2495), .A2(n2483), .ZN(n3097) );
  OR2_X1 U3159 ( .A1(n2421), .A2(n3097), .ZN(n2486) );
  INV_X1 U3160 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2484) );
  OR2_X1 U3161 ( .A1(n2423), .A2(n2484), .ZN(n2485) );
  NAND4_X1 U3162 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n3691)
         );
  NAND2_X1 U3163 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  XNOR2_X1 U3164 ( .A(n2490), .B(IR_REG_8__SCAN_IN), .ZN(n3763) );
  MUX2_X1 U3165 ( .A(n3763), .B(DATAI_8_), .S(n3526), .Z(n3088) );
  AND2_X1 U3166 ( .A1(n3691), .A2(n3088), .ZN(n2492) );
  NAND2_X1 U3167 ( .A1(n3080), .A2(n3095), .ZN(n2491) );
  NAND2_X1 U3168 ( .A1(n2407), .A2(REG2_REG_9__SCAN_IN), .ZN(n2500) );
  INV_X1 U3169 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2493) );
  OR2_X1 U3170 ( .A1(n3290), .A2(n2493), .ZN(n2499) );
  INV_X1 U3171 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3740) );
  OR2_X1 U3172 ( .A1(n2423), .A2(n3740), .ZN(n2498) );
  NAND2_X1 U3173 ( .A1(n2495), .A2(n2494), .ZN(n2496) );
  NAND2_X1 U3174 ( .A1(n2512), .A2(n2496), .ZN(n3085) );
  OR2_X1 U3175 ( .A1(n2421), .A2(n3085), .ZN(n2497) );
  NAND4_X1 U3176 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n3690)
         );
  INV_X1 U3177 ( .A(IR_REG_6__SCAN_IN), .ZN(n2503) );
  INV_X1 U3178 ( .A(IR_REG_8__SCAN_IN), .ZN(n2501) );
  NAND3_X1 U3179 ( .A1(n2503), .A2(n2502), .A3(n2501), .ZN(n2504) );
  NOR2_X1 U3180 ( .A1(n2507), .A2(n2767), .ZN(n2506) );
  MUX2_X1 U3181 ( .A(n2767), .B(n2506), .S(IR_REG_9__SCAN_IN), .Z(n2509) );
  NAND2_X1 U3182 ( .A1(n2507), .A2(n4313), .ZN(n2528) );
  INV_X1 U3183 ( .A(n2528), .ZN(n2508) );
  MUX2_X1 U3184 ( .A(n4486), .B(DATAI_9_), .S(n3526), .Z(n3082) );
  NAND2_X1 U3185 ( .A1(n2407), .A2(REG2_REG_10__SCAN_IN), .ZN(n2518) );
  INV_X1 U3186 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2511) );
  OR2_X1 U3187 ( .A1(n3290), .A2(n2511), .ZN(n2517) );
  NAND2_X1 U3188 ( .A1(n2512), .A2(n4215), .ZN(n2513) );
  NAND2_X1 U3189 ( .A1(n2521), .A2(n2513), .ZN(n3131) );
  OR2_X1 U3190 ( .A1(n2421), .A2(n3131), .ZN(n2516) );
  INV_X1 U3191 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2514) );
  OR2_X1 U3192 ( .A1(n2423), .A2(n2514), .ZN(n2515) );
  NAND4_X1 U3193 ( .A1(n2518), .A2(n2517), .A3(n2516), .A4(n2515), .ZN(n4656)
         );
  NAND2_X1 U3194 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  XNOR2_X1 U3195 ( .A(n2519), .B(IR_REG_10__SCAN_IN), .ZN(n3767) );
  MUX2_X1 U3196 ( .A(n3767), .B(DATAI_10_), .S(n3526), .Z(n3121) );
  INV_X1 U3197 ( .A(n4656), .ZN(n3164) );
  INV_X1 U3198 ( .A(n3121), .ZN(n3129) );
  NAND2_X1 U3199 ( .A1(n2407), .A2(REG2_REG_11__SCAN_IN), .ZN(n2527) );
  INV_X1 U3200 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2520) );
  OR2_X1 U3201 ( .A1(n3290), .A2(n2520), .ZN(n2526) );
  AND2_X1 U3202 ( .A1(n2521), .A2(n3163), .ZN(n2522) );
  NOR2_X1 U3203 ( .A1(n2541), .A2(n2522), .ZN(n4664) );
  INV_X1 U3204 ( .A(n4664), .ZN(n3168) );
  OR2_X1 U3205 ( .A1(n2421), .A2(n3168), .ZN(n2525) );
  INV_X1 U3206 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2523) );
  OR2_X1 U3207 ( .A1(n2423), .A2(n2523), .ZN(n2524) );
  NAND2_X1 U3208 ( .A1(n2529), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U3209 ( .A(n2537), .B(IR_REG_11__SCAN_IN), .ZN(n4741) );
  MUX2_X1 U32100 ( .A(n4741), .B(DATAI_11_), .S(n3526), .Z(n4667) );
  NAND2_X1 U32110 ( .A1(n3158), .A2(n4667), .ZN(n3609) );
  INV_X1 U32120 ( .A(n4667), .ZN(n3156) );
  NAND2_X1 U32130 ( .A1(n3689), .A2(n3156), .ZN(n3600) );
  NAND2_X1 U32140 ( .A1(n3609), .A2(n3600), .ZN(n4659) );
  NAND2_X1 U32150 ( .A1(n2407), .A2(REG2_REG_12__SCAN_IN), .ZN(n2535) );
  INV_X1 U32160 ( .A(REG0_REG_12__SCAN_IN), .ZN(n2530) );
  OR2_X1 U32170 ( .A1(n3290), .A2(n2530), .ZN(n2534) );
  INV_X1 U32180 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2531) );
  OR2_X1 U32190 ( .A1(n2423), .A2(n2531), .ZN(n2533) );
  XNOR2_X1 U32200 ( .A(n2541), .B(REG3_REG_12__SCAN_IN), .ZN(n3145) );
  OR2_X1 U32210 ( .A1(n2421), .A2(n3145), .ZN(n2532) );
  NAND4_X1 U32220 ( .A1(n2535), .A2(n2534), .A3(n2533), .A4(n2532), .ZN(n3688)
         );
  INV_X1 U32230 ( .A(IR_REG_11__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32240 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  NAND2_X1 U32250 ( .A1(n2538), .A2(IR_REG_31__SCAN_IN), .ZN(n2539) );
  XNOR2_X1 U32260 ( .A(n2539), .B(IR_REG_12__SCAN_IN), .ZN(n3772) );
  MUX2_X1 U32270 ( .A(n3772), .B(DATAI_12_), .S(n3526), .Z(n3172) );
  NOR2_X1 U32280 ( .A1(n3688), .A2(n3172), .ZN(n2540) );
  INV_X1 U32290 ( .A(n3688), .ZN(n4658) );
  NAND2_X1 U32300 ( .A1(n2407), .A2(REG2_REG_13__SCAN_IN), .ZN(n2546) );
  INV_X1 U32310 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4476) );
  OR2_X1 U32320 ( .A1(n3290), .A2(n4476), .ZN(n2545) );
  AOI21_X1 U32330 ( .B1(n2541), .B2(REG3_REG_12__SCAN_IN), .A(
        REG3_REG_13__SCAN_IN), .ZN(n2542) );
  OR2_X1 U32340 ( .A1(n2552), .A2(n2542), .ZN(n3223) );
  OR2_X1 U32350 ( .A1(n2421), .A2(n3223), .ZN(n2544) );
  INV_X1 U32360 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4271) );
  OR2_X1 U32370 ( .A1(n2423), .A2(n4271), .ZN(n2543) );
  NAND4_X1 U32380 ( .A1(n2546), .A2(n2545), .A3(n2544), .A4(n2543), .ZN(n3687)
         );
  NAND2_X1 U32390 ( .A1(n2547), .A2(IR_REG_31__SCAN_IN), .ZN(n2548) );
  XNOR2_X1 U32400 ( .A(n2548), .B(IR_REG_13__SCAN_IN), .ZN(n3774) );
  MUX2_X1 U32410 ( .A(n3774), .B(DATAI_13_), .S(n3526), .Z(n3216) );
  AND2_X1 U32420 ( .A1(n3687), .A2(n3216), .ZN(n2550) );
  NAND2_X1 U32430 ( .A1(n3263), .A2(n3221), .ZN(n2549) );
  NAND2_X1 U32440 ( .A1(n2407), .A2(REG2_REG_14__SCAN_IN), .ZN(n2557) );
  INV_X1 U32450 ( .A(REG0_REG_14__SCAN_IN), .ZN(n2551) );
  OR2_X1 U32460 ( .A1(n3290), .A2(n2551), .ZN(n2556) );
  OR2_X1 U32470 ( .A1(n2552), .A2(REG3_REG_14__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32480 ( .A1(n2563), .A2(n2553), .ZN(n3270) );
  OR2_X1 U32490 ( .A1(n2421), .A2(n3270), .ZN(n2555) );
  INV_X1 U32500 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4367) );
  OR2_X1 U32510 ( .A1(n2423), .A2(n4367), .ZN(n2554) );
  OR2_X1 U32520 ( .A1(n2558), .A2(n2767), .ZN(n2559) );
  XNOR2_X1 U32530 ( .A(n2559), .B(IR_REG_14__SCAN_IN), .ZN(n4736) );
  MUX2_X1 U32540 ( .A(n4736), .B(DATAI_14_), .S(n3526), .Z(n3268) );
  NAND2_X1 U32550 ( .A1(n4505), .A2(n3268), .ZN(n3605) );
  INV_X1 U32560 ( .A(n4505), .ZN(n3686) );
  INV_X1 U32570 ( .A(n3268), .ZN(n3244) );
  NAND2_X1 U32580 ( .A1(n3686), .A2(n3244), .ZN(n3536) );
  NAND2_X1 U32590 ( .A1(n3605), .A2(n3536), .ZN(n2701) );
  NAND2_X1 U32600 ( .A1(n3264), .A2(n2701), .ZN(n2561) );
  NAND2_X1 U32610 ( .A1(n4505), .A2(n3244), .ZN(n2560) );
  NAND2_X1 U32620 ( .A1(n2561), .A2(n2560), .ZN(n3232) );
  NAND2_X1 U32630 ( .A1(n2407), .A2(REG2_REG_15__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32640 ( .A1(n2563), .A2(n2562), .ZN(n2564) );
  NAND2_X1 U32650 ( .A1(n2572), .A2(n2564), .ZN(n4518) );
  OR2_X1 U32660 ( .A1(n2421), .A2(n4518), .ZN(n2567) );
  INV_X1 U32670 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4119) );
  OR2_X1 U32680 ( .A1(n2423), .A2(n4119), .ZN(n2566) );
  INV_X1 U32690 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4471) );
  OR2_X1 U32700 ( .A1(n3290), .A2(n4471), .ZN(n2565) );
  NAND2_X1 U32710 ( .A1(n2569), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U32720 ( .A(n2580), .B(IR_REG_15__SCAN_IN), .ZN(n3778) );
  MUX2_X1 U32730 ( .A(n3778), .B(DATAI_15_), .S(n3526), .Z(n4508) );
  NOR2_X1 U32740 ( .A1(n3685), .A2(n4508), .ZN(n2571) );
  NAND2_X1 U32750 ( .A1(n3685), .A2(n4508), .ZN(n2570) );
  NAND2_X1 U32760 ( .A1(n2407), .A2(REG2_REG_16__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32770 ( .A1(n2572), .A2(n4361), .ZN(n2574) );
  INV_X1 U32780 ( .A(n2573), .ZN(n2583) );
  NAND2_X1 U32790 ( .A1(n2574), .A2(n2583), .ZN(n4501) );
  OR2_X1 U32800 ( .A1(n2421), .A2(n4501), .ZN(n2577) );
  INV_X1 U32810 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4115) );
  OR2_X1 U32820 ( .A1(n2423), .A2(n4115), .ZN(n2576) );
  INV_X1 U32830 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4466) );
  OR2_X1 U32840 ( .A1(n3290), .A2(n4466), .ZN(n2575) );
  NAND2_X1 U32850 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND2_X1 U32860 ( .A1(n2581), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  XNOR2_X1 U32870 ( .A(n2582), .B(IR_REG_16__SCAN_IN), .ZN(n4485) );
  MUX2_X1 U32880 ( .A(n4485), .B(DATAI_16_), .S(n3526), .Z(n4495) );
  NAND2_X1 U32890 ( .A1(n4502), .A2(n4495), .ZN(n3651) );
  INV_X1 U32900 ( .A(n4502), .ZN(n4013) );
  NAND2_X1 U32910 ( .A1(n2407), .A2(REG2_REG_17__SCAN_IN), .ZN(n2590) );
  INV_X1 U32920 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4463) );
  OR2_X1 U32930 ( .A1(n3290), .A2(n4463), .ZN(n2589) );
  INV_X1 U32940 ( .A(n2594), .ZN(n2586) );
  INV_X1 U32950 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32960 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  NAND2_X1 U32970 ( .A1(n2586), .A2(n2585), .ZN(n4021) );
  OR2_X1 U32980 ( .A1(n2421), .A2(n4021), .ZN(n2588) );
  INV_X1 U32990 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4274) );
  OR2_X1 U33000 ( .A1(n2423), .A2(n4274), .ZN(n2587) );
  INV_X1 U33010 ( .A(n4491), .ZN(n3684) );
  NAND2_X1 U33020 ( .A1(n2591), .A2(IR_REG_31__SCAN_IN), .ZN(n2592) );
  XNOR2_X1 U33030 ( .A(n2592), .B(IR_REG_17__SCAN_IN), .ZN(n4732) );
  MUX2_X1 U33040 ( .A(n4732), .B(DATAI_17_), .S(n3526), .Z(n3464) );
  NAND2_X1 U33050 ( .A1(n3684), .A2(n3464), .ZN(n2593) );
  NAND2_X1 U33060 ( .A1(n2407), .A2(REG2_REG_18__SCAN_IN), .ZN(n2599) );
  INV_X1 U33070 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4230) );
  OR2_X1 U33080 ( .A1(n3290), .A2(n4230), .ZN(n2598) );
  OAI21_X1 U33090 ( .B1(n2594), .B2(REG3_REG_18__SCAN_IN), .A(n2604), .ZN(
        n4004) );
  OR2_X1 U33100 ( .A1(n2421), .A2(n4004), .ZN(n2597) );
  INV_X1 U33110 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2595) );
  OR2_X1 U33120 ( .A1(n2423), .A2(n2595), .ZN(n2596) );
  NOR2_X1 U33130 ( .A1(n2600), .A2(n2767), .ZN(n2601) );
  MUX2_X1 U33140 ( .A(n2767), .B(n2601), .S(IR_REG_18__SCAN_IN), .Z(n2603) );
  OR2_X1 U33150 ( .A1(n2603), .A2(n2602), .ZN(n3799) );
  MUX2_X1 U33160 ( .A(n3807), .B(DATAI_18_), .S(n3526), .Z(n3994) );
  NAND2_X1 U33170 ( .A1(n4011), .A2(n3994), .ZN(n3972) );
  INV_X1 U33180 ( .A(n3994), .ZN(n4002) );
  NAND2_X1 U33190 ( .A1(n3979), .A2(n4002), .ZN(n3973) );
  NAND2_X1 U33200 ( .A1(n2407), .A2(REG2_REG_19__SCAN_IN), .ZN(n2609) );
  INV_X1 U33210 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4458) );
  OR2_X1 U33220 ( .A1(n3290), .A2(n4458), .ZN(n2608) );
  INV_X1 U33230 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4104) );
  OR2_X1 U33240 ( .A1(n2423), .A2(n4104), .ZN(n2607) );
  AND2_X1 U33250 ( .A1(n2604), .A2(n4420), .ZN(n2605) );
  OR2_X1 U33260 ( .A1(n2605), .A2(n2615), .ZN(n3987) );
  OR2_X1 U33270 ( .A1(n2421), .A2(n3987), .ZN(n2606) );
  NAND4_X1 U33280 ( .A1(n2609), .A2(n2608), .A3(n2607), .A4(n2606), .ZN(n3995)
         );
  INV_X1 U33290 ( .A(n2602), .ZN(n2610) );
  NAND2_X1 U33300 ( .A1(n2612), .A2(IR_REG_19__SCAN_IN), .ZN(n2613) );
  INV_X1 U33310 ( .A(DATAI_19_), .ZN(n4202) );
  MUX2_X1 U33320 ( .A(n3811), .B(n4202), .S(n3526), .Z(n3986) );
  NAND2_X1 U33330 ( .A1(n2407), .A2(REG2_REG_20__SCAN_IN), .ZN(n2620) );
  INV_X1 U33340 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4454) );
  OR2_X1 U33350 ( .A1(n3290), .A2(n4454), .ZN(n2619) );
  INV_X1 U33360 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4289) );
  OR2_X1 U33370 ( .A1(n2423), .A2(n4289), .ZN(n2618) );
  OR2_X1 U33380 ( .A1(n2615), .A2(REG3_REG_20__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U33390 ( .A1(n2635), .A2(n2616), .ZN(n3482) );
  OR2_X1 U33400 ( .A1(n2421), .A2(n3482), .ZN(n2617) );
  NAND4_X1 U33410 ( .A1(n2620), .A2(n2619), .A3(n2618), .A4(n2617), .ZN(n3939)
         );
  INV_X1 U33420 ( .A(n3962), .ZN(n3328) );
  NAND2_X1 U33430 ( .A1(n3939), .A2(n3328), .ZN(n3564) );
  NOR2_X1 U33440 ( .A1(n3939), .A2(n3328), .ZN(n3566) );
  NAND2_X1 U33450 ( .A1(n2407), .A2(REG2_REG_21__SCAN_IN), .ZN(n2624) );
  INV_X1 U33460 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4450) );
  OR2_X1 U33470 ( .A1(n3290), .A2(n4450), .ZN(n2623) );
  INV_X1 U33480 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4280) );
  OR2_X1 U33490 ( .A1(n2423), .A2(n4280), .ZN(n2622) );
  INV_X1 U33500 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3441) );
  XNOR2_X1 U33510 ( .A(n2635), .B(n3441), .ZN(n3440) );
  OR2_X1 U33520 ( .A1(n2421), .A2(n3440), .ZN(n2621) );
  NAND2_X1 U3353 ( .A1(n3956), .A2(n3944), .ZN(n2626) );
  NOR2_X1 U33540 ( .A1(n3956), .A2(n3944), .ZN(n2625) );
  NAND2_X1 U3355 ( .A1(n2407), .A2(REG2_REG_23__SCAN_IN), .ZN(n2631) );
  INV_X1 U3356 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4445) );
  OR2_X1 U3357 ( .A1(n3290), .A2(n4445), .ZN(n2630) );
  NAND2_X1 U3358 ( .A1(n2636), .A2(n3414), .ZN(n2627) );
  NAND2_X1 U3359 ( .A1(n2644), .A2(n2627), .ZN(n3413) );
  OR2_X1 U3360 ( .A1(n2421), .A2(n3413), .ZN(n2629) );
  INV_X1 U3361 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4418) );
  OR2_X1 U3362 ( .A1(n2423), .A2(n4418), .ZN(n2628) );
  NAND4_X1 U3363 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n3922)
         );
  NOR2_X1 U3364 ( .A1(n3922), .A2(n3903), .ZN(n2642) );
  NAND2_X1 U3365 ( .A1(n2407), .A2(REG2_REG_22__SCAN_IN), .ZN(n2641) );
  INV_X1 U3366 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2632) );
  OR2_X1 U3367 ( .A1(n3290), .A2(n2632), .ZN(n2640) );
  INV_X1 U3368 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2633) );
  OR2_X1 U3369 ( .A1(n2423), .A2(n2633), .ZN(n2639) );
  INV_X1 U3370 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2634) );
  OAI21_X1 U3371 ( .B1(n2635), .B2(n3441), .A(n2634), .ZN(n2637) );
  NAND2_X1 U3372 ( .A1(n2637), .A2(n2636), .ZN(n3927) );
  OR2_X1 U3373 ( .A1(n2421), .A2(n3927), .ZN(n2638) );
  NAND2_X1 U3374 ( .A1(n3442), .A2(n3929), .ZN(n3899) );
  INV_X1 U3375 ( .A(n3929), .ZN(n3492) );
  NAND2_X1 U3376 ( .A1(n3938), .A2(n3492), .ZN(n2710) );
  NAND2_X1 U3377 ( .A1(n3938), .A2(n3929), .ZN(n3895) );
  INV_X1 U3378 ( .A(n3903), .ZN(n3908) );
  OAI22_X1 U3379 ( .A1(n2642), .A2(n3895), .B1(n3885), .B2(n3908), .ZN(n2643)
         );
  NAND2_X1 U3380 ( .A1(n2407), .A2(REG2_REG_24__SCAN_IN), .ZN(n2650) );
  INV_X1 U3381 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4441) );
  OR2_X1 U3382 ( .A1(n3290), .A2(n4441), .ZN(n2649) );
  INV_X1 U3383 ( .A(n2653), .ZN(n2646) );
  NAND2_X1 U3384 ( .A1(n2644), .A2(n3471), .ZN(n2645) );
  NAND2_X1 U3385 ( .A1(n2646), .A2(n2645), .ZN(n3470) );
  OR2_X1 U3386 ( .A1(n2421), .A2(n3470), .ZN(n2648) );
  INV_X1 U3387 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4217) );
  OR2_X1 U3388 ( .A1(n2423), .A2(n4217), .ZN(n2647) );
  INV_X1 U3389 ( .A(n3906), .ZN(n3683) );
  NAND2_X1 U3390 ( .A1(n3683), .A2(n3881), .ZN(n2652) );
  NAND2_X1 U3391 ( .A1(n2407), .A2(REG2_REG_25__SCAN_IN), .ZN(n2659) );
  INV_X1 U3392 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4437) );
  OR2_X1 U3393 ( .A1(n3290), .A2(n4437), .ZN(n2658) );
  OR2_X1 U3394 ( .A1(n2653), .A2(REG3_REG_25__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3395 ( .A1(n2655), .A2(n2654), .ZN(n3452) );
  INV_X1 U3396 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4366) );
  OR2_X1 U3397 ( .A1(n2423), .A2(n4366), .ZN(n2656) );
  AOI21_X1 U3398 ( .B1(n3857), .B2(n2368), .A(n2660), .ZN(n2661) );
  NAND2_X1 U3399 ( .A1(n2407), .A2(REG2_REG_27__SCAN_IN), .ZN(n2668) );
  INV_X1 U3400 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4244) );
  OR2_X1 U3401 ( .A1(n3290), .A2(n4244), .ZN(n2667) );
  INV_X1 U3402 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4287) );
  OR2_X1 U3403 ( .A1(n2423), .A2(n4287), .ZN(n2666) );
  INV_X1 U3404 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4394) );
  INV_X1 U3405 ( .A(n2672), .ZN(n2664) );
  NAND2_X1 U3406 ( .A1(n2662), .A2(n4394), .ZN(n2663) );
  NAND2_X1 U3407 ( .A1(n2664), .A2(n2663), .ZN(n3825) );
  OR2_X1 U3408 ( .A1(n2421), .A2(n3825), .ZN(n2665) );
  NAND2_X1 U3409 ( .A1(n2407), .A2(REG2_REG_28__SCAN_IN), .ZN(n2677) );
  INV_X1 U3410 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4296) );
  OR2_X1 U3411 ( .A1(n3290), .A2(n4296), .ZN(n2676) );
  INV_X1 U3412 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4304) );
  OR2_X1 U3413 ( .A1(n2423), .A2(n4304), .ZN(n2675) );
  NAND2_X1 U3414 ( .A1(n2672), .A2(REG3_REG_28__SCAN_IN), .ZN(n3294) );
  OR2_X1 U3415 ( .A1(n2672), .A2(REG3_REG_28__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3416 ( .A1(n3294), .A2(n2673), .ZN(n3816) );
  OR2_X1 U3417 ( .A1(n2421), .A2(n3816), .ZN(n2674) );
  NAND2_X1 U3418 ( .A1(n3404), .A2(n3392), .ZN(n3532) );
  INV_X1 U3419 ( .A(n3392), .ZN(n3385) );
  NAND2_X1 U3420 ( .A1(n3832), .A2(n3385), .ZN(n3523) );
  XNOR2_X1 U3421 ( .A(n3278), .B(n3572), .ZN(n3815) );
  OAI21_X1 U3422 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U3423 ( .A1(n2682), .A2(n2681), .ZN(n2684) );
  XNOR2_X2 U3424 ( .A(n2684), .B(n2683), .ZN(n2720) );
  NAND2_X1 U3425 ( .A1(n2165), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  XNOR2_X1 U3426 ( .A(n2930), .B(n4482), .ZN(n2686) );
  NAND2_X1 U3427 ( .A1(n2686), .A2(n3811), .ZN(n4684) );
  AND2_X1 U3428 ( .A1(n2687), .A2(n4484), .ZN(n4710) );
  INV_X1 U3429 ( .A(n4482), .ZN(n2721) );
  NAND2_X1 U3430 ( .A1(n2391), .A2(n2688), .ZN(n2689) );
  INV_X1 U3431 ( .A(n3697), .ZN(n4679) );
  NAND2_X1 U3432 ( .A1(n4679), .A2(n4689), .ZN(n3613) );
  NAND2_X1 U3433 ( .A1(n4671), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U3434 ( .A1(n4045), .A2(n3616), .ZN(n2979) );
  XNOR2_X1 U3435 ( .A(n4046), .B(n3620), .ZN(n3584) );
  INV_X1 U3436 ( .A(n4046), .ZN(n3621) );
  NAND2_X1 U3437 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  INV_X1 U3438 ( .A(n3623), .ZN(n2693) );
  AND2_X1 U3439 ( .A1(n3694), .A2(n3010), .ZN(n3004) );
  INV_X1 U3440 ( .A(n3694), .ZN(n2973) );
  NAND2_X1 U3441 ( .A1(n2973), .A2(n2946), .ZN(n3634) );
  NAND2_X1 U3442 ( .A1(n3693), .A2(n2306), .ZN(n3635) );
  NAND2_X1 U3443 ( .A1(n2989), .A2(n3635), .ZN(n2694) );
  INV_X1 U3444 ( .A(n3693), .ZN(n3027) );
  NAND2_X1 U3445 ( .A1(n3027), .A2(n2993), .ZN(n3628) );
  INV_X1 U3446 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U3447 ( .A1(n3080), .A2(n3088), .ZN(n3631) );
  NAND2_X1 U3448 ( .A1(n3691), .A2(n3095), .ZN(n3636) );
  INV_X1 U3449 ( .A(n3062), .ZN(n2697) );
  NAND2_X1 U3450 ( .A1(n3123), .A2(n3082), .ZN(n3632) );
  NAND2_X1 U3451 ( .A1(n4656), .A2(n3129), .ZN(n3599) );
  NAND2_X1 U3452 ( .A1(n3120), .A2(n3599), .ZN(n2699) );
  NAND2_X1 U3453 ( .A1(n3164), .A2(n3121), .ZN(n3602) );
  NAND2_X1 U3454 ( .A1(n2699), .A2(n3602), .ZN(n4654) );
  NAND2_X1 U3455 ( .A1(n4654), .A2(n3600), .ZN(n2700) );
  NOR2_X1 U3456 ( .A1(n3688), .A2(n3185), .ZN(n3606) );
  NAND2_X1 U3457 ( .A1(n3688), .A2(n3185), .ZN(n3598) );
  NAND2_X1 U34580 ( .A1(n3263), .A2(n3216), .ZN(n3603) );
  NAND2_X1 U34590 ( .A1(n4492), .A2(n4508), .ZN(n3604) );
  INV_X1 U3460 ( .A(n4508), .ZN(n3300) );
  NAND2_X1 U3461 ( .A1(n3685), .A2(n3300), .ZN(n3537) );
  NAND2_X1 U3462 ( .A1(n3995), .A2(n3986), .ZN(n2702) );
  AND2_X1 U3463 ( .A1(n3973), .A2(n2702), .ZN(n2703) );
  OR2_X1 U3464 ( .A1(n4491), .A2(n3464), .ZN(n3969) );
  NAND2_X1 U3465 ( .A1(n2703), .A2(n3969), .ZN(n3648) );
  AND2_X1 U3466 ( .A1(n3939), .A2(n3962), .ZN(n3649) );
  NAND2_X1 U34670 ( .A1(n4491), .A2(n3464), .ZN(n3970) );
  NAND2_X1 U3468 ( .A1(n3972), .A2(n3970), .ZN(n2704) );
  NAND2_X1 U34690 ( .A1(n2704), .A2(n2703), .ZN(n2706) );
  NAND2_X1 U3470 ( .A1(n3502), .A2(n3424), .ZN(n2705) );
  NAND2_X1 U34710 ( .A1(n2706), .A2(n2705), .ZN(n3951) );
  NOR2_X1 U3472 ( .A1(n3939), .A2(n3962), .ZN(n2707) );
  OR2_X1 U34730 ( .A1(n3951), .A2(n2707), .ZN(n3542) );
  INV_X1 U3474 ( .A(n3649), .ZN(n3541) );
  INV_X1 U34750 ( .A(n3652), .ZN(n2708) );
  NAND2_X1 U3476 ( .A1(n3956), .A2(n3937), .ZN(n3897) );
  AND2_X1 U34770 ( .A1(n3899), .A2(n3897), .ZN(n3654) );
  NOR2_X1 U3478 ( .A1(n3956), .A2(n3937), .ZN(n3898) );
  INV_X1 U34790 ( .A(n3898), .ZN(n2713) );
  INV_X1 U3480 ( .A(n3899), .ZN(n2712) );
  NOR2_X1 U34810 ( .A1(n3885), .A2(n3903), .ZN(n3558) );
  INV_X1 U3482 ( .A(n2710), .ZN(n2711) );
  NOR2_X1 U34830 ( .A1(n3558), .A2(n2711), .ZN(n3658) );
  OAI21_X1 U3484 ( .B1(n2713), .B2(n2712), .A(n3658), .ZN(n3544) );
  NAND2_X1 U34850 ( .A1(n3885), .A2(n3903), .ZN(n3557) );
  NAND2_X1 U3486 ( .A1(n3906), .A2(n3881), .ZN(n3560) );
  NAND2_X1 U34870 ( .A1(n3557), .A2(n3560), .ZN(n3656) );
  NAND2_X1 U3488 ( .A1(n3847), .A2(n3863), .ZN(n3840) );
  NAND2_X1 U34890 ( .A1(n3835), .A2(n3844), .ZN(n3575) );
  NAND2_X1 U3490 ( .A1(n3840), .A2(n3575), .ZN(n3657) );
  INV_X1 U34910 ( .A(n3657), .ZN(n3548) );
  NAND2_X1 U3492 ( .A1(n3683), .A2(n3888), .ZN(n3859) );
  NAND2_X1 U34930 ( .A1(n3882), .A2(n3869), .ZN(n3559) );
  AND2_X1 U3494 ( .A1(n3859), .A2(n3559), .ZN(n3839) );
  NAND2_X1 U34950 ( .A1(n3864), .A2(n3850), .ZN(n3574) );
  OAI21_X1 U3496 ( .B1(n3657), .B2(n3839), .A(n3574), .ZN(n3662) );
  NAND2_X1 U34970 ( .A1(n3514), .A2(n3831), .ZN(n3531) );
  NAND2_X1 U3498 ( .A1(n3845), .A2(n3403), .ZN(n3660) );
  XNOR2_X1 U34990 ( .A(n3282), .B(n3572), .ZN(n2715) );
  INV_X1 U3500 ( .A(n2687), .ZN(n4483) );
  NAND2_X1 U35010 ( .A1(n4483), .A2(n2720), .ZN(n3554) );
  NAND2_X1 U3502 ( .A1(n4482), .A2(n4484), .ZN(n2714) );
  NAND2_X1 U35030 ( .A1(n2715), .A2(n4702), .ZN(n2723) );
  NAND2_X1 U3504 ( .A1(n2407), .A2(REG2_REG_29__SCAN_IN), .ZN(n2719) );
  INV_X1 U35050 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4303) );
  OR2_X1 U35060 ( .A1(n3290), .A2(n4303), .ZN(n2718) );
  OR2_X1 U35070 ( .A1(n2421), .A2(n3294), .ZN(n2717) );
  INV_X1 U35080 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4301) );
  OR2_X1 U35090 ( .A1(n2423), .A2(n4301), .ZN(n2716) );
  NAND4_X1 U35100 ( .A1(n2719), .A2(n2718), .A3(n2717), .A4(n2716), .ZN(n3682)
         );
  NAND2_X1 U35110 ( .A1(n2875), .A2(n2791), .ZN(n4705) );
  INV_X1 U35120 ( .A(n2720), .ZN(n2751) );
  AND2_X2 U35130 ( .A1(n4707), .A2(n4483), .ZN(n4674) );
  AOI22_X1 U35140 ( .A1(n3682), .A2(n4675), .B1(n3392), .B2(n4674), .ZN(n2722)
         );
  OAI211_X1 U35150 ( .C1(n3514), .C2(n4678), .A(n2723), .B(n2722), .ZN(n3821)
         );
  AOI21_X1 U35160 ( .B1(n3815), .B2(n4797), .A(n3821), .ZN(n2761) );
  OAI21_X2 U35170 ( .B1(n2165), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U35180 ( .A1(n2749), .A2(n4319), .ZN(n2748) );
  INV_X1 U35190 ( .A(IR_REG_24__SCAN_IN), .ZN(n2724) );
  OR2_X1 U35200 ( .A1(n2726), .A2(n2767), .ZN(n2727) );
  NAND2_X1 U35210 ( .A1(n2749), .A2(n2727), .ZN(n2728) );
  NAND2_X1 U35220 ( .A1(n2744), .A2(n2745), .ZN(n2729) );
  MUX2_X1 U35230 ( .A(n2744), .B(n2729), .S(B_REG_SCAN_IN), .Z(n2733) );
  INV_X1 U35240 ( .A(n2730), .ZN(n2731) );
  NOR4_X1 U35250 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2742) );
  NOR4_X1 U35260 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2741) );
  INV_X1 U35270 ( .A(D_REG_27__SCAN_IN), .ZN(n4719) );
  INV_X1 U35280 ( .A(D_REG_6__SCAN_IN), .ZN(n4726) );
  INV_X1 U35290 ( .A(D_REG_28__SCAN_IN), .ZN(n4718) );
  INV_X1 U35300 ( .A(D_REG_10__SCAN_IN), .ZN(n4725) );
  NAND4_X1 U35310 ( .A1(n4719), .A2(n4726), .A3(n4718), .A4(n4725), .ZN(n2739)
         );
  NOR4_X1 U35320 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2737) );
  NOR4_X1 U35330 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2736) );
  NOR4_X1 U35340 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2735) );
  NOR4_X1 U35350 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2734) );
  NAND4_X1 U35360 ( .A1(n2737), .A2(n2736), .A3(n2735), .A4(n2734), .ZN(n2738)
         );
  NOR4_X1 U35370 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(n2739), 
        .A4(n2738), .ZN(n2740) );
  NAND3_X1 U35380 ( .A1(n2742), .A2(n2741), .A3(n2740), .ZN(n2743) );
  INV_X1 U35390 ( .A(n2744), .ZN(n2747) );
  INV_X1 U35400 ( .A(n2745), .ZN(n2746) );
  OR2_X1 U35410 ( .A1(n2749), .A2(n4319), .ZN(n2750) );
  NAND2_X1 U35420 ( .A1(n2748), .A2(n2750), .ZN(n2777) );
  NAND2_X1 U35430 ( .A1(n2687), .A2(n3811), .ZN(n2792) );
  AND2_X1 U35440 ( .A1(n2791), .A2(n2792), .ZN(n2822) );
  NOR2_X1 U35450 ( .A1(n2796), .A2(n2822), .ZN(n2926) );
  NAND2_X1 U35460 ( .A1(n4803), .A2(n2751), .ZN(n2808) );
  NAND2_X1 U35470 ( .A1(n2926), .A2(n2808), .ZN(n2752) );
  NOR2_X1 U35480 ( .A1(n2924), .A2(n2752), .ZN(n2755) );
  INV_X1 U35490 ( .A(D_REG_1__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U35500 ( .A1(n2772), .A2(n4258), .ZN(n2754) );
  NAND2_X1 U35510 ( .A1(n2745), .A2(n3399), .ZN(n2753) );
  NAND2_X1 U35520 ( .A1(n2754), .A2(n2753), .ZN(n2923) );
  INV_X1 U35530 ( .A(D_REG_0__SCAN_IN), .ZN(n4362) );
  INV_X1 U35540 ( .A(n2790), .ZN(n2928) );
  MUX2_X1 U35550 ( .A(n2761), .B(n4296), .S(n4812), .Z(n2759) );
  INV_X1 U35560 ( .A(n4689), .ZN(n4709) );
  NAND2_X1 U35570 ( .A1(n2756), .A2(n4709), .ZN(n4692) );
  INV_X1 U35580 ( .A(n4495), .ZN(n4036) );
  OAI21_X1 U35590 ( .B1(n2308), .B2(n3385), .A(n3280), .ZN(n3819) );
  NAND2_X2 U35600 ( .A1(n2687), .A2(n4707), .ZN(n4798) );
  NAND2_X1 U35610 ( .A1(n2759), .A2(n2758), .ZN(U3514) );
  MUX2_X1 U35620 ( .A(n4304), .B(n2761), .S(n4828), .Z(n2763) );
  NAND2_X1 U35630 ( .A1(n2763), .A2(n2762), .ZN(U3546) );
  INV_X2 U35640 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X4 U35650 ( .A1(n2798), .A2(n2806), .ZN(U4043) );
  INV_X1 U35660 ( .A(DATAI_18_), .ZN(n4221) );
  NAND2_X1 U35670 ( .A1(n3807), .A2(STATE_REG_SCAN_IN), .ZN(n2764) );
  OAI21_X1 U35680 ( .B1(STATE_REG_SCAN_IN), .B2(n4221), .A(n2764), .ZN(U3334)
         );
  INV_X1 U35690 ( .A(DATAI_26_), .ZN(n4421) );
  NAND2_X1 U35700 ( .A1(n2765), .A2(STATE_REG_SCAN_IN), .ZN(n2766) );
  OAI21_X1 U35710 ( .B1(STATE_REG_SCAN_IN), .B2(n4421), .A(n2766), .ZN(U3326)
         );
  INV_X1 U35720 ( .A(DATAI_31_), .ZN(n2769) );
  OR4_X1 U35730 ( .A1(n2185), .A2(IR_REG_30__SCAN_IN), .A3(n2767), .A4(U3149), 
        .ZN(n2768) );
  OAI21_X1 U35740 ( .B1(STATE_REG_SCAN_IN), .B2(n2769), .A(n2768), .ZN(U3321)
         );
  INV_X1 U35750 ( .A(DATAI_24_), .ZN(n2770) );
  MUX2_X1 U35760 ( .A(n2770), .B(n2744), .S(STATE_REG_SCAN_IN), .Z(n2771) );
  INV_X1 U35770 ( .A(n2771), .ZN(U3328) );
  INV_X1 U35780 ( .A(n2772), .ZN(n2773) );
  AOI22_X1 U35790 ( .A1(n4729), .A2(n4362), .B1(n2774), .B2(n4730), .ZN(U3458)
         );
  INV_X1 U35800 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4259) );
  MUX2_X1 U35810 ( .A(REG2_REG_2__SCAN_IN), .B(n4259), .S(n4489), .Z(n3719) );
  INV_X1 U3582 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2775) );
  AND2_X1 U3583 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3709)
         );
  NAND2_X1 U3584 ( .A1(n4490), .A2(REG2_REG_1__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3585 ( .A1(n3707), .A2(n2776), .ZN(n3718) );
  NAND2_X1 U3586 ( .A1(n3719), .A2(n3718), .ZN(n3717) );
  OAI21_X1 U3587 ( .B1(n4259), .B2(n2417), .A(n3717), .ZN(n2879) );
  XOR2_X1 U3588 ( .A(n4488), .B(n2879), .Z(n2880) );
  XNOR2_X1 U3589 ( .A(n2880), .B(REG2_REG_3__SCAN_IN), .ZN(n2788) );
  INV_X1 U3590 ( .A(n2777), .ZN(n2821) );
  NAND2_X1 U3591 ( .A1(n2821), .A2(STATE_REG_SCAN_IN), .ZN(n3679) );
  NAND2_X1 U3592 ( .A1(n2796), .A2(n3679), .ZN(n2780) );
  NAND2_X1 U3593 ( .A1(n2791), .A2(n2777), .ZN(n2778) );
  AND2_X1 U3594 ( .A1(n3526), .A2(n2778), .ZN(n2779) );
  XNOR2_X1 U3595 ( .A(n2391), .B(IR_REG_27__SCAN_IN), .ZN(n4481) );
  INV_X1 U3596 ( .A(n4481), .ZN(n3698) );
  NOR2_X1 U3597 ( .A1(n3698), .A2(n2875), .ZN(n3675) );
  INV_X1 U3598 ( .A(n2779), .ZN(n2781) );
  INV_X1 U3599 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4205) );
  NOR2_X1 U3600 ( .A1(STATE_REG_SCAN_IN), .A2(n4205), .ZN(n2863) );
  NOR2_X1 U3601 ( .A1(n4653), .A2(n2434), .ZN(n2782) );
  AOI211_X1 U3602 ( .C1(n4645), .C2(ADDR_REG_3__SCAN_IN), .A(n2863), .B(n2782), 
        .ZN(n2787) );
  INV_X1 U3603 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4817) );
  MUX2_X1 U3604 ( .A(REG1_REG_2__SCAN_IN), .B(n4817), .S(n4489), .Z(n3722) );
  INV_X1 U3605 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4815) );
  MUX2_X1 U3606 ( .A(REG1_REG_1__SCAN_IN), .B(n4815), .S(n4490), .Z(n3712) );
  AND2_X1 U3607 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3711)
         );
  NAND2_X1 U3608 ( .A1(n3712), .A2(n3711), .ZN(n3710) );
  NAND2_X1 U3609 ( .A1(n4490), .A2(REG1_REG_1__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U3610 ( .A1(n3710), .A2(n2783), .ZN(n3721) );
  NAND2_X1 U3611 ( .A1(n4489), .A2(REG1_REG_2__SCAN_IN), .ZN(n2784) );
  OAI211_X1 U3612 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2785), .A(n4646), .B(n2883), 
        .ZN(n2786) );
  OAI211_X1 U3613 ( .C1(n2788), .C2(n4639), .A(n2787), .B(n2786), .ZN(U3243)
         );
  NOR2_X1 U3614 ( .A1(n2924), .A2(n2923), .ZN(n2789) );
  NAND2_X1 U3615 ( .A1(n2790), .A2(n2789), .ZN(n2812) );
  INV_X1 U3616 ( .A(n2791), .ZN(n2794) );
  NAND2_X1 U3617 ( .A1(n4707), .A2(n2792), .ZN(n2793) );
  NAND2_X1 U3618 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  INV_X1 U3619 ( .A(n2930), .ZN(n2797) );
  NAND2_X1 U3620 ( .A1(n3697), .A2(n2839), .ZN(n2799) );
  AND2_X4 U3621 ( .A1(n2798), .A2(n2930), .ZN(n2841) );
  NAND2_X1 U3622 ( .A1(n4689), .A2(n2841), .ZN(n2846) );
  OAI211_X1 U3623 ( .C1(n2800), .C2(n2798), .A(n2799), .B(n2846), .ZN(n2805)
         );
  INV_X1 U3624 ( .A(n2798), .ZN(n2801) );
  AOI22_X1 U3625 ( .A1(n4689), .A2(n2839), .B1(n2801), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2803) );
  NAND2_X1 U3626 ( .A1(n3697), .A2(n2830), .ZN(n2802) );
  NAND2_X1 U3627 ( .A1(n2803), .A2(n2802), .ZN(n2804) );
  NAND2_X1 U3628 ( .A1(n2805), .A2(n2804), .ZN(n2848) );
  OAI21_X1 U3629 ( .B1(n2805), .B2(n2804), .A(n2848), .ZN(n2873) );
  INV_X1 U3630 ( .A(n2812), .ZN(n2807) );
  NAND2_X1 U3631 ( .A1(n4482), .A2(n3811), .ZN(n2828) );
  NOR3_X1 U3632 ( .A1(n2838), .A2(n2828), .A3(n2806), .ZN(n3676) );
  NAND2_X1 U3633 ( .A1(n2807), .A2(n3676), .ZN(n2861) );
  NOR2_X1 U3634 ( .A1(n2861), .A2(n4480), .ZN(n3431) );
  NAND2_X1 U3635 ( .A1(n2812), .A2(n2808), .ZN(n2824) );
  NAND2_X1 U3636 ( .A1(n2824), .A2(n2926), .ZN(n3430) );
  AOI22_X1 U3637 ( .A1(n3431), .A2(n2840), .B1(REG3_REG_0__SCAN_IN), .B2(n3430), .ZN(n2814) );
  NAND2_X1 U3638 ( .A1(n2810), .A2(n4674), .ZN(n2811) );
  INV_X1 U3639 ( .A(n2808), .ZN(n2809) );
  NAND2_X1 U3640 ( .A1(n2153), .A2(n4689), .ZN(n2813) );
  OAI211_X1 U3641 ( .C1(n3519), .C2(n2873), .A(n2814), .B(n2813), .ZN(U3229)
         );
  NOR2_X1 U3642 ( .A1(n4645), .A2(U4043), .ZN(U3148) );
  INV_X1 U3643 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n2820) );
  INV_X1 U3644 ( .A(REG0_REG_31__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U3645 ( .A1(n2407), .A2(REG2_REG_31__SCAN_IN), .ZN(n2817) );
  INV_X1 U3646 ( .A(REG1_REG_31__SCAN_IN), .ZN(n2815) );
  OR2_X1 U3647 ( .A1(n2423), .A2(n2815), .ZN(n2816) );
  OAI211_X1 U3648 ( .C1(n3290), .C2(n2818), .A(n2817), .B(n2816), .ZN(n4061)
         );
  NAND2_X1 U3649 ( .A1(n4061), .A2(U4043), .ZN(n2819) );
  OAI21_X1 U3650 ( .B1(U4043), .B2(n2820), .A(n2819), .ZN(U3581) );
  NOR2_X1 U3651 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  NAND3_X1 U3652 ( .A1(n2824), .A2(n2823), .A3(n2798), .ZN(n2825) );
  NAND2_X1 U3653 ( .A1(n4046), .A2(n2839), .ZN(n2827) );
  NAND2_X1 U3654 ( .A1(n2827), .A2(n2826), .ZN(n2829) );
  AOI22_X1 U3655 ( .A1(n4046), .A2(n2830), .B1(n2832), .B2(n3620), .ZN(n2895)
         );
  XNOR2_X1 U3656 ( .A(n2894), .B(n2895), .ZN(n2892) );
  NAND2_X1 U3657 ( .A1(n2841), .A2(n4055), .ZN(n2834) );
  NAND2_X1 U3658 ( .A1(n4676), .A2(n2839), .ZN(n2833) );
  OR2_X1 U3659 ( .A1(n2418), .A2(n3384), .ZN(n2837) );
  NAND2_X1 U3660 ( .A1(n4055), .A2(n2839), .ZN(n2836) );
  NAND2_X1 U3661 ( .A1(n2837), .A2(n2836), .ZN(n2856) );
  XNOR2_X1 U3662 ( .A(n2855), .B(n2856), .ZN(n2866) );
  INV_X1 U3663 ( .A(n2866), .ZN(n2854) );
  NAND2_X1 U3664 ( .A1(n2840), .A2(n2832), .ZN(n2843) );
  NAND2_X1 U3665 ( .A1(n2843), .A2(n2842), .ZN(n2844) );
  NAND2_X1 U3666 ( .A1(n4690), .A2(n2839), .ZN(n2845) );
  NAND2_X1 U3667 ( .A1(n2846), .A2(n3335), .ZN(n2847) );
  NAND2_X1 U3668 ( .A1(n2848), .A2(n2847), .ZN(n3428) );
  NAND2_X1 U3669 ( .A1(n3429), .A2(n3428), .ZN(n3427) );
  INV_X1 U3670 ( .A(n2849), .ZN(n2851) );
  NAND2_X1 U3671 ( .A1(n2851), .A2(n2850), .ZN(n2852) );
  NAND2_X1 U3672 ( .A1(n3427), .A2(n2852), .ZN(n2867) );
  INV_X1 U3673 ( .A(n2867), .ZN(n2853) );
  NAND2_X1 U3674 ( .A1(n2854), .A2(n2853), .ZN(n2868) );
  INV_X1 U3675 ( .A(n2855), .ZN(n2858) );
  INV_X1 U3676 ( .A(n2856), .ZN(n2857) );
  NAND2_X1 U3677 ( .A1(n2858), .A2(n2857), .ZN(n2859) );
  NAND2_X1 U3678 ( .A1(n2868), .A2(n2859), .ZN(n2893) );
  XNOR2_X1 U3679 ( .A(n2892), .B(n2893), .ZN(n2860) );
  NAND2_X1 U3680 ( .A1(n2860), .A2(n4514), .ZN(n2865) );
  NOR2_X1 U3681 ( .A1(n2861), .A2(n2875), .ZN(n3432) );
  OAI22_X1 U3682 ( .A1(n2418), .A2(n4504), .B1(n4503), .B2(n2944), .ZN(n2862)
         );
  AOI211_X1 U3683 ( .C1(n3620), .C2(n2153), .A(n2863), .B(n2862), .ZN(n2864)
         );
  OAI211_X1 U3684 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4519), .A(n2865), .B(n2864), 
        .ZN(U3215) );
  INV_X1 U3685 ( .A(n2868), .ZN(n2869) );
  AOI21_X1 U3686 ( .B1(n2866), .B2(n2867), .A(n2869), .ZN(n2872) );
  AOI22_X1 U3687 ( .A1(n2153), .A2(n4055), .B1(n3430), .B2(REG3_REG_2__SCAN_IN), .ZN(n2871) );
  AOI22_X1 U3688 ( .A1(n3431), .A2(n4046), .B1(n3432), .B2(n2840), .ZN(n2870)
         );
  OAI211_X1 U3689 ( .C1(n2872), .C2(n3519), .A(n2871), .B(n2870), .ZN(U3234)
         );
  NAND3_X1 U3690 ( .A1(n2873), .A2(n4480), .A3(n3698), .ZN(n2878) );
  INV_X1 U3691 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2874) );
  AND2_X1 U3692 ( .A1(n4481), .A2(n2874), .ZN(n2876) );
  OR2_X1 U3693 ( .A1(n2876), .A2(n2875), .ZN(n3701) );
  INV_X1 U3694 ( .A(IR_REG_0__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U3695 ( .A1(n3675), .A2(n3709), .B1(n3701), .B2(n3699), .ZN(n2877)
         );
  NAND3_X1 U3696 ( .A1(n2878), .A2(U4043), .A3(n2877), .ZN(n3728) );
  AOI22_X1 U3697 ( .A1(n2880), .A2(REG2_REG_3__SCAN_IN), .B1(n4488), .B2(n2879), .ZN(n3757) );
  XNOR2_X1 U3698 ( .A(n3757), .B(n4487), .ZN(n3754) );
  XOR2_X1 U3699 ( .A(REG2_REG_4__SCAN_IN), .B(n3754), .Z(n2890) );
  INV_X1 U3700 ( .A(n4487), .ZN(n3756) );
  NAND2_X1 U3701 ( .A1(n2881), .A2(n4488), .ZN(n2882) );
  NAND2_X1 U3702 ( .A1(n2883), .A2(n2882), .ZN(n3729) );
  INV_X1 U3703 ( .A(n2884), .ZN(n2885) );
  NAND2_X1 U3704 ( .A1(n2885), .A2(n2438), .ZN(n2886) );
  NAND3_X1 U3705 ( .A1(n4646), .A2(n3731), .A3(n2886), .ZN(n2888) );
  AND2_X1 U3706 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2906) );
  AOI21_X1 U3707 ( .B1(n4645), .B2(ADDR_REG_4__SCAN_IN), .A(n2906), .ZN(n2887)
         );
  OAI211_X1 U3708 ( .C1(n4653), .C2(n3756), .A(n2888), .B(n2887), .ZN(n2889)
         );
  AOI21_X1 U3709 ( .B1(n4610), .B2(n2890), .A(n2889), .ZN(n2891) );
  NAND2_X1 U3710 ( .A1(n3728), .A2(n2891), .ZN(U3244) );
  NAND2_X1 U3711 ( .A1(n2893), .A2(n2892), .ZN(n2898) );
  INV_X1 U3712 ( .A(n2894), .ZN(n2896) );
  NAND2_X1 U3713 ( .A1(n2896), .A2(n2895), .ZN(n2897) );
  OAI22_X1 U3714 ( .A1(n2944), .A2(n2838), .B1(n2831), .B2(n2915), .ZN(n2899)
         );
  XNOR2_X1 U3715 ( .A(n2899), .B(n3386), .ZN(n2936) );
  OR2_X1 U3716 ( .A1(n2944), .A2(n3384), .ZN(n2901) );
  NAND2_X1 U3717 ( .A1(n2907), .A2(n2839), .ZN(n2900) );
  NAND2_X1 U3718 ( .A1(n2901), .A2(n2900), .ZN(n2935) );
  AOI21_X1 U3719 ( .B1(n2902), .B2(n2903), .A(n3519), .ZN(n2904) );
  NAND2_X1 U3720 ( .A1(n2904), .A2(n2938), .ZN(n2909) );
  OAI22_X1 U3721 ( .A1(n2973), .A2(n4503), .B1(n4504), .B2(n3621), .ZN(n2905)
         );
  AOI211_X1 U3722 ( .C1(n2907), .C2(n2153), .A(n2906), .B(n2905), .ZN(n2908)
         );
  OAI211_X1 U3723 ( .C1(n4519), .C2(n2911), .A(n2909), .B(n2908), .ZN(U3227)
         );
  OAI21_X1 U3724 ( .B1(n2984), .B2(n2915), .A(n4811), .ZN(n2910) );
  NOR2_X1 U3725 ( .A1(n2910), .A2(n3011), .ZN(n4772) );
  NOR2_X1 U3726 ( .A1(n4716), .A2(n2911), .ZN(n2922) );
  INV_X1 U3727 ( .A(n3589), .ZN(n2919) );
  XNOR2_X1 U3728 ( .A(n2912), .B(n2919), .ZN(n2917) );
  INV_X1 U3729 ( .A(n4674), .ZN(n4010) );
  NAND2_X1 U3730 ( .A1(n4046), .A2(n4655), .ZN(n2914) );
  NAND2_X1 U3731 ( .A1(n3694), .A2(n4675), .ZN(n2913) );
  OAI211_X1 U3732 ( .C1(n4010), .C2(n2915), .A(n2914), .B(n2913), .ZN(n2916)
         );
  AOI21_X1 U3733 ( .B1(n2917), .B2(n4702), .A(n2916), .ZN(n2921) );
  XNOR2_X1 U3734 ( .A(n2918), .B(n2919), .ZN(n4771) );
  INV_X1 U3735 ( .A(n4684), .ZN(n4703) );
  NAND2_X1 U3736 ( .A1(n4771), .A2(n4703), .ZN(n2920) );
  NAND2_X1 U3737 ( .A1(n2921), .A2(n2920), .ZN(n4776) );
  AOI211_X1 U3738 ( .C1(n4772), .C2(n3811), .A(n2922), .B(n4776), .ZN(n2933)
         );
  INV_X1 U3739 ( .A(n2923), .ZN(n2927) );
  INV_X1 U3740 ( .A(n2924), .ZN(n2925) );
  NAND4_X1 U3741 ( .A1(n2928), .A2(n2927), .A3(n2926), .A4(n2925), .ZN(n2929)
         );
  OR2_X1 U3742 ( .A1(n2930), .A2(n3811), .ZN(n2931) );
  INV_X1 U3743 ( .A(n4693), .ZN(n4701) );
  AOI22_X1 U3744 ( .A1(n4771), .A2(n4701), .B1(REG2_REG_4__SCAN_IN), .B2(n4700), .ZN(n2932) );
  OAI21_X1 U3745 ( .B1(n2933), .B2(n4700), .A(n2932), .ZN(U3286) );
  NAND2_X1 U3746 ( .A1(n3696), .A2(DATAO_REG_21__SCAN_IN), .ZN(n2934) );
  OAI21_X1 U3747 ( .B1(n3956), .B2(n3696), .A(n2934), .ZN(U3571) );
  NAND2_X1 U3748 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3749 ( .A1(n3694), .A2(n2839), .ZN(n2940) );
  NAND2_X1 U3750 ( .A1(n2946), .A2(n2841), .ZN(n2939) );
  NAND2_X1 U3751 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  XNOR2_X1 U3752 ( .A(n2941), .B(n3386), .ZN(n2962) );
  AOI22_X1 U3753 ( .A1(n3694), .A2(n2830), .B1(n2839), .B2(n2946), .ZN(n2960)
         );
  XNOR2_X1 U3754 ( .A(n2962), .B(n2960), .ZN(n2942) );
  NAND2_X1 U3755 ( .A1(n2943), .A2(n2942), .ZN(n2964) );
  OAI211_X1 U3756 ( .C1(n2943), .C2(n2942), .A(n2964), .B(n4514), .ZN(n2948)
         );
  AND2_X1 U3757 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4531) );
  OAI22_X1 U3758 ( .A1(n2944), .A2(n4504), .B1(n4503), .B2(n3027), .ZN(n2945)
         );
  AOI211_X1 U3759 ( .C1(n2946), .C2(n2153), .A(n4531), .B(n2945), .ZN(n2947)
         );
  OAI211_X1 U3760 ( .C1(n4519), .C2(n3012), .A(n2948), .B(n2947), .ZN(U3224)
         );
  XNOR2_X1 U3761 ( .A(n2949), .B(n2175), .ZN(n2952) );
  AOI22_X1 U3762 ( .A1(n3691), .A2(n4675), .B1(n4674), .B2(n3029), .ZN(n2950)
         );
  OAI21_X1 U3763 ( .B1(n3027), .B2(n4678), .A(n2950), .ZN(n2951) );
  AOI21_X1 U3764 ( .B1(n2952), .B2(n4702), .A(n2951), .ZN(n4783) );
  XNOR2_X1 U3765 ( .A(n2953), .B(n2175), .ZN(n4786) );
  OR2_X1 U3766 ( .A1(n4700), .A2(n4684), .ZN(n2954) );
  INV_X1 U3767 ( .A(n2995), .ZN(n2956) );
  INV_X1 U3768 ( .A(n3096), .ZN(n2955) );
  OAI211_X1 U3769 ( .C1(n2956), .C2(n3022), .A(n2955), .B(n4811), .ZN(n4782)
         );
  OR2_X1 U3770 ( .A1(n4700), .A2(n4484), .ZN(n4003) );
  NOR2_X1 U3771 ( .A1(n4782), .A2(n4003), .ZN(n2958) );
  INV_X1 U3772 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3752) );
  OAI22_X1 U3773 ( .A1(n4712), .A2(n3752), .B1(n3032), .B2(n4716), .ZN(n2957)
         );
  AOI211_X1 U3774 ( .C1(n4786), .C2(n4042), .A(n2958), .B(n2957), .ZN(n2959)
         );
  OAI21_X1 U3775 ( .B1(n4783), .B2(n4700), .A(n2959), .ZN(U3283) );
  INV_X1 U3776 ( .A(n2960), .ZN(n2961) );
  NAND2_X1 U3777 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  NAND2_X1 U3778 ( .A1(n2964), .A2(n2963), .ZN(n3019) );
  NAND2_X1 U3779 ( .A1(n3693), .A2(n2832), .ZN(n2966) );
  NAND2_X1 U3780 ( .A1(n2993), .A2(n2841), .ZN(n2965) );
  NAND2_X1 U3781 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  XNOR2_X1 U3782 ( .A(n2967), .B(n3386), .ZN(n3017) );
  NAND2_X1 U3783 ( .A1(n3693), .A2(n2830), .ZN(n2969) );
  NAND2_X1 U3784 ( .A1(n2993), .A2(n2839), .ZN(n2968) );
  NAND2_X1 U3785 ( .A1(n2969), .A2(n2968), .ZN(n3018) );
  XNOR2_X1 U3786 ( .A(n3017), .B(n3018), .ZN(n2970) );
  XNOR2_X1 U3787 ( .A(n3019), .B(n2970), .ZN(n2971) );
  NAND2_X1 U3788 ( .A1(n2971), .A2(n4514), .ZN(n2976) );
  INV_X1 U3789 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2972) );
  NOR2_X1 U3790 ( .A1(STATE_REG_SCAN_IN), .A2(n2972), .ZN(n4541) );
  OAI22_X1 U3791 ( .A1(n3090), .A2(n4503), .B1(n4504), .B2(n2973), .ZN(n2974)
         );
  AOI211_X1 U3792 ( .C1(n2993), .C2(n2153), .A(n4541), .B(n2974), .ZN(n2975)
         );
  OAI211_X1 U3793 ( .C1(n4519), .C2(n2996), .A(n2976), .B(n2975), .ZN(U3236)
         );
  XNOR2_X1 U3794 ( .A(n2977), .B(n3584), .ZN(n4767) );
  OAI21_X1 U3795 ( .B1(n3584), .B2(n2979), .A(n2978), .ZN(n2982) );
  AOI22_X1 U3796 ( .A1(n3695), .A2(n4675), .B1(n4674), .B2(n3620), .ZN(n2980)
         );
  OAI21_X1 U3797 ( .B1(n2418), .B2(n4678), .A(n2980), .ZN(n2981) );
  AOI21_X1 U3798 ( .B1(n2982), .B2(n4702), .A(n2981), .ZN(n2983) );
  OAI21_X1 U3799 ( .B1(n4767), .B2(n4684), .A(n2983), .ZN(n4768) );
  NAND2_X1 U3800 ( .A1(n4768), .A2(n4712), .ZN(n2988) );
  AOI21_X1 U3801 ( .B1(n3620), .B2(n4762), .A(n2984), .ZN(n4770) );
  INV_X1 U3802 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2985) );
  OAI22_X1 U3803 ( .A1(n4712), .A2(n2985), .B1(n4716), .B2(REG3_REG_3__SCAN_IN), .ZN(n2986) );
  AOI21_X1 U3804 ( .B1(n4696), .B2(n4770), .A(n2986), .ZN(n2987) );
  OAI211_X1 U3805 ( .C1(n4767), .C2(n4693), .A(n2988), .B(n2987), .ZN(U3287)
         );
  OAI22_X1 U3806 ( .A1(n3090), .A2(n4705), .B1(n2306), .B2(n4010), .ZN(n2992)
         );
  NAND2_X1 U3807 ( .A1(n3628), .A2(n3635), .ZN(n3588) );
  XNOR2_X1 U3808 ( .A(n2989), .B(n3588), .ZN(n2990) );
  NOR2_X1 U3809 ( .A1(n2990), .A2(n4015), .ZN(n2991) );
  AOI211_X1 U3810 ( .C1(n4655), .C2(n3694), .A(n2992), .B(n2991), .ZN(n3033)
         );
  NAND2_X1 U3811 ( .A1(n3009), .A2(n2993), .ZN(n2994) );
  INV_X1 U3812 ( .A(n3037), .ZN(n3001) );
  INV_X1 U3813 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2997) );
  OAI22_X1 U3814 ( .A1(n4712), .A2(n2997), .B1(n2996), .B2(n4716), .ZN(n3000)
         );
  XOR2_X1 U3815 ( .A(n3588), .B(n2998), .Z(n3034) );
  NOR2_X1 U3816 ( .A1(n3034), .A2(n3967), .ZN(n2999) );
  AOI211_X1 U3817 ( .C1(n3001), .C2(n4696), .A(n3000), .B(n2999), .ZN(n3002)
         );
  OAI21_X1 U3818 ( .B1(n4700), .B2(n3033), .A(n3002), .ZN(U3284) );
  INV_X1 U3819 ( .A(n3004), .ZN(n3625) );
  NAND2_X1 U3820 ( .A1(n3625), .A2(n3634), .ZN(n3586) );
  XNOR2_X1 U3821 ( .A(n3003), .B(n3586), .ZN(n4779) );
  XOR2_X1 U3822 ( .A(n3586), .B(n3005), .Z(n3008) );
  OAI22_X1 U3823 ( .A1(n3027), .A2(n4705), .B1(n4010), .B2(n3010), .ZN(n3006)
         );
  AOI21_X1 U3824 ( .B1(n4655), .B2(n3695), .A(n3006), .ZN(n3007) );
  OAI21_X1 U3825 ( .B1(n3008), .B2(n4015), .A(n3007), .ZN(n4781) );
  NAND2_X1 U3826 ( .A1(n4781), .A2(n4712), .ZN(n3016) );
  OAI21_X1 U3827 ( .B1(n3011), .B2(n3010), .A(n3009), .ZN(n4777) );
  INV_X1 U3828 ( .A(n4777), .ZN(n3014) );
  INV_X1 U3829 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3758) );
  OAI22_X1 U3830 ( .A1(n4712), .A2(n3758), .B1(n3012), .B2(n4716), .ZN(n3013)
         );
  AOI21_X1 U3831 ( .B1(n3014), .B2(n4696), .A(n3013), .ZN(n3015) );
  OAI211_X1 U3832 ( .C1(n3967), .C2(n4779), .A(n3016), .B(n3015), .ZN(U3285)
         );
  OAI21_X1 U3833 ( .B1(n3019), .B2(n3018), .A(n3017), .ZN(n3021) );
  NAND2_X1 U3834 ( .A1(n3019), .A2(n3018), .ZN(n3020) );
  NAND2_X1 U3835 ( .A1(n3021), .A2(n3020), .ZN(n3042) );
  OAI22_X1 U3836 ( .A1(n3090), .A2(n2838), .B1(n2831), .B2(n3022), .ZN(n3023)
         );
  XNOR2_X1 U3837 ( .A(n3023), .B(n3335), .ZN(n3043) );
  OR2_X1 U3838 ( .A1(n3090), .A2(n3384), .ZN(n3025) );
  NAND2_X1 U3839 ( .A1(n3029), .A2(n2839), .ZN(n3024) );
  NAND2_X1 U3840 ( .A1(n3025), .A2(n3024), .ZN(n3044) );
  XNOR2_X1 U3841 ( .A(n3043), .B(n3044), .ZN(n3041) );
  XOR2_X1 U3842 ( .A(n3042), .B(n3041), .Z(n3026) );
  NAND2_X1 U3843 ( .A1(n3026), .A2(n4514), .ZN(n3031) );
  AND2_X1 U3844 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n4551) );
  OAI22_X1 U3845 ( .A1(n3027), .A2(n4504), .B1(n4503), .B2(n3080), .ZN(n3028)
         );
  AOI211_X1 U3846 ( .C1(n3029), .C2(n2153), .A(n4551), .B(n3028), .ZN(n3030)
         );
  OAI211_X1 U3847 ( .C1(n4519), .C2(n3032), .A(n3031), .B(n3030), .ZN(U3210)
         );
  OAI21_X1 U3848 ( .B1(n4778), .B2(n3034), .A(n3033), .ZN(n3039) );
  OAI22_X1 U3849 ( .A1(n3037), .A2(n4130), .B1(n4828), .B2(n2461), .ZN(n3035)
         );
  AOI21_X1 U3850 ( .B1(n3039), .B2(n4828), .A(n3035), .ZN(n3036) );
  INV_X1 U3851 ( .A(n3036), .ZN(U3524) );
  OAI22_X1 U3852 ( .A1(n3037), .A2(n4478), .B1(n4813), .B2(n2460), .ZN(n3038)
         );
  AOI21_X1 U3853 ( .B1(n3039), .B2(n4813), .A(n3038), .ZN(n3040) );
  INV_X1 U3854 ( .A(n3040), .ZN(U3479) );
  INV_X1 U3855 ( .A(n3043), .ZN(n3045) );
  NAND2_X1 U3856 ( .A1(n3045), .A2(n3044), .ZN(n3046) );
  NAND2_X1 U3857 ( .A1(n3691), .A2(n2839), .ZN(n3048) );
  NAND2_X1 U3858 ( .A1(n3088), .A2(n2841), .ZN(n3047) );
  NAND2_X1 U3859 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XNOR2_X1 U3860 ( .A(n3049), .B(n3386), .ZN(n3052) );
  NAND2_X1 U3861 ( .A1(n3691), .A2(n2830), .ZN(n3051) );
  NAND2_X1 U3862 ( .A1(n3088), .A2(n2839), .ZN(n3050) );
  NAND2_X1 U3863 ( .A1(n3051), .A2(n3050), .ZN(n3053) );
  AND2_X1 U3864 ( .A1(n3052), .A2(n3053), .ZN(n3073) );
  INV_X1 U3865 ( .A(n3073), .ZN(n3056) );
  INV_X1 U3866 ( .A(n3052), .ZN(n3055) );
  INV_X1 U3867 ( .A(n3053), .ZN(n3054) );
  NAND2_X1 U3868 ( .A1(n3055), .A2(n3054), .ZN(n3074) );
  NAND2_X1 U3869 ( .A1(n3056), .A2(n3074), .ZN(n3057) );
  XNOR2_X1 U3870 ( .A(n3072), .B(n3057), .ZN(n3058) );
  NAND2_X1 U3871 ( .A1(n3058), .A2(n4514), .ZN(n3061) );
  INV_X1 U3872 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4229) );
  NOR2_X1 U3873 ( .A1(STATE_REG_SCAN_IN), .A2(n4229), .ZN(n4564) );
  OAI22_X1 U3874 ( .A1(n3123), .A2(n4503), .B1(n4504), .B2(n3090), .ZN(n3059)
         );
  AOI211_X1 U3875 ( .C1(n3088), .C2(n2153), .A(n4564), .B(n3059), .ZN(n3060)
         );
  OAI211_X1 U3876 ( .C1(n4519), .C2(n3097), .A(n3061), .B(n3060), .ZN(U3218)
         );
  NAND2_X1 U3877 ( .A1(n2176), .A2(n3632), .ZN(n3561) );
  XNOR2_X1 U3878 ( .A(n3062), .B(n3561), .ZN(n3065) );
  AOI22_X1 U3879 ( .A1(n4656), .A2(n4675), .B1(n4674), .B2(n3082), .ZN(n3063)
         );
  OAI21_X1 U3880 ( .B1(n3080), .B2(n4678), .A(n3063), .ZN(n3064) );
  AOI21_X1 U3881 ( .B1(n3065), .B2(n4702), .A(n3064), .ZN(n4793) );
  XNOR2_X1 U3882 ( .A(n3066), .B(n3561), .ZN(n4796) );
  OAI21_X1 U3883 ( .B1(n4787), .B2(n3067), .A(n3128), .ZN(n4792) );
  NOR2_X1 U3884 ( .A1(n4792), .A2(n4040), .ZN(n3070) );
  INV_X1 U3885 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3068) );
  OAI22_X1 U3886 ( .A1(n4712), .A2(n3068), .B1(n3085), .B2(n4716), .ZN(n3069)
         );
  AOI211_X1 U3887 ( .C1(n4796), .C2(n4042), .A(n3070), .B(n3069), .ZN(n3071)
         );
  OAI21_X1 U3888 ( .B1(n4793), .B2(n4700), .A(n3071), .ZN(U3281) );
  NAND2_X1 U3889 ( .A1(n3075), .A2(n3074), .ZN(n3104) );
  NAND2_X1 U3890 ( .A1(n3690), .A2(n2839), .ZN(n3077) );
  NAND2_X1 U3891 ( .A1(n3082), .A2(n2841), .ZN(n3076) );
  NAND2_X1 U3892 ( .A1(n3077), .A2(n3076), .ZN(n3078) );
  XNOR2_X1 U3893 ( .A(n3078), .B(n3386), .ZN(n3105) );
  AOI22_X1 U3894 ( .A1(n3690), .A2(n2830), .B1(n2839), .B2(n3082), .ZN(n3106)
         );
  XNOR2_X1 U3895 ( .A(n3105), .B(n3106), .ZN(n3103) );
  XNOR2_X1 U3896 ( .A(n3104), .B(n3103), .ZN(n3079) );
  NAND2_X1 U3897 ( .A1(n3079), .A2(n4514), .ZN(n3084) );
  NOR2_X1 U3898 ( .A1(STATE_REG_SCAN_IN), .A2(n2494), .ZN(n4576) );
  OAI22_X1 U3899 ( .A1(n3080), .A2(n4504), .B1(n4503), .B2(n3164), .ZN(n3081)
         );
  AOI211_X1 U3900 ( .C1(n3082), .C2(n2153), .A(n4576), .B(n3081), .ZN(n3083)
         );
  OAI211_X1 U3901 ( .C1(n4519), .C2(n3085), .A(n3084), .B(n3083), .ZN(U3228)
         );
  NAND2_X1 U3902 ( .A1(n3631), .A2(n3636), .ZN(n3587) );
  XNOR2_X1 U3903 ( .A(n3086), .B(n3587), .ZN(n3094) );
  XNOR2_X1 U3904 ( .A(n3087), .B(n3587), .ZN(n3092) );
  AOI22_X1 U3905 ( .A1(n3690), .A2(n4675), .B1(n3088), .B2(n4674), .ZN(n3089)
         );
  OAI21_X1 U3906 ( .B1(n3090), .B2(n4678), .A(n3089), .ZN(n3091) );
  AOI21_X1 U3907 ( .B1(n3092), .B2(n4702), .A(n3091), .ZN(n3093) );
  OAI21_X1 U3908 ( .B1(n3094), .B2(n4684), .A(n3093), .ZN(n4789) );
  INV_X1 U3909 ( .A(n4789), .ZN(n3102) );
  INV_X1 U3910 ( .A(n3094), .ZN(n4791) );
  NOR2_X1 U3911 ( .A1(n3096), .A2(n3095), .ZN(n4788) );
  NOR3_X1 U3912 ( .A1(n4788), .A2(n4787), .A3(n4040), .ZN(n3100) );
  INV_X1 U3913 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3098) );
  OAI22_X1 U3914 ( .A1(n4712), .A2(n3098), .B1(n3097), .B2(n4716), .ZN(n3099)
         );
  AOI211_X1 U3915 ( .C1(n4791), .C2(n4701), .A(n3100), .B(n3099), .ZN(n3101)
         );
  OAI21_X1 U3916 ( .B1(n3102), .B2(n4700), .A(n3101), .ZN(U3282) );
  INV_X1 U3917 ( .A(n3105), .ZN(n3107) );
  NAND2_X1 U3918 ( .A1(n3107), .A2(n3106), .ZN(n3108) );
  NAND2_X1 U3919 ( .A1(n4656), .A2(n2839), .ZN(n3110) );
  NAND2_X1 U3920 ( .A1(n3121), .A2(n2841), .ZN(n3109) );
  NAND2_X1 U3921 ( .A1(n3110), .A2(n3109), .ZN(n3111) );
  XNOR2_X1 U3922 ( .A(n3111), .B(n3335), .ZN(n3150) );
  AOI22_X1 U3923 ( .A1(n4656), .A2(n2830), .B1(n2839), .B2(n3121), .ZN(n3151)
         );
  XNOR2_X1 U3924 ( .A(n3150), .B(n3151), .ZN(n3113) );
  AOI21_X1 U3925 ( .B1(n3112), .B2(n3113), .A(n3519), .ZN(n3115) );
  NAND2_X1 U3926 ( .A1(n3115), .A2(n3155), .ZN(n3118) );
  NOR2_X1 U3927 ( .A1(STATE_REG_SCAN_IN), .A2(n4215), .ZN(n4585) );
  OAI22_X1 U3928 ( .A1(n3158), .A2(n4503), .B1(n4504), .B2(n3123), .ZN(n3116)
         );
  AOI211_X1 U3929 ( .C1(n3121), .C2(n2153), .A(n4585), .B(n3116), .ZN(n3117)
         );
  OAI211_X1 U3930 ( .C1(n4519), .C2(n3131), .A(n3118), .B(n3117), .ZN(U3214)
         );
  AND2_X1 U3931 ( .A1(n3602), .A2(n3599), .ZN(n3568) );
  XOR2_X1 U3932 ( .A(n3568), .B(n3119), .Z(n3127) );
  XNOR2_X1 U3933 ( .A(n3120), .B(n3568), .ZN(n3125) );
  AOI22_X1 U3934 ( .A1(n3689), .A2(n4675), .B1(n3121), .B2(n4674), .ZN(n3122)
         );
  OAI21_X1 U3935 ( .B1(n3123), .B2(n4678), .A(n3122), .ZN(n3124) );
  AOI21_X1 U3936 ( .B1(n3125), .B2(n4702), .A(n3124), .ZN(n3126) );
  OAI21_X1 U3937 ( .B1(n3127), .B2(n4684), .A(n3126), .ZN(n4801) );
  INV_X1 U3938 ( .A(n4801), .ZN(n3136) );
  INV_X1 U3939 ( .A(n3127), .ZN(n4804) );
  INV_X1 U3940 ( .A(n3128), .ZN(n3130) );
  NOR2_X1 U3941 ( .A1(n3130), .A2(n3129), .ZN(n4800) );
  INV_X1 U3942 ( .A(n4666), .ZN(n4799) );
  NOR3_X1 U3943 ( .A1(n4800), .A2(n4799), .A3(n4040), .ZN(n3134) );
  INV_X1 U3944 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3132) );
  OAI22_X1 U3945 ( .A1(n4712), .A2(n3132), .B1(n3131), .B2(n4716), .ZN(n3133)
         );
  AOI211_X1 U3946 ( .C1(n4804), .C2(n4701), .A(n3134), .B(n3133), .ZN(n3135)
         );
  OAI21_X1 U3947 ( .B1(n3136), .B2(n4700), .A(n3135), .ZN(U3280) );
  INV_X1 U3948 ( .A(n3598), .ZN(n3137) );
  OR2_X1 U3949 ( .A1(n3137), .A2(n3606), .ZN(n3567) );
  XNOR2_X1 U3950 ( .A(n3138), .B(n3567), .ZN(n3141) );
  OAI22_X1 U3951 ( .A1(n3263), .A2(n4705), .B1(n4010), .B2(n3185), .ZN(n3139)
         );
  AOI21_X1 U3952 ( .B1(n4655), .B2(n3689), .A(n3139), .ZN(n3140) );
  OAI21_X1 U3953 ( .B1(n3141), .B2(n4015), .A(n3140), .ZN(n3190) );
  INV_X1 U3954 ( .A(n3190), .ZN(n3149) );
  XNOR2_X1 U3955 ( .A(n3142), .B(n3567), .ZN(n3191) );
  INV_X1 U3956 ( .A(n3143), .ZN(n4665) );
  INV_X1 U3957 ( .A(n3222), .ZN(n3144) );
  OAI21_X1 U3958 ( .B1(n4665), .B2(n3185), .A(n3144), .ZN(n3195) );
  INV_X1 U3959 ( .A(n3145), .ZN(n3187) );
  INV_X1 U3960 ( .A(n4716), .ZN(n4688) );
  AOI22_X1 U3961 ( .A1(n4700), .A2(REG2_REG_12__SCAN_IN), .B1(n3187), .B2(
        n4688), .ZN(n3146) );
  OAI21_X1 U3962 ( .B1(n3195), .B2(n4040), .A(n3146), .ZN(n3147) );
  AOI21_X1 U3963 ( .B1(n3191), .B2(n4042), .A(n3147), .ZN(n3148) );
  OAI21_X1 U3964 ( .B1(n3149), .B2(n4700), .A(n3148), .ZN(U3278) );
  INV_X1 U3965 ( .A(n3150), .ZN(n3153) );
  INV_X1 U3966 ( .A(n3151), .ZN(n3152) );
  NAND2_X1 U3967 ( .A1(n3153), .A2(n3152), .ZN(n3154) );
  NAND2_X1 U3968 ( .A1(n3155), .A2(n3154), .ZN(n3203) );
  OAI22_X1 U3969 ( .A1(n3158), .A2(n2838), .B1(n2831), .B2(n3156), .ZN(n3157)
         );
  XNOR2_X1 U3970 ( .A(n3157), .B(n3335), .ZN(n3198) );
  OR2_X1 U3971 ( .A1(n3158), .A2(n3384), .ZN(n3160) );
  NAND2_X1 U3972 ( .A1(n4667), .A2(n2839), .ZN(n3159) );
  XNOR2_X1 U3973 ( .A(n3198), .B(n3197), .ZN(n3161) );
  XNOR2_X1 U3974 ( .A(n3203), .B(n3161), .ZN(n3162) );
  NAND2_X1 U3975 ( .A1(n3162), .A2(n4514), .ZN(n3167) );
  NOR2_X1 U3976 ( .A1(STATE_REG_SCAN_IN), .A2(n3163), .ZN(n4597) );
  OAI22_X1 U3977 ( .A1(n4658), .A2(n4503), .B1(n4504), .B2(n3164), .ZN(n3165)
         );
  AOI211_X1 U3978 ( .C1(n4667), .C2(n2153), .A(n4597), .B(n3165), .ZN(n3166)
         );
  OAI211_X1 U3979 ( .C1(n4519), .C2(n3168), .A(n3167), .B(n3166), .ZN(U3233)
         );
  NAND2_X1 U3980 ( .A1(n3688), .A2(n2832), .ZN(n3170) );
  NAND2_X1 U3981 ( .A1(n3172), .A2(n2841), .ZN(n3169) );
  NAND2_X1 U3982 ( .A1(n3170), .A2(n3169), .ZN(n3171) );
  XNOR2_X1 U3983 ( .A(n3171), .B(n3386), .ZN(n3175) );
  NAND2_X1 U3984 ( .A1(n3688), .A2(n2830), .ZN(n3174) );
  NAND2_X1 U3985 ( .A1(n3172), .A2(n2839), .ZN(n3173) );
  NAND2_X1 U3986 ( .A1(n3174), .A2(n3173), .ZN(n3176) );
  NAND2_X1 U3987 ( .A1(n3175), .A2(n3176), .ZN(n3196) );
  INV_X1 U3988 ( .A(n3175), .ZN(n3178) );
  INV_X1 U3989 ( .A(n3176), .ZN(n3177) );
  NAND2_X1 U3990 ( .A1(n3178), .A2(n3177), .ZN(n3199) );
  NAND2_X1 U3991 ( .A1(n3196), .A2(n3199), .ZN(n3183) );
  INV_X1 U3992 ( .A(n3197), .ZN(n3179) );
  NOR2_X1 U3993 ( .A1(n3203), .A2(n3179), .ZN(n3181) );
  INV_X1 U3994 ( .A(n3203), .ZN(n3180) );
  OAI22_X1 U3995 ( .A1(n3181), .A2(n3198), .B1(n3180), .B2(n3197), .ZN(n3182)
         );
  XOR2_X1 U3996 ( .A(n3183), .B(n3182), .Z(n3189) );
  INV_X1 U3997 ( .A(n2153), .ZN(n3513) );
  AOI22_X1 U3998 ( .A1(n3432), .A2(n3689), .B1(n3431), .B2(n3687), .ZN(n3184)
         );
  NAND2_X1 U3999 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4602) );
  OAI211_X1 U4000 ( .C1(n3513), .C2(n3185), .A(n3184), .B(n4602), .ZN(n3186)
         );
  AOI21_X1 U4001 ( .B1(n3187), .B2(n3517), .A(n3186), .ZN(n3188) );
  OAI21_X1 U4002 ( .B1(n3189), .B2(n3519), .A(n3188), .ZN(U3221) );
  AOI21_X1 U4003 ( .B1(n4797), .B2(n3191), .A(n3190), .ZN(n3193) );
  MUX2_X1 U4004 ( .A(n2531), .B(n3193), .S(n4828), .Z(n3192) );
  OAI21_X1 U4005 ( .B1(n3195), .B2(n4130), .A(n3192), .ZN(U3530) );
  INV_X2 U4006 ( .A(n4812), .ZN(n4813) );
  MUX2_X1 U4007 ( .A(n2530), .B(n3193), .S(n4813), .Z(n3194) );
  OAI21_X1 U4008 ( .B1(n3195), .B2(n4478), .A(n3194), .ZN(U3491) );
  OAI21_X1 U4009 ( .B1(n3198), .B2(n3197), .A(n3196), .ZN(n3202) );
  NAND3_X1 U4010 ( .A1(n3198), .A2(n3197), .A3(n3196), .ZN(n3200) );
  AND2_X1 U4011 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  NAND2_X1 U4012 ( .A1(n3687), .A2(n2839), .ZN(n3205) );
  NAND2_X1 U4013 ( .A1(n3216), .A2(n2841), .ZN(n3204) );
  NAND2_X1 U4014 ( .A1(n3205), .A2(n3204), .ZN(n3206) );
  NAND2_X1 U4015 ( .A1(n3687), .A2(n2830), .ZN(n3208) );
  NAND2_X1 U4016 ( .A1(n3216), .A2(n2832), .ZN(n3207) );
  NAND2_X1 U4017 ( .A1(n3208), .A2(n3207), .ZN(n3241) );
  XNOR2_X1 U4018 ( .A(n3243), .B(n3241), .ZN(n3209) );
  XNOR2_X1 U4019 ( .A(n3242), .B(n3209), .ZN(n3210) );
  NAND2_X1 U4020 ( .A1(n3210), .A2(n4514), .ZN(n3213) );
  AND2_X1 U4021 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4615) );
  OAI22_X1 U4022 ( .A1(n4658), .A2(n4504), .B1(n4503), .B2(n4505), .ZN(n3211)
         );
  AOI211_X1 U4023 ( .C1(n3216), .C2(n2153), .A(n4615), .B(n3211), .ZN(n3212)
         );
  OAI211_X1 U4024 ( .C1(n4519), .C2(n3223), .A(n3213), .B(n3212), .ZN(U3231)
         );
  AND2_X1 U4025 ( .A1(n2182), .A2(n3603), .ZN(n3570) );
  XOR2_X1 U4026 ( .A(n3570), .B(n3214), .Z(n4126) );
  XOR2_X1 U4027 ( .A(n3570), .B(n3215), .Z(n3219) );
  AOI22_X1 U4028 ( .A1(n3686), .A2(n4675), .B1(n4674), .B2(n3216), .ZN(n3217)
         );
  OAI21_X1 U4029 ( .B1(n4658), .B2(n4678), .A(n3217), .ZN(n3218) );
  AOI21_X1 U4030 ( .B1(n3219), .B2(n4702), .A(n3218), .ZN(n3220) );
  OAI21_X1 U4031 ( .B1(n4126), .B2(n4684), .A(n3220), .ZN(n4127) );
  NAND2_X1 U4032 ( .A1(n4127), .A2(n4712), .ZN(n3227) );
  OAI21_X1 U4033 ( .B1(n3222), .B2(n3221), .A(n3269), .ZN(n4479) );
  INV_X1 U4034 ( .A(n4479), .ZN(n3225) );
  INV_X1 U4035 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4609) );
  OAI22_X1 U4036 ( .A1(n4712), .A2(n4609), .B1(n3223), .B2(n4716), .ZN(n3224)
         );
  AOI21_X1 U4037 ( .B1(n3225), .B2(n4696), .A(n3224), .ZN(n3226) );
  OAI211_X1 U4038 ( .C1(n4126), .C2(n4693), .A(n3227), .B(n3226), .ZN(U3277)
         );
  XNOR2_X1 U4039 ( .A(n3228), .B(n3233), .ZN(n3231) );
  OAI22_X1 U4040 ( .A1(n4502), .A2(n4705), .B1(n4010), .B2(n3300), .ZN(n3229)
         );
  AOI21_X1 U4041 ( .B1(n4655), .B2(n3686), .A(n3229), .ZN(n3230) );
  OAI21_X1 U4042 ( .B1(n3231), .B2(n4015), .A(n3230), .ZN(n4117) );
  INV_X1 U40430 ( .A(n4117), .ZN(n3240) );
  XNOR2_X1 U4044 ( .A(n3232), .B(n3233), .ZN(n4118) );
  INV_X1 U4045 ( .A(n4122), .ZN(n3235) );
  INV_X1 U4046 ( .A(n4037), .ZN(n3234) );
  OAI21_X1 U4047 ( .B1(n3235), .B2(n3300), .A(n3234), .ZN(n4473) );
  NOR2_X1 U4048 ( .A1(n4473), .A2(n4040), .ZN(n3238) );
  INV_X1 U4049 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3236) );
  OAI22_X1 U4050 ( .A1(n4712), .A2(n3236), .B1(n4518), .B2(n4716), .ZN(n3237)
         );
  AOI211_X1 U4051 ( .C1(n4118), .C2(n4042), .A(n3238), .B(n3237), .ZN(n3239)
         );
  OAI21_X1 U4052 ( .B1(n3240), .B2(n4700), .A(n3239), .ZN(U3275) );
  OAI22_X1 U4053 ( .A1(n4505), .A2(n2838), .B1(n2831), .B2(n3244), .ZN(n3245)
         );
  XNOR2_X1 U4054 ( .A(n3245), .B(n3386), .ZN(n3248) );
  OR2_X1 U4055 ( .A1(n4505), .A2(n3384), .ZN(n3247) );
  NAND2_X1 U4056 ( .A1(n3268), .A2(n2839), .ZN(n3246) );
  NAND2_X1 U4057 ( .A1(n3247), .A2(n3246), .ZN(n3249) );
  NAND2_X1 U4058 ( .A1(n3248), .A2(n3249), .ZN(n3254) );
  NAND2_X1 U4059 ( .A1(n3253), .A2(n3254), .ZN(n3299) );
  INV_X1 U4060 ( .A(n3248), .ZN(n3251) );
  INV_X1 U4061 ( .A(n3249), .ZN(n3250) );
  NAND2_X1 U4062 ( .A1(n3251), .A2(n3250), .ZN(n3298) );
  INV_X1 U4063 ( .A(n3298), .ZN(n3252) );
  NOR2_X1 U4064 ( .A1(n3299), .A2(n3252), .ZN(n3256) );
  AOI21_X1 U4065 ( .B1(n3298), .B2(n3254), .A(n3253), .ZN(n3255) );
  OAI21_X1 U4066 ( .B1(n3256), .B2(n3255), .A(n4514), .ZN(n3260) );
  INV_X1 U4067 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3257) );
  NOR2_X1 U4068 ( .A1(STATE_REG_SCAN_IN), .A2(n3257), .ZN(n4624) );
  OAI22_X1 U4069 ( .A1(n4492), .A2(n4503), .B1(n4504), .B2(n3263), .ZN(n3258)
         );
  AOI211_X1 U4070 ( .C1(n3268), .C2(n2153), .A(n4624), .B(n3258), .ZN(n3259)
         );
  OAI211_X1 U4071 ( .C1(n4519), .C2(n3270), .A(n3260), .B(n3259), .ZN(U3212)
         );
  OAI21_X1 U4072 ( .B1(n3592), .B2(n3539), .A(n3261), .ZN(n3267) );
  AOI22_X1 U4073 ( .A1(n3685), .A2(n4675), .B1(n3268), .B2(n4674), .ZN(n3262)
         );
  OAI21_X1 U4074 ( .B1(n3263), .B2(n4678), .A(n3262), .ZN(n3266) );
  XNOR2_X1 U4075 ( .A(n3264), .B(n3592), .ZN(n4125) );
  NOR2_X1 U4076 ( .A1(n4125), .A2(n4684), .ZN(n3265) );
  AOI211_X1 U4077 ( .C1(n4702), .C2(n3267), .A(n3266), .B(n3265), .ZN(n4124)
         );
  INV_X1 U4078 ( .A(n4125), .ZN(n3274) );
  NAND2_X1 U4079 ( .A1(n3269), .A2(n3268), .ZN(n4121) );
  AND3_X1 U4080 ( .A1(n4122), .A2(n4696), .A3(n4121), .ZN(n3273) );
  INV_X1 U4081 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3271) );
  OAI22_X1 U4082 ( .A1(n4712), .A2(n3271), .B1(n3270), .B2(n4716), .ZN(n3272)
         );
  AOI211_X1 U4083 ( .C1(n3274), .C2(n4701), .A(n3273), .B(n3272), .ZN(n3275)
         );
  OAI21_X1 U4084 ( .B1(n4124), .B2(n4700), .A(n3275), .ZN(U3276) );
  INV_X1 U4085 ( .A(n3572), .ZN(n3277) );
  NAND2_X1 U4086 ( .A1(n3526), .A2(DATAI_29_), .ZN(n3521) );
  XOR2_X1 U4087 ( .A(n3521), .B(n3682), .Z(n3573) );
  XNOR2_X1 U4088 ( .A(n3279), .B(n3573), .ZN(n4072) );
  NOR2_X2 U4089 ( .A1(n3280), .A2(n3528), .ZN(n4066) );
  AOI21_X1 U4090 ( .B1(n3528), .B2(n3280), .A(n4066), .ZN(n4071) );
  AOI22_X1 U4091 ( .A1(n4071), .A2(n4696), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4700), .ZN(n3297) );
  INV_X1 U4092 ( .A(n3532), .ZN(n3281) );
  INV_X1 U4093 ( .A(n3283), .ZN(n3284) );
  XNOR2_X1 U4094 ( .A(n3284), .B(n3573), .ZN(n3285) );
  INV_X1 U4095 ( .A(REG0_REG_30__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4096 ( .A1(n2407), .A2(REG2_REG_30__SCAN_IN), .ZN(n3288) );
  INV_X1 U4097 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3286) );
  OR2_X1 U4098 ( .A1(n2423), .A2(n3286), .ZN(n3287) );
  OAI211_X1 U4099 ( .C1(n3290), .C2(n3289), .A(n3288), .B(n3287), .ZN(n3681)
         );
  AOI21_X1 U4100 ( .B1(B_REG_SCAN_IN), .B2(n4481), .A(n4705), .ZN(n4060) );
  AOI22_X1 U4101 ( .A1(n3681), .A2(n4060), .B1(n4674), .B2(n3528), .ZN(n3291)
         );
  NOR2_X1 U4102 ( .A1(n4716), .A2(n3294), .ZN(n3295) );
  OAI21_X1 U4103 ( .B1(n4070), .B2(n3295), .A(n4712), .ZN(n3296) );
  OAI211_X1 U4104 ( .C1(n4072), .C2(n3967), .A(n3297), .B(n3296), .ZN(U3354)
         );
  OAI22_X1 U4105 ( .A1(n4492), .A2(n2838), .B1(n2831), .B2(n3300), .ZN(n3301)
         );
  XNOR2_X1 U4106 ( .A(n3301), .B(n3386), .ZN(n3309) );
  OR2_X1 U4107 ( .A1(n4492), .A2(n3384), .ZN(n3303) );
  NAND2_X1 U4108 ( .A1(n4508), .A2(n2839), .ZN(n3302) );
  OAI22_X1 U4109 ( .A1(n4502), .A2(n2838), .B1(n2831), .B2(n4036), .ZN(n3304)
         );
  XNOR2_X1 U4110 ( .A(n3304), .B(n3386), .ZN(n3308) );
  OR2_X1 U4111 ( .A1(n4502), .A2(n3384), .ZN(n3306) );
  NAND2_X1 U4112 ( .A1(n4495), .A2(n2839), .ZN(n3305) );
  NAND2_X1 U4113 ( .A1(n3306), .A2(n3305), .ZN(n3307) );
  NOR2_X1 U4114 ( .A1(n3308), .A2(n3307), .ZN(n3310) );
  AOI21_X1 U4115 ( .B1(n3308), .B2(n3307), .A(n3310), .ZN(n4497) );
  OAI22_X1 U4116 ( .A1(n4491), .A2(n2838), .B1(n2831), .B2(n4020), .ZN(n3311)
         );
  XNOR2_X1 U4117 ( .A(n3311), .B(n3386), .ZN(n3315) );
  OR2_X1 U4118 ( .A1(n4491), .A2(n3384), .ZN(n3313) );
  NAND2_X1 U4119 ( .A1(n3464), .A2(n2839), .ZN(n3312) );
  NAND2_X1 U4120 ( .A1(n3313), .A2(n3312), .ZN(n3314) );
  NAND2_X1 U4121 ( .A1(n3315), .A2(n3314), .ZN(n3458) );
  NOR2_X1 U4122 ( .A1(n3315), .A2(n3314), .ZN(n3460) );
  AOI21_X1 U4123 ( .B1(n3457), .B2(n3458), .A(n3460), .ZN(n3500) );
  INV_X1 U4124 ( .A(n3500), .ZN(n3321) );
  OR2_X1 U4125 ( .A1(n4011), .A2(n3384), .ZN(n3317) );
  NAND2_X1 U4126 ( .A1(n3994), .A2(n2839), .ZN(n3316) );
  NAND2_X1 U4127 ( .A1(n3317), .A2(n3316), .ZN(n3497) );
  OAI22_X1 U4128 ( .A1(n4011), .A2(n2838), .B1(n2831), .B2(n4002), .ZN(n3318)
         );
  XNOR2_X1 U4129 ( .A(n3318), .B(n3386), .ZN(n3498) );
  NAND2_X1 U4130 ( .A1(n3497), .A2(n3498), .ZN(n3320) );
  AOI21_X1 U4131 ( .B1(n3321), .B2(n3320), .A(n3319), .ZN(n3421) );
  NAND2_X1 U4132 ( .A1(n3995), .A2(n2839), .ZN(n3323) );
  OR2_X1 U4133 ( .A1(n3986), .A2(n2831), .ZN(n3322) );
  NAND2_X1 U4134 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  XNOR2_X1 U4135 ( .A(n3324), .B(n3386), .ZN(n3326) );
  OAI22_X1 U4136 ( .A1(n3502), .A2(n3384), .B1(n2838), .B2(n3986), .ZN(n3325)
         );
  XNOR2_X1 U4137 ( .A(n3326), .B(n3325), .ZN(n3420) );
  NAND2_X1 U4138 ( .A1(n3939), .A2(n2839), .ZN(n3330) );
  NAND2_X1 U4139 ( .A1(n3328), .A2(n2841), .ZN(n3329) );
  NAND2_X1 U4140 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  XNOR2_X1 U4141 ( .A(n3331), .B(n3335), .ZN(n3334) );
  NOR2_X1 U4142 ( .A1(n3962), .A2(n2838), .ZN(n3332) );
  AOI21_X1 U4143 ( .B1(n3939), .B2(n2830), .A(n3332), .ZN(n3333) );
  OR2_X1 U4144 ( .A1(n3334), .A2(n3333), .ZN(n3478) );
  NAND2_X1 U4145 ( .A1(n3477), .A2(n3478), .ZN(n3476) );
  NAND2_X1 U4146 ( .A1(n3334), .A2(n3333), .ZN(n3480) );
  NAND2_X1 U4147 ( .A1(n3476), .A2(n3480), .ZN(n3439) );
  INV_X1 U4148 ( .A(n3439), .ZN(n3342) );
  OAI22_X1 U4149 ( .A1(n3956), .A2(n2838), .B1(n2831), .B2(n3944), .ZN(n3336)
         );
  XNOR2_X1 U4150 ( .A(n3336), .B(n3335), .ZN(n3437) );
  OR2_X1 U4151 ( .A1(n3956), .A2(n3384), .ZN(n3338) );
  NAND2_X1 U4152 ( .A1(n2839), .A2(n3937), .ZN(n3337) );
  INV_X1 U4153 ( .A(n3437), .ZN(n3340) );
  INV_X1 U4154 ( .A(n3436), .ZN(n3339) );
  AOI21_X2 U4155 ( .B1(n3342), .B2(n3341), .A(n2365), .ZN(n3489) );
  OAI22_X1 U4156 ( .A1(n3442), .A2(n3384), .B1(n2838), .B2(n3492), .ZN(n3349)
         );
  OAI22_X1 U4157 ( .A1(n3442), .A2(n2838), .B1(n2831), .B2(n3492), .ZN(n3343)
         );
  XNOR2_X1 U4158 ( .A(n3343), .B(n3386), .ZN(n3348) );
  XOR2_X1 U4159 ( .A(n3349), .B(n3348), .Z(n3490) );
  NAND2_X1 U4160 ( .A1(n3922), .A2(n2839), .ZN(n3345) );
  NAND2_X1 U4161 ( .A1(n2841), .A2(n3903), .ZN(n3344) );
  NAND2_X1 U4162 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  XNOR2_X1 U4163 ( .A(n3346), .B(n3386), .ZN(n3357) );
  AND2_X1 U4164 ( .A1(n2839), .A2(n3903), .ZN(n3347) );
  AOI21_X1 U4165 ( .B1(n3922), .B2(n2830), .A(n3347), .ZN(n3355) );
  XNOR2_X1 U4166 ( .A(n3357), .B(n3355), .ZN(n3411) );
  INV_X1 U4167 ( .A(n3348), .ZN(n3351) );
  INV_X1 U4168 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4169 ( .A1(n3351), .A2(n3350), .ZN(n3412) );
  OR2_X1 U4170 ( .A1(n3906), .A2(n3384), .ZN(n3354) );
  NAND2_X1 U4171 ( .A1(n2839), .A2(n3881), .ZN(n3353) );
  AND2_X1 U4172 ( .A1(n3354), .A2(n3353), .ZN(n3359) );
  INV_X1 U4173 ( .A(n3355), .ZN(n3356) );
  NAND2_X1 U4174 ( .A1(n3357), .A2(n3356), .ZN(n3360) );
  OAI22_X1 U4175 ( .A1(n3906), .A2(n2838), .B1(n2831), .B2(n3888), .ZN(n3358)
         );
  XNOR2_X1 U4176 ( .A(n3358), .B(n3386), .ZN(n3468) );
  NAND2_X1 U4177 ( .A1(n3882), .A2(n2839), .ZN(n3362) );
  NAND2_X1 U4178 ( .A1(n2841), .A2(n3863), .ZN(n3361) );
  NAND2_X1 U4179 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  XNOR2_X1 U4180 ( .A(n3363), .B(n3386), .ZN(n3367) );
  NAND2_X1 U4181 ( .A1(n3882), .A2(n2830), .ZN(n3365) );
  NAND2_X1 U4182 ( .A1(n2839), .A2(n3863), .ZN(n3364) );
  NAND2_X1 U4183 ( .A1(n3365), .A2(n3364), .ZN(n3366) );
  NOR2_X1 U4184 ( .A1(n3367), .A2(n3366), .ZN(n3448) );
  NAND2_X1 U4185 ( .A1(n3367), .A2(n3366), .ZN(n3449) );
  NAND2_X1 U4186 ( .A1(n3864), .A2(n2832), .ZN(n3369) );
  NAND2_X1 U4187 ( .A1(n2841), .A2(n3844), .ZN(n3368) );
  NAND2_X1 U4188 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  XNOR2_X1 U4189 ( .A(n3370), .B(n3386), .ZN(n3373) );
  NAND2_X1 U4190 ( .A1(n3864), .A2(n2830), .ZN(n3372) );
  NAND2_X1 U4191 ( .A1(n2839), .A2(n3844), .ZN(n3371) );
  NAND2_X1 U4192 ( .A1(n3372), .A2(n3371), .ZN(n3374) );
  AND2_X1 U4193 ( .A1(n3373), .A2(n3374), .ZN(n3507) );
  INV_X1 U4194 ( .A(n3373), .ZN(n3376) );
  INV_X1 U4195 ( .A(n3374), .ZN(n3375) );
  NAND2_X1 U4196 ( .A1(n3376), .A2(n3375), .ZN(n3506) );
  OAI22_X1 U4197 ( .A1(n3514), .A2(n2838), .B1(n3403), .B2(n2831), .ZN(n3377)
         );
  XNOR2_X1 U4198 ( .A(n3377), .B(n3386), .ZN(n3381) );
  OR2_X1 U4199 ( .A1(n3514), .A2(n3384), .ZN(n3379) );
  NAND2_X1 U4200 ( .A1(n2832), .A2(n3831), .ZN(n3378) );
  NAND2_X1 U4201 ( .A1(n3379), .A2(n3378), .ZN(n3380) );
  XNOR2_X1 U4202 ( .A(n3381), .B(n3380), .ZN(n3402) );
  INV_X1 U4203 ( .A(n3380), .ZN(n3383) );
  INV_X1 U4204 ( .A(n3381), .ZN(n3382) );
  OAI22_X1 U4205 ( .A1(n3401), .A2(n3402), .B1(n3383), .B2(n3382), .ZN(n3391)
         );
  OAI22_X1 U4206 ( .A1(n3404), .A2(n3384), .B1(n2838), .B2(n3385), .ZN(n3389)
         );
  OAI22_X1 U4207 ( .A1(n3404), .A2(n2838), .B1(n2831), .B2(n3385), .ZN(n3387)
         );
  XNOR2_X1 U4208 ( .A(n3387), .B(n3386), .ZN(n3388) );
  XOR2_X1 U4209 ( .A(n3389), .B(n3388), .Z(n3390) );
  XNOR2_X1 U4210 ( .A(n3391), .B(n3390), .ZN(n3397) );
  AOI22_X1 U4211 ( .A1(n3431), .A2(n3682), .B1(n3432), .B2(n3845), .ZN(n3394)
         );
  AOI22_X1 U4212 ( .A1(n2153), .A2(n3392), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3393) );
  OAI211_X1 U4213 ( .C1(n3816), .C2(n4519), .A(n3394), .B(n3393), .ZN(n3395)
         );
  INV_X1 U4214 ( .A(n3395), .ZN(n3396) );
  OAI21_X1 U4215 ( .B1(n3397), .B2(n3519), .A(n3396), .ZN(U3217) );
  NAND2_X1 U4216 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3398) );
  OAI21_X1 U4217 ( .B1(n2745), .B2(U3149), .A(n3398), .ZN(U3327) );
  AND2_X1 U4218 ( .A1(n4730), .A2(n3399), .ZN(n3400) );
  AOI22_X1 U4219 ( .A1(n4729), .A2(n4258), .B1(n2745), .B2(n3400), .ZN(U3459)
         );
  XNOR2_X1 U4220 ( .A(n3401), .B(n3402), .ZN(n3409) );
  INV_X1 U4221 ( .A(n3825), .ZN(n3407) );
  OAI22_X1 U4222 ( .A1(n3513), .A2(n3403), .B1(STATE_REG_SCAN_IN), .B2(n4394), 
        .ZN(n3406) );
  OAI22_X1 U4223 ( .A1(n3404), .A2(n4503), .B1(n4504), .B2(n3835), .ZN(n3405)
         );
  AOI211_X1 U4224 ( .C1(n3407), .C2(n3517), .A(n3406), .B(n3405), .ZN(n3408)
         );
  OAI21_X1 U4225 ( .B1(n3409), .B2(n3519), .A(n3408), .ZN(U3211) );
  NAND2_X1 U4226 ( .A1(n3410), .A2(n4514), .ZN(n3419) );
  AOI21_X1 U4227 ( .B1(n3488), .B2(n3412), .A(n3411), .ZN(n3418) );
  INV_X1 U4228 ( .A(n3413), .ZN(n3910) );
  OAI22_X1 U4229 ( .A1(n3513), .A2(n3908), .B1(STATE_REG_SCAN_IN), .B2(n3414), 
        .ZN(n3416) );
  OAI22_X1 U4230 ( .A1(n3906), .A2(n4503), .B1(n4504), .B2(n3442), .ZN(n3415)
         );
  AOI211_X1 U4231 ( .C1(n3910), .C2(n3517), .A(n3416), .B(n3415), .ZN(n3417)
         );
  OAI21_X1 U4232 ( .B1(n3419), .B2(n3418), .A(n3417), .ZN(U3213) );
  XNOR2_X1 U4233 ( .A(n3421), .B(n3420), .ZN(n3422) );
  NAND2_X1 U4234 ( .A1(n3422), .A2(n4514), .ZN(n3426) );
  NOR2_X1 U4235 ( .A1(n4420), .A2(STATE_REG_SCAN_IN), .ZN(n3809) );
  INV_X1 U4236 ( .A(n3939), .ZN(n3977) );
  OAI22_X1 U4237 ( .A1(n4011), .A2(n4504), .B1(n4503), .B2(n3977), .ZN(n3423)
         );
  AOI211_X1 U4238 ( .C1(n3424), .C2(n2153), .A(n3809), .B(n3423), .ZN(n3425)
         );
  OAI211_X1 U4239 ( .C1(n4519), .C2(n3987), .A(n3426), .B(n3425), .ZN(U3216)
         );
  OAI211_X1 U4240 ( .C1(n3429), .C2(n3428), .A(n3427), .B(n4514), .ZN(n3435)
         );
  AOI22_X1 U4241 ( .A1(n2153), .A2(n4690), .B1(n3430), .B2(REG3_REG_1__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4242 ( .A1(n3432), .A2(n3697), .B1(n3431), .B2(n4676), .ZN(n3433)
         );
  NAND3_X1 U4243 ( .A1(n3435), .A2(n3434), .A3(n3433), .ZN(U3219) );
  XNOR2_X1 U4244 ( .A(n3437), .B(n3436), .ZN(n3438) );
  XNOR2_X1 U4245 ( .A(n3439), .B(n3438), .ZN(n3446) );
  INV_X1 U4246 ( .A(n3440), .ZN(n3945) );
  OAI22_X1 U4247 ( .A1(n3513), .A2(n3944), .B1(STATE_REG_SCAN_IN), .B2(n3441), 
        .ZN(n3444) );
  OAI22_X1 U4248 ( .A1(n3977), .A2(n4504), .B1(n4503), .B2(n3442), .ZN(n3443)
         );
  AOI211_X1 U4249 ( .C1(n3945), .C2(n3517), .A(n3444), .B(n3443), .ZN(n3445)
         );
  OAI21_X1 U4250 ( .B1(n3446), .B2(n3519), .A(n3445), .ZN(U3220) );
  INV_X1 U4251 ( .A(n3448), .ZN(n3450) );
  NAND2_X1 U4252 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  XNOR2_X1 U4253 ( .A(n3447), .B(n3451), .ZN(n3456) );
  INV_X1 U4254 ( .A(n3452), .ZN(n3870) );
  INV_X1 U4255 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4220) );
  OAI22_X1 U4256 ( .A1(n3513), .A2(n3869), .B1(STATE_REG_SCAN_IN), .B2(n4220), 
        .ZN(n3454) );
  OAI22_X1 U4257 ( .A1(n3906), .A2(n4504), .B1(n4503), .B2(n3835), .ZN(n3453)
         );
  AOI211_X1 U4258 ( .C1(n3870), .C2(n3517), .A(n3454), .B(n3453), .ZN(n3455)
         );
  OAI21_X1 U4259 ( .B1(n3456), .B2(n3519), .A(n3455), .ZN(U3222) );
  INV_X1 U4260 ( .A(n3458), .ZN(n3459) );
  NOR2_X1 U4261 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  XNOR2_X1 U4262 ( .A(n3457), .B(n3461), .ZN(n3462) );
  NAND2_X1 U4263 ( .A1(n3462), .A2(n4514), .ZN(n3466) );
  AND2_X1 U4264 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4644) );
  OAI22_X1 U4265 ( .A1(n4011), .A2(n4503), .B1(n4504), .B2(n4502), .ZN(n3463)
         );
  AOI211_X1 U4266 ( .C1(n3464), .C2(n2153), .A(n4644), .B(n3463), .ZN(n3465)
         );
  OAI211_X1 U4267 ( .C1(n4519), .C2(n4021), .A(n3466), .B(n3465), .ZN(U3225)
         );
  NOR2_X1 U4268 ( .A1(n3467), .A2(n2167), .ZN(n3469) );
  XNOR2_X1 U4269 ( .A(n3469), .B(n3468), .ZN(n3475) );
  INV_X1 U4270 ( .A(n3470), .ZN(n3890) );
  OAI22_X1 U4271 ( .A1(n3513), .A2(n3888), .B1(STATE_REG_SCAN_IN), .B2(n3471), 
        .ZN(n3473) );
  OAI22_X1 U4272 ( .A1(n3885), .A2(n4504), .B1(n4503), .B2(n3847), .ZN(n3472)
         );
  AOI211_X1 U4273 ( .C1(n3890), .C2(n3517), .A(n3473), .B(n3472), .ZN(n3474)
         );
  OAI21_X1 U4274 ( .B1(n3475), .B2(n3519), .A(n3474), .ZN(U3226) );
  INV_X1 U4275 ( .A(n3476), .ZN(n3481) );
  AOI21_X1 U4276 ( .B1(n3480), .B2(n3478), .A(n3477), .ZN(n3479) );
  AOI21_X1 U4277 ( .B1(n3481), .B2(n3480), .A(n3479), .ZN(n3487) );
  INV_X1 U4278 ( .A(n3482), .ZN(n3963) );
  INV_X1 U4279 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3483) );
  OAI22_X1 U4280 ( .A1(n3513), .A2(n3962), .B1(STATE_REG_SCAN_IN), .B2(n3483), 
        .ZN(n3485) );
  OAI22_X1 U4281 ( .A1(n3502), .A2(n4504), .B1(n4503), .B2(n3956), .ZN(n3484)
         );
  AOI211_X1 U4282 ( .C1(n3963), .C2(n3517), .A(n3485), .B(n3484), .ZN(n3486)
         );
  OAI21_X1 U4283 ( .B1(n3487), .B2(n3519), .A(n3486), .ZN(U3230) );
  OAI21_X1 U4284 ( .B1(n3490), .B2(n3489), .A(n3488), .ZN(n3491) );
  NAND2_X1 U4285 ( .A1(n3491), .A2(n4514), .ZN(n3496) );
  NOR2_X1 U4286 ( .A1(n3513), .A2(n3492), .ZN(n3494) );
  OAI22_X1 U4287 ( .A1(n3885), .A2(n4503), .B1(n4504), .B2(n3956), .ZN(n3493)
         );
  AOI211_X1 U4288 ( .C1(REG3_REG_22__SCAN_IN), .C2(U3149), .A(n3494), .B(n3493), .ZN(n3495) );
  OAI211_X1 U4289 ( .C1(n4519), .C2(n3927), .A(n3496), .B(n3495), .ZN(U3232)
         );
  XNOR2_X1 U4290 ( .A(n3498), .B(n3497), .ZN(n3499) );
  XNOR2_X1 U4291 ( .A(n3500), .B(n3499), .ZN(n3501) );
  NAND2_X1 U4292 ( .A1(n3501), .A2(n4514), .ZN(n3505) );
  INV_X1 U4293 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4417) );
  NOR2_X1 U4294 ( .A1(STATE_REG_SCAN_IN), .A2(n4417), .ZN(n3797) );
  OAI22_X1 U4295 ( .A1(n3502), .A2(n4503), .B1(n4504), .B2(n4491), .ZN(n3503)
         );
  AOI211_X1 U4296 ( .C1(n3994), .C2(n2153), .A(n3797), .B(n3503), .ZN(n3504)
         );
  OAI211_X1 U4297 ( .C1(n4519), .C2(n4004), .A(n3505), .B(n3504), .ZN(U3235)
         );
  INV_X1 U4298 ( .A(n3506), .ZN(n3508) );
  NOR2_X1 U4299 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  XNOR2_X1 U4300 ( .A(n3510), .B(n3509), .ZN(n3520) );
  INV_X1 U4301 ( .A(n3511), .ZN(n3851) );
  OAI22_X1 U4302 ( .A1(n3513), .A2(n3850), .B1(STATE_REG_SCAN_IN), .B2(n3512), 
        .ZN(n3516) );
  OAI22_X1 U4303 ( .A1(n3847), .A2(n4504), .B1(n4503), .B2(n3514), .ZN(n3515)
         );
  AOI211_X1 U4304 ( .C1(n3851), .C2(n3517), .A(n3516), .B(n3515), .ZN(n3518)
         );
  OAI21_X1 U4305 ( .B1(n3520), .B2(n3519), .A(n3518), .ZN(U3237) );
  NAND2_X1 U4306 ( .A1(n3526), .A2(DATAI_30_), .ZN(n4065) );
  INV_X1 U4307 ( .A(n3829), .ZN(n3525) );
  INV_X1 U4308 ( .A(n3574), .ZN(n3524) );
  NAND2_X1 U4309 ( .A1(n3682), .A2(n3521), .ZN(n3522) );
  NAND2_X1 U4310 ( .A1(n3523), .A2(n3522), .ZN(n3661) );
  NOR3_X1 U4311 ( .A1(n3525), .A2(n3524), .A3(n3661), .ZN(n3551) );
  OR2_X1 U4312 ( .A1(n3681), .A2(n4065), .ZN(n3527) );
  NAND2_X1 U4313 ( .A1(n3526), .A2(DATAI_31_), .ZN(n4059) );
  NAND2_X1 U4314 ( .A1(n4061), .A2(n4059), .ZN(n3665) );
  AND2_X1 U4315 ( .A1(n3527), .A2(n3665), .ZN(n3578) );
  INV_X1 U4316 ( .A(n3682), .ZN(n3529) );
  NAND2_X1 U4317 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  NAND2_X1 U4318 ( .A1(n3578), .A2(n3530), .ZN(n3534) );
  INV_X1 U4319 ( .A(n3534), .ZN(n3535) );
  NAND2_X1 U4320 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  NOR2_X1 U4321 ( .A1(n3534), .A2(n3533), .ZN(n3547) );
  AOI21_X1 U4322 ( .B1(n3535), .B2(n3661), .A(n3547), .ZN(n3668) );
  NAND2_X1 U4323 ( .A1(n3605), .A2(n3604), .ZN(n3538) );
  NAND2_X1 U4324 ( .A1(n3537), .A2(n3536), .ZN(n3639) );
  NAND2_X1 U4325 ( .A1(n3639), .A2(n3604), .ZN(n3597) );
  OAI21_X1 U4326 ( .B1(n3539), .B2(n3538), .A(n3597), .ZN(n3540) );
  AOI211_X1 U4327 ( .C1(n3540), .C2(n3651), .A(n2222), .B(n3648), .ZN(n3543)
         );
  OAI21_X1 U4328 ( .B1(n3543), .B2(n3542), .A(n3541), .ZN(n3545) );
  AOI21_X1 U4329 ( .B1(n3545), .B2(n3654), .A(n3544), .ZN(n3546) );
  OAI21_X1 U4330 ( .B1(n3546), .B2(n3656), .A(n3839), .ZN(n3549) );
  NAND3_X1 U4331 ( .A1(n3549), .A2(n3548), .A3(n3547), .ZN(n3550) );
  OAI21_X1 U4332 ( .B1(n3551), .B2(n3668), .A(n3550), .ZN(n3552) );
  OAI21_X1 U4333 ( .B1(n4065), .B2(n4061), .A(n3552), .ZN(n3556) );
  INV_X1 U4334 ( .A(n3681), .ZN(n3553) );
  INV_X1 U4335 ( .A(n4065), .ZN(n4068) );
  NOR2_X1 U4336 ( .A1(n3553), .A2(n4068), .ZN(n3576) );
  INV_X1 U4337 ( .A(n4061), .ZN(n3577) );
  INV_X1 U4338 ( .A(n4059), .ZN(n4062) );
  OAI21_X1 U4339 ( .B1(n3576), .B2(n3577), .A(n4062), .ZN(n3555) );
  AOI21_X1 U4340 ( .B1(n3556), .B2(n3555), .A(n3554), .ZN(n3673) );
  INV_X1 U4341 ( .A(n3557), .ZN(n3876) );
  NOR2_X1 U4342 ( .A1(n3558), .A2(n3876), .ZN(n3900) );
  INV_X1 U4343 ( .A(n3900), .ZN(n3562) );
  NAND2_X1 U4344 ( .A1(n3840), .A2(n3559), .ZN(n3860) );
  NAND2_X1 U4345 ( .A1(n3560), .A2(n3859), .ZN(n3878) );
  NOR4_X1 U4346 ( .A1(n3562), .A2(n3860), .A3(n3878), .A4(n3561), .ZN(n3585)
         );
  INV_X1 U4347 ( .A(n3897), .ZN(n3563) );
  OR2_X1 U4348 ( .A1(n3898), .A2(n3563), .ZN(n3935) );
  INV_X1 U4349 ( .A(n3935), .ZN(n3583) );
  INV_X1 U4350 ( .A(n3564), .ZN(n3565) );
  NOR2_X1 U4351 ( .A1(n3566), .A2(n3565), .ZN(n3954) );
  INV_X1 U4352 ( .A(n3567), .ZN(n3569) );
  NAND4_X1 U4353 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3581)
         );
  NAND4_X1 U4354 ( .A1(n3573), .A2(n3572), .A3(n4000), .A4(n4033), .ZN(n3580)
         );
  AOI21_X1 U4355 ( .B1(n3577), .B2(n4062), .A(n3576), .ZN(n3666) );
  NAND4_X1 U4356 ( .A1(n3829), .A2(n3842), .A3(n3578), .A4(n3666), .ZN(n3579)
         );
  NOR4_X1 U4357 ( .A1(n3954), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3582)
         );
  NAND4_X1 U4358 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3595)
         );
  NAND2_X1 U4359 ( .A1(n3969), .A2(n3970), .ZN(n4017) );
  NOR4_X1 U4360 ( .A1(n2691), .A2(n3586), .A3(n4017), .A4(n4659), .ZN(n3591)
         );
  INV_X1 U4361 ( .A(n3918), .ZN(n3917) );
  NOR4_X1 U4362 ( .A1(n3917), .A2(n3589), .A3(n3588), .A4(n3587), .ZN(n3590)
         );
  NAND2_X1 U4363 ( .A1(n3591), .A2(n3590), .ZN(n3594) );
  XNOR2_X1 U4364 ( .A(n3995), .B(n3986), .ZN(n3983) );
  INV_X1 U4365 ( .A(n4681), .ZN(n4673) );
  NAND2_X1 U4366 ( .A1(n3697), .A2(n4709), .ZN(n3614) );
  AND2_X1 U4367 ( .A1(n3613), .A2(n3614), .ZN(n4699) );
  NAND4_X1 U4368 ( .A1(n3592), .A2(n4673), .A3(n2175), .A4(n4699), .ZN(n3593)
         );
  NOR2_X1 U4369 ( .A1(n3596), .A2(n2720), .ZN(n3671) );
  INV_X1 U4370 ( .A(n3597), .ZN(n3645) );
  NAND2_X1 U4371 ( .A1(n2182), .A2(n3598), .ZN(n3607) );
  NAND2_X1 U4372 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  NOR2_X1 U4373 ( .A1(n3607), .A2(n3601), .ZN(n3641) );
  INV_X1 U4374 ( .A(n3602), .ZN(n3612) );
  NAND3_X1 U4375 ( .A1(n3605), .A2(n3604), .A3(n3603), .ZN(n3611) );
  INV_X1 U4376 ( .A(n3606), .ZN(n3608) );
  AOI21_X1 U4377 ( .B1(n3609), .B2(n3608), .A(n3607), .ZN(n3610) );
  AOI211_X1 U4378 ( .C1(n3641), .C2(n3612), .A(n3611), .B(n3610), .ZN(n3644)
         );
  INV_X1 U4379 ( .A(n3613), .ZN(n4672) );
  OAI211_X1 U4380 ( .C1(n4672), .C2(n2720), .A(n3615), .B(n3614), .ZN(n3617)
         );
  NAND3_X1 U4381 ( .A1(n3617), .A2(n3616), .A3(n2690), .ZN(n3619) );
  OAI211_X1 U4382 ( .C1(n3621), .C2(n3620), .A(n3619), .B(n3618), .ZN(n3624)
         );
  NAND3_X1 U4383 ( .A1(n3624), .A2(n3623), .A3(n3622), .ZN(n3626) );
  NAND4_X1 U4384 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3635), .ZN(n3629)
         );
  NAND3_X1 U4385 ( .A1(n3629), .A2(n2175), .A3(n3628), .ZN(n3630) );
  NAND3_X1 U4386 ( .A1(n3630), .A2(n3637), .A3(n3636), .ZN(n3633) );
  AND3_X1 U4387 ( .A1(n3633), .A2(n3632), .A3(n3631), .ZN(n3640) );
  NAND4_X1 U4388 ( .A1(n2211), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3638)
         );
  OAI22_X1 U4389 ( .A1(n3640), .A2(n3639), .B1(n3645), .B2(n3638), .ZN(n3642)
         );
  NAND3_X1 U4390 ( .A1(n3642), .A2(n3641), .A3(n2176), .ZN(n3643) );
  OAI21_X1 U4391 ( .B1(n3645), .B2(n3644), .A(n3643), .ZN(n3646) );
  NAND2_X1 U4392 ( .A1(n3647), .A2(n3646), .ZN(n3650) );
  AOI211_X1 U4393 ( .C1(n3651), .C2(n3650), .A(n3649), .B(n3648), .ZN(n3653)
         );
  NOR2_X1 U4394 ( .A1(n3653), .A2(n3652), .ZN(n3655) );
  OAI21_X1 U4395 ( .B1(n3898), .B2(n3655), .A(n3654), .ZN(n3659) );
  AOI211_X1 U4396 ( .C1(n3659), .C2(n3658), .A(n3657), .B(n3656), .ZN(n3664)
         );
  INV_X1 U4397 ( .A(n3660), .ZN(n3663) );
  NOR4_X1 U4398 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3669)
         );
  INV_X1 U4399 ( .A(n3665), .ZN(n3667) );
  OAI22_X1 U4400 ( .A1(n3669), .A2(n3668), .B1(n3667), .B2(n3666), .ZN(n3670)
         );
  MUX2_X1 U4401 ( .A(n3671), .B(n3670), .S(n2687), .Z(n3672) );
  NOR2_X1 U4402 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  XNOR2_X1 U4403 ( .A(n3674), .B(n4484), .ZN(n3680) );
  NAND2_X1 U4404 ( .A1(n3676), .A2(n3675), .ZN(n3677) );
  OAI211_X1 U4405 ( .C1(n4482), .C2(n3679), .A(n3677), .B(B_REG_SCAN_IN), .ZN(
        n3678) );
  OAI21_X1 U4406 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(U3239) );
  MUX2_X1 U4407 ( .A(n3681), .B(DATAO_REG_30__SCAN_IN), .S(n3696), .Z(U3580)
         );
  MUX2_X1 U4408 ( .A(n3682), .B(DATAO_REG_29__SCAN_IN), .S(n3696), .Z(U3579)
         );
  MUX2_X1 U4409 ( .A(DATAO_REG_28__SCAN_IN), .B(n3832), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4410 ( .A(DATAO_REG_27__SCAN_IN), .B(n3845), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4411 ( .A(n3864), .B(DATAO_REG_26__SCAN_IN), .S(n3696), .Z(U3576)
         );
  MUX2_X1 U4412 ( .A(n3882), .B(DATAO_REG_25__SCAN_IN), .S(n3696), .Z(U3575)
         );
  MUX2_X1 U4413 ( .A(DATAO_REG_24__SCAN_IN), .B(n3683), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4414 ( .A(DATAO_REG_23__SCAN_IN), .B(n3922), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4415 ( .A(DATAO_REG_22__SCAN_IN), .B(n3938), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4416 ( .A(n3939), .B(DATAO_REG_20__SCAN_IN), .S(n3696), .Z(U3570)
         );
  MUX2_X1 U4417 ( .A(n3995), .B(DATAO_REG_19__SCAN_IN), .S(n3696), .Z(U3569)
         );
  MUX2_X1 U4418 ( .A(DATAO_REG_18__SCAN_IN), .B(n3979), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4419 ( .A(DATAO_REG_17__SCAN_IN), .B(n3684), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4420 ( .A(DATAO_REG_16__SCAN_IN), .B(n4013), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4421 ( .A(DATAO_REG_15__SCAN_IN), .B(n3685), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4422 ( .A(DATAO_REG_14__SCAN_IN), .B(n3686), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4423 ( .A(n3687), .B(DATAO_REG_13__SCAN_IN), .S(n3696), .Z(U3563)
         );
  MUX2_X1 U4424 ( .A(n3688), .B(DATAO_REG_12__SCAN_IN), .S(n3696), .Z(U3562)
         );
  MUX2_X1 U4425 ( .A(DATAO_REG_11__SCAN_IN), .B(n3689), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4426 ( .A(n4656), .B(DATAO_REG_10__SCAN_IN), .S(n3696), .Z(U3560)
         );
  MUX2_X1 U4427 ( .A(n3690), .B(DATAO_REG_9__SCAN_IN), .S(n3696), .Z(U3559) );
  MUX2_X1 U4428 ( .A(n3691), .B(DATAO_REG_8__SCAN_IN), .S(n3696), .Z(U3558) );
  MUX2_X1 U4429 ( .A(DATAO_REG_7__SCAN_IN), .B(n3692), .S(U4043), .Z(U3557) );
  MUX2_X1 U4430 ( .A(n3693), .B(DATAO_REG_6__SCAN_IN), .S(n3696), .Z(U3556) );
  MUX2_X1 U4431 ( .A(n3694), .B(DATAO_REG_5__SCAN_IN), .S(n3696), .Z(U3555) );
  MUX2_X1 U4432 ( .A(DATAO_REG_4__SCAN_IN), .B(n3695), .S(U4043), .Z(U3554) );
  MUX2_X1 U4433 ( .A(n4046), .B(DATAO_REG_3__SCAN_IN), .S(n3696), .Z(U3553) );
  MUX2_X1 U4434 ( .A(DATAO_REG_2__SCAN_IN), .B(n4676), .S(U4043), .Z(U3552) );
  MUX2_X1 U4435 ( .A(DATAO_REG_1__SCAN_IN), .B(n2840), .S(U4043), .Z(U3551) );
  MUX2_X1 U4436 ( .A(DATAO_REG_0__SCAN_IN), .B(n3697), .S(U4043), .Z(U3550) );
  NAND3_X1 U4437 ( .A1(n4646), .A2(IR_REG_0__SCAN_IN), .A3(n2800), .ZN(n3706)
         );
  AOI22_X1 U4438 ( .A1(n4645), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3705) );
  AOI21_X1 U4439 ( .B1(n2800), .B2(n3698), .A(n3701), .ZN(n3700) );
  MUX2_X1 U4440 ( .A(n3701), .B(n3700), .S(n3699), .Z(n3703) );
  NAND2_X1 U4441 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  NAND3_X1 U4442 ( .A1(n3706), .A2(n3705), .A3(n3704), .ZN(U3240) );
  OAI211_X1 U4443 ( .C1(n3709), .C2(n3708), .A(n4610), .B(n3707), .ZN(n3716)
         );
  OAI211_X1 U4444 ( .C1(n3712), .C2(n3711), .A(n4646), .B(n3710), .ZN(n3715)
         );
  INV_X1 U4445 ( .A(n4653), .ZN(n3783) );
  NAND2_X1 U4446 ( .A1(n3783), .A2(n4490), .ZN(n3714) );
  AOI22_X1 U4447 ( .A1(n4645), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3713) );
  NAND4_X1 U4448 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(U3241)
         );
  AOI22_X1 U4449 ( .A1(n4645), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3727) );
  OAI211_X1 U4450 ( .C1(n3719), .C2(n3718), .A(n4610), .B(n3717), .ZN(n3724)
         );
  OAI211_X1 U4451 ( .C1(n3722), .C2(n3721), .A(n4646), .B(n3720), .ZN(n3723)
         );
  AND2_X1 U4452 ( .A1(n3724), .A2(n3723), .ZN(n3726) );
  NAND2_X1 U4453 ( .A1(n3783), .A2(n4489), .ZN(n3725) );
  NAND4_X1 U4454 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(U3242)
         );
  INV_X1 U4455 ( .A(n3778), .ZN(n4735) );
  AOI22_X1 U4456 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3778), .B1(n4735), .B2(
        n4119), .ZN(n4636) );
  INV_X1 U4457 ( .A(n3774), .ZN(n4739) );
  AOI22_X1 U4458 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3774), .B1(n4739), .B2(
        n4271), .ZN(n4618) );
  INV_X1 U4459 ( .A(n4741), .ZN(n4595) );
  AOI22_X1 U4460 ( .A1(n4741), .A2(REG1_REG_11__SCAN_IN), .B1(n2523), .B2(
        n4595), .ZN(n4589) );
  INV_X1 U4461 ( .A(n4486), .ZN(n4574) );
  NAND2_X1 U4462 ( .A1(n3729), .A2(n4487), .ZN(n3730) );
  INV_X1 U4463 ( .A(n3753), .ZN(n4751) );
  AOI22_X1 U4464 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4751), .B1(n3753), .B2(n2452), .ZN(n4528) );
  NOR2_X1 U4465 ( .A1(n3733), .A2(n2304), .ZN(n3734) );
  NAND2_X1 U4466 ( .A1(n3763), .A2(n3738), .ZN(n3739) );
  INV_X1 U4467 ( .A(n3763), .ZN(n4746) );
  NAND2_X1 U4468 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U4469 ( .A1(n3739), .A2(n4557), .ZN(n4568) );
  MUX2_X1 U4470 ( .A(REG1_REG_9__SCAN_IN), .B(n3740), .S(n4486), .Z(n4567) );
  NAND2_X1 U4471 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OAI21_X1 U4472 ( .B1(n3740), .B2(n4574), .A(n4566), .ZN(n3741) );
  NAND2_X1 U4473 ( .A1(n3767), .A2(n3741), .ZN(n3742) );
  INV_X1 U4474 ( .A(n3767), .ZN(n4744) );
  XNOR2_X1 U4475 ( .A(n3741), .B(n4744), .ZN(n4579) );
  NAND2_X1 U4476 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U4477 ( .A1(n3772), .A2(n3743), .ZN(n3744) );
  NAND2_X1 U4478 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U4479 ( .A1(n4736), .A2(n3745), .ZN(n3746) );
  NAND2_X1 U4480 ( .A1(n3746), .A2(n4625), .ZN(n4635) );
  NAND2_X1 U4481 ( .A1(n4636), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U4482 ( .A1(n3778), .A2(REG1_REG_15__SCAN_IN), .ZN(n3747) );
  INV_X1 U4483 ( .A(n4485), .ZN(n3791) );
  AOI21_X1 U4484 ( .B1(n3748), .B2(REG1_REG_16__SCAN_IN), .A(n3787), .ZN(n3785) );
  INV_X1 U4485 ( .A(n4646), .ZN(n4537) );
  INV_X1 U4486 ( .A(n4645), .ZN(n3751) );
  INV_X1 U4487 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n3750) );
  NOR2_X1 U4488 ( .A1(STATE_REG_SCAN_IN), .A2(n4361), .ZN(n4494) );
  INV_X1 U4489 ( .A(n4494), .ZN(n3749) );
  OAI21_X1 U4490 ( .B1(n3751), .B2(n3750), .A(n3749), .ZN(n3782) );
  NOR2_X1 U4491 ( .A1(n4609), .A2(n4739), .ZN(n4608) );
  INV_X1 U4492 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4493 ( .A1(n4741), .A2(REG2_REG_11__SCAN_IN), .B1(n3770), .B2(
        n4595), .ZN(n4592) );
  NAND2_X1 U4494 ( .A1(n4486), .A2(REG2_REG_9__SCAN_IN), .ZN(n3766) );
  MUX2_X1 U4495 ( .A(REG2_REG_9__SCAN_IN), .B(n3068), .S(n4486), .Z(n4570) );
  NAND2_X1 U4496 ( .A1(n4546), .A2(REG2_REG_7__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4497 ( .A1(n4546), .A2(REG2_REG_7__SCAN_IN), .B1(n3752), .B2(n4748), .ZN(n4554) );
  AOI22_X1 U4498 ( .A1(REG2_REG_5__SCAN_IN), .A2(n3753), .B1(n4751), .B2(n3758), .ZN(n4534) );
  NAND2_X1 U4499 ( .A1(n3754), .A2(REG2_REG_4__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4500 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  NAND2_X1 U4501 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4543), .ZN(n4542) );
  NAND2_X1 U4502 ( .A1(n3761), .A2(n4542), .ZN(n4553) );
  NAND2_X1 U4503 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  NAND2_X1 U4504 ( .A1(n3762), .A2(n4552), .ZN(n3764) );
  NAND2_X1 U4505 ( .A1(n3763), .A2(n3764), .ZN(n3765) );
  XNOR2_X1 U4506 ( .A(n3764), .B(n4746), .ZN(n4560) );
  NAND2_X1 U4507 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U4508 ( .A1(n3765), .A2(n4559), .ZN(n4571) );
  NAND2_X1 U4509 ( .A1(n4570), .A2(n4571), .ZN(n4569) );
  NAND2_X1 U4510 ( .A1(n3766), .A2(n4569), .ZN(n3768) );
  NAND2_X1 U4511 ( .A1(n3767), .A2(n3768), .ZN(n3769) );
  XNOR2_X1 U4512 ( .A(n3768), .B(n4744), .ZN(n4581) );
  NAND2_X1 U4513 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U4514 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  NAND2_X1 U4515 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4600), .ZN(n4599) );
  NOR2_X1 U4516 ( .A1(n2293), .A2(n3775), .ZN(n3776) );
  NOR2_X1 U4517 ( .A1(n3776), .A2(n4621), .ZN(n4631) );
  NAND2_X1 U4518 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3778), .ZN(n3777) );
  OAI21_X1 U4519 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3778), .A(n3777), .ZN(n4630) );
  NOR2_X1 U4520 ( .A1(n4631), .A2(n4630), .ZN(n4629) );
  AND2_X1 U4521 ( .A1(n3778), .A2(REG2_REG_15__SCAN_IN), .ZN(n3779) );
  NOR2_X1 U4522 ( .A1(n4629), .A2(n3779), .ZN(n3792) );
  XNOR2_X1 U4523 ( .A(n3792), .B(n4485), .ZN(n3780) );
  INV_X1 U4524 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4227) );
  NAND2_X1 U4525 ( .A1(n3780), .A2(n4227), .ZN(n3793) );
  AOI221_X1 U4526 ( .B1(n3780), .B2(n3793), .C1(n4227), .C2(n3793), .A(n4639), 
        .ZN(n3781) );
  AOI211_X1 U4527 ( .C1(n3783), .C2(n4485), .A(n3782), .B(n3781), .ZN(n3784)
         );
  OAI21_X1 U4528 ( .B1(n3785), .B2(n4537), .A(n3784), .ZN(U3256) );
  XNOR2_X1 U4529 ( .A(n3799), .B(REG1_REG_18__SCAN_IN), .ZN(n3802) );
  INV_X1 U4530 ( .A(n4732), .ZN(n4652) );
  INV_X1 U4531 ( .A(n3786), .ZN(n3788) );
  AOI22_X1 U4532 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4652), .B1(n4732), .B2(
        n4274), .ZN(n4647) );
  INV_X1 U4533 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3790) );
  NOR2_X1 U4534 ( .A1(n3807), .A2(n3790), .ZN(n3789) );
  AOI21_X1 U4535 ( .B1(n3807), .B2(n3790), .A(n3789), .ZN(n3796) );
  INV_X1 U4536 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4537 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4732), .B1(n4652), .B2(
        n4406), .ZN(n4642) );
  NAND2_X1 U4538 ( .A1(n3792), .A2(n3791), .ZN(n3794) );
  NAND2_X1 U4539 ( .A1(n3794), .A2(n3793), .ZN(n4640) );
  NAND2_X1 U4540 ( .A1(n4642), .A2(n4640), .ZN(n4641) );
  OAI21_X1 U4541 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4732), .A(n4641), .ZN(n3795) );
  AOI211_X1 U4542 ( .C1(n3796), .C2(n3795), .A(n3806), .B(n4639), .ZN(n3801)
         );
  AOI21_X1 U4543 ( .B1(n4645), .B2(ADDR_REG_18__SCAN_IN), .A(n3797), .ZN(n3798) );
  OAI21_X1 U4544 ( .B1(n3799), .B2(n4653), .A(n3798), .ZN(n3800) );
  AOI22_X1 U4545 ( .A1(n3803), .A2(n3802), .B1(REG1_REG_18__SCAN_IN), .B2(
        n3807), .ZN(n3805) );
  XNOR2_X1 U4546 ( .A(n3811), .B(n4104), .ZN(n3804) );
  XNOR2_X1 U4547 ( .A(n3805), .B(n3804), .ZN(n3814) );
  XNOR2_X1 U4548 ( .A(n3811), .B(REG2_REG_19__SCAN_IN), .ZN(n3808) );
  AOI21_X1 U4549 ( .B1(n4645), .B2(ADDR_REG_19__SCAN_IN), .A(n3809), .ZN(n3810) );
  OAI21_X1 U4550 ( .B1(n3811), .B2(n4653), .A(n3810), .ZN(n3812) );
  OAI21_X1 U4551 ( .B1(n3814), .B2(n4537), .A(n3813), .ZN(U3259) );
  INV_X1 U4552 ( .A(n3815), .ZN(n3823) );
  INV_X1 U4553 ( .A(n3816), .ZN(n3817) );
  AOI22_X1 U4554 ( .A1(n4700), .A2(REG2_REG_28__SCAN_IN), .B1(n3817), .B2(
        n4688), .ZN(n3818) );
  OAI21_X1 U4555 ( .B1(n3819), .B2(n4040), .A(n3818), .ZN(n3820) );
  AOI21_X1 U4556 ( .B1(n3821), .B2(n4712), .A(n3820), .ZN(n3822) );
  OAI21_X1 U4557 ( .B1(n3823), .B2(n3967), .A(n3822), .ZN(U3262) );
  XOR2_X1 U4558 ( .A(n3829), .B(n3824), .Z(n4076) );
  AOI21_X1 U4559 ( .B1(n3831), .B2(n2155), .A(n2308), .ZN(n4074) );
  INV_X1 U4560 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3826) );
  OAI22_X1 U4561 ( .A1(n4712), .A2(n3826), .B1(n3825), .B2(n4716), .ZN(n3827)
         );
  AOI21_X1 U4562 ( .B1(n4074), .B2(n4696), .A(n3827), .ZN(n3837) );
  OAI21_X1 U4563 ( .B1(n2174), .B2(n3829), .A(n3828), .ZN(n3830) );
  NAND2_X1 U4564 ( .A1(n3830), .A2(n4702), .ZN(n3834) );
  AOI22_X1 U4565 ( .A1(n3832), .A2(n4675), .B1(n3831), .B2(n4674), .ZN(n3833)
         );
  OAI211_X1 U4566 ( .C1(n3835), .C2(n4678), .A(n3834), .B(n3833), .ZN(n4073)
         );
  NAND2_X1 U4567 ( .A1(n4073), .A2(n4712), .ZN(n3836) );
  OAI211_X1 U4568 ( .C1(n4076), .C2(n3967), .A(n3837), .B(n3836), .ZN(U3263)
         );
  XNOR2_X1 U4569 ( .A(n3838), .B(n3842), .ZN(n4080) );
  INV_X1 U4570 ( .A(n4080), .ZN(n3856) );
  INV_X1 U4571 ( .A(n3839), .ZN(n3841) );
  OAI21_X1 U4572 ( .B1(n3858), .B2(n3841), .A(n3840), .ZN(n3843) );
  XNOR2_X1 U4573 ( .A(n3843), .B(n3842), .ZN(n3849) );
  AOI22_X1 U4574 ( .A1(n3845), .A2(n4675), .B1(n4674), .B2(n3844), .ZN(n3846)
         );
  OAI21_X1 U4575 ( .B1(n3847), .B2(n4678), .A(n3846), .ZN(n3848) );
  AOI21_X1 U4576 ( .B1(n3849), .B2(n4702), .A(n3848), .ZN(n4077) );
  INV_X1 U4577 ( .A(n4077), .ZN(n3854) );
  OAI21_X1 U4578 ( .B1(n3867), .B2(n3850), .A(n2155), .ZN(n4078) );
  AOI22_X1 U4579 ( .A1(n4700), .A2(REG2_REG_26__SCAN_IN), .B1(n3851), .B2(
        n4688), .ZN(n3852) );
  OAI21_X1 U4580 ( .B1(n4078), .B2(n4040), .A(n3852), .ZN(n3853) );
  AOI21_X1 U4581 ( .B1(n3854), .B2(n4712), .A(n3853), .ZN(n3855) );
  OAI21_X1 U4582 ( .B1(n3856), .B2(n3967), .A(n3855), .ZN(U3264) );
  XOR2_X1 U4583 ( .A(n3860), .B(n3857), .Z(n4083) );
  INV_X1 U4584 ( .A(n4083), .ZN(n3874) );
  NAND2_X1 U4585 ( .A1(n2203), .A2(n3859), .ZN(n3861) );
  XNOR2_X1 U4586 ( .A(n3861), .B(n3860), .ZN(n3862) );
  NAND2_X1 U4587 ( .A1(n3862), .A2(n4702), .ZN(n3866) );
  AOI22_X1 U4588 ( .A1(n3864), .A2(n4675), .B1(n4674), .B2(n3863), .ZN(n3865)
         );
  OAI211_X1 U4589 ( .C1(n3906), .C2(n4678), .A(n3866), .B(n3865), .ZN(n4082)
         );
  INV_X1 U4590 ( .A(n3867), .ZN(n3868) );
  OAI21_X1 U4591 ( .B1(n3886), .B2(n3869), .A(n3868), .ZN(n4439) );
  AOI22_X1 U4592 ( .A1(n4700), .A2(REG2_REG_25__SCAN_IN), .B1(n3870), .B2(
        n4688), .ZN(n3871) );
  OAI21_X1 U4593 ( .B1(n4439), .B2(n4040), .A(n3871), .ZN(n3872) );
  AOI21_X1 U4594 ( .B1(n4082), .B2(n4712), .A(n3872), .ZN(n3873) );
  OAI21_X1 U4595 ( .B1(n3874), .B2(n3967), .A(n3873), .ZN(U3265) );
  XNOR2_X1 U4596 ( .A(n3875), .B(n3878), .ZN(n4086) );
  INV_X1 U4597 ( .A(n4086), .ZN(n3894) );
  NOR2_X1 U4598 ( .A1(n3877), .A2(n3876), .ZN(n3879) );
  XNOR2_X1 U4599 ( .A(n3879), .B(n3878), .ZN(n3880) );
  NAND2_X1 U4600 ( .A1(n3880), .A2(n4702), .ZN(n3884) );
  AOI22_X1 U4601 ( .A1(n3882), .A2(n4675), .B1(n4674), .B2(n3881), .ZN(n3883)
         );
  OAI211_X1 U4602 ( .C1(n3885), .C2(n4678), .A(n3884), .B(n3883), .ZN(n4085)
         );
  INV_X1 U4603 ( .A(n3907), .ZN(n3889) );
  INV_X1 U4604 ( .A(n3886), .ZN(n3887) );
  OAI21_X1 U4605 ( .B1(n3889), .B2(n3888), .A(n3887), .ZN(n4443) );
  AOI22_X1 U4606 ( .A1(n4700), .A2(REG2_REG_24__SCAN_IN), .B1(n3890), .B2(
        n4688), .ZN(n3891) );
  OAI21_X1 U4607 ( .B1(n4443), .B2(n4040), .A(n3891), .ZN(n3892) );
  AOI21_X1 U4608 ( .B1(n4085), .B2(n4712), .A(n3892), .ZN(n3893) );
  OAI21_X1 U4609 ( .B1(n3894), .B2(n3967), .A(n3893), .ZN(U3266) );
  OR2_X1 U4610 ( .A1(n3915), .A2(n3918), .ZN(n3916) );
  NAND2_X1 U4611 ( .A1(n3916), .A2(n3895), .ZN(n3896) );
  XNOR2_X1 U4612 ( .A(n3896), .B(n3900), .ZN(n4089) );
  INV_X1 U4613 ( .A(n4089), .ZN(n3914) );
  OAI21_X1 U4614 ( .B1(n3936), .B2(n3898), .A(n3897), .ZN(n3919) );
  NAND2_X1 U4615 ( .A1(n3919), .A2(n3918), .ZN(n3921) );
  NAND2_X1 U4616 ( .A1(n3921), .A2(n3899), .ZN(n3901) );
  XNOR2_X1 U4617 ( .A(n3901), .B(n3900), .ZN(n3902) );
  NAND2_X1 U4618 ( .A1(n3902), .A2(n4702), .ZN(n3905) );
  AOI22_X1 U4619 ( .A1(n3938), .A2(n4655), .B1(n4674), .B2(n3903), .ZN(n3904)
         );
  OAI211_X1 U4620 ( .C1(n3906), .C2(n4705), .A(n3905), .B(n3904), .ZN(n4088)
         );
  INV_X1 U4621 ( .A(n4092), .ZN(n3909) );
  OAI21_X1 U4622 ( .B1(n3909), .B2(n3908), .A(n3907), .ZN(n4447) );
  AOI22_X1 U4623 ( .A1(n4700), .A2(REG2_REG_23__SCAN_IN), .B1(n3910), .B2(
        n4688), .ZN(n3911) );
  OAI21_X1 U4624 ( .B1(n4447), .B2(n4040), .A(n3911), .ZN(n3912) );
  AOI21_X1 U4625 ( .B1(n4088), .B2(n4712), .A(n3912), .ZN(n3913) );
  OAI21_X1 U4626 ( .B1(n3914), .B2(n3967), .A(n3913), .ZN(U3267) );
  OAI21_X1 U4627 ( .B1(n2242), .B2(n3917), .A(n3916), .ZN(n4095) );
  OR2_X1 U4628 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  NAND2_X1 U4629 ( .A1(n3921), .A2(n3920), .ZN(n3926) );
  NAND2_X1 U4630 ( .A1(n3929), .A2(n4674), .ZN(n3924) );
  NAND2_X1 U4631 ( .A1(n3922), .A2(n4675), .ZN(n3923) );
  OAI211_X1 U4632 ( .C1(n3956), .C2(n4678), .A(n3924), .B(n3923), .ZN(n3925)
         );
  AOI21_X1 U4633 ( .B1(n3926), .B2(n4702), .A(n3925), .ZN(n4094) );
  NOR2_X1 U4634 ( .A1(n4716), .A2(n3927), .ZN(n3928) );
  AOI21_X1 U4635 ( .B1(n4700), .B2(REG2_REG_22__SCAN_IN), .A(n3928), .ZN(n3931) );
  NAND2_X1 U4636 ( .A1(n3943), .A2(n3929), .ZN(n4091) );
  NAND3_X1 U4637 ( .A1(n4092), .A2(n4696), .A3(n4091), .ZN(n3930) );
  OAI211_X1 U4638 ( .C1(n4094), .C2(n4700), .A(n3931), .B(n3930), .ZN(n3932)
         );
  INV_X1 U4639 ( .A(n3932), .ZN(n3933) );
  OAI21_X1 U4640 ( .B1(n4095), .B2(n3967), .A(n3933), .ZN(U3268) );
  XOR2_X1 U4641 ( .A(n3935), .B(n3934), .Z(n4097) );
  INV_X1 U4642 ( .A(n4097), .ZN(n3949) );
  XOR2_X1 U4643 ( .A(n3936), .B(n3935), .Z(n3942) );
  AOI22_X1 U4644 ( .A1(n3938), .A2(n4675), .B1(n4674), .B2(n3937), .ZN(n3941)
         );
  NAND2_X1 U4645 ( .A1(n3939), .A2(n4655), .ZN(n3940) );
  OAI211_X1 U4646 ( .C1(n3942), .C2(n4015), .A(n3941), .B(n3940), .ZN(n4096)
         );
  OAI21_X1 U4647 ( .B1(n3960), .B2(n3944), .A(n3943), .ZN(n4452) );
  AOI22_X1 U4648 ( .A1(n4700), .A2(REG2_REG_21__SCAN_IN), .B1(n3945), .B2(
        n4688), .ZN(n3946) );
  OAI21_X1 U4649 ( .B1(n4452), .B2(n4040), .A(n3946), .ZN(n3947) );
  AOI21_X1 U4650 ( .B1(n4096), .B2(n4712), .A(n3947), .ZN(n3948) );
  OAI21_X1 U4651 ( .B1(n3949), .B2(n3967), .A(n3948), .ZN(U3269) );
  XNOR2_X1 U4652 ( .A(n3950), .B(n3954), .ZN(n4100) );
  INV_X1 U4653 ( .A(n4100), .ZN(n3968) );
  INV_X1 U4654 ( .A(n3951), .ZN(n3952) );
  NAND2_X1 U4655 ( .A1(n3953), .A2(n3952), .ZN(n3955) );
  XNOR2_X1 U4656 ( .A(n3955), .B(n3954), .ZN(n3959) );
  OAI22_X1 U4657 ( .A1(n3956), .A2(n4705), .B1(n4010), .B2(n3962), .ZN(n3957)
         );
  AOI21_X1 U4658 ( .B1(n4655), .B2(n3995), .A(n3957), .ZN(n3958) );
  OAI21_X1 U4659 ( .B1(n3959), .B2(n4015), .A(n3958), .ZN(n4099) );
  INV_X1 U4660 ( .A(n3960), .ZN(n3961) );
  OAI21_X1 U4661 ( .B1(n3984), .B2(n3962), .A(n3961), .ZN(n4456) );
  AOI22_X1 U4662 ( .A1(n4700), .A2(REG2_REG_20__SCAN_IN), .B1(n3963), .B2(
        n4688), .ZN(n3964) );
  OAI21_X1 U4663 ( .B1(n4456), .B2(n4040), .A(n3964), .ZN(n3965) );
  AOI21_X1 U4664 ( .B1(n4099), .B2(n4712), .A(n3965), .ZN(n3966) );
  OAI21_X1 U4665 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(U3270) );
  INV_X1 U4666 ( .A(n3969), .ZN(n3971) );
  OAI21_X1 U4667 ( .B1(n4009), .B2(n3971), .A(n3970), .ZN(n3993) );
  INV_X1 U4668 ( .A(n3972), .ZN(n3974) );
  OAI21_X1 U4669 ( .B1(n3993), .B2(n3974), .A(n3973), .ZN(n3976) );
  INV_X1 U4670 ( .A(n3983), .ZN(n3975) );
  XNOR2_X1 U4671 ( .A(n3976), .B(n3975), .ZN(n3981) );
  OAI22_X1 U4672 ( .A1(n3977), .A2(n4705), .B1(n4010), .B2(n3986), .ZN(n3978)
         );
  AOI21_X1 U4673 ( .B1(n4655), .B2(n3979), .A(n3978), .ZN(n3980) );
  OAI21_X1 U4674 ( .B1(n3981), .B2(n4015), .A(n3980), .ZN(n4102) );
  INV_X1 U4675 ( .A(n4102), .ZN(n3992) );
  XNOR2_X1 U4676 ( .A(n3982), .B(n3983), .ZN(n4103) );
  INV_X1 U4677 ( .A(n3984), .ZN(n3985) );
  OAI21_X1 U4678 ( .B1(n2321), .B2(n3986), .A(n3985), .ZN(n4460) );
  INV_X1 U4679 ( .A(n3987), .ZN(n3988) );
  AOI22_X1 U4680 ( .A1(n4700), .A2(REG2_REG_19__SCAN_IN), .B1(n3988), .B2(
        n4688), .ZN(n3989) );
  OAI21_X1 U4681 ( .B1(n4460), .B2(n4040), .A(n3989), .ZN(n3990) );
  AOI21_X1 U4682 ( .B1(n4103), .B2(n4042), .A(n3990), .ZN(n3991) );
  OAI21_X1 U4683 ( .B1(n3992), .B2(n4700), .A(n3991), .ZN(U3271) );
  XNOR2_X1 U4684 ( .A(n3993), .B(n4000), .ZN(n3998) );
  AOI22_X1 U4685 ( .A1(n3995), .A2(n4675), .B1(n3994), .B2(n4674), .ZN(n3996)
         );
  OAI21_X1 U4686 ( .B1(n4491), .B2(n4678), .A(n3996), .ZN(n3997) );
  AOI21_X1 U4687 ( .B1(n3998), .B2(n4702), .A(n3997), .ZN(n4107) );
  XOR2_X1 U4688 ( .A(n4000), .B(n3999), .Z(n4108) );
  INV_X1 U4689 ( .A(n4108), .ZN(n4007) );
  OAI211_X1 U4690 ( .C1(n2316), .C2(n4002), .A(n4001), .B(n4811), .ZN(n4106)
         );
  NOR2_X1 U4691 ( .A1(n4106), .A2(n4003), .ZN(n4006) );
  OAI22_X1 U4692 ( .A1(n4712), .A2(n3790), .B1(n4004), .B2(n4716), .ZN(n4005)
         );
  AOI211_X1 U4693 ( .C1(n4007), .C2(n4042), .A(n4006), .B(n4005), .ZN(n4008)
         );
  OAI21_X1 U4694 ( .B1(n4700), .B2(n4107), .A(n4008), .ZN(U3272) );
  XOR2_X1 U4695 ( .A(n4017), .B(n4009), .Z(n4016) );
  OAI22_X1 U4696 ( .A1(n4011), .A2(n4705), .B1(n4020), .B2(n4010), .ZN(n4012)
         );
  AOI21_X1 U4697 ( .B1(n4655), .B2(n4013), .A(n4012), .ZN(n4014) );
  OAI21_X1 U4698 ( .B1(n4016), .B2(n4015), .A(n4014), .ZN(n4109) );
  INV_X1 U4699 ( .A(n4109), .ZN(n4025) );
  XNOR2_X1 U4700 ( .A(n4018), .B(n4017), .ZN(n4110) );
  OAI21_X1 U4701 ( .B1(n4034), .B2(n4020), .A(n4019), .ZN(n4465) );
  NOR2_X1 U4702 ( .A1(n4465), .A2(n4040), .ZN(n4023) );
  OAI22_X1 U4703 ( .A1(n4712), .A2(n4406), .B1(n4021), .B2(n4716), .ZN(n4022)
         );
  AOI211_X1 U4704 ( .C1(n4110), .C2(n4042), .A(n4023), .B(n4022), .ZN(n4024)
         );
  OAI21_X1 U4705 ( .B1(n4025), .B2(n4700), .A(n4024), .ZN(U3273) );
  XNOR2_X1 U4706 ( .A(n4027), .B(n4026), .ZN(n4031) );
  OR2_X1 U4707 ( .A1(n4492), .A2(n4678), .ZN(n4029) );
  NAND2_X1 U4708 ( .A1(n4495), .A2(n4674), .ZN(n4028) );
  OAI211_X1 U4709 ( .C1(n4491), .C2(n4705), .A(n4029), .B(n4028), .ZN(n4030)
         );
  AOI21_X1 U4710 ( .B1(n4031), .B2(n4702), .A(n4030), .ZN(n4114) );
  XNOR2_X1 U4711 ( .A(n4032), .B(n4033), .ZN(n4112) );
  INV_X1 U4712 ( .A(n4034), .ZN(n4035) );
  OAI21_X1 U4713 ( .B1(n4037), .B2(n4036), .A(n4035), .ZN(n4469) );
  INV_X1 U4714 ( .A(n4501), .ZN(n4038) );
  AOI22_X1 U4715 ( .A1(n4700), .A2(REG2_REG_16__SCAN_IN), .B1(n4038), .B2(
        n4688), .ZN(n4039) );
  OAI21_X1 U4716 ( .B1(n4469), .B2(n4040), .A(n4039), .ZN(n4041) );
  AOI21_X1 U4717 ( .B1(n4112), .B2(n4042), .A(n4041), .ZN(n4043) );
  OAI21_X1 U4718 ( .B1(n4114), .B2(n4700), .A(n4043), .ZN(U3274) );
  NAND3_X1 U4719 ( .A1(n2691), .A2(n2690), .A3(n4671), .ZN(n4044) );
  NAND2_X1 U4720 ( .A1(n4045), .A2(n4044), .ZN(n4049) );
  AOI22_X1 U4721 ( .A1(n4046), .A2(n4675), .B1(n4055), .B2(n4674), .ZN(n4047)
         );
  OAI21_X1 U4722 ( .B1(n4706), .B2(n4678), .A(n4047), .ZN(n4048) );
  AOI21_X1 U4723 ( .B1(n4049), .B2(n4702), .A(n4048), .ZN(n4054) );
  NAND2_X1 U4724 ( .A1(n4051), .A2(n2154), .ZN(n4052) );
  NAND2_X1 U4725 ( .A1(n4050), .A2(n4052), .ZN(n4766) );
  NAND2_X1 U4726 ( .A1(n4766), .A2(n4703), .ZN(n4053) );
  AND2_X1 U4727 ( .A1(n4054), .A2(n4053), .ZN(n4763) );
  MUX2_X1 U4728 ( .A(n4763), .B(n4259), .S(n4700), .Z(n4058) );
  AOI22_X1 U4729 ( .A1(n4766), .A2(n4701), .B1(REG3_REG_2__SCAN_IN), .B2(n4688), .ZN(n4057) );
  NAND2_X1 U4730 ( .A1(n4692), .A2(n4055), .ZN(n4761) );
  NAND3_X1 U4731 ( .A1(n4696), .A2(n4762), .A3(n4761), .ZN(n4056) );
  NAND3_X1 U4732 ( .A1(n4058), .A2(n4057), .A3(n4056), .ZN(U3288) );
  NAND2_X1 U4733 ( .A1(n4066), .A2(n4065), .ZN(n4064) );
  XNOR2_X1 U4734 ( .A(n4064), .B(n4059), .ZN(n4520) );
  INV_X1 U4735 ( .A(n4520), .ZN(n4132) );
  AND2_X1 U4736 ( .A1(n4061), .A2(n4060), .ZN(n4067) );
  AOI21_X1 U4737 ( .B1(n4062), .B2(n4674), .A(n4067), .ZN(n4522) );
  MUX2_X1 U4738 ( .A(n2815), .B(n4522), .S(n4828), .Z(n4063) );
  OAI21_X1 U4739 ( .B1(n4132), .B2(n4130), .A(n4063), .ZN(U3549) );
  OAI21_X1 U4740 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4523) );
  AOI21_X1 U4741 ( .B1(n4068), .B2(n4674), .A(n4067), .ZN(n4526) );
  MUX2_X1 U4742 ( .A(n3286), .B(n4526), .S(n4828), .Z(n4069) );
  OAI21_X1 U4743 ( .B1(n4523), .B2(n4130), .A(n4069), .ZN(U3548) );
  MUX2_X1 U4744 ( .A(REG1_REG_29__SCAN_IN), .B(n4134), .S(n4828), .Z(U3547) );
  AOI21_X1 U4745 ( .B1(n4811), .B2(n4074), .A(n4073), .ZN(n4075) );
  OAI21_X1 U4746 ( .B1(n4076), .B2(n4778), .A(n4075), .ZN(n4135) );
  MUX2_X1 U4747 ( .A(REG1_REG_27__SCAN_IN), .B(n4135), .S(n4828), .Z(U3545) );
  OAI21_X1 U4748 ( .B1(n4798), .B2(n4078), .A(n4077), .ZN(n4079) );
  AOI21_X1 U4749 ( .B1(n4080), .B2(n4797), .A(n4079), .ZN(n4136) );
  INV_X1 U4750 ( .A(n4136), .ZN(n4081) );
  MUX2_X1 U4751 ( .A(REG1_REG_26__SCAN_IN), .B(n4081), .S(n4828), .Z(U3544) );
  AOI21_X1 U4752 ( .B1(n4083), .B2(n4797), .A(n4082), .ZN(n4436) );
  MUX2_X1 U4753 ( .A(n4366), .B(n4436), .S(n4828), .Z(n4084) );
  OAI21_X1 U4754 ( .B1(n4130), .B2(n4439), .A(n4084), .ZN(U3543) );
  AOI21_X1 U4755 ( .B1(n4086), .B2(n4797), .A(n4085), .ZN(n4440) );
  MUX2_X1 U4756 ( .A(n4217), .B(n4440), .S(n4828), .Z(n4087) );
  OAI21_X1 U4757 ( .B1(n4130), .B2(n4443), .A(n4087), .ZN(U3542) );
  AOI21_X1 U4758 ( .B1(n4089), .B2(n4797), .A(n4088), .ZN(n4444) );
  MUX2_X1 U4759 ( .A(n4418), .B(n4444), .S(n4828), .Z(n4090) );
  OAI21_X1 U4760 ( .B1(n4130), .B2(n4447), .A(n4090), .ZN(U3541) );
  NAND3_X1 U4761 ( .A1(n4092), .A2(n4811), .A3(n4091), .ZN(n4093) );
  OAI211_X1 U4762 ( .C1(n4095), .C2(n4778), .A(n4094), .B(n4093), .ZN(n4448)
         );
  MUX2_X1 U4763 ( .A(REG1_REG_22__SCAN_IN), .B(n4448), .S(n4828), .Z(U3540) );
  AOI21_X1 U4764 ( .B1(n4097), .B2(n4797), .A(n4096), .ZN(n4449) );
  MUX2_X1 U4765 ( .A(n4280), .B(n4449), .S(n4828), .Z(n4098) );
  OAI21_X1 U4766 ( .B1(n4130), .B2(n4452), .A(n4098), .ZN(U3539) );
  AOI21_X1 U4767 ( .B1(n4100), .B2(n4797), .A(n4099), .ZN(n4453) );
  MUX2_X1 U4768 ( .A(n4289), .B(n4453), .S(n4828), .Z(n4101) );
  OAI21_X1 U4769 ( .B1(n4130), .B2(n4456), .A(n4101), .ZN(U3538) );
  AOI21_X1 U4770 ( .B1(n4797), .B2(n4103), .A(n4102), .ZN(n4457) );
  MUX2_X1 U4771 ( .A(n4104), .B(n4457), .S(n4828), .Z(n4105) );
  OAI21_X1 U4772 ( .B1(n4130), .B2(n4460), .A(n4105), .ZN(U3537) );
  OAI211_X1 U4773 ( .C1(n4108), .C2(n4778), .A(n4107), .B(n4106), .ZN(n4461)
         );
  MUX2_X1 U4774 ( .A(REG1_REG_18__SCAN_IN), .B(n4461), .S(n4828), .Z(U3536) );
  AOI21_X1 U4775 ( .B1(n4110), .B2(n4797), .A(n4109), .ZN(n4462) );
  MUX2_X1 U4776 ( .A(n4274), .B(n4462), .S(n4828), .Z(n4111) );
  OAI21_X1 U4777 ( .B1(n4130), .B2(n4465), .A(n4111), .ZN(U3535) );
  NAND2_X1 U4778 ( .A1(n4112), .A2(n4797), .ZN(n4113) );
  AND2_X1 U4779 ( .A1(n4114), .A2(n4113), .ZN(n4467) );
  MUX2_X1 U4780 ( .A(n4467), .B(n4115), .S(n4826), .Z(n4116) );
  OAI21_X1 U4781 ( .B1(n4130), .B2(n4469), .A(n4116), .ZN(U3534) );
  AOI21_X1 U4782 ( .B1(n4797), .B2(n4118), .A(n4117), .ZN(n4470) );
  MUX2_X1 U4783 ( .A(n4119), .B(n4470), .S(n4828), .Z(n4120) );
  OAI21_X1 U4784 ( .B1(n4130), .B2(n4473), .A(n4120), .ZN(U3533) );
  NAND3_X1 U4785 ( .A1(n4122), .A2(n4811), .A3(n4121), .ZN(n4123) );
  OAI211_X1 U4786 ( .C1(n4125), .C2(n4805), .A(n4124), .B(n4123), .ZN(n4474)
         );
  MUX2_X1 U4787 ( .A(REG1_REG_14__SCAN_IN), .B(n4474), .S(n4828), .Z(U3532) );
  INV_X1 U4788 ( .A(n4126), .ZN(n4128) );
  AOI21_X1 U4789 ( .B1(n4803), .B2(n4128), .A(n4127), .ZN(n4475) );
  MUX2_X1 U4790 ( .A(n4271), .B(n4475), .S(n4828), .Z(n4129) );
  OAI21_X1 U4791 ( .B1(n4130), .B2(n4479), .A(n4129), .ZN(U3531) );
  MUX2_X1 U4792 ( .A(n2818), .B(n4522), .S(n4813), .Z(n4131) );
  OAI21_X1 U4793 ( .B1(n4132), .B2(n4478), .A(n4131), .ZN(U3517) );
  MUX2_X1 U4794 ( .A(n3289), .B(n4526), .S(n4813), .Z(n4133) );
  OAI21_X1 U4795 ( .B1(n4523), .B2(n4478), .A(n4133), .ZN(U3516) );
  MUX2_X1 U4796 ( .A(REG0_REG_29__SCAN_IN), .B(n4134), .S(n4813), .Z(U3515) );
  MUX2_X1 U4797 ( .A(REG0_REG_27__SCAN_IN), .B(n4135), .S(n4813), .Z(U3513) );
  MUX2_X1 U4798 ( .A(n4137), .B(n4136), .S(n4813), .Z(n4435) );
  INV_X1 U4799 ( .A(keyinput118), .ZN(n4138) );
  NOR4_X1 U4800 ( .A1(keyinput97), .A2(keyinput88), .A3(keyinput2), .A4(n4138), 
        .ZN(n4143) );
  NOR4_X1 U4801 ( .A1(keyinput53), .A2(keyinput96), .A3(keyinput69), .A4(
        keyinput29), .ZN(n4142) );
  INV_X1 U4802 ( .A(keyinput14), .ZN(n4354) );
  NOR4_X1 U4803 ( .A1(keyinput59), .A2(keyinput33), .A3(keyinput22), .A4(n4354), .ZN(n4141) );
  NAND2_X1 U4804 ( .A1(keyinput61), .A2(keyinput109), .ZN(n4139) );
  NOR3_X1 U4805 ( .A1(keyinput115), .A2(keyinput125), .A3(n4139), .ZN(n4140)
         );
  NAND4_X1 U4806 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4182)
         );
  INV_X1 U4807 ( .A(keyinput5), .ZN(n4145) );
  NAND4_X1 U4808 ( .A1(keyinput107), .A2(keyinput62), .A3(keyinput108), .A4(
        keyinput121), .ZN(n4144) );
  NOR3_X1 U4809 ( .A1(keyinput7), .A2(n4145), .A3(n4144), .ZN(n4148) );
  INV_X1 U4810 ( .A(keyinput13), .ZN(n4390) );
  INV_X1 U4811 ( .A(keyinput30), .ZN(n4388) );
  INV_X1 U4812 ( .A(keyinput12), .ZN(n4387) );
  INV_X1 U4813 ( .A(keyinput93), .ZN(n4397) );
  NOR4_X1 U4814 ( .A1(n4390), .A2(n4388), .A3(n4387), .A4(n4397), .ZN(n4147)
         );
  INV_X1 U4815 ( .A(keyinput40), .ZN(n4393) );
  NOR4_X1 U4816 ( .A1(keyinput68), .A2(keyinput78), .A3(keyinput80), .A4(n4393), .ZN(n4146) );
  NAND4_X1 U4817 ( .A1(keyinput16), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(
        n4181) );
  NAND2_X1 U4818 ( .A1(keyinput122), .A2(keyinput75), .ZN(n4149) );
  NOR3_X1 U4819 ( .A1(keyinput126), .A2(keyinput119), .A3(n4149), .ZN(n4165)
         );
  INV_X1 U4820 ( .A(keyinput67), .ZN(n4150) );
  NOR4_X1 U4821 ( .A1(keyinput70), .A2(keyinput71), .A3(keyinput79), .A4(n4150), .ZN(n4164) );
  NAND2_X1 U4822 ( .A1(keyinput19), .A2(keyinput102), .ZN(n4151) );
  NOR3_X1 U4823 ( .A1(keyinput123), .A2(keyinput18), .A3(n4151), .ZN(n4152) );
  NAND3_X1 U4824 ( .A1(keyinput31), .A2(keyinput26), .A3(n4152), .ZN(n4153) );
  NOR3_X1 U4825 ( .A1(keyinput111), .A2(keyinput23), .A3(n4153), .ZN(n4163) );
  INV_X1 U4826 ( .A(keyinput63), .ZN(n4154) );
  NAND4_X1 U4827 ( .A1(keyinput50), .A2(keyinput55), .A3(keyinput51), .A4(
        n4154), .ZN(n4161) );
  NOR2_X1 U4828 ( .A1(keyinput6), .A2(keyinput54), .ZN(n4155) );
  NAND3_X1 U4829 ( .A1(keyinput27), .A2(keyinput10), .A3(n4155), .ZN(n4160) );
  NOR2_X1 U4830 ( .A1(keyinput46), .A2(keyinput42), .ZN(n4156) );
  NAND3_X1 U4831 ( .A1(keyinput35), .A2(keyinput47), .A3(n4156), .ZN(n4159) );
  INV_X1 U4832 ( .A(keyinput34), .ZN(n4157) );
  NAND4_X1 U4833 ( .A1(keyinput38), .A2(keyinput58), .A3(keyinput39), .A4(
        n4157), .ZN(n4158) );
  NOR4_X1 U4834 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4162)
         );
  NAND4_X1 U4835 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4180)
         );
  NOR2_X1 U4836 ( .A1(keyinput1), .A2(keyinput25), .ZN(n4166) );
  NAND3_X1 U4837 ( .A1(keyinput37), .A2(keyinput9), .A3(n4166), .ZN(n4167) );
  NOR3_X1 U4838 ( .A1(keyinput57), .A2(keyinput49), .A3(n4167), .ZN(n4178) );
  NAND2_X1 U4839 ( .A1(keyinput20), .A2(keyinput0), .ZN(n4168) );
  NOR3_X1 U4840 ( .A1(keyinput44), .A2(keyinput4), .A3(n4168), .ZN(n4169) );
  NAND3_X1 U4841 ( .A1(keyinput120), .A2(keyinput76), .A3(n4169), .ZN(n4176)
         );
  AND4_X1 U4842 ( .A1(keyinput117), .A2(keyinput101), .A3(keyinput89), .A4(
        keyinput85), .ZN(n4174) );
  INV_X1 U4843 ( .A(keyinput81), .ZN(n4170) );
  NOR4_X1 U4844 ( .A1(keyinput43), .A2(keyinput113), .A3(keyinput73), .A4(
        n4170), .ZN(n4173) );
  NOR4_X1 U4845 ( .A1(keyinput36), .A2(keyinput32), .A3(keyinput28), .A4(
        keyinput24), .ZN(n4172) );
  NOR4_X1 U4846 ( .A1(keyinput92), .A2(keyinput72), .A3(keyinput64), .A4(
        keyinput124), .ZN(n4171) );
  NAND4_X1 U4847 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4175)
         );
  NOR4_X1 U4848 ( .A1(keyinput8), .A2(keyinput56), .A3(n4176), .A4(n4175), 
        .ZN(n4177) );
  NAND4_X1 U4849 ( .A1(keyinput77), .A2(keyinput65), .A3(n4178), .A4(n4177), 
        .ZN(n4179) );
  NOR4_X1 U4850 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4199)
         );
  NAND2_X1 U4851 ( .A1(keyinput95), .A2(keyinput17), .ZN(n4183) );
  NOR3_X1 U4852 ( .A1(keyinput86), .A2(keyinput90), .A3(n4183), .ZN(n4184) );
  NAND3_X1 U4853 ( .A1(keyinput3), .A2(keyinput84), .A3(n4184), .ZN(n4193) );
  NAND2_X1 U4854 ( .A1(keyinput98), .A2(keyinput74), .ZN(n4185) );
  NOR3_X1 U4855 ( .A1(keyinput106), .A2(keyinput114), .A3(n4185), .ZN(n4191)
         );
  INV_X1 U4856 ( .A(keyinput83), .ZN(n4186) );
  NOR4_X1 U4857 ( .A1(keyinput104), .A2(keyinput60), .A3(keyinput110), .A4(
        n4186), .ZN(n4190) );
  NAND2_X1 U4858 ( .A1(keyinput15), .A2(keyinput21), .ZN(n4187) );
  NOR3_X1 U4859 ( .A1(keyinput103), .A2(keyinput91), .A3(n4187), .ZN(n4189) );
  INV_X1 U4860 ( .A(keyinput45), .ZN(n4255) );
  NOR4_X1 U4861 ( .A1(keyinput52), .A2(keyinput82), .A3(keyinput116), .A4(
        n4255), .ZN(n4188) );
  NAND4_X1 U4862 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4192)
         );
  NOR4_X1 U4863 ( .A1(keyinput87), .A2(keyinput94), .A3(n4193), .A4(n4192), 
        .ZN(n4198) );
  NAND3_X1 U4864 ( .A1(keyinput11), .A2(keyinput112), .A3(keyinput99), .ZN(
        n4194) );
  NOR2_X1 U4865 ( .A1(keyinput100), .A2(n4194), .ZN(n4197) );
  NAND2_X1 U4866 ( .A1(keyinput105), .A2(keyinput66), .ZN(n4195) );
  NOR3_X1 U4867 ( .A1(keyinput41), .A2(keyinput127), .A3(n4195), .ZN(n4196) );
  NAND4_X1 U4868 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4200)
         );
  INV_X1 U4869 ( .A(DATAI_29_), .ZN(n4402) );
  AOI21_X1 U4870 ( .B1(n4200), .B2(keyinput48), .A(n4402), .ZN(n4433) );
  INV_X1 U4871 ( .A(D_REG_3__SCAN_IN), .ZN(n4727) );
  AOI22_X1 U4872 ( .A1(n4202), .A2(keyinput19), .B1(n4727), .B2(keyinput31), 
        .ZN(n4201) );
  OAI221_X1 U4873 ( .B1(n4202), .B2(keyinput19), .C1(n4727), .C2(keyinput31), 
        .A(n4201), .ZN(n4212) );
  INV_X1 U4874 ( .A(keyinput2), .ZN(n4204) );
  AOI22_X1 U4875 ( .A1(n4205), .A2(keyinput88), .B1(ADDR_REG_0__SCAN_IN), .B2(
        n4204), .ZN(n4203) );
  OAI221_X1 U4876 ( .B1(n4205), .B2(keyinput88), .C1(n4204), .C2(
        ADDR_REG_0__SCAN_IN), .A(n4203), .ZN(n4211) );
  INV_X1 U4877 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4878 ( .A1(n3826), .A2(keyinput29), .B1(keyinput97), .B2(n4207), 
        .ZN(n4206) );
  OAI221_X1 U4879 ( .B1(n3826), .B2(keyinput29), .C1(n4207), .C2(keyinput97), 
        .A(n4206), .ZN(n4210) );
  AOI22_X1 U4880 ( .A1(n4476), .A2(keyinput25), .B1(n2874), .B2(keyinput1), 
        .ZN(n4208) );
  OAI221_X1 U4881 ( .B1(n4476), .B2(keyinput25), .C1(n2874), .C2(keyinput1), 
        .A(n4208), .ZN(n4209) );
  OR4_X1 U4882 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4344) );
  INV_X1 U4883 ( .A(D_REG_20__SCAN_IN), .ZN(n4721) );
  INV_X1 U4884 ( .A(DATAI_7_), .ZN(n4747) );
  AOI22_X1 U4885 ( .A1(n4721), .A2(keyinput76), .B1(keyinput4), .B2(n4747), 
        .ZN(n4213) );
  OAI221_X1 U4886 ( .B1(n4721), .B2(keyinput76), .C1(n4747), .C2(keyinput4), 
        .A(n4213), .ZN(n4225) );
  INV_X1 U4887 ( .A(D_REG_30__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U4888 ( .A1(n4717), .A2(keyinput49), .B1(keyinput37), .B2(n4215), 
        .ZN(n4214) );
  OAI221_X1 U4889 ( .B1(n4717), .B2(keyinput49), .C1(n4215), .C2(keyinput37), 
        .A(n4214), .ZN(n4224) );
  INV_X1 U4890 ( .A(DATAI_0_), .ZN(n4218) );
  AOI22_X1 U4891 ( .A1(n4218), .A2(keyinput65), .B1(n4217), .B2(keyinput57), 
        .ZN(n4216) );
  OAI221_X1 U4892 ( .B1(n4218), .B2(keyinput65), .C1(n4217), .C2(keyinput57), 
        .A(n4216), .ZN(n4223) );
  AOI22_X1 U4893 ( .A1(n4221), .A2(keyinput38), .B1(n4220), .B2(keyinput39), 
        .ZN(n4219) );
  OAI221_X1 U4894 ( .B1(n4221), .B2(keyinput38), .C1(n4220), .C2(keyinput39), 
        .A(n4219), .ZN(n4222) );
  NOR4_X1 U4895 ( .A1(n4225), .A2(n4224), .A3(n4223), .A4(n4222), .ZN(n4251)
         );
  AOI22_X1 U4896 ( .A1(n4227), .A2(keyinput42), .B1(keyinput43), .B2(n2530), 
        .ZN(n4226) );
  OAI221_X1 U4897 ( .B1(n4227), .B2(keyinput42), .C1(n2530), .C2(keyinput43), 
        .A(n4226), .ZN(n4234) );
  AOI22_X1 U4898 ( .A1(n4230), .A2(keyinput102), .B1(n4229), .B2(keyinput111), 
        .ZN(n4228) );
  OAI221_X1 U4899 ( .B1(n4230), .B2(keyinput102), .C1(n4229), .C2(keyinput111), 
        .A(n4228), .ZN(n4233) );
  XNOR2_X1 U4900 ( .A(keyinput9), .B(n4137), .ZN(n4232) );
  XNOR2_X1 U4901 ( .A(keyinput26), .B(n2520), .ZN(n4231) );
  NOR4_X1 U4902 ( .A1(n4234), .A2(n4233), .A3(n4232), .A4(n4231), .ZN(n4250)
         );
  AOI22_X1 U4903 ( .A1(n2494), .A2(keyinput63), .B1(keyinput58), .B2(n2447), 
        .ZN(n4235) );
  OAI221_X1 U4904 ( .B1(n2494), .B2(keyinput63), .C1(n2447), .C2(keyinput58), 
        .A(n4235), .ZN(n4238) );
  INV_X1 U4905 ( .A(DATAI_15_), .ZN(n4734) );
  AOI22_X1 U4906 ( .A1(n4734), .A2(keyinput6), .B1(keyinput10), .B2(n2460), 
        .ZN(n4236) );
  OAI221_X1 U4907 ( .B1(n4734), .B2(keyinput6), .C1(n2460), .C2(keyinput10), 
        .A(n4236), .ZN(n4237) );
  NOR2_X1 U4908 ( .A1(n4238), .A2(n4237), .ZN(n4249) );
  INV_X1 U4909 ( .A(D_REG_19__SCAN_IN), .ZN(n4722) );
  INV_X1 U4910 ( .A(D_REG_16__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U4911 ( .A1(n4722), .A2(keyinput50), .B1(keyinput51), .B2(n4723), 
        .ZN(n4239) );
  OAI221_X1 U4912 ( .B1(n4722), .B2(keyinput50), .C1(n4723), .C2(keyinput51), 
        .A(n4239), .ZN(n4247) );
  INV_X1 U4913 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4242) );
  INV_X1 U4914 ( .A(B_REG_SCAN_IN), .ZN(n4241) );
  AOI22_X1 U4915 ( .A1(n4242), .A2(keyinput96), .B1(n4241), .B2(keyinput69), 
        .ZN(n4240) );
  OAI221_X1 U4916 ( .B1(n4242), .B2(keyinput96), .C1(n4241), .C2(keyinput69), 
        .A(n4240), .ZN(n4246) );
  INV_X1 U4917 ( .A(DATAI_23_), .ZN(n4731) );
  AOI22_X1 U4918 ( .A1(n4731), .A2(keyinput34), .B1(n4244), .B2(keyinput35), 
        .ZN(n4243) );
  OAI221_X1 U4919 ( .B1(n4731), .B2(keyinput34), .C1(n4244), .C2(keyinput35), 
        .A(n4243), .ZN(n4245) );
  NOR3_X1 U4920 ( .A1(n4247), .A2(n4246), .A3(n4245), .ZN(n4248) );
  NAND4_X1 U4921 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4343)
         );
  AOI22_X1 U4922 ( .A1(n2452), .A2(keyinput110), .B1(keyinput74), .B2(n2775), 
        .ZN(n4252) );
  OAI221_X1 U4923 ( .B1(n2452), .B2(keyinput110), .C1(n2775), .C2(keyinput74), 
        .A(n4252), .ZN(n4263) );
  AOI22_X1 U4924 ( .A1(n3740), .A2(keyinput60), .B1(keyinput83), .B2(n2470), 
        .ZN(n4253) );
  OAI221_X1 U4925 ( .B1(n3740), .B2(keyinput60), .C1(n2470), .C2(keyinput83), 
        .A(n4253), .ZN(n4262) );
  INV_X1 U4926 ( .A(keyinput98), .ZN(n4256) );
  AOI22_X1 U4927 ( .A1(n4256), .A2(DATAO_REG_17__SCAN_IN), .B1(
        DATAO_REG_20__SCAN_IN), .B2(n4255), .ZN(n4254) );
  OAI221_X1 U4928 ( .B1(n4256), .B2(DATAO_REG_17__SCAN_IN), .C1(n4255), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4254), .ZN(n4261) );
  AOI22_X1 U4929 ( .A1(n4259), .A2(keyinput114), .B1(n4258), .B2(keyinput106), 
        .ZN(n4257) );
  OAI221_X1 U4930 ( .B1(n4259), .B2(keyinput114), .C1(n4258), .C2(keyinput106), 
        .A(n4257), .ZN(n4260) );
  NOR4_X1 U4931 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4312)
         );
  INV_X1 U4932 ( .A(keyinput11), .ZN(n4266) );
  INV_X1 U4933 ( .A(keyinput66), .ZN(n4265) );
  AOI22_X1 U4934 ( .A1(n4266), .A2(ADDR_REG_15__SCAN_IN), .B1(
        ADDR_REG_16__SCAN_IN), .B2(n4265), .ZN(n4264) );
  OAI221_X1 U4935 ( .B1(n4266), .B2(ADDR_REG_15__SCAN_IN), .C1(n4265), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4264), .ZN(n4278) );
  INV_X1 U4936 ( .A(keyinput99), .ZN(n4269) );
  INV_X1 U4937 ( .A(keyinput100), .ZN(n4268) );
  AOI22_X1 U4938 ( .A1(n4269), .A2(ADDR_REG_12__SCAN_IN), .B1(
        ADDR_REG_13__SCAN_IN), .B2(n4268), .ZN(n4267) );
  OAI221_X1 U4939 ( .B1(n4269), .B2(ADDR_REG_12__SCAN_IN), .C1(n4268), .C2(
        ADDR_REG_13__SCAN_IN), .A(n4267), .ZN(n4277) );
  AOI22_X1 U4940 ( .A1(n4271), .A2(keyinput105), .B1(n2523), .B2(keyinput104), 
        .ZN(n4270) );
  OAI221_X1 U4941 ( .B1(n4271), .B2(keyinput105), .C1(n2523), .C2(keyinput104), 
        .A(n4270), .ZN(n4276) );
  INV_X1 U4942 ( .A(keyinput127), .ZN(n4273) );
  AOI22_X1 U4943 ( .A1(n4274), .A2(keyinput41), .B1(ADDR_REG_17__SCAN_IN), 
        .B2(n4273), .ZN(n4272) );
  OAI221_X1 U4944 ( .B1(n4274), .B2(keyinput41), .C1(n4273), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4272), .ZN(n4275) );
  NOR4_X1 U4945 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(n4311)
         );
  INV_X1 U4946 ( .A(DATAI_1_), .ZN(n4281) );
  AOI22_X1 U4947 ( .A1(n4281), .A2(keyinput86), .B1(keyinput87), .B2(n4280), 
        .ZN(n4279) );
  OAI221_X1 U4948 ( .B1(n4281), .B2(keyinput86), .C1(n4280), .C2(keyinput87), 
        .A(n4279), .ZN(n4293) );
  INV_X1 U4949 ( .A(keyinput84), .ZN(n4284) );
  INV_X1 U4950 ( .A(keyinput17), .ZN(n4283) );
  AOI22_X1 U4951 ( .A1(n4284), .A2(DATAO_REG_31__SCAN_IN), .B1(
        REG1_REG_31__SCAN_IN), .B2(n4283), .ZN(n4282) );
  OAI221_X1 U4952 ( .B1(n4284), .B2(DATAO_REG_31__SCAN_IN), .C1(n4283), .C2(
        REG1_REG_31__SCAN_IN), .A(n4282), .ZN(n4292) );
  AOI22_X1 U4953 ( .A1(n4287), .A2(keyinput90), .B1(n4286), .B2(keyinput70), 
        .ZN(n4285) );
  OAI221_X1 U4954 ( .B1(n4287), .B2(keyinput90), .C1(n4286), .C2(keyinput70), 
        .A(n4285), .ZN(n4291) );
  INV_X1 U4955 ( .A(DATAI_5_), .ZN(n4750) );
  AOI22_X1 U4956 ( .A1(n4750), .A2(keyinput94), .B1(n4289), .B2(keyinput95), 
        .ZN(n4288) );
  OAI221_X1 U4957 ( .B1(n4750), .B2(keyinput94), .C1(n4289), .C2(keyinput95), 
        .A(n4288), .ZN(n4290) );
  NOR4_X1 U4958 ( .A1(n4293), .A2(n4292), .A3(n4291), .A4(n4290), .ZN(n4310)
         );
  INV_X1 U4959 ( .A(keyinput116), .ZN(n4295) );
  AOI22_X1 U4960 ( .A1(n4296), .A2(keyinput21), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4295), .ZN(n4294) );
  OAI221_X1 U4961 ( .B1(n4296), .B2(keyinput21), .C1(n4295), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4294), .ZN(n4308) );
  INV_X1 U4962 ( .A(keyinput82), .ZN(n4299) );
  INV_X1 U4963 ( .A(keyinput52), .ZN(n4298) );
  AOI22_X1 U4964 ( .A1(n4299), .A2(DATAO_REG_23__SCAN_IN), .B1(
        DATAO_REG_24__SCAN_IN), .B2(n4298), .ZN(n4297) );
  OAI221_X1 U4965 ( .B1(n4299), .B2(DATAO_REG_23__SCAN_IN), .C1(n4298), .C2(
        DATAO_REG_24__SCAN_IN), .A(n4297), .ZN(n4307) );
  AOI22_X1 U4966 ( .A1(n4301), .A2(keyinput15), .B1(keyinput3), .B2(n3289), 
        .ZN(n4300) );
  OAI221_X1 U4967 ( .B1(n4301), .B2(keyinput15), .C1(n3289), .C2(keyinput3), 
        .A(n4300), .ZN(n4306) );
  AOI22_X1 U4968 ( .A1(n4304), .A2(keyinput91), .B1(n4303), .B2(keyinput103), 
        .ZN(n4302) );
  OAI221_X1 U4969 ( .B1(n4304), .B2(keyinput91), .C1(n4303), .C2(keyinput103), 
        .A(n4302), .ZN(n4305) );
  NOR4_X1 U4970 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), .ZN(n4309)
         );
  NAND4_X1 U4971 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4342)
         );
  XOR2_X1 U4972 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput56), .Z(n4317) );
  XOR2_X1 U4973 ( .A(IR_REG_0__SCAN_IN), .B(keyinput115), .Z(n4316) );
  XOR2_X1 U4974 ( .A(IR_REG_1__SCAN_IN), .B(keyinput92), .Z(n4315) );
  XNOR2_X1 U4975 ( .A(n4313), .B(keyinput16), .ZN(n4314) );
  NOR4_X1 U4976 ( .A1(n4317), .A2(n4316), .A3(n4315), .A4(n4314), .ZN(n4340)
         );
  XNOR2_X1 U4977 ( .A(n4318), .B(keyinput0), .ZN(n4325) );
  XNOR2_X1 U4978 ( .A(n4319), .B(keyinput44), .ZN(n4324) );
  XNOR2_X1 U4979 ( .A(n4320), .B(keyinput27), .ZN(n4323) );
  XNOR2_X1 U4980 ( .A(n4321), .B(keyinput20), .ZN(n4322) );
  NOR4_X1 U4981 ( .A1(n4325), .A2(n4324), .A3(n4323), .A4(n4322), .ZN(n4339)
         );
  XNOR2_X1 U4982 ( .A(n4326), .B(keyinput47), .ZN(n4332) );
  XNOR2_X1 U4983 ( .A(n4327), .B(keyinput23), .ZN(n4331) );
  XNOR2_X1 U4984 ( .A(n4328), .B(keyinput54), .ZN(n4330) );
  XNOR2_X1 U4985 ( .A(n4441), .B(keyinput18), .ZN(n4329) );
  NOR4_X1 U4986 ( .A1(n4332), .A2(n4331), .A3(n4330), .A4(n4329), .ZN(n4338)
         );
  XOR2_X1 U4987 ( .A(REG2_REG_24__SCAN_IN), .B(keyinput55), .Z(n4336) );
  XOR2_X1 U4988 ( .A(REG1_REG_16__SCAN_IN), .B(keyinput120), .Z(n4335) );
  XNOR2_X1 U4989 ( .A(keyinput118), .B(n2800), .ZN(n4334) );
  XNOR2_X1 U4990 ( .A(keyinput46), .B(n2404), .ZN(n4333) );
  NOR4_X1 U4991 ( .A1(n4336), .A2(n4335), .A3(n4334), .A4(n4333), .ZN(n4337)
         );
  NAND4_X1 U4992 ( .A1(n4340), .A2(n4339), .A3(n4338), .A4(n4337), .ZN(n4341)
         );
  NOR4_X1 U4993 ( .A1(n4344), .A2(n4343), .A3(n4342), .A4(n4341), .ZN(n4376)
         );
  INV_X1 U4994 ( .A(keyinput61), .ZN(n4346) );
  AOI22_X1 U4995 ( .A1(n2461), .A2(keyinput59), .B1(ADDR_REG_6__SCAN_IN), .B2(
        n4346), .ZN(n4345) );
  OAI221_X1 U4996 ( .B1(n2461), .B2(keyinput59), .C1(n4346), .C2(
        ADDR_REG_6__SCAN_IN), .A(n4345), .ZN(n4359) );
  INV_X1 U4997 ( .A(keyinput109), .ZN(n4349) );
  INV_X1 U4998 ( .A(keyinput125), .ZN(n4348) );
  AOI22_X1 U4999 ( .A1(n4349), .A2(ADDR_REG_4__SCAN_IN), .B1(
        ADDR_REG_5__SCAN_IN), .B2(n4348), .ZN(n4347) );
  OAI221_X1 U5000 ( .B1(n4349), .B2(ADDR_REG_4__SCAN_IN), .C1(n4348), .C2(
        ADDR_REG_5__SCAN_IN), .A(n4347), .ZN(n4358) );
  INV_X1 U5001 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4352) );
  INV_X1 U5002 ( .A(keyinput22), .ZN(n4351) );
  AOI22_X1 U5003 ( .A1(n4352), .A2(keyinput112), .B1(ADDR_REG_11__SCAN_IN), 
        .B2(n4351), .ZN(n4350) );
  OAI221_X1 U5004 ( .B1(n4352), .B2(keyinput112), .C1(n4351), .C2(
        ADDR_REG_11__SCAN_IN), .A(n4350), .ZN(n4357) );
  INV_X1 U5005 ( .A(keyinput33), .ZN(n4355) );
  AOI22_X1 U5006 ( .A1(n4355), .A2(ADDR_REG_7__SCAN_IN), .B1(
        ADDR_REG_10__SCAN_IN), .B2(n4354), .ZN(n4353) );
  OAI221_X1 U5007 ( .B1(n4355), .B2(ADDR_REG_7__SCAN_IN), .C1(n4354), .C2(
        ADDR_REG_10__SCAN_IN), .A(n4353), .ZN(n4356) );
  NOR4_X1 U5008 ( .A1(n4359), .A2(n4358), .A3(n4357), .A4(n4356), .ZN(n4375)
         );
  AOI22_X1 U5009 ( .A1(n4362), .A2(keyinput113), .B1(keyinput117), .B2(n4361), 
        .ZN(n4360) );
  OAI221_X1 U5010 ( .B1(n4362), .B2(keyinput113), .C1(n4361), .C2(keyinput117), 
        .A(n4360), .ZN(n4373) );
  INV_X1 U5011 ( .A(keyinput89), .ZN(n4364) );
  AOI22_X1 U5012 ( .A1(n4437), .A2(keyinput101), .B1(DATAO_REG_21__SCAN_IN), 
        .B2(n4364), .ZN(n4363) );
  OAI221_X1 U5013 ( .B1(n4437), .B2(keyinput101), .C1(n4364), .C2(
        DATAO_REG_21__SCAN_IN), .A(n4363), .ZN(n4372) );
  AOI22_X1 U5014 ( .A1(n4367), .A2(keyinput85), .B1(keyinput81), .B2(n4366), 
        .ZN(n4365) );
  OAI221_X1 U5015 ( .B1(n4367), .B2(keyinput85), .C1(n4366), .C2(keyinput81), 
        .A(n4365), .ZN(n4371) );
  INV_X1 U5016 ( .A(DATAI_13_), .ZN(n4738) );
  AOI22_X1 U5017 ( .A1(n4738), .A2(keyinput73), .B1(n4369), .B2(keyinput77), 
        .ZN(n4368) );
  OAI221_X1 U5018 ( .B1(n4738), .B2(keyinput73), .C1(n4369), .C2(keyinput77), 
        .A(n4368), .ZN(n4370) );
  NOR4_X1 U5019 ( .A1(n4373), .A2(n4372), .A3(n4371), .A4(n4370), .ZN(n4374)
         );
  NAND3_X1 U5020 ( .A1(n4376), .A2(n4375), .A3(n4374), .ZN(n4432) );
  AOI22_X1 U5021 ( .A1(n4719), .A2(keyinput71), .B1(keyinput67), .B2(n4726), 
        .ZN(n4377) );
  OAI221_X1 U5022 ( .B1(n4719), .B2(keyinput71), .C1(n4726), .C2(keyinput67), 
        .A(n4377), .ZN(n4385) );
  AOI22_X1 U5023 ( .A1(n4718), .A2(keyinput79), .B1(keyinput75), .B2(n4725), 
        .ZN(n4378) );
  OAI221_X1 U5024 ( .B1(n4718), .B2(keyinput79), .C1(n4725), .C2(keyinput75), 
        .A(n4378), .ZN(n4384) );
  INV_X1 U5025 ( .A(D_REG_15__SCAN_IN), .ZN(n4724) );
  INV_X1 U5026 ( .A(DATAI_4_), .ZN(n4380) );
  AOI22_X1 U5027 ( .A1(n4724), .A2(keyinput119), .B1(keyinput126), .B2(n4380), 
        .ZN(n4379) );
  OAI221_X1 U5028 ( .B1(n4724), .B2(keyinput119), .C1(n4380), .C2(keyinput126), 
        .A(n4379), .ZN(n4383) );
  INV_X1 U5029 ( .A(D_REG_26__SCAN_IN), .ZN(n4720) );
  AOI22_X1 U5030 ( .A1(n4720), .A2(keyinput122), .B1(keyinput123), .B2(n4445), 
        .ZN(n4381) );
  OAI221_X1 U5031 ( .B1(n4720), .B2(keyinput122), .C1(n4445), .C2(keyinput123), 
        .A(n4381), .ZN(n4382) );
  NOR4_X1 U5032 ( .A1(n4385), .A2(n4384), .A3(n4383), .A4(n4382), .ZN(n4430)
         );
  AOI22_X1 U5033 ( .A1(n4388), .A2(DATAO_REG_8__SCAN_IN), .B1(
        DATAO_REG_12__SCAN_IN), .B2(n4387), .ZN(n4386) );
  OAI221_X1 U5034 ( .B1(n4388), .B2(DATAO_REG_8__SCAN_IN), .C1(n4387), .C2(
        DATAO_REG_12__SCAN_IN), .A(n4386), .ZN(n4401) );
  INV_X1 U5035 ( .A(keyinput78), .ZN(n4391) );
  AOI22_X1 U5036 ( .A1(n4391), .A2(DATAO_REG_4__SCAN_IN), .B1(
        DATAO_REG_10__SCAN_IN), .B2(n4390), .ZN(n4389) );
  OAI221_X1 U5037 ( .B1(n4391), .B2(DATAO_REG_4__SCAN_IN), .C1(n4390), .C2(
        DATAO_REG_10__SCAN_IN), .A(n4389), .ZN(n4400) );
  AOI22_X1 U5038 ( .A1(n4394), .A2(keyinput53), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n4393), .ZN(n4392) );
  OAI221_X1 U5039 ( .B1(n4394), .B2(keyinput53), .C1(n4393), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4392), .ZN(n4399) );
  INV_X1 U5040 ( .A(keyinput80), .ZN(n4396) );
  AOI22_X1 U5041 ( .A1(n4397), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n4396), .ZN(n4395) );
  OAI221_X1 U5042 ( .B1(n4397), .B2(DATAO_REG_6__SCAN_IN), .C1(n4396), .C2(
        DATAO_REG_13__SCAN_IN), .A(n4395), .ZN(n4398) );
  NOR4_X1 U5043 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .ZN(n4429)
         );
  INV_X1 U5044 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U5045 ( .A1(keyinput107), .A2(n4404), .B1(keyinput48), .B2(n4402), 
        .ZN(n4403) );
  OAI21_X1 U5046 ( .B1(n4404), .B2(keyinput107), .A(n4403), .ZN(n4414) );
  AOI22_X1 U5047 ( .A1(U3149), .A2(keyinput5), .B1(keyinput7), .B2(n4406), 
        .ZN(n4405) );
  OAI221_X1 U5048 ( .B1(U3149), .B2(keyinput5), .C1(n4406), .C2(keyinput7), 
        .A(n4405), .ZN(n4413) );
  AOI22_X1 U5049 ( .A1(n2422), .A2(keyinput121), .B1(n2398), .B2(keyinput68), 
        .ZN(n4407) );
  OAI221_X1 U5050 ( .B1(n2422), .B2(keyinput121), .C1(n2398), .C2(keyinput68), 
        .A(n4407), .ZN(n4412) );
  INV_X1 U5051 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4410) );
  INV_X1 U5052 ( .A(keyinput108), .ZN(n4409) );
  AOI22_X1 U5053 ( .A1(n4410), .A2(keyinput62), .B1(ADDR_REG_3__SCAN_IN), .B2(
        n4409), .ZN(n4408) );
  OAI221_X1 U5054 ( .B1(n4410), .B2(keyinput62), .C1(n4409), .C2(
        ADDR_REG_3__SCAN_IN), .A(n4408), .ZN(n4411) );
  NOR4_X1 U5055 ( .A1(n4414), .A2(n4413), .A3(n4412), .A4(n4411), .ZN(n4428)
         );
  AOI22_X1 U5056 ( .A1(n2437), .A2(keyinput72), .B1(keyinput64), .B2(n4450), 
        .ZN(n4415) );
  OAI221_X1 U5057 ( .B1(n2437), .B2(keyinput72), .C1(n4450), .C2(keyinput64), 
        .A(n4415), .ZN(n4426) );
  AOI22_X1 U5058 ( .A1(n4418), .A2(keyinput124), .B1(n4417), .B2(keyinput36), 
        .ZN(n4416) );
  OAI221_X1 U5059 ( .B1(n4418), .B2(keyinput124), .C1(n4417), .C2(keyinput36), 
        .A(n4416), .ZN(n4425) );
  AOI22_X1 U5060 ( .A1(n4421), .A2(keyinput32), .B1(n4420), .B2(keyinput28), 
        .ZN(n4419) );
  OAI221_X1 U5061 ( .B1(n4421), .B2(keyinput32), .C1(n4420), .C2(keyinput28), 
        .A(n4419), .ZN(n4424) );
  INV_X1 U5062 ( .A(DATAI_8_), .ZN(n4745) );
  AOI22_X1 U5063 ( .A1(n4745), .A2(keyinput24), .B1(n2493), .B2(keyinput8), 
        .ZN(n4422) );
  OAI221_X1 U5064 ( .B1(n4745), .B2(keyinput24), .C1(n2493), .C2(keyinput8), 
        .A(n4422), .ZN(n4423) );
  NOR4_X1 U5065 ( .A1(n4426), .A2(n4425), .A3(n4424), .A4(n4423), .ZN(n4427)
         );
  NAND4_X1 U5066 ( .A1(n4430), .A2(n4429), .A3(n4428), .A4(n4427), .ZN(n4431)
         );
  NOR3_X1 U5067 ( .A1(n4433), .A2(n4432), .A3(n4431), .ZN(n4434) );
  XNOR2_X1 U5068 ( .A(n4435), .B(n4434), .ZN(U3512) );
  MUX2_X1 U5069 ( .A(n4437), .B(n4436), .S(n4813), .Z(n4438) );
  OAI21_X1 U5070 ( .B1(n4439), .B2(n4478), .A(n4438), .ZN(U3511) );
  MUX2_X1 U5071 ( .A(n4441), .B(n4440), .S(n4813), .Z(n4442) );
  OAI21_X1 U5072 ( .B1(n4443), .B2(n4478), .A(n4442), .ZN(U3510) );
  MUX2_X1 U5073 ( .A(n4445), .B(n4444), .S(n4813), .Z(n4446) );
  OAI21_X1 U5074 ( .B1(n4447), .B2(n4478), .A(n4446), .ZN(U3509) );
  MUX2_X1 U5075 ( .A(REG0_REG_22__SCAN_IN), .B(n4448), .S(n4813), .Z(U3508) );
  MUX2_X1 U5076 ( .A(n4450), .B(n4449), .S(n4813), .Z(n4451) );
  OAI21_X1 U5077 ( .B1(n4452), .B2(n4478), .A(n4451), .ZN(U3507) );
  MUX2_X1 U5078 ( .A(n4454), .B(n4453), .S(n4813), .Z(n4455) );
  OAI21_X1 U5079 ( .B1(n4456), .B2(n4478), .A(n4455), .ZN(U3506) );
  MUX2_X1 U5080 ( .A(n4458), .B(n4457), .S(n4813), .Z(n4459) );
  OAI21_X1 U5081 ( .B1(n4460), .B2(n4478), .A(n4459), .ZN(U3505) );
  MUX2_X1 U5082 ( .A(REG0_REG_18__SCAN_IN), .B(n4461), .S(n4813), .Z(U3503) );
  MUX2_X1 U5083 ( .A(n4463), .B(n4462), .S(n4813), .Z(n4464) );
  OAI21_X1 U5084 ( .B1(n4465), .B2(n4478), .A(n4464), .ZN(U3501) );
  MUX2_X1 U5085 ( .A(n4467), .B(n4466), .S(n4812), .Z(n4468) );
  OAI21_X1 U5086 ( .B1(n4469), .B2(n4478), .A(n4468), .ZN(U3499) );
  MUX2_X1 U5087 ( .A(n4471), .B(n4470), .S(n4813), .Z(n4472) );
  OAI21_X1 U5088 ( .B1(n4473), .B2(n4478), .A(n4472), .ZN(U3497) );
  MUX2_X1 U5089 ( .A(REG0_REG_14__SCAN_IN), .B(n4474), .S(n4813), .Z(U3495) );
  MUX2_X1 U5090 ( .A(n4476), .B(n4475), .S(n4813), .Z(n4477) );
  OAI21_X1 U5091 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(U3493) );
  MUX2_X1 U5092 ( .A(n2384), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5093 ( .A(DATAI_29_), .B(n2193), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5094 ( .A(DATAI_28_), .B(n4480), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5095 ( .A(n4481), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5096 ( .A(DATAI_22_), .B(n4482), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5097 ( .A(DATAI_21_), .B(n2720), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5098 ( .A(DATAI_20_), .B(n4483), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5099 ( .A(n4484), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5100 ( .A(DATAI_16_), .B(n4485), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5101 ( .A(DATAI_9_), .B(n4486), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5102 ( .A(DATAI_4_), .B(n4487), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5103 ( .A(n4488), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5104 ( .A(n4489), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5105 ( .A(n4490), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5106 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  OAI22_X1 U5107 ( .A1(n4492), .A2(n4504), .B1(n4503), .B2(n4491), .ZN(n4493)
         );
  AOI211_X1 U5108 ( .C1(n4495), .C2(n2153), .A(n4494), .B(n4493), .ZN(n4500)
         );
  AOI21_X1 U5109 ( .B1(n4512), .B2(n4509), .A(n4511), .ZN(n4496) );
  XOR2_X1 U5110 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND2_X1 U5111 ( .A1(n4498), .A2(n4514), .ZN(n4499) );
  OAI211_X1 U5112 ( .C1(n4519), .C2(n4501), .A(n4500), .B(n4499), .ZN(U3223)
         );
  AND2_X1 U5113 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4633) );
  OAI22_X1 U5114 ( .A1(n4505), .A2(n4504), .B1(n4503), .B2(n4502), .ZN(n4506)
         );
  AOI211_X1 U5115 ( .C1(n4508), .C2(n2153), .A(n4633), .B(n4506), .ZN(n4517)
         );
  INV_X1 U5116 ( .A(n4509), .ZN(n4510) );
  NOR2_X1 U5117 ( .A1(n4511), .A2(n4510), .ZN(n4513) );
  XNOR2_X1 U5118 ( .A(n4513), .B(n4512), .ZN(n4515) );
  NAND2_X1 U5119 ( .A1(n4515), .A2(n4514), .ZN(n4516) );
  OAI211_X1 U5120 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4516), .ZN(U3238)
         );
  AOI22_X1 U5121 ( .A1(n4520), .A2(n4696), .B1(n4700), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4521) );
  OAI21_X1 U5122 ( .B1(n4700), .B2(n4522), .A(n4521), .ZN(U3260) );
  INV_X1 U5123 ( .A(n4523), .ZN(n4524) );
  AOI22_X1 U5124 ( .A1(n4524), .A2(n4696), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4700), .ZN(n4525) );
  OAI21_X1 U5125 ( .B1(n4700), .B2(n4526), .A(n4525), .ZN(U3261) );
  AOI211_X1 U5126 ( .C1(n4529), .C2(n4528), .A(n4527), .B(n4537), .ZN(n4530)
         );
  AOI211_X1 U5127 ( .C1(n4645), .C2(ADDR_REG_5__SCAN_IN), .A(n4531), .B(n4530), 
        .ZN(n4536) );
  OAI211_X1 U5128 ( .C1(n4534), .C2(n4533), .A(n4610), .B(n4532), .ZN(n4535)
         );
  OAI211_X1 U5129 ( .C1(n4653), .C2(n4751), .A(n4536), .B(n4535), .ZN(U3245)
         );
  AOI211_X1 U5130 ( .C1(n2461), .C2(n4539), .A(n4538), .B(n4537), .ZN(n4540)
         );
  AOI211_X1 U5131 ( .C1(n4645), .C2(ADDR_REG_6__SCAN_IN), .A(n4541), .B(n4540), 
        .ZN(n4545) );
  OAI211_X1 U5132 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4543), .A(n4610), .B(n4542), 
        .ZN(n4544) );
  OAI211_X1 U5133 ( .C1(n4653), .C2(n2304), .A(n4545), .B(n4544), .ZN(U3246)
         );
  AOI22_X1 U5134 ( .A1(n4546), .A2(n2470), .B1(REG1_REG_7__SCAN_IN), .B2(n4748), .ZN(n4548) );
  OAI21_X1 U5135 ( .B1(n4549), .B2(n4548), .A(n4646), .ZN(n4547) );
  AOI21_X1 U5136 ( .B1(n4549), .B2(n4548), .A(n4547), .ZN(n4550) );
  AOI211_X1 U5137 ( .C1(n4645), .C2(ADDR_REG_7__SCAN_IN), .A(n4551), .B(n4550), 
        .ZN(n4556) );
  OAI211_X1 U5138 ( .C1(n4554), .C2(n4553), .A(n4610), .B(n4552), .ZN(n4555)
         );
  OAI211_X1 U5139 ( .C1(n4653), .C2(n4748), .A(n4556), .B(n4555), .ZN(U3247)
         );
  OAI211_X1 U5140 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4558), .A(n4646), .B(n4557), 
        .ZN(n4562) );
  OAI211_X1 U5141 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4560), .A(n4610), .B(n4559), 
        .ZN(n4561) );
  OAI211_X1 U5142 ( .C1(n4653), .C2(n4746), .A(n4562), .B(n4561), .ZN(n4563)
         );
  AOI211_X1 U5143 ( .C1(n4645), .C2(ADDR_REG_8__SCAN_IN), .A(n4564), .B(n4563), 
        .ZN(n4565) );
  INV_X1 U5144 ( .A(n4565), .ZN(U3248) );
  OAI211_X1 U5145 ( .C1(n4568), .C2(n4567), .A(n4566), .B(n4646), .ZN(n4573)
         );
  OAI211_X1 U5146 ( .C1(n4571), .C2(n4570), .A(n4610), .B(n4569), .ZN(n4572)
         );
  OAI211_X1 U5147 ( .C1(n4653), .C2(n4574), .A(n4573), .B(n4572), .ZN(n4575)
         );
  AOI211_X1 U5148 ( .C1(n4645), .C2(ADDR_REG_9__SCAN_IN), .A(n4576), .B(n4575), 
        .ZN(n4577) );
  INV_X1 U5149 ( .A(n4577), .ZN(U3249) );
  OAI211_X1 U5150 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4579), .A(n4646), .B(n4578), .ZN(n4583) );
  OAI211_X1 U5151 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4581), .A(n4610), .B(n4580), .ZN(n4582) );
  OAI211_X1 U5152 ( .C1(n4653), .C2(n4744), .A(n4583), .B(n4582), .ZN(n4584)
         );
  AOI211_X1 U5153 ( .C1(n4645), .C2(ADDR_REG_10__SCAN_IN), .A(n4585), .B(n4584), .ZN(n4586) );
  INV_X1 U5154 ( .A(n4586), .ZN(U3250) );
  OAI211_X1 U5155 ( .C1(n4589), .C2(n4588), .A(n4646), .B(n4587), .ZN(n4594)
         );
  OAI211_X1 U5156 ( .C1(n4592), .C2(n4591), .A(n4610), .B(n4590), .ZN(n4593)
         );
  OAI211_X1 U5157 ( .C1(n4653), .C2(n4595), .A(n4594), .B(n4593), .ZN(n4596)
         );
  AOI211_X1 U5158 ( .C1(n4645), .C2(ADDR_REG_11__SCAN_IN), .A(n4597), .B(n4596), .ZN(n4598) );
  INV_X1 U5159 ( .A(n4598), .ZN(U3251) );
  OAI211_X1 U5160 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4600), .A(n4610), .B(n4599), .ZN(n4601) );
  NAND2_X1 U5161 ( .A1(n4602), .A2(n4601), .ZN(n4603) );
  AOI21_X1 U5162 ( .B1(n4645), .B2(ADDR_REG_12__SCAN_IN), .A(n4603), .ZN(n4607) );
  OAI211_X1 U5163 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4605), .A(n4646), .B(n4604), .ZN(n4606) );
  OAI211_X1 U5164 ( .C1(n4653), .C2(n2292), .A(n4607), .B(n4606), .ZN(U3252)
         );
  AOI21_X1 U5165 ( .B1(n4609), .B2(n4739), .A(n4608), .ZN(n4613) );
  OAI21_X1 U5166 ( .B1(n4613), .B2(n4612), .A(n4610), .ZN(n4611) );
  AOI21_X1 U5167 ( .B1(n4613), .B2(n4612), .A(n4611), .ZN(n4614) );
  AOI211_X1 U5168 ( .C1(n4645), .C2(ADDR_REG_13__SCAN_IN), .A(n4615), .B(n4614), .ZN(n4620) );
  OAI211_X1 U5169 ( .C1(n4618), .C2(n4617), .A(n4646), .B(n4616), .ZN(n4619)
         );
  OAI211_X1 U5170 ( .C1(n4653), .C2(n4739), .A(n4620), .B(n4619), .ZN(U3253)
         );
  AOI211_X1 U5171 ( .C1(n3271), .C2(n4622), .A(n4621), .B(n4639), .ZN(n4623)
         );
  AOI211_X1 U5172 ( .C1(n4645), .C2(ADDR_REG_14__SCAN_IN), .A(n4624), .B(n4623), .ZN(n4628) );
  OAI211_X1 U5173 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4626), .A(n4646), .B(n4625), .ZN(n4627) );
  OAI211_X1 U5174 ( .C1(n4653), .C2(n2293), .A(n4628), .B(n4627), .ZN(U3254)
         );
  AOI211_X1 U5175 ( .C1(n4631), .C2(n4630), .A(n4629), .B(n4639), .ZN(n4632)
         );
  AOI211_X1 U5176 ( .C1(ADDR_REG_15__SCAN_IN), .C2(n4645), .A(n4633), .B(n4632), .ZN(n4638) );
  OAI211_X1 U5177 ( .C1(n4636), .C2(n4635), .A(n4646), .B(n4634), .ZN(n4637)
         );
  OAI211_X1 U5178 ( .C1(n4653), .C2(n4735), .A(n4638), .B(n4637), .ZN(U3255)
         );
  AOI221_X1 U5179 ( .B1(n4642), .B2(n4641), .C1(n4640), .C2(n4641), .A(n4639), 
        .ZN(n4643) );
  AOI211_X1 U5180 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4645), .A(n4644), .B(n4643), .ZN(n4651) );
  OAI221_X1 U5181 ( .B1(n4649), .B2(n4648), .C1(n4649), .C2(n4647), .A(n4646), 
        .ZN(n4650) );
  OAI211_X1 U5182 ( .C1(n4653), .C2(n4652), .A(n4651), .B(n4650), .ZN(U3257)
         );
  XOR2_X1 U5183 ( .A(n4654), .B(n4659), .Z(n4663) );
  AOI22_X1 U5184 ( .A1(n4656), .A2(n4655), .B1(n4674), .B2(n4667), .ZN(n4657)
         );
  OAI21_X1 U5185 ( .B1(n4658), .B2(n4705), .A(n4657), .ZN(n4662) );
  XOR2_X1 U5186 ( .A(n4660), .B(n4659), .Z(n4806) );
  NOR2_X1 U5187 ( .A1(n4806), .A2(n4684), .ZN(n4661) );
  AOI211_X1 U5188 ( .C1(n4663), .C2(n4702), .A(n4662), .B(n4661), .ZN(n4807)
         );
  AOI22_X1 U5189 ( .A1(n4664), .A2(n4688), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4700), .ZN(n4670) );
  INV_X1 U5190 ( .A(n4806), .ZN(n4668) );
  AOI21_X1 U5191 ( .B1(n4667), .B2(n4666), .A(n4665), .ZN(n4810) );
  AOI22_X1 U5192 ( .A1(n4668), .A2(n4701), .B1(n4696), .B2(n4810), .ZN(n4669)
         );
  OAI211_X1 U5193 ( .C1(n4700), .C2(n4807), .A(n4670), .B(n4669), .ZN(U3279)
         );
  OAI21_X1 U5194 ( .B1(n4673), .B2(n4672), .A(n4671), .ZN(n4687) );
  AOI22_X1 U5195 ( .A1(n4676), .A2(n4675), .B1(n4674), .B2(n4690), .ZN(n4677)
         );
  OAI21_X1 U5196 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n4686) );
  OR2_X1 U5197 ( .A1(n4681), .A2(n4680), .ZN(n4682) );
  NAND2_X1 U5198 ( .A1(n4683), .A2(n4682), .ZN(n4757) );
  NOR2_X1 U5199 ( .A1(n4757), .A2(n4684), .ZN(n4685) );
  AOI211_X1 U5200 ( .C1(n4702), .C2(n4687), .A(n4686), .B(n4685), .ZN(n4755)
         );
  AOI22_X1 U5201 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4688), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4700), .ZN(n4698) );
  NAND2_X1 U5202 ( .A1(n4690), .A2(n4689), .ZN(n4691) );
  NAND2_X1 U5203 ( .A1(n4692), .A2(n4691), .ZN(n4756) );
  INV_X1 U5204 ( .A(n4756), .ZN(n4695) );
  NOR2_X1 U5205 ( .A1(n4693), .A2(n4757), .ZN(n4694) );
  AOI21_X1 U5206 ( .B1(n4696), .B2(n4695), .A(n4694), .ZN(n4697) );
  OAI211_X1 U5207 ( .C1(n4700), .C2(n4755), .A(n4698), .B(n4697), .ZN(U3289)
         );
  INV_X1 U5208 ( .A(n4699), .ZN(n4754) );
  AOI22_X1 U5209 ( .A1(n4701), .A2(n4754), .B1(REG2_REG_0__SCAN_IN), .B2(n4700), .ZN(n4715) );
  OAI21_X1 U5210 ( .B1(n4703), .B2(n4702), .A(n4754), .ZN(n4704) );
  OAI21_X1 U5211 ( .B1(n4706), .B2(n4705), .A(n4704), .ZN(n4752) );
  INV_X1 U5212 ( .A(n4707), .ZN(n4708) );
  NOR2_X1 U5213 ( .A1(n4709), .A2(n4708), .ZN(n4753) );
  INV_X1 U5214 ( .A(n4753), .ZN(n4711) );
  NOR2_X1 U5215 ( .A1(n4711), .A2(n4710), .ZN(n4713) );
  OAI21_X1 U5216 ( .B1(n4752), .B2(n4713), .A(n4712), .ZN(n4714) );
  OAI211_X1 U5217 ( .C1(n4716), .C2(n2398), .A(n4715), .B(n4714), .ZN(U3290)
         );
  AND2_X1 U5218 ( .A1(D_REG_31__SCAN_IN), .A2(n4729), .ZN(U3291) );
  NOR2_X1 U5219 ( .A1(n4728), .A2(n4717), .ZN(U3292) );
  AND2_X1 U5220 ( .A1(D_REG_29__SCAN_IN), .A2(n4729), .ZN(U3293) );
  NOR2_X1 U5221 ( .A1(n4728), .A2(n4718), .ZN(U3294) );
  NOR2_X1 U5222 ( .A1(n4728), .A2(n4719), .ZN(U3295) );
  NOR2_X1 U5223 ( .A1(n4728), .A2(n4720), .ZN(U3296) );
  AND2_X1 U5224 ( .A1(D_REG_25__SCAN_IN), .A2(n4729), .ZN(U3297) );
  AND2_X1 U5225 ( .A1(D_REG_24__SCAN_IN), .A2(n4729), .ZN(U3298) );
  AND2_X1 U5226 ( .A1(D_REG_23__SCAN_IN), .A2(n4729), .ZN(U3299) );
  AND2_X1 U5227 ( .A1(D_REG_22__SCAN_IN), .A2(n4729), .ZN(U3300) );
  AND2_X1 U5228 ( .A1(D_REG_21__SCAN_IN), .A2(n4729), .ZN(U3301) );
  NOR2_X1 U5229 ( .A1(n4728), .A2(n4721), .ZN(U3302) );
  NOR2_X1 U5230 ( .A1(n4728), .A2(n4722), .ZN(U3303) );
  AND2_X1 U5231 ( .A1(D_REG_18__SCAN_IN), .A2(n4729), .ZN(U3304) );
  AND2_X1 U5232 ( .A1(D_REG_17__SCAN_IN), .A2(n4729), .ZN(U3305) );
  NOR2_X1 U5233 ( .A1(n4728), .A2(n4723), .ZN(U3306) );
  NOR2_X1 U5234 ( .A1(n4728), .A2(n4724), .ZN(U3307) );
  AND2_X1 U5235 ( .A1(D_REG_14__SCAN_IN), .A2(n4729), .ZN(U3308) );
  AND2_X1 U5236 ( .A1(D_REG_13__SCAN_IN), .A2(n4729), .ZN(U3309) );
  AND2_X1 U5237 ( .A1(D_REG_12__SCAN_IN), .A2(n4729), .ZN(U3310) );
  AND2_X1 U5238 ( .A1(D_REG_11__SCAN_IN), .A2(n4729), .ZN(U3311) );
  NOR2_X1 U5239 ( .A1(n4728), .A2(n4725), .ZN(U3312) );
  AND2_X1 U5240 ( .A1(D_REG_9__SCAN_IN), .A2(n4729), .ZN(U3313) );
  AND2_X1 U5241 ( .A1(D_REG_8__SCAN_IN), .A2(n4729), .ZN(U3314) );
  AND2_X1 U5242 ( .A1(D_REG_7__SCAN_IN), .A2(n4729), .ZN(U3315) );
  NOR2_X1 U5243 ( .A1(n4728), .A2(n4726), .ZN(U3316) );
  AND2_X1 U5244 ( .A1(D_REG_5__SCAN_IN), .A2(n4729), .ZN(U3317) );
  AND2_X1 U5245 ( .A1(D_REG_4__SCAN_IN), .A2(n4729), .ZN(U3318) );
  NOR2_X1 U5246 ( .A1(n4728), .A2(n4727), .ZN(U3319) );
  AND2_X1 U5247 ( .A1(D_REG_2__SCAN_IN), .A2(n4729), .ZN(U3320) );
  AOI21_X1 U5248 ( .B1(U3149), .B2(n4731), .A(n4730), .ZN(U3329) );
  OAI22_X1 U5249 ( .A1(U3149), .A2(n4732), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4733) );
  INV_X1 U5250 ( .A(n4733), .ZN(U3335) );
  AOI22_X1 U5251 ( .A1(STATE_REG_SCAN_IN), .A2(n4735), .B1(n4734), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5252 ( .A1(U3149), .A2(n4736), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4737) );
  INV_X1 U5253 ( .A(n4737), .ZN(U3338) );
  AOI22_X1 U5254 ( .A1(STATE_REG_SCAN_IN), .A2(n4739), .B1(n4738), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5255 ( .A(DATAI_12_), .ZN(n4740) );
  AOI22_X1 U5256 ( .A1(STATE_REG_SCAN_IN), .A2(n2292), .B1(n4740), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5257 ( .A1(U3149), .A2(n4741), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4742) );
  INV_X1 U5258 ( .A(n4742), .ZN(U3341) );
  INV_X1 U5259 ( .A(DATAI_10_), .ZN(n4743) );
  AOI22_X1 U5260 ( .A1(STATE_REG_SCAN_IN), .A2(n4744), .B1(n4743), .B2(U3149), 
        .ZN(U3342) );
  AOI22_X1 U5261 ( .A1(STATE_REG_SCAN_IN), .A2(n4746), .B1(n4745), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5262 ( .A1(STATE_REG_SCAN_IN), .A2(n4748), .B1(n4747), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5263 ( .A(DATAI_6_), .ZN(n4749) );
  AOI22_X1 U5264 ( .A1(STATE_REG_SCAN_IN), .A2(n2304), .B1(n4749), .B2(U3149), 
        .ZN(U3346) );
  AOI22_X1 U5265 ( .A1(STATE_REG_SCAN_IN), .A2(n4751), .B1(n4750), .B2(U3149), 
        .ZN(U3347) );
  AOI211_X1 U5266 ( .C1(n4803), .C2(n4754), .A(n4753), .B(n4752), .ZN(n4814)
         );
  AOI22_X1 U5267 ( .A1(n4813), .A2(n4814), .B1(n2397), .B2(n4812), .ZN(U3467)
         );
  INV_X1 U5268 ( .A(n4755), .ZN(n4759) );
  OAI22_X1 U5269 ( .A1(n4757), .A2(n4805), .B1(n4798), .B2(n4756), .ZN(n4758)
         );
  NOR2_X1 U5270 ( .A1(n4759), .A2(n4758), .ZN(n4816) );
  INV_X1 U5271 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5272 ( .A1(n4813), .A2(n4816), .B1(n4760), .B2(n4812), .ZN(U3469)
         );
  AND3_X1 U5273 ( .A1(n4762), .A2(n4811), .A3(n4761), .ZN(n4765) );
  INV_X1 U5274 ( .A(n4763), .ZN(n4764) );
  AOI211_X1 U5275 ( .C1(n4803), .C2(n4766), .A(n4765), .B(n4764), .ZN(n4818)
         );
  AOI22_X1 U5276 ( .A1(n4813), .A2(n4818), .B1(n2404), .B2(n4812), .ZN(U3471)
         );
  NOR2_X1 U5277 ( .A1(n4767), .A2(n4805), .ZN(n4769) );
  AOI211_X1 U5278 ( .C1(n4811), .C2(n4770), .A(n4769), .B(n4768), .ZN(n4819)
         );
  AOI22_X1 U5279 ( .A1(n4813), .A2(n4819), .B1(n2424), .B2(n4812), .ZN(U3473)
         );
  NAND2_X1 U5280 ( .A1(n4771), .A2(n4803), .ZN(n4774) );
  INV_X1 U5281 ( .A(n4772), .ZN(n4773) );
  NAND2_X1 U5282 ( .A1(n4774), .A2(n4773), .ZN(n4775) );
  NOR2_X1 U5283 ( .A1(n4776), .A2(n4775), .ZN(n4820) );
  AOI22_X1 U5284 ( .A1(n4813), .A2(n4820), .B1(n2437), .B2(n4812), .ZN(U3475)
         );
  OAI22_X1 U5285 ( .A1(n4779), .A2(n4778), .B1(n4798), .B2(n4777), .ZN(n4780)
         );
  NOR2_X1 U5286 ( .A1(n4781), .A2(n4780), .ZN(n4821) );
  AOI22_X1 U5287 ( .A1(n4813), .A2(n4821), .B1(n2447), .B2(n4812), .ZN(U3477)
         );
  INV_X1 U5288 ( .A(n4782), .ZN(n4785) );
  INV_X1 U5289 ( .A(n4783), .ZN(n4784) );
  AOI211_X1 U5290 ( .C1(n4786), .C2(n4797), .A(n4785), .B(n4784), .ZN(n4822)
         );
  AOI22_X1 U5291 ( .A1(n4813), .A2(n4822), .B1(n2469), .B2(n4812), .ZN(U3481)
         );
  NOR3_X1 U5292 ( .A1(n4788), .A2(n4787), .A3(n4798), .ZN(n4790) );
  AOI211_X1 U5293 ( .C1(n4791), .C2(n4803), .A(n4790), .B(n4789), .ZN(n4823)
         );
  AOI22_X1 U5294 ( .A1(n4813), .A2(n4823), .B1(n2481), .B2(n4812), .ZN(U3483)
         );
  NOR2_X1 U5295 ( .A1(n4792), .A2(n4798), .ZN(n4795) );
  INV_X1 U5296 ( .A(n4793), .ZN(n4794) );
  AOI211_X1 U5297 ( .C1(n4797), .C2(n4796), .A(n4795), .B(n4794), .ZN(n4824)
         );
  AOI22_X1 U5298 ( .A1(n4813), .A2(n4824), .B1(n2493), .B2(n4812), .ZN(U3485)
         );
  NOR3_X1 U5299 ( .A1(n4800), .A2(n4799), .A3(n4798), .ZN(n4802) );
  AOI211_X1 U5300 ( .C1(n4804), .C2(n4803), .A(n4802), .B(n4801), .ZN(n4825)
         );
  AOI22_X1 U5301 ( .A1(n4813), .A2(n4825), .B1(n2511), .B2(n4812), .ZN(U3487)
         );
  NOR2_X1 U5302 ( .A1(n4806), .A2(n4805), .ZN(n4809) );
  INV_X1 U5303 ( .A(n4807), .ZN(n4808) );
  AOI211_X1 U5304 ( .C1(n4811), .C2(n4810), .A(n4809), .B(n4808), .ZN(n4827)
         );
  AOI22_X1 U5305 ( .A1(n4813), .A2(n4827), .B1(n2520), .B2(n4812), .ZN(U3489)
         );
  AOI22_X1 U5306 ( .A1(n4828), .A2(n4814), .B1(n2800), .B2(n4826), .ZN(U3518)
         );
  AOI22_X1 U5307 ( .A1(n4828), .A2(n4816), .B1(n4815), .B2(n4826), .ZN(U3519)
         );
  AOI22_X1 U5308 ( .A1(n4828), .A2(n4818), .B1(n4817), .B2(n4826), .ZN(U3520)
         );
  AOI22_X1 U5309 ( .A1(n4828), .A2(n4819), .B1(n2422), .B2(n4826), .ZN(U3521)
         );
  AOI22_X1 U5310 ( .A1(n4828), .A2(n4820), .B1(n2438), .B2(n4826), .ZN(U3522)
         );
  AOI22_X1 U5311 ( .A1(n4828), .A2(n4821), .B1(n2452), .B2(n4826), .ZN(U3523)
         );
  AOI22_X1 U5312 ( .A1(n4828), .A2(n4822), .B1(n2470), .B2(n4826), .ZN(U3525)
         );
  AOI22_X1 U5313 ( .A1(n4828), .A2(n4823), .B1(n2484), .B2(n4826), .ZN(U3526)
         );
  AOI22_X1 U5314 ( .A1(n4828), .A2(n4824), .B1(n3740), .B2(n4826), .ZN(U3527)
         );
  AOI22_X1 U5315 ( .A1(n4828), .A2(n4825), .B1(n2514), .B2(n4826), .ZN(U3528)
         );
  AOI22_X1 U5316 ( .A1(n4828), .A2(n4827), .B1(n2523), .B2(n4826), .ZN(U3529)
         );
endmodule

