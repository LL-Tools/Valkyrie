

module b21_C_gen_AntiSAT_k_128_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4309, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074;

  NAND2_X1 U4813 ( .A1(n4751), .A2(n4752), .ZN(n8245) );
  INV_X1 U4814 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U4815 ( .A1(n5677), .A2(n7228), .ZN(n7233) );
  INV_X2 U4816 ( .A(n5899), .ZN(n5916) );
  OR2_X1 U4817 ( .A1(n5911), .A2(n5910), .ZN(n5913) );
  INV_X1 U4818 ( .A(n5943), .ZN(n8645) );
  INV_X2 U4819 ( .A(n6504), .ZN(n5877) );
  INV_X1 U4821 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n4309) );
  INV_X1 U4823 ( .A(n6380), .ZN(n6346) );
  INV_X1 U4824 ( .A(n5638), .ZN(n6984) );
  NAND2_X1 U4825 ( .A1(n6935), .A2(n9930), .ZN(n5447) );
  INV_X2 U4826 ( .A(n7222), .ZN(n6255) );
  INV_X1 U4827 ( .A(n5117), .ZN(n5424) );
  INV_X1 U4828 ( .A(n5927), .ZN(n8639) );
  NAND2_X1 U4829 ( .A1(n4621), .A2(n7006), .ZN(n7363) );
  CLKBUF_X2 U4830 ( .A(n4344), .Z(n8650) );
  BUF_X1 U4831 ( .A(n9986), .Z(n4315) );
  OR2_X1 U4832 ( .A1(n7566), .A2(n7570), .ZN(n7568) );
  AND4_X1 U4833 ( .A1(n5958), .A2(n5957), .A3(n5956), .A4(n5955), .ZN(n7392)
         );
  NOR2_X1 U4834 ( .A1(n7776), .A2(n8707), .ZN(n7777) );
  NAND2_X1 U4835 ( .A1(n4694), .A2(n4892), .ZN(n5116) );
  INV_X2 U4836 ( .A(n9938), .ZN(n9942) );
  NAND2_X2 U4837 ( .A1(n9821), .A2(n9819), .ZN(n9823) );
  NAND2_X2 U4838 ( .A1(n7994), .A2(n7996), .ZN(n7995) );
  NAND2_X1 U4839 ( .A1(n6506), .A2(n4401), .ZN(n4311) );
  NAND2_X2 U4840 ( .A1(n7987), .A2(n5740), .ZN(n5741) );
  NAND2_X2 U4841 ( .A1(n5736), .A2(n7983), .ZN(n7987) );
  NAND2_X1 U4842 ( .A1(n5630), .A2(n5629), .ZN(n6970) );
  INV_X1 U4843 ( .A(n5761), .ZN(n5662) );
  XNOR2_X2 U4844 ( .A(n5850), .B(n5849), .ZN(n7752) );
  CLKBUF_X2 U4845 ( .A(n9916), .Z(n4312) );
  OAI21_X2 U4846 ( .B1(n6551), .B2(n5117), .A(n4367), .ZN(n9811) );
  AOI22_X2 U4847 ( .A1(n8245), .A2(n8244), .B1(n8479), .B2(n8065), .ZN(n8229)
         );
  NAND2_X2 U4848 ( .A1(n5179), .A2(n5178), .ZN(n9827) );
  OAI21_X2 U4849 ( .B1(n5215), .B2(n4928), .A(n4927), .ZN(n5229) );
  INV_X1 U4850 ( .A(n6478), .ZN(n5629) );
  AND2_X1 U4851 ( .A1(n4317), .A2(n4401), .ZN(n4313) );
  AND2_X1 U4852 ( .A1(n4317), .A2(n4401), .ZN(n4314) );
  OAI211_X1 U4855 ( .C1(n5117), .C2(n6549), .A(n5098), .B(n5097), .ZN(n9986)
         );
  NAND2_X1 U4856 ( .A1(n8625), .A2(n6343), .ZN(n8516) );
  NAND2_X1 U4857 ( .A1(n8558), .A2(n8559), .ZN(n8625) );
  NOR2_X1 U4858 ( .A1(n9112), .A2(n8744), .ZN(n9104) );
  NAND2_X1 U4859 ( .A1(n6327), .A2(n6326), .ZN(n9283) );
  NAND2_X1 U4860 ( .A1(n7568), .A2(n4847), .ZN(n7672) );
  NAND2_X1 U4861 ( .A1(n7233), .A2(n5679), .ZN(n7415) );
  NAND2_X2 U4862 ( .A1(n8848), .A2(n8924), .ZN(n8798) );
  INV_X1 U4863 ( .A(n7287), .ZN(n9773) );
  INV_X4 U4864 ( .A(n5909), .ZN(n6378) );
  INV_X1 U4865 ( .A(n9986), .ZN(n9885) );
  NAND2_X4 U4866 ( .A1(n7026), .A2(n7025), .ZN(n7222) );
  NAND2_X1 U4867 ( .A1(n5580), .A2(n5579), .ZN(n6446) );
  CLKBUF_X3 U4868 ( .A(n5893), .Z(n6356) );
  NAND2_X1 U4869 ( .A1(n6447), .A2(n9958), .ZN(n5579) );
  INV_X1 U4870 ( .A(n6952), .ZN(n9761) );
  INV_X1 U4871 ( .A(n6380), .ZN(n5880) );
  INV_X1 U4872 ( .A(n6379), .ZN(n4316) );
  INV_X1 U4873 ( .A(n9930), .ZN(n9968) );
  NAND2_X1 U4874 ( .A1(n6506), .A2(n4401), .ZN(n5943) );
  INV_X4 U4875 ( .A(n6506), .ZN(n5921) );
  CLKBUF_X2 U4876 ( .A(n5074), .Z(n4324) );
  CLKBUF_X2 U4877 ( .A(n5074), .Z(n4323) );
  NOR2_X1 U4878 ( .A1(n6388), .A2(n7752), .ZN(n5851) );
  AND2_X1 U4879 ( .A1(n8501), .A2(n8503), .ZN(n5074) );
  NOR2_X1 U4880 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4565) );
  INV_X2 U4881 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AOI211_X1 U4882 ( .C1(n9272), .C2(n9240), .A(n9078), .B(n9077), .ZN(n9079)
         );
  NOR2_X1 U4883 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U4884 ( .A1(n4571), .A2(n4569), .ZN(n9269) );
  NOR2_X1 U4885 ( .A1(n7962), .A2(n7961), .ZN(n8017) );
  NOR3_X1 U4886 ( .A1(n8788), .A2(n8905), .A3(n6386), .ZN(n8913) );
  OR2_X1 U4887 ( .A1(n9046), .A2(n9246), .ZN(n4571) );
  AOI21_X1 U4888 ( .B1(n9076), .B2(n9237), .A(n9075), .ZN(n9270) );
  AOI211_X1 U4889 ( .C1(n9347), .C2(n9290), .A(n9289), .B(n9288), .ZN(n9291)
         );
  AOI21_X1 U4890 ( .B1(n9092), .B2(n9237), .A(n4402), .ZN(n9286) );
  XOR2_X1 U4891 ( .A(n9105), .B(n9104), .Z(n9106) );
  AOI21_X1 U4892 ( .B1(n9150), .B2(n8794), .A(n8793), .ZN(n9135) );
  NAND2_X1 U4893 ( .A1(n4764), .A2(n4761), .ZN(n8365) );
  NAND2_X1 U4894 ( .A1(n8232), .A2(n5433), .ZN(n8244) );
  NAND2_X1 U4895 ( .A1(n7733), .A2(n4762), .ZN(n4764) );
  NAND2_X1 U4896 ( .A1(n5369), .A2(n5368), .ZN(n8406) );
  NAND2_X1 U4897 ( .A1(n7415), .A2(n4830), .ZN(n7423) );
  NAND2_X1 U4898 ( .A1(n4745), .A2(n4748), .ZN(n7519) );
  CLKBUF_X1 U4899 ( .A(n7508), .Z(n4406) );
  NAND2_X1 U4900 ( .A1(n7387), .A2(n7386), .ZN(n7508) );
  NAND2_X1 U4901 ( .A1(n5167), .A2(n5166), .ZN(n9877) );
  AND2_X1 U4902 ( .A1(n5463), .A2(n5462), .ZN(n7070) );
  NOR2_X1 U4903 ( .A1(n7274), .A2(n7287), .ZN(n7396) );
  INV_X1 U4904 ( .A(n7385), .ZN(n9780) );
  AOI21_X1 U4905 ( .B1(n6566), .B2(n8645), .A(n4429), .ZN(n7583) );
  AND2_X1 U4906 ( .A1(n4728), .A2(n5121), .ZN(n7264) );
  AND4_X1 U4907 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n7369)
         );
  AND4_X1 U4908 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n7302)
         );
  INV_X1 U4909 ( .A(n6915), .ZN(n8104) );
  INV_X1 U4910 ( .A(n5048), .ZN(n6447) );
  INV_X1 U4911 ( .A(n6379), .ZN(n5893) );
  NAND4_X1 U4912 ( .A1(n5042), .A2(n5041), .A3(n5040), .A4(n5039), .ZN(n5048)
         );
  CLKBUF_X3 U4913 ( .A(n5914), .Z(n6298) );
  OAI211_X1 U4914 ( .C1(n8655), .C2(n6676), .A(n5929), .B(n5928), .ZN(n6952)
         );
  CLKBUF_X1 U4915 ( .A(n5875), .Z(n7025) );
  AND2_X1 U4916 ( .A1(n5827), .A2(n5826), .ZN(n5914) );
  NAND2_X2 U4917 ( .A1(n5631), .A2(n6970), .ZN(n5761) );
  OR2_X1 U4918 ( .A1(n10004), .A2(n8254), .ZN(n5638) );
  OAI211_X1 U4919 ( .C1(n5117), .C2(n6546), .A(n5058), .B(n5057), .ZN(n9930)
         );
  BUF_X2 U4920 ( .A(n5068), .Z(n4319) );
  XNOR2_X1 U4921 ( .A(n5842), .B(n5841), .ZN(n8947) );
  NAND2_X4 U4922 ( .A1(n6423), .A2(n8951), .ZN(n6506) );
  CLKBUF_X1 U4923 ( .A(n5067), .Z(n5409) );
  NAND2_X1 U4924 ( .A1(n5825), .A2(n5824), .ZN(n7912) );
  OAI21_X1 U4925 ( .B1(n5873), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5867) );
  AND2_X1 U4926 ( .A1(n5874), .A2(n5873), .ZN(n9018) );
  MUX2_X1 U4927 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5823), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5825) );
  NAND2_X1 U4928 ( .A1(n5572), .A2(n7463), .ZN(n6972) );
  NAND2_X1 U4929 ( .A1(n5848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U4930 ( .A1(n4864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4865) );
  CLKBUF_X1 U4931 ( .A(n5429), .Z(n7343) );
  INV_X1 U4932 ( .A(n5024), .ZN(n8503) );
  NAND2_X1 U4933 ( .A1(n5863), .A2(n5862), .ZN(n8951) );
  XNOR2_X1 U4934 ( .A(n4862), .B(n5000), .ZN(n7463) );
  CLKBUF_X1 U4935 ( .A(n5822), .Z(n5858) );
  XNOR2_X1 U4936 ( .A(n5607), .B(n5608), .ZN(n5572) );
  NAND2_X1 U4937 ( .A1(n5021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5022) );
  XNOR2_X1 U4938 ( .A(n5013), .B(n5012), .ZN(n6703) );
  OR2_X1 U4939 ( .A1(n4863), .A2(n8498), .ZN(n4866) );
  NAND2_X1 U4940 ( .A1(n5010), .A2(n5016), .ZN(n5622) );
  AND2_X1 U4941 ( .A1(n4860), .A2(n4826), .ZN(n4863) );
  MUX2_X1 U4942 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5007), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5010) );
  NOR2_X1 U4943 ( .A1(n5618), .A2(n4768), .ZN(n4766) );
  NAND2_X2 U4944 ( .A1(n4401), .A2(P1_U3084), .ZN(n9378) );
  NAND2_X1 U4945 ( .A1(n5006), .A2(n4769), .ZN(n4768) );
  AND2_X1 U4946 ( .A1(n4856), .A2(n4855), .ZN(n4840) );
  INV_X1 U4947 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5834) );
  INV_X1 U4948 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5991) );
  INV_X1 U4949 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4998) );
  INV_X1 U4950 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U4951 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4564) );
  NOR2_X1 U4952 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4566) );
  NOR2_X1 U4953 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4855) );
  INV_X1 U4954 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5849) );
  NOR2_X1 U4955 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4857) );
  INV_X1 U4956 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5002) );
  NOR2_X1 U4957 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6151) );
  NOR2_X1 U4958 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9596) );
  AND2_X1 U4959 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9595) );
  NAND2_X1 U4960 ( .A1(n5622), .A2(n6703), .ZN(n4317) );
  NAND2_X2 U4961 ( .A1(n5622), .A2(n6703), .ZN(n6700) );
  INV_X1 U4962 ( .A(n7963), .ZN(n7962) );
  XNOR2_X1 U4963 ( .A(n4824), .B(n5747), .ZN(n7963) );
  NAND2_X1 U4964 ( .A1(n6461), .A2(n5129), .ZN(n6463) );
  OAI21_X2 U4966 ( .B1(n9826), .B2(n4834), .A(n4833), .ZN(n9637) );
  NAND2_X2 U4967 ( .A1(n9823), .A2(n9820), .ZN(n9826) );
  AND2_X1 U4968 ( .A1(n8503), .A2(n5023), .ZN(n4318) );
  BUF_X2 U4969 ( .A(n5068), .Z(n4320) );
  NAND2_X2 U4970 ( .A1(n5833), .A2(n5814), .ZN(n6411) );
  NOR2_X4 U4971 ( .A1(n6075), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U4972 ( .A1(n5631), .A2(n6970), .ZN(n4321) );
  NAND2_X1 U4973 ( .A1(n5631), .A2(n6970), .ZN(n4322) );
  XNOR2_X2 U4974 ( .A(n5844), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6393) );
  OAI22_X2 U4975 ( .A1(n8296), .A2(n8297), .B1(n8083), .B2(n8299), .ZN(n8282)
         );
  AOI22_X2 U4976 ( .A1(n8308), .A2(n6472), .B1(n6471), .B2(n8318), .ZN(n8296)
         );
  AOI21_X2 U4977 ( .B1(n8602), .B2(n8605), .A(n8604), .ZN(n8531) );
  NOR2_X2 U4978 ( .A1(n6276), .A2(n6275), .ZN(n8604) );
  INV_X1 U4979 ( .A(n5899), .ZN(n4325) );
  INV_X1 U4980 ( .A(n4325), .ZN(n4326) );
  XNOR2_X2 U4982 ( .A(n7041), .B(n7032), .ZN(n7028) );
  NAND4_X4 U4983 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n7041)
         );
  OAI222_X1 U4984 ( .A1(n9378), .A2(n9371), .B1(P1_U3084), .B2(n5828), .C1(
        n9370), .C2(n9369), .ZN(P1_U3323) );
  XNOR2_X2 U4985 ( .A(n5821), .B(n5820), .ZN(n5828) );
  OR2_X1 U4986 ( .A1(n8329), .A2(n7985), .ZN(n5522) );
  INV_X1 U4987 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4867) );
  NAND2_X1 U4988 ( .A1(n9595), .A2(n4868), .ZN(n4869) );
  INV_X1 U4989 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4868) );
  AOI21_X1 U4990 ( .B1(n7915), .B2(n7914), .A(n4425), .ZN(n4424) );
  OR2_X1 U4991 ( .A1(n9339), .A2(n8965), .ZN(n7914) );
  NOR2_X1 U4992 ( .A1(n7916), .A2(n9247), .ZN(n4425) );
  NAND2_X1 U4993 ( .A1(n5160), .A2(n5159), .ZN(n4912) );
  AND2_X1 U4994 ( .A1(n6745), .A2(n6423), .ZN(n9234) );
  NAND2_X1 U4995 ( .A1(n6506), .A2(n4574), .ZN(n4573) );
  INV_X1 U4996 ( .A(n4690), .ZN(n4689) );
  OAI21_X1 U4997 ( .B1(n5380), .B2(n4691), .A(n5390), .ZN(n4690) );
  INV_X1 U4998 ( .A(n4650), .ZN(n4649) );
  AOI21_X1 U4999 ( .B1(n4539), .B2(n5568), .A(n4369), .ZN(n4538) );
  OR2_X1 U5000 ( .A1(n8271), .A2(n8020), .ZN(n5532) );
  OR2_X1 U5001 ( .A1(n8299), .A2(n7964), .ZN(n5525) );
  OR2_X1 U5002 ( .A1(n7743), .A2(n7744), .ZN(n7834) );
  INV_X1 U5003 ( .A(n4768), .ZN(n4767) );
  NOR2_X1 U5004 ( .A1(n9626), .A2(n4643), .ZN(n8782) );
  AND2_X1 U5005 ( .A1(n8790), .A2(n9027), .ZN(n4643) );
  OR2_X1 U5006 ( .A1(n9290), .A2(n9116), .ZN(n9086) );
  INV_X1 U5007 ( .A(n4780), .ZN(n4423) );
  OAI21_X1 U5008 ( .B1(n4781), .B2(n4331), .A(n4366), .ZN(n4780) );
  NAND2_X1 U5009 ( .A1(n9132), .A2(n9153), .ZN(n4790) );
  AND2_X1 U5010 ( .A1(n9305), .A2(n9161), .ZN(n4791) );
  AND2_X1 U5011 ( .A1(n9305), .A2(n8553), .ZN(n8793) );
  OR2_X1 U5012 ( .A1(n9305), .A2(n8553), .ZN(n8794) );
  NAND2_X1 U5013 ( .A1(n4455), .A2(n9249), .ZN(n4778) );
  OR2_X1 U5014 ( .A1(n8707), .A2(n9607), .ZN(n7756) );
  INV_X1 U5015 ( .A(n7388), .ZN(n7387) );
  AND2_X1 U5016 ( .A1(n5878), .A2(n9018), .ZN(n8781) );
  INV_X1 U5017 ( .A(n9208), .ZN(n9202) );
  NAND2_X1 U5018 ( .A1(n4995), .A2(n4994), .ZN(n5420) );
  OAI21_X1 U5019 ( .B1(n5318), .B2(n5317), .A(n4961), .ZN(n5331) );
  AND2_X1 U5020 ( .A1(n4968), .A2(n4967), .ZN(n5330) );
  INV_X1 U5021 ( .A(SI_21_), .ZN(n4954) );
  NAND2_X1 U5022 ( .A1(n4953), .A2(n4952), .ZN(n5305) );
  NAND2_X1 U5023 ( .A1(n5296), .A2(n5295), .ZN(n4953) );
  AOI21_X1 U5024 ( .B1(n4670), .B2(n4346), .A(n4669), .ZN(n4668) );
  AND2_X1 U5025 ( .A1(n4924), .A2(n4923), .ZN(n5201) );
  INV_X1 U5026 ( .A(n4671), .ZN(n4670) );
  OAI21_X1 U5027 ( .B1(n4674), .B2(n4346), .A(n4919), .ZN(n4671) );
  AOI21_X1 U5028 ( .B1(n4679), .B2(n4682), .A(n4678), .ZN(n4677) );
  OR2_X1 U5029 ( .A1(n6017), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6056) );
  AND2_X1 U5030 ( .A1(n4871), .A2(n4872), .ZN(n4696) );
  INV_X1 U5031 ( .A(n4822), .ZN(n4821) );
  AOI22_X1 U5032 ( .A1(n5746), .A2(n4823), .B1(n5748), .B2(n5747), .ZN(n4822)
         );
  AOI21_X1 U5033 ( .B1(n4328), .B2(n8281), .A(n4372), .ZN(n4752) );
  AND2_X1 U5034 ( .A1(n8421), .A2(n8082), .ZN(n6473) );
  OR2_X1 U5035 ( .A1(n8278), .A2(n4558), .ZN(n4440) );
  INV_X1 U5036 ( .A(n4735), .ZN(n8308) );
  NAND2_X1 U5037 ( .A1(n4743), .A2(n8322), .ZN(n4739) );
  INV_X1 U5038 ( .A(n4737), .ZN(n4736) );
  NOR2_X1 U5039 ( .A1(n7827), .A2(n4763), .ZN(n4762) );
  INV_X1 U5040 ( .A(n4765), .ZN(n4763) );
  INV_X1 U5041 ( .A(n4851), .ZN(n4757) );
  NAND2_X1 U5042 ( .A1(n7114), .A2(n5130), .ZN(n7069) );
  NAND2_X1 U5043 ( .A1(n8101), .A2(n9885), .ZN(n7113) );
  NAND3_X1 U5044 ( .A1(n4870), .A2(n4869), .A3(n4873), .ZN(n5038) );
  INV_X1 U5045 ( .A(n6298), .ZN(n6425) );
  AND2_X1 U5046 ( .A1(n4795), .A2(n9070), .ZN(n4794) );
  NAND2_X1 U5047 ( .A1(n4796), .A2(n4800), .ZN(n4795) );
  AND2_X1 U5048 ( .A1(n4602), .A2(n8792), .ZN(n9089) );
  OR2_X1 U5049 ( .A1(n8557), .A2(n9183), .ZN(n4845) );
  NAND2_X1 U5050 ( .A1(n9178), .A2(n7918), .ZN(n4422) );
  AND4_X1 U5051 ( .A1(n6221), .A2(n6220), .A3(n6219), .A4(n6218), .ZN(n9182)
         );
  INV_X1 U5052 ( .A(n4775), .ZN(n4774) );
  AND2_X1 U5053 ( .A1(n9346), .A2(n8966), .ZN(n7863) );
  INV_X1 U5054 ( .A(n9248), .ZN(n9232) );
  NAND2_X1 U5055 ( .A1(n8641), .A2(n8640), .ZN(n9267) );
  INV_X1 U5056 ( .A(n9269), .ZN(n4431) );
  INV_X1 U5057 ( .A(n9380), .ZN(n4464) );
  NAND2_X1 U5058 ( .A1(n4556), .A2(n4889), .ZN(n5109) );
  INV_X1 U5059 ( .A(n4553), .ZN(n4552) );
  INV_X1 U5060 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U5061 ( .B1(n8168), .B2(n9869), .A(n4533), .ZN(n4532) );
  AOI21_X1 U5062 ( .B1(n8170), .B2(n9864), .A(n8169), .ZN(n4533) );
  AND2_X1 U5063 ( .A1(n6368), .A2(n6329), .ZN(n9083) );
  NAND2_X1 U5064 ( .A1(n5817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5856) );
  AOI211_X1 U5065 ( .C1(n5510), .C2(n4559), .A(n4558), .B(n4557), .ZN(n5531)
         );
  NOR2_X1 U5066 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  OAI22_X1 U5067 ( .A1(n5525), .A2(n5559), .B1(n5511), .B2(n5570), .ZN(n4557)
         );
  OAI22_X1 U5068 ( .A1(n4542), .A2(n5542), .B1(n5541), .B2(n5570), .ZN(n4541)
         );
  AOI21_X1 U5069 ( .B1(n4544), .B2(n4543), .A(n4412), .ZN(n4542) );
  NOR2_X1 U5070 ( .A1(n8406), .A2(n8253), .ZN(n4486) );
  INV_X1 U5071 ( .A(n4988), .ZN(n4691) );
  NAND2_X1 U5072 ( .A1(n4653), .A2(n5258), .ZN(n4647) );
  NOR2_X1 U5073 ( .A1(n4649), .A2(n4940), .ZN(n4648) );
  AOI21_X1 U5074 ( .B1(n5228), .B2(n4932), .A(n4655), .ZN(n4654) );
  INV_X1 U5075 ( .A(n5245), .ZN(n4655) );
  NOR2_X1 U5076 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4562) );
  NOR2_X1 U5077 ( .A1(n5131), .A2(n4684), .ZN(n4683) );
  INV_X1 U5078 ( .A(n4895), .ZN(n4684) );
  NAND2_X1 U5079 ( .A1(n4700), .A2(n4360), .ZN(n4704) );
  NAND2_X1 U5080 ( .A1(n4708), .A2(n4710), .ZN(n4700) );
  INV_X1 U5081 ( .A(n4711), .ZN(n4710) );
  NOR2_X1 U5082 ( .A1(n8378), .A2(n4443), .ZN(n4442) );
  INV_X1 U5083 ( .A(n5501), .ZN(n4443) );
  OR2_X1 U5084 ( .A1(n7663), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U5085 ( .A1(n7732), .A2(n4480), .ZN(n4479) );
  OR2_X1 U5086 ( .A1(n5429), .A2(n5572), .ZN(n5628) );
  NAND2_X1 U5087 ( .A1(n4859), .A2(n4829), .ZN(n4828) );
  INV_X1 U5088 ( .A(n8616), .ZN(n4632) );
  OAI22_X1 U5089 ( .A1(n7392), .A2(n6379), .B1(n9773), .B2(n6380), .ZN(n5964)
         );
  NAND2_X1 U5090 ( .A1(n4371), .A2(n4811), .ZN(n4810) );
  OR2_X1 U5091 ( .A1(n9280), .A2(n8631), .ZN(n9040) );
  INV_X1 U5092 ( .A(n4506), .ZN(n4503) );
  NAND2_X1 U5093 ( .A1(n8527), .A2(n4462), .ZN(n4461) );
  NAND2_X1 U5094 ( .A1(n4602), .A2(n4603), .ZN(n4601) );
  INV_X1 U5095 ( .A(n4601), .ZN(n4599) );
  NAND2_X1 U5096 ( .A1(n9040), .A2(n8898), .ZN(n9035) );
  NOR2_X1 U5097 ( .A1(n8744), .A2(n4604), .ZN(n4603) );
  INV_X1 U5098 ( .A(n8758), .ZN(n4604) );
  OR2_X1 U5099 ( .A1(n9298), .A2(n9153), .ZN(n8862) );
  NOR2_X1 U5100 ( .A1(n4585), .A2(n9194), .ZN(n4584) );
  NOR2_X1 U5101 ( .A1(n7923), .A2(n8867), .ZN(n4585) );
  NOR2_X1 U5102 ( .A1(n9336), .A2(n9339), .ZN(n4456) );
  OR2_X1 U5103 ( .A1(n6041), .A2(n6040), .ZN(n6061) );
  OR2_X1 U5104 ( .A1(n4806), .A2(n8805), .ZN(n4416) );
  NAND2_X1 U5105 ( .A1(n5423), .A2(n4664), .ZN(n4663) );
  INV_X1 U5106 ( .A(n4666), .ZN(n4664) );
  NOR2_X1 U5107 ( .A1(n5423), .A2(n4662), .ZN(n4661) );
  INV_X1 U5108 ( .A(n4665), .ZN(n4662) );
  NAND2_X1 U5109 ( .A1(n5423), .A2(n4665), .ZN(n4659) );
  AND2_X1 U5110 ( .A1(n4666), .A2(n4665), .ZN(n4660) );
  AND2_X1 U5111 ( .A1(n4988), .A2(n4987), .ZN(n5380) );
  NAND2_X1 U5112 ( .A1(n4982), .A2(n4981), .ZN(n5379) );
  OAI21_X1 U5113 ( .B1(n5355), .B2(n5354), .A(n4976), .ZN(n5367) );
  AND2_X1 U5114 ( .A1(n4812), .A2(n5849), .ZN(n4811) );
  INV_X1 U5115 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4812) );
  OAI21_X1 U5116 ( .B1(n5305), .B2(n4955), .A(n4957), .ZN(n5318) );
  NAND2_X1 U5117 ( .A1(n4944), .A2(n4943), .ZN(n5287) );
  AND2_X1 U5118 ( .A1(n5836), .A2(n5834), .ZN(n4639) );
  AOI21_X1 U5119 ( .B1(n4654), .B2(n4652), .A(n4651), .ZN(n4650) );
  INV_X1 U5120 ( .A(n4937), .ZN(n4651) );
  INV_X1 U5121 ( .A(n4932), .ZN(n4652) );
  INV_X1 U5122 ( .A(n4654), .ZN(n4653) );
  NOR2_X1 U5123 ( .A1(n4915), .A2(n4675), .ZN(n4674) );
  INV_X1 U5124 ( .A(n4911), .ZN(n4675) );
  AND2_X1 U5125 ( .A1(n4905), .A2(n4904), .ZN(n5144) );
  AOI21_X1 U5126 ( .B1(n4683), .B2(n4681), .A(n4680), .ZN(n4679) );
  INV_X1 U5127 ( .A(n4900), .ZN(n4680) );
  INV_X1 U5128 ( .A(n5115), .ZN(n4681) );
  INV_X1 U5129 ( .A(n4683), .ZN(n4682) );
  INV_X1 U5130 ( .A(SI_17_), .ZN(n9502) );
  XNOR2_X1 U5132 ( .A(n4321), .B(n9958), .ZN(n5633) );
  NAND2_X1 U5133 ( .A1(n5745), .A2(n5744), .ZN(n4824) );
  NAND2_X1 U5134 ( .A1(n5279), .A2(n5278), .ZN(n5290) );
  AOI21_X1 U5135 ( .B1(n4538), .B2(n4536), .A(n6478), .ZN(n4535) );
  INV_X1 U5136 ( .A(n4539), .ZN(n4536) );
  OR2_X1 U5137 ( .A1(n5569), .A2(n4537), .ZN(n4534) );
  INV_X1 U5138 ( .A(n4538), .ZN(n4537) );
  INV_X1 U5139 ( .A(n4702), .ZN(n4701) );
  OAI21_X1 U5140 ( .B1(n4705), .B2(n4704), .A(n5600), .ZN(n4702) );
  NAND2_X1 U5141 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  INV_X1 U5142 ( .A(n4712), .ZN(n4706) );
  INV_X1 U5143 ( .A(n4319), .ZN(n5412) );
  NOR2_X2 U5144 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5055) );
  NOR2_X1 U5145 ( .A1(n7188), .A2(n4526), .ZN(n8132) );
  AND2_X1 U5146 ( .A1(n7189), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4526) );
  OR2_X1 U5147 ( .A1(n6487), .A2(n8196), .ZN(n8181) );
  OR2_X1 U5148 ( .A1(n5370), .A2(n9527), .ZN(n5395) );
  OR2_X1 U5149 ( .A1(n8253), .A2(n8065), .ZN(n8232) );
  AND2_X1 U5150 ( .A1(n5539), .A2(n8218), .ZN(n8231) );
  INV_X1 U5151 ( .A(n6473), .ZN(n4754) );
  OR2_X1 U5152 ( .A1(n8298), .A2(n8299), .ZN(n8300) );
  NAND2_X1 U5153 ( .A1(n4723), .A2(n4724), .ZN(n8278) );
  AOI21_X1 U5154 ( .B1(n4726), .B2(n8310), .A(n4725), .ZN(n4724) );
  INV_X1 U5155 ( .A(n5525), .ZN(n4725) );
  AND2_X1 U5156 ( .A1(n5525), .A2(n5511), .ZN(n8297) );
  NOR2_X1 U5157 ( .A1(n8291), .A2(n5521), .ZN(n4726) );
  OR2_X1 U5158 ( .A1(n8309), .A2(n8310), .ZN(n4727) );
  AOI21_X1 U5159 ( .B1(n4743), .B2(n4741), .A(n4365), .ZN(n4740) );
  INV_X1 U5160 ( .A(n6469), .ZN(n4741) );
  NAND2_X1 U5161 ( .A1(n8338), .A2(n8337), .ZN(n4720) );
  AND2_X1 U5162 ( .A1(n5514), .A2(n5515), .ZN(n8337) );
  NOR2_X1 U5163 ( .A1(n7834), .A2(n8459), .ZN(n8368) );
  AND2_X1 U5164 ( .A1(n8378), .A2(n4341), .ZN(n4761) );
  NAND2_X1 U5165 ( .A1(n7736), .A2(n4721), .ZN(n7829) );
  NOR2_X1 U5166 ( .A1(n7832), .A2(n4722), .ZN(n4721) );
  INV_X1 U5167 ( .A(n5497), .ZN(n4722) );
  NAND2_X1 U5168 ( .A1(n7738), .A2(n7737), .ZN(n7736) );
  AND2_X1 U5169 ( .A1(n5490), .A2(n5489), .ZN(n7570) );
  NOR2_X1 U5170 ( .A1(n7596), .A2(n9827), .ZN(n7528) );
  NOR3_X1 U5171 ( .A1(n7596), .A2(n7663), .A3(n9827), .ZN(n7574) );
  NAND2_X1 U5172 ( .A1(n4718), .A2(n5473), .ZN(n4716) );
  AOI21_X1 U5173 ( .B1(n6466), .B2(n4749), .A(n4353), .ZN(n4748) );
  NAND2_X1 U5174 ( .A1(n7593), .A2(n4746), .ZN(n4745) );
  INV_X1 U5175 ( .A(n6465), .ZN(n4749) );
  NAND2_X1 U5176 ( .A1(n4719), .A2(n4717), .ZN(n7598) );
  INV_X1 U5177 ( .A(n4718), .ZN(n4717) );
  NAND2_X1 U5178 ( .A1(n7177), .A2(n5467), .ZN(n7317) );
  NOR2_X1 U5179 ( .A1(n7178), .A2(n4760), .ZN(n4759) );
  INV_X1 U5180 ( .A(n6462), .ZN(n4760) );
  NAND2_X1 U5181 ( .A1(n7264), .A2(n8099), .ZN(n5463) );
  NAND2_X1 U5182 ( .A1(n4441), .A2(n7069), .ZN(n7177) );
  AND2_X1 U5183 ( .A1(n7178), .A2(n5463), .ZN(n4441) );
  NAND2_X1 U5184 ( .A1(n9891), .A2(n5114), .ZN(n7114) );
  NAND2_X1 U5185 ( .A1(n4335), .A2(n6457), .ZN(n4732) );
  NAND2_X1 U5186 ( .A1(n7071), .A2(n5460), .ZN(n7117) );
  OR2_X1 U5187 ( .A1(n6477), .A2(n8254), .ZN(n7602) );
  NAND2_X1 U5188 ( .A1(n8102), .A2(n9979), .ZN(n9889) );
  AND2_X1 U5189 ( .A1(n5438), .A2(n7113), .ZN(n9887) );
  INV_X1 U5190 ( .A(n9922), .ZN(n9907) );
  NAND2_X1 U5191 ( .A1(n5628), .A2(n6482), .ZN(n9922) );
  NOR2_X1 U5192 ( .A1(n9958), .A2(n9951), .ZN(n9924) );
  NAND2_X1 U5193 ( .A1(n5427), .A2(n5426), .ZN(n8175) );
  NAND2_X1 U5194 ( .A1(n5307), .A2(n5306), .ZN(n8433) );
  NAND2_X1 U5195 ( .A1(n5275), .A2(n5274), .ZN(n8357) );
  NAND2_X1 U5196 ( .A1(n5235), .A2(n5234), .ZN(n7744) );
  INV_X1 U5197 ( .A(n9811), .ZN(n9979) );
  OR2_X1 U5198 ( .A1(n9946), .A2(n5785), .ZN(n6966) );
  AND2_X1 U5199 ( .A1(n6489), .A2(n6904), .ZN(n6968) );
  NAND2_X1 U5200 ( .A1(n5021), .A2(n5020), .ZN(n5024) );
  NAND2_X1 U5201 ( .A1(n5609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U5202 ( .A1(n5607), .A2(n5608), .ZN(n5609) );
  OAI211_X1 U5203 ( .C1(n8655), .C2(n6619), .A(n5994), .B(n5993), .ZN(n7385)
         );
  OAI21_X1 U5204 ( .B1(n8595), .B2(n8549), .A(n8548), .ZN(n8547) );
  OR2_X1 U5205 ( .A1(n6136), .A2(n6135), .ZN(n6158) );
  NAND2_X1 U5206 ( .A1(n4636), .A2(n4634), .ZN(n7465) );
  NOR2_X1 U5207 ( .A1(n4635), .A2(n7467), .ZN(n4634) );
  INV_X1 U5208 ( .A(n4637), .ZN(n4635) );
  INV_X1 U5209 ( .A(n8591), .ZN(n4626) );
  OR2_X1 U5210 ( .A1(n6211), .A2(n4632), .ZN(n4630) );
  AND2_X1 U5211 ( .A1(n8538), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U5212 ( .A1(n4631), .A2(n4630), .ZN(n4629) );
  AND2_X1 U5213 ( .A1(n6211), .A2(n4632), .ZN(n4631) );
  AND2_X1 U5214 ( .A1(n8947), .A2(n9168), .ZN(n6418) );
  AOI21_X1 U5215 ( .B1(n8658), .B2(n8908), .A(n8657), .ZN(n8785) );
  NAND2_X1 U5216 ( .A1(n6619), .A2(n6514), .ZN(n4504) );
  INV_X1 U5217 ( .A(n4504), .ZN(n4502) );
  INV_X1 U5218 ( .A(n4500), .ZN(n4499) );
  OAI21_X1 U5219 ( .B1(n4348), .B2(n4502), .A(n4501), .ZN(n4500) );
  INV_X1 U5220 ( .A(n6605), .ZN(n4501) );
  NOR2_X1 U5221 ( .A1(n6687), .A2(n4385), .ZN(n6691) );
  OAI21_X1 U5222 ( .B1(n9705), .B2(n4491), .A(n4490), .ZN(n9716) );
  NAND2_X1 U5223 ( .A1(n4494), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5224 ( .A1(n8985), .A2(n4494), .ZN(n4490) );
  INV_X1 U5225 ( .A(n9717), .ZN(n4494) );
  OR2_X1 U5226 ( .A1(n9705), .A2(n9704), .ZN(n4493) );
  NOR2_X1 U5227 ( .A1(n9727), .A2(n4400), .ZN(n9743) );
  NOR2_X1 U5228 ( .A1(n9743), .A2(n9744), .ZN(n9742) );
  NAND2_X1 U5229 ( .A1(n8648), .A2(n8647), .ZN(n9031) );
  INV_X1 U5230 ( .A(n9035), .ZN(n8827) );
  NOR3_X1 U5231 ( .A1(n9117), .A2(n9283), .A3(n9290), .ZN(n9081) );
  AND2_X1 U5232 ( .A1(n6304), .A2(n6303), .ZN(n9107) );
  NAND2_X1 U5233 ( .A1(n4782), .A2(n4790), .ZN(n4781) );
  INV_X1 U5234 ( .A(n4785), .ZN(n4782) );
  AOI21_X1 U5235 ( .B1(n4787), .B2(n4786), .A(n4361), .ZN(n4785) );
  NAND2_X1 U5236 ( .A1(n4787), .A2(n4790), .ZN(n4783) );
  NOR2_X1 U5237 ( .A1(n4791), .A2(n4789), .ZN(n4788) );
  INV_X1 U5238 ( .A(n4845), .ZN(n4789) );
  AND2_X1 U5239 ( .A1(n8862), .A2(n8746), .ZN(n9134) );
  AND2_X1 U5240 ( .A1(n8795), .A2(n8794), .ZN(n9151) );
  AND3_X1 U5241 ( .A1(n6252), .A2(n6251), .A3(n6250), .ZN(n9183) );
  NAND2_X1 U5242 ( .A1(n4582), .A2(n8726), .ZN(n4581) );
  INV_X1 U5243 ( .A(n4584), .ZN(n4582) );
  NAND2_X1 U5244 ( .A1(n8726), .A2(n8869), .ZN(n4583) );
  AND2_X1 U5245 ( .A1(n9156), .A2(n8796), .ZN(n9179) );
  AOI22_X1 U5246 ( .A1(n9192), .A2(n7917), .B1(n9221), .B2(n9202), .ZN(n9178)
         );
  AND4_X1 U5247 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n9197)
         );
  OAI21_X1 U5248 ( .B1(n9218), .B2(n7923), .A(n4584), .ZN(n4586) );
  NAND2_X1 U5249 ( .A1(n4373), .A2(n4778), .ZN(n4775) );
  AND2_X1 U5250 ( .A1(n9336), .A2(n9233), .ZN(n4779) );
  NOR2_X1 U5251 ( .A1(n4428), .A2(n4383), .ZN(n4427) );
  NAND2_X1 U5252 ( .A1(n4350), .A2(n4329), .ZN(n4587) );
  OAI22_X1 U5253 ( .A1(n7537), .A2(n7536), .B1(n7535), .B2(n8970), .ZN(n7614)
         );
  AND2_X1 U5254 ( .A1(n8679), .A2(n8681), .ZN(n8809) );
  INV_X1 U5255 ( .A(n8809), .ZN(n7554) );
  OAI21_X1 U5256 ( .B1(n7394), .B2(n8803), .A(n7393), .ZN(n7395) );
  AND4_X1 U5257 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n7504)
         );
  AND2_X1 U5258 ( .A1(n8664), .A2(n8853), .ZN(n8801) );
  NAND2_X1 U5259 ( .A1(n7136), .A2(n8797), .ZN(n7219) );
  NAND2_X1 U5260 ( .A1(n8663), .A2(n8854), .ZN(n8797) );
  AND4_X2 U5261 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n7303)
         );
  NAND2_X1 U5262 ( .A1(n7045), .A2(n7044), .ZN(n7134) );
  OR2_X1 U5263 ( .A1(n7030), .A2(n6423), .ZN(n9248) );
  AND2_X1 U5264 ( .A1(n8787), .A2(n8906), .ZN(n9246) );
  NAND2_X1 U5265 ( .A1(n8956), .A2(n9168), .ZN(n7026) );
  INV_X1 U5266 ( .A(n9234), .ZN(n9250) );
  INV_X1 U5267 ( .A(n9122), .ZN(n9295) );
  NAND2_X1 U5268 ( .A1(n6227), .A2(n6226), .ZN(n9316) );
  NOR2_X1 U5269 ( .A1(n6772), .A2(n6771), .ZN(n7097) );
  INV_X1 U5270 ( .A(n9790), .ZN(n9653) );
  INV_X1 U5271 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5866) );
  INV_X1 U5272 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5839) );
  INV_X1 U5273 ( .A(n5871), .ZN(n5840) );
  INV_X1 U5274 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6174) );
  OAI21_X1 U5275 ( .B1(n5229), .B2(n5228), .A(n4932), .ZN(n5246) );
  OAI21_X1 U5276 ( .B1(n4912), .B2(n4346), .A(n4670), .ZN(n5202) );
  XNOR2_X1 U5277 ( .A(n4545), .B(n5175), .ZN(n6596) );
  NAND2_X1 U5278 ( .A1(n4912), .A2(n4911), .ZN(n4545) );
  NAND2_X1 U5279 ( .A1(n4685), .A2(n4895), .ZN(n5132) );
  NAND2_X1 U5280 ( .A1(n5116), .A2(n5115), .ZN(n4685) );
  NAND2_X1 U5281 ( .A1(n4409), .A2(n4883), .ZN(n5080) );
  NOR2_X1 U5282 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5807) );
  AND2_X1 U5283 ( .A1(n4465), .A2(n4496), .ZN(n5904) );
  INV_X1 U5284 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4496) );
  OAI211_X1 U5285 ( .C1(n4699), .C2(n4696), .A(n4697), .B(n4695), .ZN(n5044)
         );
  NAND2_X1 U5286 ( .A1(n4698), .A2(n4874), .ZN(n4695) );
  NAND2_X1 U5287 ( .A1(n4871), .A2(n4336), .ZN(n4697) );
  NAND2_X2 U5288 ( .A1(n5333), .A2(n5332), .ZN(n8421) );
  NAND2_X1 U5289 ( .A1(n4816), .A2(n9859), .ZN(n4815) );
  AND2_X1 U5290 ( .A1(n8207), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5291 ( .A1(n5795), .A2(n9854), .ZN(n4817) );
  NAND2_X1 U5292 ( .A1(n6908), .A2(n6909), .ZN(n6907) );
  XNOR2_X1 U5293 ( .A(n4519), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U5294 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4519) );
  INV_X1 U5295 ( .A(n4515), .ZN(n8160) );
  NOR2_X1 U5296 ( .A1(n9869), .A2(n5622), .ZN(n9865) );
  AND2_X1 U5297 ( .A1(n6704), .A2(n6703), .ZN(n9864) );
  OAI21_X1 U5298 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n4530) );
  INV_X1 U5299 ( .A(n7264), .ZN(n7080) );
  AOI21_X1 U5300 ( .B1(n9617), .B2(n4608), .A(n4364), .ZN(n4607) );
  NOR2_X1 U5301 ( .A1(n4614), .A2(n9618), .ZN(n4612) );
  NOR2_X1 U5302 ( .A1(n4617), .A2(n4615), .ZN(n4614) );
  INV_X1 U5303 ( .A(n4618), .ZN(n4615) );
  NAND2_X1 U5304 ( .A1(n4618), .A2(n4619), .ZN(n4616) );
  OAI21_X1 U5305 ( .B1(n9067), .B2(n8637), .A(n6442), .ZN(n6443) );
  AND2_X1 U5306 ( .A1(n8517), .A2(n8518), .ZN(n6364) );
  INV_X1 U5307 ( .A(n7583), .ZN(n7559) );
  INV_X1 U5308 ( .A(n7292), .ZN(n7217) );
  NAND2_X1 U5309 ( .A1(n4576), .A2(n4575), .ZN(n5863) );
  NAND2_X1 U5310 ( .A1(n5816), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4575) );
  INV_X1 U5311 ( .A(n5878), .ZN(n8956) );
  AND2_X1 U5312 ( .A1(n6377), .A2(n6376), .ZN(n9049) );
  OR2_X1 U5313 ( .A1(n9064), .A2(n6425), .ZN(n6377) );
  NAND2_X1 U5314 ( .A1(n6335), .A2(n6334), .ZN(n8962) );
  INV_X1 U5315 ( .A(n7504), .ZN(n8972) );
  NAND2_X1 U5316 ( .A1(n5914), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U5317 ( .A1(n6796), .A2(n4386), .ZN(n6631) );
  NAND2_X1 U5318 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  NAND2_X1 U5319 ( .A1(n9059), .A2(n9061), .ZN(n9277) );
  NAND2_X1 U5320 ( .A1(n4793), .A2(n4796), .ZN(n9060) );
  NAND2_X1 U5321 ( .A1(n4801), .A2(n4799), .ZN(n4793) );
  NAND2_X1 U5322 ( .A1(n4404), .A2(n4403), .ZN(n4402) );
  NAND2_X1 U5323 ( .A1(n9090), .A2(n9232), .ZN(n4403) );
  NAND2_X1 U5324 ( .A1(n9263), .A2(n7224), .ZN(n9260) );
  AND2_X1 U5325 ( .A1(n9203), .A2(n9646), .ZN(n9240) );
  INV_X1 U5326 ( .A(n9268), .ZN(n4466) );
  NAND2_X1 U5327 ( .A1(n9266), .A2(n9790), .ZN(n4430) );
  AOI211_X1 U5328 ( .C1(n5493), .C2(n7570), .A(n5492), .B(n5591), .ZN(n4551)
         );
  INV_X1 U5329 ( .A(n5505), .ZN(n4547) );
  INV_X1 U5330 ( .A(n5503), .ZN(n4549) );
  AOI21_X1 U5331 ( .B1(n4550), .B2(n4548), .A(n4546), .ZN(n5517) );
  NOR2_X1 U5332 ( .A1(n4549), .A2(n8378), .ZN(n4548) );
  NAND2_X1 U5333 ( .A1(n4547), .A2(n5513), .ZN(n4546) );
  OAI21_X1 U5334 ( .B1(n4551), .B2(n5500), .A(n4363), .ZN(n4550) );
  INV_X1 U5335 ( .A(n5511), .ZN(n4561) );
  NAND2_X1 U5336 ( .A1(n5518), .A2(n5570), .ZN(n4560) );
  AOI21_X1 U5337 ( .B1(n8231), .B2(n4413), .A(n5559), .ZN(n4412) );
  INV_X1 U5338 ( .A(n4414), .ZN(n4413) );
  OAI21_X1 U5339 ( .B1(n8244), .B2(n5535), .A(n5433), .ZN(n4414) );
  NAND2_X1 U5340 ( .A1(n5538), .A2(n5537), .ZN(n4544) );
  NOR2_X1 U5341 ( .A1(n8244), .A2(n5536), .ZN(n4543) );
  NAND2_X1 U5342 ( .A1(n5554), .A2(n5553), .ZN(n5557) );
  NOR2_X1 U5343 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  NAND2_X1 U5344 ( .A1(n4541), .A2(n5544), .ZN(n5554) );
  AOI21_X1 U5345 ( .B1(n5557), .B2(n6484), .A(n6475), .ZN(n5558) );
  AOI21_X1 U5346 ( .B1(n5417), .B2(n5561), .A(n4393), .ZN(n4711) );
  AOI21_X1 U5347 ( .B1(n4711), .B2(n4709), .A(n8182), .ZN(n4708) );
  INV_X1 U5348 ( .A(n5561), .ZN(n4709) );
  AND2_X1 U5349 ( .A1(n4474), .A2(n4473), .ZN(n4472) );
  NOR2_X1 U5350 ( .A1(n8453), .A2(n8357), .ZN(n4474) );
  INV_X1 U5351 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U5352 ( .A1(n5419), .A2(SI_30_), .ZN(n4666) );
  NAND2_X1 U5353 ( .A1(n5419), .A2(SI_30_), .ZN(n4665) );
  INV_X1 U5354 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5811) );
  INV_X1 U5355 ( .A(n5201), .ZN(n4669) );
  INV_X1 U5356 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4920) );
  INV_X1 U5357 ( .A(n5144), .ZN(n4678) );
  INV_X1 U5358 ( .A(SI_11_), .ZN(n9429) );
  NAND3_X1 U5359 ( .A1(n5628), .A2(n6972), .A3(n7463), .ZN(n5631) );
  NAND2_X1 U5360 ( .A1(n4540), .A2(n5559), .ZN(n4539) );
  AND2_X1 U5361 ( .A1(n5561), .A2(n4713), .ZN(n4712) );
  INV_X1 U5362 ( .A(n5418), .ZN(n4713) );
  INV_X1 U5363 ( .A(n4708), .ZN(n4707) );
  OR2_X1 U5364 ( .A1(n8196), .A2(n5416), .ZN(n5560) );
  NAND2_X1 U5365 ( .A1(n8207), .A2(n6484), .ZN(n5547) );
  OR2_X1 U5366 ( .A1(n8207), .A2(n6484), .ZN(n5550) );
  NOR2_X1 U5367 ( .A1(n8207), .A2(n4484), .ZN(n4482) );
  OR2_X1 U5368 ( .A1(n8401), .A2(n6474), .ZN(n5545) );
  OR2_X1 U5369 ( .A1(n8406), .A2(n7953), .ZN(n5539) );
  OAI21_X1 U5370 ( .B1(n4740), .B2(n4738), .A(n4370), .ZN(n4737) );
  INV_X1 U5371 ( .A(n5575), .ZN(n4436) );
  INV_X1 U5372 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5192) );
  NOR2_X1 U5373 ( .A1(n4750), .A2(n4747), .ZN(n4746) );
  NAND2_X1 U5374 ( .A1(n4747), .A2(n5158), .ZN(n4718) );
  NAND2_X1 U5375 ( .A1(n8269), .A2(n4486), .ZN(n8237) );
  NAND2_X1 U5376 ( .A1(n8269), .A2(n8479), .ZN(n8250) );
  AND2_X1 U5377 ( .A1(n8368), .A2(n4470), .ZN(n8328) );
  NOR2_X1 U5378 ( .A1(n4471), .A2(n8329), .ZN(n4470) );
  INV_X1 U5379 ( .A(n4472), .ZN(n4471) );
  NAND2_X1 U5380 ( .A1(n8368), .A2(n4474), .ZN(n8355) );
  NOR2_X1 U5381 ( .A1(n4478), .A2(n9638), .ZN(n4477) );
  NOR2_X1 U5382 ( .A1(n7080), .A2(n7111), .ZN(n7182) );
  NAND2_X1 U5383 ( .A1(n4467), .A2(n7152), .ZN(n7111) );
  INV_X1 U5384 ( .A(n9884), .ZN(n4467) );
  OAI21_X1 U5385 ( .B1(n5784), .B2(n5783), .A(n9943), .ZN(n6489) );
  INV_X1 U5386 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4997) );
  INV_X1 U5387 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5118) );
  INV_X1 U5388 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4854) );
  INV_X1 U5389 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4838) );
  INV_X1 U5390 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5216) );
  INV_X1 U5391 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4858) );
  INV_X1 U5392 ( .A(n5081), .ZN(n4839) );
  INV_X1 U5393 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5230) );
  NOR2_X1 U5394 ( .A1(n5146), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5162) );
  OR2_X1 U5395 ( .A1(n5133), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U5396 ( .A1(n4642), .A2(n4641), .ZN(n8657) );
  NAND2_X1 U5397 ( .A1(n9072), .A2(n8781), .ZN(n4641) );
  OR2_X1 U5398 ( .A1(n8782), .A2(n4375), .ZN(n4642) );
  NOR2_X1 U5399 ( .A1(n9675), .A2(n4508), .ZN(n8982) );
  NOR2_X1 U5400 ( .A1(n4510), .A2(n4509), .ZN(n4508) );
  INV_X1 U5401 ( .A(n9674), .ZN(n4510) );
  OR2_X1 U5402 ( .A1(n9271), .A2(n9049), .ZN(n8832) );
  INV_X1 U5403 ( .A(n4788), .ZN(n4786) );
  NOR2_X1 U5404 ( .A1(n4804), .A2(n4802), .ZN(n4428) );
  NOR2_X1 U5405 ( .A1(n7753), .A2(n4803), .ZN(n4802) );
  INV_X1 U5406 ( .A(n7627), .ZN(n4803) );
  INV_X1 U5407 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6098) );
  INV_X1 U5408 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6060) );
  NOR2_X1 U5409 ( .A1(n7511), .A2(n4451), .ZN(n4453) );
  NAND2_X1 U5410 ( .A1(n4452), .A2(n9660), .ZN(n4451) );
  NOR2_X1 U5411 ( .A1(n7613), .A2(n7535), .ZN(n4452) );
  INV_X1 U5412 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6040) );
  INV_X1 U5413 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6021) );
  OR2_X1 U5414 ( .A1(n6022), .A2(n6021), .ZN(n6041) );
  OR2_X1 U5415 ( .A1(n7558), .A2(n7559), .ZN(n7511) );
  NAND2_X1 U5416 ( .A1(n7047), .A2(n4407), .ZN(n8922) );
  NAND2_X1 U5417 ( .A1(n7046), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U5418 ( .A1(n6385), .A2(n8956), .ZN(n7030) );
  AOI21_X1 U5419 ( .B1(n4689), .B2(n4691), .A(n4397), .ZN(n4686) );
  INV_X1 U5420 ( .A(n5343), .ZN(n4692) );
  OAI21_X1 U5421 ( .B1(n5287), .B2(n5286), .A(n4948), .ZN(n5296) );
  AND2_X1 U5422 ( .A1(n4952), .A2(n4951), .ZN(n5295) );
  INV_X1 U5423 ( .A(n4646), .ZN(n4645) );
  OAI21_X1 U5424 ( .B1(n4649), .B2(n4647), .A(n4939), .ZN(n4646) );
  INV_X1 U5425 ( .A(n4914), .ZN(n4672) );
  INV_X1 U5426 ( .A(n5959), .ZN(n4405) );
  NOR2_X1 U5427 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4563) );
  INV_X1 U5428 ( .A(n4886), .ZN(n4555) );
  OAI21_X1 U5429 ( .B1(n5079), .B2(n4555), .A(n5091), .ZN(n4553) );
  INV_X1 U5430 ( .A(SI_13_), .ZN(n9469) );
  INV_X1 U5431 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9481) );
  INV_X1 U5432 ( .A(SI_16_), .ZN(n9525) );
  INV_X1 U5433 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9441) );
  OR2_X1 U5434 ( .A1(n7657), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U5435 ( .A1(n4836), .A2(n5700), .ZN(n4833) );
  INV_X1 U5436 ( .A(n5700), .ZN(n4835) );
  NAND2_X1 U5437 ( .A1(n9637), .A2(n9636), .ZN(n9635) );
  OR2_X1 U5438 ( .A1(n5347), .A2(n9504), .ZN(n5359) );
  AND2_X1 U5439 ( .A1(n7125), .A2(n5667), .ZN(n4832) );
  NAND2_X1 U5440 ( .A1(n7700), .A2(n4837), .ZN(n4836) );
  INV_X1 U5441 ( .A(n4853), .ZN(n4837) );
  NOR2_X1 U5442 ( .A1(n5193), .A2(n5192), .ZN(n5207) );
  OR2_X1 U5443 ( .A1(n5180), .A2(n9816), .ZN(n5193) );
  NOR2_X1 U5444 ( .A1(n5801), .A2(n5800), .ZN(n6488) );
  INV_X1 U5445 ( .A(n8080), .ZN(n8065) );
  NOR2_X1 U5446 ( .A1(n5793), .A2(n9944), .ZN(n5796) );
  OR2_X1 U5447 ( .A1(n5221), .A2(n9441), .ZN(n5237) );
  NAND2_X1 U5448 ( .A1(n5236), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5252) );
  INV_X1 U5449 ( .A(n5237), .ZN(n5236) );
  NAND2_X1 U5450 ( .A1(n8107), .A2(n8106), .ZN(n8105) );
  OR2_X1 U5451 ( .A1(n6818), .A2(n6817), .ZN(n4523) );
  OR2_X1 U5452 ( .A1(n6841), .A2(n6840), .ZN(n4521) );
  OR3_X1 U5453 ( .A1(n5188), .A2(P2_IR_REG_10__SCAN_IN), .A3(
        P2_IR_REG_11__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U5454 ( .A1(n8132), .A2(n8133), .ZN(n8131) );
  NOR2_X1 U5455 ( .A1(n7351), .A2(n4525), .ZN(n7355) );
  AND2_X1 U5456 ( .A1(n7352), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5457 ( .A1(n7355), .A2(n7354), .ZN(n7451) );
  NAND2_X1 U5458 ( .A1(n7451), .A2(n4524), .ZN(n7453) );
  OR2_X1 U5459 ( .A1(n7452), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5460 ( .A1(n7453), .A2(n7454), .ZN(n7643) );
  XNOR2_X1 U5461 ( .A(n4515), .B(n8165), .ZN(n8153) );
  OR2_X1 U5462 ( .A1(n8149), .A2(n4516), .ZN(n4515) );
  NOR2_X1 U5463 ( .A1(n8145), .A2(n4517), .ZN(n4516) );
  INV_X1 U5464 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n4517) );
  NOR2_X1 U5465 ( .A1(n8182), .A2(n8181), .ZN(n8185) );
  AND2_X1 U5466 ( .A1(n5550), .A2(n5547), .ZN(n8204) );
  NAND2_X1 U5467 ( .A1(n5545), .A2(n5546), .ZN(n8216) );
  AND2_X1 U5468 ( .A1(n5395), .A2(n5371), .ZN(n8070) );
  NAND2_X1 U5469 ( .A1(n4693), .A2(n5378), .ZN(n8230) );
  INV_X1 U5470 ( .A(n8231), .ZN(n8228) );
  AOI21_X1 U5471 ( .B1(n4330), .B2(n4558), .A(n4439), .ZN(n4438) );
  INV_X1 U5472 ( .A(n5532), .ZN(n4439) );
  INV_X1 U5473 ( .A(n8244), .ZN(n8247) );
  AND2_X1 U5474 ( .A1(n8283), .A2(n4756), .ZN(n8269) );
  NOR2_X1 U5475 ( .A1(n8300), .A2(n8421), .ZN(n8283) );
  NAND2_X1 U5476 ( .A1(n5320), .A2(n5319), .ZN(n8299) );
  OR2_X1 U5477 ( .A1(n5309), .A2(n5308), .ZN(n5322) );
  OR2_X1 U5478 ( .A1(n8443), .A2(n8086), .ZN(n6470) );
  NAND2_X1 U5479 ( .A1(n8368), .A2(n8375), .ZN(n8369) );
  OAI22_X1 U5480 ( .A1(n7521), .A2(n4432), .B1(n4434), .B2(n5213), .ZN(n7675)
         );
  OR2_X1 U5481 ( .A1(n5213), .A2(n4436), .ZN(n4432) );
  INV_X1 U5482 ( .A(n4435), .ZN(n4434) );
  OAI21_X1 U5483 ( .B1(n5483), .B2(n4436), .A(n7570), .ZN(n4435) );
  NAND2_X1 U5484 ( .A1(n7675), .A2(n7674), .ZN(n7673) );
  OR2_X1 U5485 ( .A1(n7595), .A2(n9877), .ZN(n7596) );
  AND2_X1 U5486 ( .A1(n9995), .A2(n7182), .ZN(n7321) );
  NAND2_X1 U5487 ( .A1(n7321), .A2(n7327), .ZN(n7595) );
  OR2_X1 U5488 ( .A1(n5137), .A2(n9471), .ZN(n5151) );
  OR2_X1 U5489 ( .A1(n10004), .A2(n7343), .ZN(n6969) );
  NAND2_X1 U5490 ( .A1(n5100), .A2(n9887), .ZN(n9891) );
  NOR2_X1 U5491 ( .A1(n9912), .A2(n9811), .ZN(n9886) );
  NAND3_X1 U5492 ( .A1(n9924), .A2(n9968), .A3(n9973), .ZN(n9912) );
  NAND2_X1 U5493 ( .A1(n9924), .A2(n9968), .ZN(n9925) );
  NAND2_X1 U5494 ( .A1(n5206), .A2(n5205), .ZN(n7575) );
  INV_X1 U5495 ( .A(n10008), .ZN(n9962) );
  INV_X1 U5496 ( .A(n10002), .ZN(n9987) );
  XNOR2_X1 U5497 ( .A(n5613), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6507) );
  OR2_X1 U5498 ( .A1(n5801), .A2(P2_U3152), .ZN(n9944) );
  NOR2_X1 U5499 ( .A1(n4362), .A2(n4828), .ZN(n4827) );
  AND2_X1 U5500 ( .A1(n5176), .A2(n5165), .ZN(n7189) );
  INV_X1 U5501 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5984) );
  NOR2_X1 U5502 ( .A1(n5985), .A2(n5984), .ZN(n6002) );
  INV_X1 U5503 ( .A(n6094), .ZN(n4609) );
  NAND2_X1 U5504 ( .A1(n8566), .A2(n6172), .ZN(n8575) );
  NAND2_X1 U5505 ( .A1(n6156), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6180) );
  AOI22_X1 U5506 ( .A1(n6292), .A2(n8528), .B1(n6291), .B2(n8529), .ZN(n8585)
         );
  NAND2_X1 U5507 ( .A1(n7247), .A2(n7248), .ZN(n4637) );
  OR2_X1 U5508 ( .A1(n7247), .A2(n7248), .ZN(n4638) );
  AOI22_X1 U5509 ( .A1(n7270), .A2(n4316), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5877), .ZN(n5882) );
  NAND2_X1 U5510 ( .A1(n4624), .A2(n4628), .ZN(n8593) );
  NAND2_X1 U5511 ( .A1(n6210), .A2(n4630), .ZN(n4624) );
  INV_X1 U5512 ( .A(n9616), .ZN(n4610) );
  NAND2_X1 U5513 ( .A1(n7487), .A2(n7485), .ZN(n4633) );
  NOR2_X1 U5514 ( .A1(n6210), .A2(n6211), .ZN(n8614) );
  OR2_X1 U5515 ( .A1(n6180), .A2(n6179), .ZN(n6200) );
  NAND2_X1 U5516 ( .A1(n6948), .A2(n4622), .ZN(n4621) );
  INV_X1 U5517 ( .A(n5934), .ZN(n4620) );
  NAND2_X1 U5518 ( .A1(n4808), .A2(n5816), .ZN(n4807) );
  INV_X1 U5519 ( .A(n4810), .ZN(n4808) );
  OAI21_X1 U5520 ( .B1(n4577), .B2(n5860), .A(P1_IR_REG_27__SCAN_IN), .ZN(
        n4576) );
  NOR2_X1 U5521 ( .A1(n6411), .A2(n4810), .ZN(n4577) );
  AND2_X1 U5522 ( .A1(n9626), .A2(n9027), .ZN(n8905) );
  AND2_X1 U5523 ( .A1(n6352), .A2(n6351), .ZN(n8631) );
  OR2_X1 U5524 ( .A1(n6679), .A2(n6678), .ZN(n4489) );
  NAND2_X1 U5525 ( .A1(n4507), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5526 ( .A1(n6661), .A2(n4348), .ZN(n4505) );
  NOR2_X1 U5527 ( .A1(n6691), .A2(n6690), .ZN(n6723) );
  NOR2_X1 U5528 ( .A1(n8979), .A2(n4511), .ZN(n9676) );
  AND2_X1 U5529 ( .A1(n8992), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4511) );
  NOR2_X1 U5530 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  XNOR2_X1 U5531 ( .A(n8982), .B(n9002), .ZN(n9692) );
  NOR2_X1 U5532 ( .A1(n9062), .A2(n9267), .ZN(n9050) );
  NAND2_X1 U5533 ( .A1(n4460), .A2(n4459), .ZN(n4458) );
  INV_X1 U5534 ( .A(n4461), .ZN(n4460) );
  NOR2_X1 U5535 ( .A1(n9283), .A2(n9271), .ZN(n4459) );
  NAND2_X1 U5536 ( .A1(n9091), .A2(n9232), .ZN(n9074) );
  NAND2_X1 U5537 ( .A1(n9035), .A2(n4798), .ZN(n4797) );
  INV_X1 U5538 ( .A(n4849), .ZN(n4798) );
  NAND2_X1 U5539 ( .A1(n8832), .A2(n9042), .ZN(n9070) );
  OR2_X1 U5540 ( .A1(n6328), .A2(n8629), .ZN(n6368) );
  NAND2_X1 U5541 ( .A1(n4598), .A2(n4596), .ZN(n7924) );
  INV_X1 U5542 ( .A(n4597), .ZN(n4596) );
  OAI22_X1 U5543 ( .A1(n4601), .A2(n4605), .B1(n8935), .B2(n8896), .ZN(n4597)
         );
  NAND2_X1 U5544 ( .A1(n9091), .A2(n9234), .ZN(n4404) );
  OR2_X1 U5545 ( .A1(n9126), .A2(n9295), .ZN(n9117) );
  NOR2_X1 U5546 ( .A1(n9117), .A2(n9290), .ZN(n9099) );
  NAND2_X1 U5547 ( .A1(n4374), .A2(n4423), .ZN(n4418) );
  NAND2_X1 U5548 ( .A1(n9178), .A2(n4358), .ZN(n4419) );
  OR2_X1 U5549 ( .A1(n6248), .A2(n6247), .ZN(n6267) );
  INV_X1 U5550 ( .A(n8963), .ZN(n9153) );
  NAND2_X1 U5551 ( .A1(n9164), .A2(n8557), .ZN(n9165) );
  AND2_X1 U5552 ( .A1(n6265), .A2(n6264), .ZN(n9144) );
  AOI21_X1 U5553 ( .B1(n4581), .B2(n4583), .A(n4580), .ZN(n4579) );
  NAND2_X1 U5554 ( .A1(n6198), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6216) );
  INV_X1 U5555 ( .A(n6200), .ZN(n6198) );
  OAI21_X1 U5556 ( .B1(n4424), .B2(n4773), .A(n4770), .ZN(n9192) );
  AOI21_X1 U5557 ( .B1(n4772), .B2(n4774), .A(n4388), .ZN(n4770) );
  AND2_X1 U5558 ( .A1(n7866), .A2(n4454), .ZN(n9213) );
  AND2_X1 U5559 ( .A1(n4333), .A2(n9216), .ZN(n4454) );
  NAND2_X1 U5560 ( .A1(n7866), .A2(n4456), .ZN(n9251) );
  NAND2_X1 U5561 ( .A1(n7866), .A2(n7916), .ZN(n9253) );
  AND2_X1 U5562 ( .A1(n7777), .A2(n8712), .ZN(n7866) );
  OR2_X1 U5563 ( .A1(n8883), .A2(n8714), .ZN(n8818) );
  OR2_X1 U5564 ( .A1(n6099), .A2(n6098), .ZN(n6114) );
  NAND2_X1 U5565 ( .A1(n6113), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6136) );
  INV_X1 U5566 ( .A(n6114), .ZN(n6113) );
  NAND2_X1 U5567 ( .A1(n4453), .A2(n9614), .ZN(n7776) );
  AND2_X1 U5568 ( .A1(n8690), .A2(n8876), .ZN(n8815) );
  NAND2_X1 U5569 ( .A1(n7755), .A2(n7754), .ZN(n7779) );
  NAND2_X1 U5570 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  NAND2_X1 U5571 ( .A1(n7629), .A2(n7633), .ZN(n7755) );
  INV_X1 U5572 ( .A(n4453), .ZN(n7636) );
  AND4_X1 U5573 ( .A1(n6086), .A2(n6085), .A3(n6084), .A4(n6083), .ZN(n7782)
         );
  AOI21_X1 U5574 ( .B1(n7614), .B2(n8807), .A(n4382), .ZN(n7616) );
  OAI211_X1 U5575 ( .C1(n4593), .C2(n4329), .A(n4590), .B(n8840), .ZN(n7632)
         );
  OR2_X1 U5576 ( .A1(n4329), .A2(n4406), .ZN(n4590) );
  NOR2_X1 U5577 ( .A1(n7511), .A2(n4450), .ZN(n7611) );
  INV_X1 U5578 ( .A(n4452), .ZN(n4450) );
  NOR2_X1 U5579 ( .A1(n7511), .A2(n7535), .ZN(n7546) );
  NAND2_X1 U5580 ( .A1(n4592), .A2(n8681), .ZN(n7617) );
  NAND2_X1 U5581 ( .A1(n4593), .A2(n4406), .ZN(n4592) );
  AND2_X1 U5582 ( .A1(n4416), .A2(n4392), .ZN(n4415) );
  OR2_X1 U5583 ( .A1(n4806), .A2(n7395), .ZN(n4417) );
  AND4_X1 U5584 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(n7510)
         );
  AND3_X1 U5585 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5586 ( .A1(n4449), .A2(n9768), .ZN(n7274) );
  INV_X1 U5587 ( .A(n7208), .ZN(n4449) );
  OR2_X1 U5588 ( .A1(n7298), .A2(n7292), .ZN(n7208) );
  NAND2_X1 U5589 ( .A1(n7296), .A2(n9761), .ZN(n7298) );
  NOR2_X1 U5590 ( .A1(n5907), .A2(n7052), .ZN(n7296) );
  AND2_X1 U5591 ( .A1(n7043), .A2(n7042), .ZN(n7045) );
  NOR2_X1 U5592 ( .A1(n6744), .A2(n7034), .ZN(n7046) );
  AND2_X1 U5593 ( .A1(n6744), .A2(n7270), .ZN(n7029) );
  NAND2_X1 U5594 ( .A1(n6432), .A2(n7098), .ZN(n6772) );
  NAND2_X1 U5595 ( .A1(n6345), .A2(n6344), .ZN(n9280) );
  AOI21_X1 U5596 ( .B1(n6386), .B2(n7100), .A(n7096), .ZN(n6773) );
  OR2_X1 U5597 ( .A1(n7033), .A2(n8911), .ZN(n9786) );
  INV_X1 U5598 ( .A(n9347), .ZN(n9784) );
  INV_X1 U5599 ( .A(n7032), .ZN(n7101) );
  AND2_X1 U5600 ( .A1(n6387), .A2(n8949), .ZN(n9347) );
  AND2_X1 U5601 ( .A1(n6394), .A2(n6393), .ZN(n6768) );
  NAND3_X1 U5602 ( .A1(n4657), .A2(n4656), .A3(n4658), .ZN(n8654) );
  OAI21_X1 U5603 ( .B1(n4660), .B2(n5423), .A(n4659), .ZN(n4658) );
  OR2_X1 U5604 ( .A1(n5420), .A2(n4663), .ZN(n4657) );
  XNOR2_X1 U5605 ( .A(n5420), .B(n4996), .ZN(n8646) );
  XNOR2_X1 U5606 ( .A(n5404), .B(n5405), .ZN(n8638) );
  XNOR2_X1 U5607 ( .A(n5391), .B(n5390), .ZN(n8506) );
  NAND2_X1 U5608 ( .A1(n4688), .A2(n4988), .ZN(n5391) );
  XNOR2_X1 U5609 ( .A(n5379), .B(n5380), .ZN(n8509) );
  XNOR2_X1 U5610 ( .A(n5367), .B(n5366), .ZN(n7857) );
  NAND2_X1 U5611 ( .A1(n5843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  INV_X1 U5612 ( .A(n4811), .ZN(n4809) );
  INV_X1 U5613 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5845) );
  OAI21_X1 U5614 ( .B1(n5229), .B2(n4653), .A(n4650), .ZN(n5259) );
  AND2_X1 U5615 ( .A1(n5833), .A2(n5834), .ZN(n6110) );
  NAND2_X1 U5616 ( .A1(n4673), .A2(n4914), .ZN(n5187) );
  NAND2_X1 U5617 ( .A1(n4912), .A2(n4674), .ZN(n4673) );
  AND2_X1 U5618 ( .A1(n6018), .A2(n6056), .ZN(n6688) );
  OAI21_X1 U5619 ( .B1(n5116), .B2(n4682), .A(n4679), .ZN(n5145) );
  NAND2_X1 U5620 ( .A1(n4640), .A2(n5038), .ZN(n4875) );
  NAND2_X1 U5621 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5923) );
  INV_X1 U5622 ( .A(n5904), .ZN(n4495) );
  XNOR2_X1 U5623 ( .A(n5888), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6553) );
  CLKBUF_X1 U5624 ( .A(n7124), .Z(n7230) );
  NOR2_X1 U5625 ( .A1(n7421), .A2(n4831), .ZN(n4830) );
  INV_X1 U5626 ( .A(n5683), .ZN(n4831) );
  NAND2_X1 U5627 ( .A1(n7415), .A2(n5683), .ZN(n7422) );
  INV_X1 U5628 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9471) );
  NOR2_X1 U5629 ( .A1(n9826), .A2(n7657), .ZN(n7656) );
  INV_X1 U5630 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U5631 ( .B1(n5744), .B2(n4332), .A(n5749), .ZN(n4819) );
  INV_X1 U5632 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U5633 ( .A1(n9808), .A2(n4359), .ZN(n7016) );
  AND2_X1 U5634 ( .A1(n9808), .A2(n5655), .ZN(n7018) );
  AND2_X1 U5635 ( .A1(n5717), .A2(n5711), .ZN(n4843) );
  NAND2_X1 U5636 ( .A1(n5712), .A2(n5711), .ZN(n7893) );
  NOR2_X1 U5637 ( .A1(n4824), .A2(n4823), .ZN(n8016) );
  NAND2_X1 U5638 ( .A1(n6940), .A2(n4841), .ZN(n9808) );
  AND2_X1 U5639 ( .A1(n9809), .A2(n5651), .ZN(n4841) );
  AND2_X1 U5640 ( .A1(n6940), .A2(n5651), .ZN(n9810) );
  AND2_X1 U5641 ( .A1(n5734), .A2(n5729), .ZN(n4842) );
  INV_X1 U5642 ( .A(n8028), .ZN(n5734) );
  NAND2_X1 U5643 ( .A1(n7976), .A2(n5729), .ZN(n8029) );
  NOR2_X1 U5644 ( .A1(n7656), .A2(n4853), .ZN(n7701) );
  OR2_X1 U5645 ( .A1(n7656), .A2(n4836), .ZN(n7699) );
  NAND2_X1 U5646 ( .A1(n6907), .A2(n5636), .ZN(n9839) );
  INV_X1 U5647 ( .A(n9863), .ZN(n8046) );
  NAND2_X1 U5648 ( .A1(n4534), .A2(n4334), .ZN(n5606) );
  NAND2_X1 U5649 ( .A1(n4714), .A2(n5571), .ZN(n5430) );
  OR2_X1 U5650 ( .A1(n5797), .A2(n5408), .ZN(n5403) );
  NAND4_X1 U5651 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n8102)
         );
  INV_X2 U5652 ( .A(P2_U3966), .ZN(n8103) );
  NAND2_X1 U5653 ( .A1(n6713), .A2(n6714), .ZN(n6810) );
  NOR2_X1 U5654 ( .A1(n6881), .A2(n6880), .ZN(n6879) );
  AND2_X1 U5655 ( .A1(n6810), .A2(n4528), .ZN(n6881) );
  NAND2_X1 U5656 ( .A1(n6824), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4528) );
  INV_X1 U5657 ( .A(n4523), .ZN(n6838) );
  AND2_X1 U5658 ( .A1(n4523), .A2(n4522), .ZN(n6841) );
  NAND2_X1 U5659 ( .A1(n6843), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4522) );
  INV_X1 U5660 ( .A(n4521), .ZN(n6853) );
  AND2_X1 U5661 ( .A1(n4521), .A2(n4520), .ZN(n6857) );
  NAND2_X1 U5662 ( .A1(n6854), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4520) );
  NOR2_X1 U5663 ( .A1(n6920), .A2(n4527), .ZN(n6924) );
  AND2_X1 U5664 ( .A1(n6921), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5665 ( .A1(n6924), .A2(n6923), .ZN(n7188) );
  NOR2_X1 U5666 ( .A1(n7876), .A2(n4518), .ZN(n7881) );
  AND2_X1 U5667 ( .A1(n7877), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4518) );
  NOR2_X1 U5668 ( .A1(n7881), .A2(n7880), .ZN(n8149) );
  INV_X1 U5669 ( .A(n9865), .ZN(n7879) );
  NAND2_X1 U5670 ( .A1(n4755), .A2(n4328), .ZN(n8266) );
  NAND2_X1 U5671 ( .A1(n4440), .A2(n4330), .ZN(n8261) );
  AND2_X1 U5672 ( .A1(n4440), .A2(n5512), .ZN(n8263) );
  NAND2_X1 U5673 ( .A1(n4727), .A2(n4726), .ZN(n8294) );
  NAND2_X1 U5674 ( .A1(n4727), .A2(n5518), .ZN(n8292) );
  INV_X1 U5675 ( .A(n8433), .ZN(n8318) );
  NAND2_X1 U5676 ( .A1(n4720), .A2(n5515), .ZN(n8323) );
  AND2_X1 U5677 ( .A1(n4744), .A2(n4354), .ZN(n8336) );
  NAND2_X1 U5678 ( .A1(n8347), .A2(n6469), .ZN(n4744) );
  NAND2_X1 U5679 ( .A1(n7829), .A2(n5501), .ZN(n8377) );
  AND2_X1 U5680 ( .A1(n4764), .A2(n4341), .ZN(n8366) );
  NAND2_X1 U5681 ( .A1(n5251), .A2(n5250), .ZN(n8459) );
  NAND2_X1 U5682 ( .A1(n7736), .A2(n5497), .ZN(n7831) );
  NAND2_X1 U5683 ( .A1(n7733), .A2(n4765), .ZN(n7826) );
  NAND2_X1 U5684 ( .A1(n4433), .A2(n5575), .ZN(n7569) );
  NAND2_X1 U5685 ( .A1(n7521), .A2(n5483), .ZN(n4433) );
  NAND2_X1 U5686 ( .A1(n7598), .A2(n5473), .ZN(n7434) );
  NAND2_X1 U5687 ( .A1(n7591), .A2(n6465), .ZN(n7433) );
  AND2_X1 U5688 ( .A1(n4719), .A2(n5158), .ZN(n7599) );
  NOR2_X1 U5689 ( .A1(n7170), .A2(n4851), .ZN(n7313) );
  AND2_X1 U5690 ( .A1(n7069), .A2(n5463), .ZN(n4844) );
  INV_X1 U5691 ( .A(n9931), .ZN(n8374) );
  NAND2_X1 U5692 ( .A1(n4731), .A2(n6458), .ZN(n7110) );
  NAND2_X1 U5693 ( .A1(n4734), .A2(n4733), .ZN(n4731) );
  INV_X1 U5694 ( .A(n4732), .ZN(n4733) );
  NAND2_X1 U5695 ( .A1(n4734), .A2(n6457), .ZN(n9883) );
  AND2_X1 U5696 ( .A1(n9938), .A2(n9900), .ZN(n9934) );
  OR2_X1 U5697 ( .A1(n6700), .A2(n5045), .ZN(n5046) );
  INV_X1 U5698 ( .A(n8192), .ZN(n9929) );
  AND2_X2 U5699 ( .A1(n6968), .A2(n6490), .ZN(n10026) );
  INV_X1 U5700 ( .A(n8175), .ZN(n8465) );
  NAND2_X1 U5701 ( .A1(n8199), .A2(n4447), .ZN(n4446) );
  INV_X1 U5702 ( .A(n8193), .ZN(n4448) );
  INV_X1 U5703 ( .A(n7575), .ZN(n7732) );
  NAND2_X1 U5704 ( .A1(n6596), .A2(n5424), .ZN(n5179) );
  OR2_X1 U5705 ( .A1(n6561), .A2(n5117), .ZN(n4728) );
  AND2_X2 U5706 ( .A1(n6968), .A2(n6496), .ZN(n10012) );
  NOR2_X1 U5707 ( .A1(P2_U3152), .A2(n6507), .ZN(n9949) );
  INV_X1 U5708 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8498) );
  INV_X1 U5709 ( .A(n5786), .ZN(n7858) );
  XNOR2_X1 U5710 ( .A(n5615), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U5711 ( .A1(n5614), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5615) );
  INV_X1 U5712 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5612) );
  INV_X1 U5713 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7946) );
  CLKBUF_X1 U5714 ( .A(n5572), .Z(n7944) );
  INV_X1 U5715 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7432) );
  INV_X1 U5716 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7344) );
  INV_X1 U5717 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7067) );
  INV_X1 U5718 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6960) );
  INV_X1 U5719 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6734) );
  INV_X1 U5720 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6670) );
  NOR2_X1 U5721 ( .A1(n6539), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8510) );
  INV_X1 U5722 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6579) );
  INV_X1 U5723 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6570) );
  NOR2_X1 U5724 ( .A1(n6504), .A2(n6503), .ZN(n6535) );
  INV_X1 U5725 ( .A(n8962), .ZN(n9108) );
  INV_X1 U5726 ( .A(n8965), .ZN(n9247) );
  NAND2_X1 U5727 ( .A1(n6112), .A2(n6111), .ZN(n9346) );
  NAND2_X1 U5728 ( .A1(n6278), .A2(n6277), .ZN(n9298) );
  AND2_X1 U5730 ( .A1(n6273), .A2(n6272), .ZN(n8553) );
  AND4_X1 U5731 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n9612)
         );
  NAND2_X1 U5732 ( .A1(n6948), .A2(n5934), .ZN(n4623) );
  AND4_X1 U5733 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n7618)
         );
  AND2_X1 U5734 ( .A1(n6424), .A2(n6423), .ZN(n9608) );
  OAI21_X1 U5735 ( .B1(n4628), .B2(n4627), .A(n4626), .ZN(n4625) );
  INV_X1 U5736 ( .A(n8592), .ZN(n4627) );
  NAND2_X1 U5737 ( .A1(n9615), .A2(n6094), .ZN(n7715) );
  INV_X1 U5738 ( .A(n9144), .ZN(n9305) );
  NAND2_X1 U5739 ( .A1(n4633), .A2(n7484), .ZN(n7693) );
  INV_X1 U5740 ( .A(n9222), .ZN(n9249) );
  NAND2_X1 U5741 ( .A1(n9621), .A2(n9347), .ZN(n8637) );
  INV_X1 U5742 ( .A(n9625), .ZN(n8634) );
  INV_X1 U5743 ( .A(n8966), .ZN(n8703) );
  OR2_X1 U5744 ( .A1(n6439), .A2(n6423), .ZN(n9611) );
  INV_X1 U5745 ( .A(n8637), .ZN(n8611) );
  INV_X1 U5746 ( .A(n8631), .ZN(n9091) );
  INV_X1 U5747 ( .A(n9116), .ZN(n9090) );
  INV_X1 U5748 ( .A(n8553), .ZN(n9161) );
  INV_X1 U5749 ( .A(n9182), .ZN(n9221) );
  INV_X1 U5750 ( .A(n7510), .ZN(n8971) );
  INV_X1 U5751 ( .A(n7303), .ZN(n8977) );
  INV_X1 U5752 ( .A(n4489), .ZN(n6677) );
  NAND2_X1 U5753 ( .A1(n6798), .A2(n6797), .ZN(n6796) );
  AND2_X1 U5754 ( .A1(n4489), .A2(n4488), .ZN(n6798) );
  NAND2_X1 U5755 ( .A1(n6525), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5756 ( .A1(n6661), .A2(n4506), .ZN(n6617) );
  AND2_X1 U5757 ( .A1(n4505), .A2(n4504), .ZN(n6604) );
  NAND2_X1 U5758 ( .A1(n4498), .A2(n4497), .ZN(n6515) );
  AOI21_X1 U5759 ( .B1(n4499), .B2(n4502), .A(n4387), .ZN(n4497) );
  NOR2_X1 U5760 ( .A1(n6723), .A2(n4512), .ZN(n6725) );
  AND2_X1 U5761 ( .A1(n6724), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5762 ( .A1(n6725), .A2(n6726), .ZN(n6995) );
  INV_X1 U5763 ( .A(n4493), .ZN(n9703) );
  INV_X1 U5764 ( .A(n8985), .ZN(n4492) );
  XNOR2_X1 U5765 ( .A(n4513), .B(n8991), .ZN(n9015) );
  OR2_X1 U5766 ( .A1(n9742), .A2(n4514), .ZN(n4513) );
  AND2_X1 U5767 ( .A1(n9747), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4514) );
  AND2_X1 U5768 ( .A1(n6518), .A2(n6517), .ZN(n9736) );
  NAND2_X1 U5769 ( .A1(n8656), .A2(n8655), .ZN(n9626) );
  MUX2_X1 U5770 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8654), .S(n4401), .Z(n8656) );
  INV_X1 U5771 ( .A(n9031), .ZN(n9644) );
  INV_X1 U5772 ( .A(n4570), .ZN(n4569) );
  OAI22_X1 U5773 ( .A1(n9049), .A2(n9248), .B1(n9048), .B2(n9047), .ZN(n4570)
         );
  NAND2_X1 U5774 ( .A1(n9271), .A2(n9037), .ZN(n9038) );
  AOI21_X1 U5775 ( .B1(n4801), .B2(n4850), .A(n4849), .ZN(n9036) );
  AND2_X1 U5776 ( .A1(n6294), .A2(n6293), .ZN(n9122) );
  OAI21_X1 U5777 ( .B1(n9172), .B2(n4783), .A(n4781), .ZN(n9111) );
  NAND2_X1 U5778 ( .A1(n4784), .A2(n4787), .ZN(n9125) );
  NAND2_X1 U5779 ( .A1(n9172), .A2(n4788), .ZN(n4784) );
  NAND2_X1 U5780 ( .A1(n9172), .A2(n4845), .ZN(n9142) );
  AND2_X1 U5781 ( .A1(n4422), .A2(n4349), .ZN(n9171) );
  NAND2_X1 U5782 ( .A1(n6246), .A2(n6245), .ZN(n9310) );
  OAI21_X1 U5783 ( .B1(n9218), .B2(n4583), .A(n4581), .ZN(n9180) );
  AND2_X1 U5784 ( .A1(n6213), .A2(n6212), .ZN(n9208) );
  AOI21_X1 U5785 ( .B1(n9218), .B2(n8867), .A(n7923), .ZN(n9195) );
  NAND2_X1 U5786 ( .A1(n4771), .A2(n4775), .ZN(n9212) );
  OAI21_X1 U5787 ( .B1(n9242), .B2(n4774), .A(n4772), .ZN(n9211) );
  NAND2_X1 U5788 ( .A1(n9242), .A2(n4347), .ZN(n4771) );
  INV_X1 U5789 ( .A(n4779), .ZN(n4776) );
  NAND2_X1 U5790 ( .A1(n9242), .A2(n9243), .ZN(n4777) );
  NAND2_X1 U5791 ( .A1(n6155), .A2(n6154), .ZN(n9336) );
  INV_X1 U5792 ( .A(n9346), .ZN(n8712) );
  NAND2_X1 U5793 ( .A1(n6097), .A2(n6096), .ZN(n8707) );
  INV_X1 U5794 ( .A(n6010), .ZN(n4429) );
  NAND2_X1 U5795 ( .A1(n4406), .A2(n8839), .ZN(n7555) );
  NAND2_X1 U5796 ( .A1(n7506), .A2(n4805), .ZN(n7553) );
  OR2_X1 U5797 ( .A1(n5943), .A2(n6557), .ZN(n5962) );
  NAND2_X1 U5798 ( .A1(n7219), .A2(n7218), .ZN(n7221) );
  NAND2_X1 U5799 ( .A1(n7100), .A2(n7099), .ZN(n9145) );
  INV_X1 U5800 ( .A(n9145), .ZN(n9255) );
  INV_X1 U5801 ( .A(n9273), .ZN(n9274) );
  NAND2_X1 U5802 ( .A1(n5824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5821) );
  INV_X1 U5803 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7610) );
  INV_X1 U5804 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5869) );
  INV_X1 U5805 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7445) );
  NAND2_X1 U5806 ( .A1(n5873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5842) );
  INV_X1 U5807 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7346) );
  INV_X1 U5808 ( .A(n9018), .ZN(n9168) );
  AND2_X1 U5809 ( .A1(n6176), .A2(n6194), .ZN(n9731) );
  INV_X1 U5810 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6668) );
  INV_X1 U5811 ( .A(n6996), .ZN(n6990) );
  INV_X1 U5812 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6593) );
  INV_X1 U5813 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U5814 ( .A1(n4554), .A2(n4886), .ZN(n5092) );
  XNOR2_X1 U5815 ( .A(n5080), .B(n5079), .ZN(n6551) );
  AND2_X1 U5816 ( .A1(n5807), .A2(n5904), .ZN(n5940) );
  XNOR2_X1 U5817 ( .A(n5923), .B(n5922), .ZN(n6777) );
  AND2_X1 U5818 ( .A1(n5854), .A2(n4640), .ZN(n9380) );
  NOR2_X1 U5819 ( .A1(n9405), .A2(n10056), .ZN(n10055) );
  AOI21_X1 U5820 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10053), .ZN(n10052) );
  NOR2_X1 U5821 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  AOI21_X1 U5822 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10050), .ZN(n10049) );
  OAI21_X1 U5823 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10047), .ZN(n10045) );
  NAND2_X1 U5824 ( .A1(n4815), .A2(n5805), .ZN(n4814) );
  OAI211_X1 U5825 ( .C1(n8171), .C2(n8254), .A(n4531), .B(n4529), .ZN(P2_U3264) );
  INV_X1 U5826 ( .A(n4530), .ZN(n4529) );
  NAND2_X1 U5827 ( .A1(n4532), .A2(n8254), .ZN(n4531) );
  NAND2_X1 U5828 ( .A1(n4616), .A2(n8626), .ZN(n4613) );
  AND3_X1 U5829 ( .A1(n9751), .A2(n9750), .A3(n9749), .ZN(n9758) );
  NOR2_X1 U5830 ( .A1(n9286), .A2(n9257), .ZN(n9093) );
  NAND2_X1 U5831 ( .A1(n4568), .A2(n4394), .ZN(P1_U3520) );
  NAND2_X1 U5832 ( .A1(n9350), .A2(n9794), .ZN(n4568) );
  INV_X1 U5833 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5834 ( .B1(n7633), .B2(n7753), .A(n7756), .ZN(n4804) );
  AND2_X1 U5835 ( .A1(n8267), .A2(n4754), .ZN(n4328) );
  OR2_X1 U5836 ( .A1(n8875), .A2(n4591), .ZN(n4329) );
  AND2_X1 U5837 ( .A1(n8262), .A2(n5512), .ZN(n4330) );
  AND2_X1 U5838 ( .A1(n9122), .A2(n9107), .ZN(n4331) );
  INV_X1 U5839 ( .A(n7592), .ZN(n4747) );
  INV_X1 U5840 ( .A(n8322), .ZN(n4738) );
  NAND2_X1 U5841 ( .A1(n5746), .A2(n5747), .ZN(n4332) );
  AND2_X1 U5842 ( .A1(n4456), .A2(n4455), .ZN(n4333) );
  AND2_X1 U5843 ( .A1(n4535), .A2(n4399), .ZN(n4334) );
  OR2_X1 U5844 ( .A1(n8101), .A2(n4315), .ZN(n4335) );
  INV_X1 U5845 ( .A(n8207), .ZN(n8473) );
  NAND2_X1 U5846 ( .A1(n5393), .A2(n5392), .ZN(n8207) );
  AND2_X1 U5847 ( .A1(n4874), .A2(n4872), .ZN(n4336) );
  AND4_X1 U5848 ( .A1(n4854), .A2(n5230), .A3(n5163), .A4(n5118), .ZN(n4337)
         );
  AND4_X1 U5849 ( .A1(n4563), .A2(n4562), .A3(n6014), .A4(n5991), .ZN(n4338)
         );
  OR2_X1 U5850 ( .A1(n4804), .A2(n8813), .ZN(n4339) );
  AND2_X1 U5851 ( .A1(n6071), .A2(n7484), .ZN(n4340) );
  NAND2_X1 U5852 ( .A1(n8459), .A2(n8089), .ZN(n4341) );
  AND2_X1 U5853 ( .A1(n5353), .A2(n5352), .ZN(n8020) );
  OR2_X1 U5854 ( .A1(n4783), .A2(n4331), .ZN(n4342) );
  INV_X1 U5855 ( .A(n5747), .ZN(n4823) );
  NAND2_X1 U5856 ( .A1(n4860), .A2(n4859), .ZN(n5262) );
  NAND2_X1 U5857 ( .A1(n4610), .A2(n6091), .ZN(n9615) );
  AND2_X1 U5858 ( .A1(n5796), .A2(n5790), .ZN(n9841) );
  INV_X1 U5859 ( .A(n5921), .ZN(n8655) );
  OR2_X1 U5860 ( .A1(n9280), .A2(n9091), .ZN(n4343) );
  AND2_X1 U5861 ( .A1(n5828), .A2(n7912), .ZN(n4344) );
  NAND4_X1 U5862 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n6744)
         );
  OR2_X1 U5863 ( .A1(n7089), .A2(n7084), .ZN(n4345) );
  INV_X1 U5864 ( .A(n8281), .ZN(n4558) );
  OR2_X1 U5865 ( .A1(n5186), .A2(n4672), .ZN(n4346) );
  AND2_X1 U5866 ( .A1(n8615), .A2(n8616), .ZN(n8537) );
  NAND2_X1 U5867 ( .A1(n4839), .A2(n4858), .ZN(n5093) );
  OAI211_X1 U5868 ( .C1(n5117), .C2(n6542), .A(n5066), .B(n5065), .ZN(n9916)
         );
  AND2_X1 U5869 ( .A1(n5495), .A2(n5494), .ZN(n7674) );
  NOR2_X1 U5870 ( .A1(n9614), .A2(n7782), .ZN(n7753) );
  AND2_X1 U5871 ( .A1(n4778), .A2(n9243), .ZN(n4347) );
  NOR2_X1 U5872 ( .A1(n6618), .A2(n4503), .ZN(n4348) );
  AND2_X1 U5873 ( .A1(n8687), .A2(n8841), .ZN(n8813) );
  NAND2_X1 U5874 ( .A1(n4792), .A2(n4794), .ZN(n9059) );
  XNOR2_X1 U5875 ( .A(n4866), .B(n4998), .ZN(n5429) );
  OR2_X1 U5876 ( .A1(n9316), .A2(n9162), .ZN(n4349) );
  NOR2_X1 U5877 ( .A1(n7631), .A2(n4589), .ZN(n4350) );
  NAND2_X1 U5878 ( .A1(n5111), .A2(n5110), .ZN(n9858) );
  NAND2_X1 U5879 ( .A1(n5265), .A2(n5264), .ZN(n8453) );
  NAND2_X1 U5880 ( .A1(n6178), .A2(n6177), .ZN(n9329) );
  INV_X1 U5881 ( .A(n9329), .ZN(n4455) );
  NAND2_X1 U5882 ( .A1(n8971), .A2(n7583), .ZN(n8681) );
  INV_X1 U5883 ( .A(n8681), .ZN(n4591) );
  INV_X1 U5884 ( .A(n6466), .ZN(n4750) );
  AND3_X1 U5885 ( .A1(n5904), .A2(n5807), .A3(n5941), .ZN(n5971) );
  OR2_X1 U5886 ( .A1(n6411), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4351) );
  INV_X1 U5887 ( .A(n4871), .ZN(n6539) );
  CLKBUF_X3 U5888 ( .A(n4871), .Z(n4401) );
  OR3_X1 U5889 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4352) );
  INV_X1 U5890 ( .A(n8796), .ZN(n4580) );
  AND2_X1 U5891 ( .A1(n9827), .A2(n8094), .ZN(n4353) );
  NAND2_X1 U5892 ( .A1(n4419), .A2(n4418), .ZN(n9096) );
  OR2_X1 U5893 ( .A1(n8357), .A2(n8087), .ZN(n4354) );
  NAND2_X1 U5894 ( .A1(n5382), .A2(n5381), .ZN(n8401) );
  INV_X1 U5895 ( .A(n8401), .ZN(n4485) );
  AND2_X1 U5896 ( .A1(n8592), .A2(n4630), .ZN(n4355) );
  AND2_X1 U5897 ( .A1(n9329), .A2(n9222), .ZN(n4356) );
  AND2_X1 U5898 ( .A1(n5744), .A2(n4821), .ZN(n4357) );
  NAND2_X1 U5899 ( .A1(n5298), .A2(n5297), .ZN(n8329) );
  INV_X1 U5900 ( .A(n8896), .ZN(n4602) );
  INV_X1 U5901 ( .A(n9339), .ZN(n7916) );
  NAND2_X1 U5902 ( .A1(n6134), .A2(n6133), .ZN(n9339) );
  NAND2_X1 U5903 ( .A1(n8269), .A2(n4483), .ZN(n4487) );
  NAND2_X1 U5904 ( .A1(n5346), .A2(n5345), .ZN(n8271) );
  INV_X1 U5905 ( .A(n8271), .ZN(n4756) );
  NAND2_X1 U5906 ( .A1(n4687), .A2(n4686), .ZN(n5404) );
  AND2_X1 U5907 ( .A1(n4423), .A2(n7918), .ZN(n4358) );
  INV_X1 U5908 ( .A(n8253), .ZN(n8479) );
  NAND2_X1 U5909 ( .A1(n5357), .A2(n5356), .ZN(n8253) );
  AND2_X1 U5910 ( .A1(n7017), .A2(n5655), .ZN(n4359) );
  OR2_X1 U5911 ( .A1(n9877), .A2(n5174), .ZN(n5473) );
  NAND2_X1 U5912 ( .A1(n5289), .A2(n5288), .ZN(n8443) );
  INV_X1 U5913 ( .A(n8443), .ZN(n4473) );
  NOR2_X1 U5914 ( .A1(n9117), .A2(n4458), .ZN(n4463) );
  AND2_X1 U5915 ( .A1(n5502), .A2(n5501), .ZN(n7827) );
  INV_X1 U5916 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5012) );
  INV_X1 U5917 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5918 ( .A1(n4712), .A2(n5417), .ZN(n4360) );
  INV_X1 U5919 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U5920 ( .A1(n4343), .A2(n4850), .ZN(n4800) );
  AND2_X1 U5921 ( .A1(n9298), .A2(n8963), .ZN(n4361) );
  OR2_X1 U5922 ( .A1(n6411), .A2(n4809), .ZN(n5843) );
  NAND2_X1 U5923 ( .A1(n5015), .A2(n5014), .ZN(n8182) );
  INV_X1 U5924 ( .A(n4773), .ZN(n4772) );
  OAI21_X1 U5925 ( .B1(n4347), .B2(n4774), .A(n9219), .ZN(n4773) );
  OR2_X1 U5926 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4362) );
  AND2_X1 U5927 ( .A1(n7827), .A2(n5499), .ZN(n4363) );
  NOR2_X1 U5928 ( .A1(n7713), .A2(n7712), .ZN(n4364) );
  NOR2_X1 U5929 ( .A1(n4473), .A2(n8058), .ZN(n4365) );
  NAND2_X1 U5930 ( .A1(n9295), .A2(n9136), .ZN(n4366) );
  AND2_X1 U5931 ( .A1(n5083), .A2(n5084), .ZN(n4367) );
  INV_X1 U5932 ( .A(n4421), .ZN(n4420) );
  NAND2_X1 U5933 ( .A1(n9170), .A2(n4349), .ZN(n4421) );
  INV_X1 U5934 ( .A(n4484), .ZN(n4483) );
  NAND2_X1 U5935 ( .A1(n4486), .A2(n4485), .ZN(n4484) );
  AND4_X1 U5936 ( .A1(n4858), .A2(n5216), .A3(n5161), .A4(n4838), .ZN(n4368)
         );
  INV_X1 U5937 ( .A(n9271), .ZN(n9067) );
  NAND2_X1 U5938 ( .A1(n6367), .A2(n6366), .ZN(n9271) );
  NOR2_X1 U5939 ( .A1(n5571), .A2(n5570), .ZN(n4369) );
  NAND2_X1 U5940 ( .A1(n8329), .A2(n8085), .ZN(n4370) );
  INV_X1 U5941 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5841) );
  AND2_X1 U5942 ( .A1(n5845), .A2(n5815), .ZN(n4371) );
  AND2_X1 U5943 ( .A1(n5567), .A2(n5428), .ZN(n5600) );
  INV_X1 U5944 ( .A(n5600), .ZN(n4540) );
  AND2_X1 U5945 ( .A1(n4756), .A2(n8020), .ZN(n4372) );
  INV_X1 U5946 ( .A(n4743), .ZN(n4742) );
  AND2_X1 U5947 ( .A1(n6470), .A2(n4354), .ZN(n4743) );
  OR2_X1 U5948 ( .A1(n4791), .A2(n7919), .ZN(n4787) );
  OR2_X1 U5949 ( .A1(n4356), .A2(n4779), .ZN(n4373) );
  OR2_X1 U5950 ( .A1(n4342), .A2(n4421), .ZN(n4374) );
  OR2_X1 U5951 ( .A1(n9055), .A2(n8781), .ZN(n4375) );
  AND2_X1 U5952 ( .A1(n7316), .A2(n4757), .ZN(n4376) );
  AND2_X1 U5953 ( .A1(n5586), .A2(n5473), .ZN(n4377) );
  AND2_X1 U5954 ( .A1(n4738), .A2(n5515), .ZN(n4378) );
  AND2_X1 U5955 ( .A1(n4827), .A2(n5000), .ZN(n4379) );
  NOR2_X1 U5956 ( .A1(n6109), .A2(n4609), .ZN(n4608) );
  AND2_X1 U5957 ( .A1(n6171), .A2(n6149), .ZN(n4380) );
  INV_X1 U5958 ( .A(n4806), .ZN(n4805) );
  NAND2_X1 U5959 ( .A1(n7554), .A2(n7505), .ZN(n4806) );
  INV_X1 U5960 ( .A(n9324), .ZN(n9216) );
  NAND2_X1 U5961 ( .A1(n6197), .A2(n6196), .ZN(n9324) );
  AND2_X1 U5962 ( .A1(n4767), .A2(n5012), .ZN(n4381) );
  NAND2_X1 U5963 ( .A1(n4797), .A2(n4343), .ZN(n4796) );
  INV_X1 U5964 ( .A(n9114), .ZN(n4605) );
  INV_X1 U5965 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4829) );
  INV_X2 U5966 ( .A(n6232), .ZN(n5954) );
  NAND2_X1 U5967 ( .A1(n7317), .A2(n5586), .ZN(n4719) );
  NAND2_X1 U5968 ( .A1(n6313), .A2(n6312), .ZN(n9290) );
  INV_X1 U5969 ( .A(n9290), .ZN(n4462) );
  NAND2_X1 U5970 ( .A1(n4422), .A2(n4420), .ZN(n9172) );
  NAND2_X1 U5971 ( .A1(n5407), .A2(n5406), .ZN(n8196) );
  NOR2_X1 U5972 ( .A1(n7613), .A2(n8969), .ZN(n4382) );
  INV_X1 U5973 ( .A(n7028), .ZN(n4408) );
  OAI21_X1 U5974 ( .B1(n8347), .B2(n4742), .A(n4740), .ZN(n8321) );
  INV_X1 U5975 ( .A(n4424), .ZN(n9242) );
  INV_X1 U5976 ( .A(n8839), .ZN(n4594) );
  NAND2_X1 U5977 ( .A1(n6210), .A2(n6211), .ZN(n8615) );
  NAND2_X1 U5978 ( .A1(n6150), .A2(n6149), .ZN(n8565) );
  NAND2_X1 U5979 ( .A1(n4338), .A2(n4405), .ZN(n6075) );
  NOR2_X1 U5980 ( .A1(n9199), .A2(n9316), .ZN(n9164) );
  NOR2_X1 U5981 ( .A1(n9649), .A2(n8699), .ZN(n4383) );
  NAND2_X1 U5982 ( .A1(n8368), .A2(n4472), .ZN(n4475) );
  NAND2_X1 U5983 ( .A1(n7866), .A2(n4333), .ZN(n4457) );
  AND2_X1 U5984 ( .A1(n4493), .A2(n4492), .ZN(n4384) );
  AND2_X1 U5985 ( .A1(n6688), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4385) );
  OR2_X1 U5986 ( .A1(n6511), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4386) );
  INV_X1 U5987 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5163) );
  NOR2_X1 U5988 ( .A1(n6612), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4387) );
  INV_X1 U5989 ( .A(n4755), .ZN(n8425) );
  NAND2_X1 U5990 ( .A1(n4753), .A2(n4558), .ZN(n4755) );
  NOR2_X1 U5991 ( .A1(n9216), .A2(n9197), .ZN(n4388) );
  AND2_X1 U5992 ( .A1(n4777), .A2(n4776), .ZN(n4389) );
  AND2_X1 U5993 ( .A1(n6493), .A2(n4444), .ZN(n4390) );
  NAND2_X1 U5994 ( .A1(n9267), .A2(n9347), .ZN(n4391) );
  NAND2_X1 U5995 ( .A1(n8971), .A2(n7559), .ZN(n4392) );
  NAND2_X1 U5996 ( .A1(n7083), .A2(n7084), .ZN(n4734) );
  NOR2_X1 U5997 ( .A1(n7554), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U5998 ( .A1(n5220), .A2(n5219), .ZN(n9638) );
  INV_X1 U5999 ( .A(n9638), .ZN(n4481) );
  NAND2_X1 U6000 ( .A1(n4825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  NOR2_X1 U6001 ( .A1(n5418), .A2(n6595), .ZN(n4393) );
  OR2_X1 U6002 ( .A1(n9794), .A2(n4567), .ZN(n4394) );
  NAND2_X1 U6003 ( .A1(n4417), .A2(n4415), .ZN(n7537) );
  NAND2_X1 U6004 ( .A1(n7395), .A2(n8805), .ZN(n7506) );
  AND2_X1 U6005 ( .A1(n7506), .A2(n7505), .ZN(n7552) );
  NAND2_X1 U6006 ( .A1(n4636), .A2(n4637), .ZN(n7464) );
  NAND2_X1 U6007 ( .A1(n7593), .A2(n7592), .ZN(n7591) );
  NAND2_X1 U6008 ( .A1(n6463), .A2(n6462), .ZN(n7171) );
  OR2_X1 U6009 ( .A1(n7596), .A2(n4478), .ZN(n4395) );
  OR2_X1 U6010 ( .A1(n5618), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4396) );
  AND2_X1 U6011 ( .A1(n4990), .A2(n9528), .ZN(n4397) );
  INV_X1 U6012 ( .A(n4758), .ZN(n7170) );
  NAND2_X1 U6013 ( .A1(n6463), .A2(n4759), .ZN(n4758) );
  AND2_X1 U6014 ( .A1(n9856), .A2(n5667), .ZN(n4398) );
  INV_X1 U6015 ( .A(n9827), .ZN(n4480) );
  NOR2_X1 U6016 ( .A1(n9952), .A2(n5573), .ZN(n4399) );
  AND2_X1 U6017 ( .A1(n9784), .A2(n6415), .ZN(n8626) );
  INV_X1 U6018 ( .A(n8626), .ZN(n9618) );
  AND2_X1 U6019 ( .A1(n9731), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4400) );
  INV_X1 U6020 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4465) );
  INV_X1 U6021 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n4509) );
  NAND2_X2 U6022 ( .A1(n5432), .A2(n7944), .ZN(n5570) );
  INV_X1 U6023 ( .A(n4696), .ZN(n4640) );
  OAI21_X2 U6024 ( .B1(n7871), .B2(n8817), .A(n8879), .ZN(n7921) );
  OAI21_X1 U6025 ( .B1(n7758), .B2(n7757), .A(n8842), .ZN(n7781) );
  INV_X1 U6026 ( .A(n4600), .ZN(n9112) );
  INV_X1 U6027 ( .A(n8840), .ZN(n4589) );
  AOI21_X2 U6028 ( .B1(n9244), .B2(n8885), .A(n7922), .ZN(n9231) );
  NAND2_X1 U6029 ( .A1(n7299), .A2(n7138), .ZN(n4572) );
  NAND2_X1 U6030 ( .A1(n4595), .A2(n4605), .ZN(n4600) );
  NAND2_X1 U6031 ( .A1(n4600), .A2(n4603), .ZN(n9087) );
  NAND2_X1 U6032 ( .A1(n4881), .A2(n4880), .ZN(n5063) );
  NAND2_X2 U6033 ( .A1(n8365), .A2(n6468), .ZN(n8347) );
  INV_X1 U6034 ( .A(n4446), .ZN(n6497) );
  AOI21_X1 U6035 ( .B1(n8189), .B2(n10008), .A(n4448), .ZN(n4447) );
  NAND2_X1 U6036 ( .A1(n5062), .A2(n5063), .ZN(n4409) );
  INV_X1 U6037 ( .A(n5557), .ZN(n5556) );
  NAND2_X1 U6038 ( .A1(n4969), .A2(n4968), .ZN(n5344) );
  NAND2_X1 U6039 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U6040 ( .A1(n5606), .A2(n5605), .ZN(n5610) );
  AOI21_X1 U6041 ( .B1(n4411), .B2(n5566), .A(n4410), .ZN(n5569) );
  AND2_X1 U6042 ( .A1(n5574), .A2(n5570), .ZN(n4410) );
  OAI21_X1 U6043 ( .B1(n5563), .B2(n5564), .A(n5562), .ZN(n4411) );
  INV_X1 U6044 ( .A(n7616), .ZN(n4426) );
  OAI21_X1 U6045 ( .B1(n4339), .B2(n4426), .A(n4427), .ZN(n7864) );
  NAND2_X1 U6046 ( .A1(n7616), .A2(n7615), .ZN(n7628) );
  NAND4_X1 U6047 ( .A1(n4431), .A2(n4430), .A3(n4391), .A4(n4466), .ZN(n9350)
         );
  NAND2_X1 U6048 ( .A1(n8278), .A2(n4330), .ZN(n4437) );
  NAND2_X1 U6049 ( .A1(n4437), .A2(n4438), .ZN(n8246) );
  NAND2_X1 U6050 ( .A1(n7829), .A2(n4442), .ZN(n8348) );
  NAND2_X1 U6051 ( .A1(n4445), .A2(n4390), .ZN(P2_U3549) );
  OR2_X1 U6052 ( .A1(n10026), .A2(n6491), .ZN(n4444) );
  NAND2_X1 U6053 ( .A1(n4446), .A2(n10026), .ZN(n4445) );
  INV_X1 U6054 ( .A(n4457), .ZN(n9227) );
  OR3_X1 U6055 ( .A1(n9117), .A2(n9283), .A3(n4461), .ZN(n9063) );
  INV_X1 U6056 ( .A(n4463), .ZN(n9062) );
  INV_X1 U6057 ( .A(n7034), .ZN(n7270) );
  MUX2_X1 U6058 ( .A(n4465), .B(n4464), .S(n6506), .Z(n7034) );
  NAND2_X2 U6059 ( .A1(n5859), .A2(n5858), .ZN(n6423) );
  AND2_X1 U6060 ( .A1(n5047), .A2(n5046), .ZN(n4468) );
  NAND2_X2 U6061 ( .A1(n4468), .A2(n4469), .ZN(n9958) );
  OR2_X1 U6062 ( .A1(n5117), .A2(n6554), .ZN(n4469) );
  INV_X1 U6063 ( .A(n4475), .ZN(n8341) );
  INV_X1 U6064 ( .A(n7596), .ZN(n4476) );
  NAND2_X1 U6065 ( .A1(n4476), .A2(n4477), .ZN(n7743) );
  NAND2_X1 U6066 ( .A1(n8269), .A2(n4482), .ZN(n6487) );
  INV_X1 U6067 ( .A(n4487), .ZN(n8222) );
  XNOR2_X1 U6068 ( .A(n8984), .B(n9004), .ZN(n9705) );
  NAND2_X1 U6069 ( .A1(n6661), .A2(n4499), .ZN(n4498) );
  INV_X1 U6070 ( .A(n4505), .ZN(n6616) );
  INV_X1 U6071 ( .A(n6658), .ZN(n4507) );
  MUX2_X1 U6072 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6710), .S(n8109), .Z(n8107)
         );
  NAND2_X1 U6073 ( .A1(n4534), .A2(n4535), .ZN(n5604) );
  NAND2_X1 U6074 ( .A1(n5080), .A2(n5079), .ZN(n4554) );
  OAI21_X1 U6075 ( .B1(n5080), .B2(n4555), .A(n4552), .ZN(n4556) );
  INV_X1 U6076 ( .A(n5038), .ZN(n4698) );
  NAND2_X2 U6077 ( .A1(n4870), .A2(n4869), .ZN(n4871) );
  NAND2_X1 U6078 ( .A1(n8800), .A2(n8922), .ZN(n7137) );
  NAND3_X1 U6079 ( .A1(n4566), .A2(n4565), .A3(n4564), .ZN(n5959) );
  OAI21_X2 U6080 ( .B1(n8665), .B2(n7211), .A(n8854), .ZN(n7382) );
  NAND2_X1 U6081 ( .A1(n4572), .A2(n8924), .ZN(n8665) );
  OAI22_X1 U6082 ( .A1(n6554), .A2(n6539), .B1(n6555), .B2(n4401), .ZN(n4574)
         );
  AND2_X2 U6083 ( .A1(n5889), .A2(n4573), .ZN(n7032) );
  NAND2_X2 U6084 ( .A1(n6506), .A2(n6539), .ZN(n5927) );
  NAND2_X1 U6085 ( .A1(n9218), .A2(n4581), .ZN(n4578) );
  NAND2_X1 U6086 ( .A1(n4578), .A2(n4579), .ZN(n9157) );
  INV_X1 U6087 ( .A(n4586), .ZN(n9193) );
  NAND3_X1 U6088 ( .A1(n4350), .A2(n4593), .A3(n7508), .ZN(n4588) );
  NAND3_X1 U6089 ( .A1(n4588), .A2(n8687), .A3(n4587), .ZN(n7758) );
  INV_X1 U6090 ( .A(n9113), .ZN(n4595) );
  NAND2_X1 U6091 ( .A1(n9113), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U6092 ( .A1(n9616), .A2(n4608), .ZN(n4606) );
  NAND2_X1 U6093 ( .A1(n4606), .A2(n4607), .ZN(n7765) );
  NAND2_X1 U6094 ( .A1(n8515), .A2(n4612), .ZN(n4611) );
  OAI211_X1 U6095 ( .C1(n8515), .C2(n4613), .A(n4611), .B(n6444), .ZN(P1_U3218) );
  NOR2_X1 U6096 ( .A1(n6384), .A2(n6365), .ZN(n4617) );
  NAND2_X1 U6097 ( .A1(n6384), .A2(n6365), .ZN(n4618) );
  INV_X1 U6098 ( .A(n6384), .ZN(n4619) );
  NAND2_X1 U6099 ( .A1(n6150), .A2(n4380), .ZN(n8566) );
  NOR2_X1 U6100 ( .A1(n4620), .A2(n7005), .ZN(n4622) );
  XNOR2_X1 U6101 ( .A(n4623), .B(n7008), .ZN(n7014) );
  AOI21_X2 U6102 ( .B1(n6210), .B2(n4355), .A(n4625), .ZN(n8595) );
  NAND2_X1 U6103 ( .A1(n4633), .A2(n4340), .ZN(n7691) );
  NAND2_X1 U6104 ( .A1(n7250), .A2(n4638), .ZN(n4636) );
  NAND2_X1 U6105 ( .A1(n5833), .A2(n4639), .ZN(n6173) );
  XNOR2_X1 U6106 ( .A(n5867), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6385) );
  AND2_X1 U6107 ( .A1(n7158), .A2(n5999), .ZN(n6001) );
  XNOR2_X1 U6108 ( .A(n5109), .B(n5108), .ZN(n6557) );
  INV_X1 U6109 ( .A(n4766), .ZN(n5011) );
  NAND2_X1 U6110 ( .A1(n5229), .A2(n4648), .ZN(n4644) );
  NAND2_X1 U6111 ( .A1(n4644), .A2(n4645), .ZN(n5272) );
  NAND2_X1 U6112 ( .A1(n5420), .A2(n4661), .ZN(n4656) );
  NAND2_X1 U6113 ( .A1(n4912), .A2(n4670), .ZN(n4667) );
  NAND2_X1 U6114 ( .A1(n4667), .A2(n4668), .ZN(n4925) );
  NAND2_X1 U6115 ( .A1(n5116), .A2(n4679), .ZN(n4676) );
  NAND2_X1 U6116 ( .A1(n4676), .A2(n4677), .ZN(n4906) );
  NAND2_X1 U6117 ( .A1(n5379), .A2(n4689), .ZN(n4687) );
  NAND2_X1 U6118 ( .A1(n5379), .A2(n5380), .ZN(n4688) );
  OAI21_X2 U6119 ( .B1(n5344), .B2(n4692), .A(n4972), .ZN(n5355) );
  NAND2_X1 U6120 ( .A1(n8246), .A2(n8247), .ZN(n4693) );
  OAI211_X1 U6121 ( .C1(n8246), .C2(n8247), .A(n4693), .B(n9922), .ZN(n8249)
         );
  AOI21_X1 U6122 ( .B1(n4693), .B2(n8232), .A(n8231), .ZN(n8233) );
  NAND2_X1 U6123 ( .A1(n5109), .A2(n5108), .ZN(n4694) );
  NAND2_X1 U6124 ( .A1(n5043), .A2(n5044), .ZN(n4877) );
  NAND2_X1 U6125 ( .A1(n5038), .A2(SI_1_), .ZN(n4699) );
  OR2_X1 U6126 ( .A1(n6480), .A2(n4704), .ZN(n4703) );
  NAND2_X1 U6127 ( .A1(n4703), .A2(n4701), .ZN(n4714) );
  NAND2_X1 U6128 ( .A1(n7317), .A2(n4377), .ZN(n4715) );
  NAND3_X1 U6129 ( .A1(n4716), .A2(n5577), .A3(n4715), .ZN(n7521) );
  NAND2_X1 U6130 ( .A1(n4720), .A2(n4378), .ZN(n8325) );
  NAND2_X1 U6131 ( .A1(n8309), .A2(n4726), .ZN(n4723) );
  NAND3_X1 U6132 ( .A1(n4730), .A2(n7117), .A3(n4729), .ZN(n6460) );
  NAND2_X1 U6133 ( .A1(n4732), .A2(n6458), .ZN(n4729) );
  NAND3_X1 U6134 ( .A1(n7083), .A2(n7084), .A3(n6458), .ZN(n4730) );
  OAI21_X2 U6135 ( .B1(n8347), .B2(n4739), .A(n4736), .ZN(n4735) );
  INV_X1 U6136 ( .A(n8282), .ZN(n4753) );
  NAND2_X1 U6137 ( .A1(n8282), .A2(n4328), .ZN(n4751) );
  NOR2_X1 U6138 ( .A1(n8425), .A2(n6473), .ZN(n8268) );
  NAND2_X1 U6139 ( .A1(n4758), .A2(n4376), .ZN(n7312) );
  INV_X1 U6140 ( .A(n4764), .ZN(n7825) );
  OR2_X1 U6141 ( .A1(n7744), .A2(n8090), .ZN(n4765) );
  NAND2_X1 U6142 ( .A1(n5247), .A2(n5005), .ZN(n5618) );
  AND3_X2 U6143 ( .A1(n5247), .A2(n5005), .A3(n4381), .ZN(n5009) );
  INV_X1 U6144 ( .A(n9080), .ZN(n4801) );
  NAND2_X1 U6145 ( .A1(n9080), .A2(n4796), .ZN(n4792) );
  NOR2_X2 U6146 ( .A1(n6411), .A2(n4807), .ZN(n5861) );
  NAND3_X1 U6147 ( .A1(n7219), .A2(n7218), .A3(n7279), .ZN(n7278) );
  INV_X1 U6148 ( .A(n5572), .ZN(n5625) );
  NAND3_X1 U6149 ( .A1(n6907), .A2(n5643), .A3(n5636), .ZN(n6937) );
  AOI21_X1 U6150 ( .B1(n5792), .B2(n4816), .A(n4814), .ZN(n4813) );
  OAI21_X1 U6151 ( .B1(n5806), .B2(n8207), .A(n4813), .ZN(P2_U3222) );
  NAND2_X1 U6152 ( .A1(n5745), .A2(n4357), .ZN(n4820) );
  OAI211_X1 U6153 ( .C1(n5745), .C2(n4332), .A(n4820), .B(n4818), .ZN(n7994)
         );
  NAND2_X1 U6154 ( .A1(n4860), .A2(n4827), .ZN(n4861) );
  NAND2_X1 U6155 ( .A1(n4860), .A2(n4379), .ZN(n4825) );
  INV_X1 U6156 ( .A(n4828), .ZN(n4826) );
  NAND2_X1 U6157 ( .A1(n9856), .A2(n4832), .ZN(n7124) );
  NAND2_X1 U6158 ( .A1(n7124), .A2(n5672), .ZN(n5677) );
  AND4_X2 U6159 ( .A1(n4839), .A2(n4840), .A3(n4368), .A4(n4337), .ZN(n5247)
         );
  NAND2_X1 U6160 ( .A1(n7982), .A2(n5735), .ZN(n5736) );
  NAND2_X1 U6161 ( .A1(n7976), .A2(n4842), .ZN(n7982) );
  NAND2_X1 U6162 ( .A1(n7894), .A2(n5718), .ZN(n5723) );
  NAND2_X1 U6163 ( .A1(n5712), .A2(n4843), .ZN(n7894) );
  NAND2_X1 U6164 ( .A1(n6950), .A2(n6947), .ZN(n6948) );
  NAND2_X1 U6165 ( .A1(n5367), .A2(n5366), .ZN(n4982) );
  AOI21_X1 U6166 ( .B1(n7921), .B2(n8838), .A(n8883), .ZN(n9244) );
  INV_X1 U6167 ( .A(n7912), .ZN(n5827) );
  AND2_X2 U6168 ( .A1(n5826), .A2(n7912), .ZN(n6232) );
  NAND2_X1 U6169 ( .A1(n4325), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U6170 ( .A1(n5861), .A2(n5817), .ZN(n5822) );
  OR2_X1 U6171 ( .A1(n5009), .A2(n8498), .ZN(n5007) );
  NAND2_X1 U6172 ( .A1(n5819), .A2(n5818), .ZN(n5824) );
  INV_X1 U6173 ( .A(n5822), .ZN(n5819) );
  CLKBUF_X1 U6174 ( .A(n5048), .Z(n9833) );
  NAND2_X1 U6175 ( .A1(n6744), .A2(n5909), .ZN(n5881) );
  NAND2_X1 U6176 ( .A1(n6973), .A2(n5579), .ZN(n5445) );
  INV_X1 U6177 ( .A(n9270), .ZN(n9275) );
  NOR2_X1 U6178 ( .A1(n9270), .A2(n9257), .ZN(n9077) );
  NAND2_X1 U6179 ( .A1(n5011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5013) );
  OR2_X1 U6180 ( .A1(n4326), .A2(n7058), .ZN(n5902) );
  NAND2_X2 U6181 ( .A1(n5759), .A2(n8062), .ZN(n7950) );
  NAND2_X1 U6182 ( .A1(n4861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4862) );
  XNOR2_X2 U6183 ( .A(n5741), .B(n5742), .ZN(n8039) );
  INV_X1 U6184 ( .A(n5489), .ZN(n5213) );
  INV_X1 U6185 ( .A(n8378), .ZN(n5270) );
  NAND2_X1 U6186 ( .A1(n5848), .A2(n5847), .ZN(n6388) );
  INV_X1 U6187 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4859) );
  INV_X1 U6188 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5150) );
  AND2_X1 U6189 ( .A1(n7161), .A2(n6000), .ZN(n4846) );
  OR2_X1 U6190 ( .A1(n7732), .A2(n6467), .ZN(n4847) );
  AND2_X1 U6191 ( .A1(n8712), .A2(n8703), .ZN(n4848) );
  INV_X1 U6192 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9816) );
  INV_X1 U6193 ( .A(n5260), .ZN(n4860) );
  AND2_X1 U6194 ( .A1(n9283), .A2(n8962), .ZN(n4849) );
  OR2_X1 U6195 ( .A1(n9283), .A2(n8962), .ZN(n4850) );
  AND2_X1 U6196 ( .A1(n7240), .A2(n8097), .ZN(n4851) );
  AND2_X1 U6197 ( .A1(n8036), .A2(n5794), .ZN(n9859) );
  INV_X1 U6198 ( .A(n9859), .ZN(n5795) );
  AND2_X1 U6199 ( .A1(n7366), .A2(n5980), .ZN(n4852) );
  NAND2_X2 U6200 ( .A1(n7397), .A2(n9145), .ZN(n9263) );
  INV_X2 U6201 ( .A(n9803), .ZN(n9802) );
  AND2_X1 U6202 ( .A1(n5694), .A2(n5693), .ZN(n4853) );
  INV_X1 U6203 ( .A(n8357), .ZN(n8495) );
  INV_X1 U6204 ( .A(n8494), .ZN(n6500) );
  INV_X1 U6205 ( .A(n8451), .ZN(n6492) );
  OR2_X1 U6206 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  AND2_X1 U6207 ( .A1(n5528), .A2(n5532), .ZN(n5529) );
  OAI21_X1 U6208 ( .B1(n5531), .B2(n5530), .A(n5529), .ZN(n5538) );
  INV_X1 U6209 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5001) );
  INV_X1 U6210 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5810) );
  INV_X1 U6211 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5008) );
  INV_X1 U6212 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5815) );
  NOR2_X1 U6213 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  INV_X1 U6214 ( .A(n9958), .ZN(n6448) );
  INV_X1 U6215 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5006) );
  INV_X1 U6216 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5161) );
  INV_X1 U6217 ( .A(n7694), .ZN(n6071) );
  INV_X1 U6218 ( .A(n9049), .ZN(n9037) );
  INV_X1 U6219 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n4933) );
  INV_X1 U6220 ( .A(n9838), .ZN(n5643) );
  INV_X1 U6221 ( .A(n5277), .ZN(n5279) );
  INV_X1 U6222 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U6223 ( .A1(n9069), .A2(n9070), .ZN(n9068) );
  INV_X1 U6224 ( .A(n6267), .ZN(n6266) );
  INV_X1 U6225 ( .A(SI_26_), .ZN(n9499) );
  INV_X1 U6226 ( .A(SI_23_), .ZN(n4964) );
  INV_X1 U6227 ( .A(SI_20_), .ZN(n9513) );
  INV_X1 U6228 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6229 ( .A1(n8018), .A2(n8022), .ZN(n5749) );
  INV_X1 U6230 ( .A(n7892), .ZN(n5717) );
  INV_X1 U6231 ( .A(n5322), .ZN(n5321) );
  INV_X1 U6232 ( .A(n9852), .ZN(n5663) );
  NAND2_X1 U6233 ( .A1(n5334), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5347) );
  INV_X1 U6234 ( .A(n8501), .ZN(n5023) );
  NAND2_X1 U6235 ( .A1(n8375), .A2(n8056), .ZN(n6468) );
  NOR2_X1 U6236 ( .A1(n5151), .A2(n5150), .ZN(n5168) );
  INV_X1 U6237 ( .A(n7463), .ZN(n5630) );
  NAND2_X1 U6238 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  NAND2_X1 U6239 ( .A1(n5857), .A2(n5856), .ZN(n5859) );
  INV_X1 U6240 ( .A(n6158), .ZN(n6156) );
  INV_X1 U6241 ( .A(n9617), .ZN(n6091) );
  AND2_X1 U6242 ( .A1(n6410), .A2(n7096), .ZN(n6433) );
  AND2_X1 U6243 ( .A1(n8627), .A2(n8624), .ZN(n6343) );
  NAND2_X1 U6244 ( .A1(n6279), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U6245 ( .A1(n6266), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6281) );
  INV_X1 U6246 ( .A(n9164), .ZN(n9184) );
  AND2_X1 U6247 ( .A1(n8850), .A2(n8659), .ZN(n8803) );
  OR2_X1 U6248 ( .A1(n7030), .A2(n6418), .ZN(n6432) );
  INV_X1 U6249 ( .A(SI_14_), .ZN(n9522) );
  OR2_X1 U6250 ( .A1(n5123), .A2(n5122), .ZN(n5137) );
  INV_X1 U6251 ( .A(n8087), .ZN(n7970) );
  XNOR2_X1 U6252 ( .A(n5633), .B(n5634), .ZN(n6908) );
  INV_X1 U6253 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9544) );
  OR2_X1 U6254 ( .A1(n5252), .A2(n9544), .ZN(n5277) );
  OR2_X1 U6255 ( .A1(n5290), .A2(n9481), .ZN(n5309) );
  NAND2_X1 U6256 ( .A1(n5321), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5335) );
  INV_X1 U6257 ( .A(n8088), .ZN(n8056) );
  NAND2_X1 U6258 ( .A1(n5796), .A2(n5798), .ZN(n9844) );
  AND3_X1 U6259 ( .A1(n5030), .A2(n5029), .A3(n5028), .ZN(n8178) );
  INV_X1 U6260 ( .A(n4323), .ZN(n5408) );
  AND2_X2 U6261 ( .A1(n5024), .A2(n5023), .ZN(n5068) );
  INV_X1 U6262 ( .A(n8077), .ZN(n6484) );
  INV_X1 U6263 ( .A(n9834), .ZN(n8057) );
  INV_X1 U6264 ( .A(n8297), .ZN(n8291) );
  OAI22_X1 U6265 ( .A1(n7519), .A2(n7522), .B1(n7663), .B2(n8093), .ZN(n7566)
         );
  NAND2_X1 U6266 ( .A1(n6915), .A2(n9951), .ZN(n6973) );
  INV_X1 U6267 ( .A(n8196), .ZN(n6499) );
  AND2_X1 U6268 ( .A1(n5576), .A2(n5575), .ZN(n7522) );
  OR2_X1 U6269 ( .A1(n5798), .A2(n6972), .ZN(n10002) );
  OR2_X1 U6270 ( .A1(n6697), .A2(n6507), .ZN(n5801) );
  INV_X1 U6271 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5608) );
  NOR2_X1 U6272 ( .A1(n6061), .A2(n6060), .ZN(n6079) );
  OR2_X1 U6273 ( .A1(n6296), .A2(n6295), .ZN(n6316) );
  OR2_X1 U6274 ( .A1(n6224), .A2(n6223), .ZN(n8592) );
  OR2_X1 U6275 ( .A1(n9101), .A2(n6425), .ZN(n6322) );
  OR2_X1 U6276 ( .A1(n6228), .A2(n8596), .ZN(n6248) );
  NAND2_X1 U6277 ( .A1(n5914), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5885) );
  AND2_X1 U6278 ( .A1(n8999), .A2(n8998), .ZN(n9697) );
  OR2_X1 U6279 ( .A1(n9290), .A2(n9090), .ZN(n7920) );
  INV_X1 U6280 ( .A(n9298), .ZN(n9132) );
  INV_X1 U6281 ( .A(n9607), .ZN(n8699) );
  AND2_X1 U6282 ( .A1(n8680), .A2(n8671), .ZN(n8808) );
  INV_X1 U6283 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5820) );
  AND2_X1 U6284 ( .A1(n4981), .A2(n4980), .ZN(n5366) );
  AND2_X1 U6285 ( .A1(n4937), .A2(n4936), .ZN(n5245) );
  AND2_X1 U6286 ( .A1(n4911), .A2(n4910), .ZN(n5159) );
  OAI21_X1 U6287 ( .B1(n8202), .B2(n9844), .A(n5803), .ZN(n5804) );
  AND2_X1 U6288 ( .A1(n6488), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6904) );
  OR2_X1 U6289 ( .A1(n7997), .A2(n5408), .ZN(n5365) );
  AND2_X1 U6290 ( .A1(n7710), .A2(n5621), .ZN(n6697) );
  INV_X1 U6291 ( .A(n7885), .ZN(n7877) );
  AND2_X1 U6292 ( .A1(n6712), .A2(n5622), .ZN(n8169) );
  INV_X1 U6293 ( .A(n5429), .ZN(n8254) );
  OR2_X1 U6294 ( .A1(n9944), .A2(n6969), .ZN(n9894) );
  INV_X1 U6295 ( .A(n9894), .ZN(n9928) );
  AND2_X1 U6296 ( .A1(n9938), .A2(n9896), .ZN(n9931) );
  NAND2_X1 U6297 ( .A1(n7602), .A2(n7594), .ZN(n10008) );
  AND2_X1 U6298 ( .A1(n7858), .A2(n5782), .ZN(n9943) );
  AND2_X1 U6299 ( .A1(n5096), .A2(n5095), .ZN(n6821) );
  AND2_X1 U6300 ( .A1(n6436), .A2(n6419), .ZN(n9621) );
  INV_X1 U6301 ( .A(n6418), .ZN(n8949) );
  AND2_X1 U6302 ( .A1(n6322), .A2(n6321), .ZN(n9116) );
  AND4_X1 U6303 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n8579)
         );
  INV_X1 U6304 ( .A(n9748), .ZN(n6994) );
  AND2_X1 U6305 ( .A1(n6534), .A2(n6582), .ZN(n9746) );
  AND2_X1 U6306 ( .A1(n6534), .A2(n6423), .ZN(n9748) );
  AND2_X1 U6307 ( .A1(n9217), .A2(n8835), .ZN(n9230) );
  INV_X1 U6308 ( .A(n9246), .ZN(n9237) );
  AND2_X1 U6309 ( .A1(n9263), .A2(n9168), .ZN(n9203) );
  NOR2_X1 U6310 ( .A1(n6772), .A2(n6742), .ZN(n6743) );
  INV_X1 U6311 ( .A(n9786), .ZN(n9646) );
  NAND2_X1 U6312 ( .A1(n7786), .A2(n7027), .ZN(n9790) );
  AND2_X1 U6313 ( .A1(n6409), .A2(n6408), .ZN(n7096) );
  INV_X1 U6314 ( .A(n6385), .ZN(n6386) );
  INV_X1 U6315 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6129) );
  NOR2_X1 U6316 ( .A1(n9392), .A2(n9391), .ZN(n10069) );
  INV_X1 U6317 ( .A(n8174), .ZN(n9866) );
  INV_X1 U6318 ( .A(n5804), .ZN(n5805) );
  INV_X1 U6319 ( .A(n9841), .ZN(n9854) );
  NAND2_X1 U6320 ( .A1(n5802), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9863) );
  AND3_X1 U6321 ( .A1(n5027), .A2(n5026), .A3(n5025), .ZN(n6595) );
  INV_X1 U6322 ( .A(n8020), .ZN(n8081) );
  NAND2_X1 U6323 ( .A1(n6697), .A2(n9949), .ZN(n8098) );
  INV_X1 U6324 ( .A(n8169), .ZN(n9867) );
  INV_X1 U6325 ( .A(n9864), .ZN(n9868) );
  AND2_X1 U6326 ( .A1(n6577), .A2(n6576), .ZN(n8174) );
  NAND2_X2 U6327 ( .A1(n6971), .A2(n9894), .ZN(n9938) );
  INV_X1 U6328 ( .A(n9934), .ZN(n8385) );
  NAND2_X1 U6329 ( .A1(n10026), .A2(n9987), .ZN(n8451) );
  INV_X1 U6330 ( .A(n10026), .ZN(n10024) );
  INV_X1 U6331 ( .A(n8182), .ZN(n8469) );
  INV_X1 U6332 ( .A(n8329), .ZN(n8489) );
  NAND2_X1 U6333 ( .A1(n10012), .A2(n9987), .ZN(n8494) );
  INV_X1 U6334 ( .A(n10012), .ZN(n10010) );
  OR2_X1 U6335 ( .A1(n9944), .A2(n9943), .ZN(n9947) );
  INV_X1 U6336 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7797) );
  OR2_X1 U6337 ( .A1(n5249), .A2(n4860), .ZN(n7885) );
  INV_X1 U6338 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6601) );
  INV_X1 U6339 ( .A(n6443), .ZN(n6444) );
  AND2_X1 U6340 ( .A1(n6437), .A2(n6436), .ZN(n9625) );
  NAND2_X1 U6341 ( .A1(n6431), .A2(n6430), .ZN(n9072) );
  INV_X1 U6342 ( .A(n9107), .ZN(n9136) );
  INV_X1 U6343 ( .A(n8579), .ZN(n9233) );
  INV_X1 U6344 ( .A(n9746), .ZN(n9715) );
  INV_X1 U6345 ( .A(n9736), .ZN(n9756) );
  AND3_X1 U6346 ( .A1(n9734), .A2(n9733), .A3(n9732), .ZN(n9740) );
  NAND2_X1 U6347 ( .A1(n9263), .A2(n7223), .ZN(n9265) );
  INV_X1 U6348 ( .A(n9263), .ZN(n9257) );
  INV_X1 U6349 ( .A(n9263), .ZN(n9205) );
  NAND2_X1 U6350 ( .A1(n6773), .A2(n6743), .ZN(n9803) );
  NAND2_X1 U6351 ( .A1(n6773), .A2(n7097), .ZN(n9792) );
  NAND2_X1 U6352 ( .A1(n7098), .A2(n6571), .ZN(n9760) );
  AND2_X1 U6353 ( .A1(n6504), .A2(n6414), .ZN(n7098) );
  INV_X1 U6354 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7860) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6962) );
  INV_X1 U6356 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U6357 ( .A1(n10055), .A2(n10054), .ZN(n10053) );
  INV_X1 U6358 ( .A(n8098), .ZN(P2_U3966) );
  AND2_X1 U6359 ( .A1(n6535), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NOR2_X1 U6360 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4856) );
  NAND2_X1 U6361 ( .A1(n5055), .A2(n4857), .ZN(n5081) );
  NAND2_X1 U6362 ( .A1(n5247), .A2(n5002), .ZN(n5260) );
  NAND2_X1 U6363 ( .A1(n4866), .A2(n4998), .ZN(n4864) );
  XNOR2_X2 U6364 ( .A(n4865), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6478) );
  OR2_X4 U6365 ( .A1(n6972), .A2(n6478), .ZN(n10004) );
  INV_X4 U6366 ( .A(n6984), .ZN(n9898) );
  NAND2_X1 U6367 ( .A1(n5630), .A2(n6478), .ZN(n6482) );
  NAND2_X1 U6368 ( .A1(n9596), .A2(n4867), .ZN(n4870) );
  AND2_X1 U6369 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4872) );
  AND2_X1 U6370 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4873) );
  INV_X1 U6371 ( .A(SI_1_), .ZN(n4874) );
  MUX2_X1 U6372 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4871), .Z(n5043) );
  NAND2_X1 U6373 ( .A1(n4875), .A2(SI_1_), .ZN(n4876) );
  NAND2_X1 U6374 ( .A1(n4877), .A2(n4876), .ZN(n5054) );
  MUX2_X1 U6375 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4871), .Z(n4879) );
  INV_X1 U6376 ( .A(SI_2_), .ZN(n4878) );
  XNOR2_X1 U6377 ( .A(n4879), .B(n4878), .ZN(n5053) );
  NAND2_X1 U6378 ( .A1(n5054), .A2(n5053), .ZN(n4881) );
  NAND2_X1 U6379 ( .A1(n4879), .A2(SI_2_), .ZN(n4880) );
  MUX2_X1 U6380 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4871), .Z(n4882) );
  INV_X1 U6381 ( .A(SI_3_), .ZN(n9482) );
  XNOR2_X1 U6382 ( .A(n4882), .B(n9482), .ZN(n5062) );
  NAND2_X1 U6383 ( .A1(n4882), .A2(SI_3_), .ZN(n4883) );
  MUX2_X1 U6384 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4871), .Z(n4885) );
  INV_X1 U6385 ( .A(SI_4_), .ZN(n4884) );
  XNOR2_X1 U6386 ( .A(n4885), .B(n4884), .ZN(n5079) );
  NAND2_X1 U6387 ( .A1(n4885), .A2(SI_4_), .ZN(n4886) );
  MUX2_X1 U6388 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4871), .Z(n4888) );
  INV_X1 U6389 ( .A(SI_5_), .ZN(n4887) );
  XNOR2_X1 U6390 ( .A(n4888), .B(n4887), .ZN(n5091) );
  NAND2_X1 U6391 ( .A1(n4888), .A2(SI_5_), .ZN(n4889) );
  INV_X1 U6392 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6558) );
  INV_X1 U6393 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6556) );
  MUX2_X1 U6394 ( .A(n6558), .B(n6556), .S(n4871), .Z(n4890) );
  XNOR2_X1 U6395 ( .A(n4890), .B(SI_6_), .ZN(n5108) );
  INV_X1 U6396 ( .A(n4890), .ZN(n4891) );
  NAND2_X1 U6397 ( .A1(n4891), .A2(SI_6_), .ZN(n4892) );
  MUX2_X1 U6398 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4871), .Z(n4894) );
  INV_X1 U6399 ( .A(SI_7_), .ZN(n4893) );
  XNOR2_X1 U6400 ( .A(n4894), .B(n4893), .ZN(n5115) );
  NAND2_X1 U6401 ( .A1(n4894), .A2(SI_7_), .ZN(n4895) );
  MUX2_X1 U6402 ( .A(n6570), .B(n6568), .S(n4871), .Z(n4897) );
  INV_X1 U6403 ( .A(SI_8_), .ZN(n4896) );
  NAND2_X1 U6404 ( .A1(n4897), .A2(n4896), .ZN(n4900) );
  INV_X1 U6405 ( .A(n4897), .ZN(n4898) );
  NAND2_X1 U6406 ( .A1(n4898), .A2(SI_8_), .ZN(n4899) );
  NAND2_X1 U6407 ( .A1(n4900), .A2(n4899), .ZN(n5131) );
  MUX2_X1 U6408 ( .A(n6579), .B(n6593), .S(n4871), .Z(n4902) );
  INV_X1 U6409 ( .A(SI_9_), .ZN(n4901) );
  NAND2_X1 U6410 ( .A1(n4902), .A2(n4901), .ZN(n4905) );
  INV_X1 U6411 ( .A(n4902), .ZN(n4903) );
  NAND2_X1 U6412 ( .A1(n4903), .A2(SI_9_), .ZN(n4904) );
  NAND2_X1 U6413 ( .A1(n4906), .A2(n4905), .ZN(n5160) );
  MUX2_X1 U6414 ( .A(n6601), .B(n6599), .S(n4401), .Z(n4908) );
  INV_X1 U6415 ( .A(SI_10_), .ZN(n4907) );
  NAND2_X1 U6416 ( .A1(n4908), .A2(n4907), .ZN(n4911) );
  INV_X1 U6417 ( .A(n4908), .ZN(n4909) );
  NAND2_X1 U6418 ( .A1(n4909), .A2(SI_10_), .ZN(n4910) );
  MUX2_X1 U6419 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4401), .Z(n4913) );
  XNOR2_X1 U6420 ( .A(n4913), .B(n9429), .ZN(n5175) );
  INV_X1 U6421 ( .A(n5175), .ZN(n4915) );
  NAND2_X1 U6422 ( .A1(n4913), .A2(SI_11_), .ZN(n4914) );
  MUX2_X1 U6423 ( .A(n6670), .B(n6668), .S(n4401), .Z(n4916) );
  NAND2_X1 U6424 ( .A1(n4916), .A2(n9439), .ZN(n4919) );
  INV_X1 U6425 ( .A(n4916), .ZN(n4917) );
  NAND2_X1 U6426 ( .A1(n4917), .A2(SI_12_), .ZN(n4918) );
  NAND2_X1 U6427 ( .A1(n4919), .A2(n4918), .ZN(n5186) );
  MUX2_X1 U6428 ( .A(n6734), .B(n4920), .S(n4401), .Z(n4921) );
  NAND2_X1 U6429 ( .A1(n4921), .A2(n9469), .ZN(n4924) );
  INV_X1 U6430 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6431 ( .A1(n4922), .A2(SI_13_), .ZN(n4923) );
  NAND2_X1 U6432 ( .A1(n4925), .A2(n4924), .ZN(n5215) );
  MUX2_X1 U6433 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4401), .Z(n4926) );
  XNOR2_X1 U6434 ( .A(n4926), .B(n9522), .ZN(n5214) );
  INV_X1 U6435 ( .A(n5214), .ZN(n4928) );
  NAND2_X1 U6436 ( .A1(n4926), .A2(SI_14_), .ZN(n4927) );
  MUX2_X1 U6437 ( .A(n6960), .B(n6962), .S(n4401), .Z(n4929) );
  NAND2_X1 U6438 ( .A1(n4929), .A2(n9523), .ZN(n4932) );
  INV_X1 U6439 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6440 ( .A1(n4930), .A2(SI_15_), .ZN(n4931) );
  NAND2_X1 U6441 ( .A1(n4932), .A2(n4931), .ZN(n5228) );
  MUX2_X1 U6442 ( .A(n7067), .B(n4933), .S(n4401), .Z(n4934) );
  NAND2_X1 U6443 ( .A1(n4934), .A2(n9525), .ZN(n4937) );
  INV_X1 U6444 ( .A(n4934), .ZN(n4935) );
  NAND2_X1 U6445 ( .A1(n4935), .A2(SI_16_), .ZN(n4936) );
  MUX2_X1 U6446 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4401), .Z(n4938) );
  XNOR2_X1 U6447 ( .A(n4938), .B(n9502), .ZN(n5258) );
  INV_X1 U6448 ( .A(n5258), .ZN(n4940) );
  NAND2_X1 U6449 ( .A1(n4938), .A2(SI_17_), .ZN(n4939) );
  MUX2_X1 U6450 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4401), .Z(n4942) );
  XNOR2_X1 U6451 ( .A(n4942), .B(SI_18_), .ZN(n5271) );
  INV_X1 U6452 ( .A(n5271), .ZN(n4941) );
  NAND2_X1 U6453 ( .A1(n5272), .A2(n4941), .ZN(n4944) );
  NAND2_X1 U6454 ( .A1(n4942), .A2(SI_18_), .ZN(n4943) );
  MUX2_X1 U6455 ( .A(n7344), .B(n7346), .S(n4401), .Z(n4945) );
  NAND2_X1 U6456 ( .A1(n4945), .A2(n9539), .ZN(n4948) );
  INV_X1 U6457 ( .A(n4945), .ZN(n4946) );
  NAND2_X1 U6458 ( .A1(n4946), .A2(SI_19_), .ZN(n4947) );
  NAND2_X1 U6459 ( .A1(n4948), .A2(n4947), .ZN(n5286) );
  MUX2_X1 U6460 ( .A(n7432), .B(n7445), .S(n4401), .Z(n4949) );
  NAND2_X1 U6461 ( .A1(n4949), .A2(n9513), .ZN(n4952) );
  INV_X1 U6462 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6463 ( .A1(n4950), .A2(SI_20_), .ZN(n4951) );
  MUX2_X1 U6464 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4401), .Z(n4956) );
  XNOR2_X1 U6465 ( .A(n4956), .B(n4954), .ZN(n5304) );
  INV_X1 U6466 ( .A(n5304), .ZN(n4955) );
  NAND2_X1 U6467 ( .A1(n4956), .A2(SI_21_), .ZN(n4957) );
  MUX2_X1 U6468 ( .A(n7946), .B(n7610), .S(n4401), .Z(n4958) );
  INV_X1 U6469 ( .A(SI_22_), .ZN(n9473) );
  NAND2_X1 U6470 ( .A1(n4958), .A2(n9473), .ZN(n4961) );
  INV_X1 U6471 ( .A(n4958), .ZN(n4959) );
  NAND2_X1 U6472 ( .A1(n4959), .A2(SI_22_), .ZN(n4960) );
  NAND2_X1 U6473 ( .A1(n4961), .A2(n4960), .ZN(n5317) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n4963) );
  INV_X1 U6475 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4962) );
  MUX2_X1 U6476 ( .A(n4963), .B(n4962), .S(n4401), .Z(n4965) );
  NAND2_X1 U6477 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  INV_X1 U6478 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6479 ( .A1(n4966), .A2(SI_23_), .ZN(n4967) );
  NAND2_X1 U6480 ( .A1(n5331), .A2(n5330), .ZN(n4969) );
  MUX2_X1 U6481 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4401), .Z(n4971) );
  INV_X1 U6482 ( .A(SI_24_), .ZN(n4970) );
  XNOR2_X1 U6483 ( .A(n4971), .B(n4970), .ZN(n5343) );
  NAND2_X1 U6484 ( .A1(n4971), .A2(SI_24_), .ZN(n4972) );
  INV_X1 U6485 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7794) );
  MUX2_X1 U6486 ( .A(n7797), .B(n7794), .S(n4401), .Z(n4973) );
  INV_X1 U6487 ( .A(SI_25_), .ZN(n9537) );
  NAND2_X1 U6488 ( .A1(n4973), .A2(n9537), .ZN(n4976) );
  INV_X1 U6489 ( .A(n4973), .ZN(n4974) );
  NAND2_X1 U6490 ( .A1(n4974), .A2(SI_25_), .ZN(n4975) );
  NAND2_X1 U6491 ( .A1(n4976), .A2(n4975), .ZN(n5354) );
  INV_X1 U6492 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n4977) );
  MUX2_X1 U6493 ( .A(n4977), .B(n7860), .S(n4401), .Z(n4978) );
  NAND2_X1 U6494 ( .A1(n4978), .A2(n9499), .ZN(n4981) );
  INV_X1 U6495 ( .A(n4978), .ZN(n4979) );
  NAND2_X1 U6496 ( .A1(n4979), .A2(SI_26_), .ZN(n4980) );
  INV_X1 U6497 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n4984) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n4983) );
  MUX2_X1 U6499 ( .A(n4984), .B(n4983), .S(n4401), .Z(n4985) );
  INV_X1 U6500 ( .A(SI_27_), .ZN(n9468) );
  NAND2_X1 U6501 ( .A1(n4985), .A2(n9468), .ZN(n4988) );
  INV_X1 U6502 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6503 ( .A1(n4986), .A2(SI_27_), .ZN(n4987) );
  MUX2_X1 U6504 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4401), .Z(n4989) );
  XNOR2_X1 U6505 ( .A(n4989), .B(n9528), .ZN(n5390) );
  INV_X1 U6506 ( .A(n4989), .ZN(n4990) );
  MUX2_X1 U6507 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4401), .Z(n4991) );
  INV_X1 U6508 ( .A(SI_29_), .ZN(n4992) );
  XNOR2_X1 U6509 ( .A(n4991), .B(n4992), .ZN(n5405) );
  NAND2_X1 U6510 ( .A1(n5404), .A2(n5405), .ZN(n4995) );
  INV_X1 U6511 ( .A(n4991), .ZN(n4993) );
  NAND2_X1 U6512 ( .A1(n4993), .A2(n4992), .ZN(n4994) );
  MUX2_X1 U6513 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4401), .Z(n5419) );
  INV_X1 U6514 ( .A(SI_30_), .ZN(n5421) );
  XNOR2_X1 U6515 ( .A(n5419), .B(n5421), .ZN(n4996) );
  NOR2_X1 U6516 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4999) );
  NAND4_X1 U6517 ( .A1(n4999), .A2(n4998), .A3(n4829), .A4(n4997), .ZN(n5004)
         );
  NAND4_X1 U6518 ( .A1(n4859), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n5003)
         );
  NOR2_X1 U6519 ( .A1(n5004), .A2(n5003), .ZN(n5005) );
  NAND2_X1 U6520 ( .A1(n5009), .A2(n5008), .ZN(n5016) );
  NAND2_X2 U6521 ( .A1(n6700), .A2(n6539), .ZN(n5117) );
  NAND2_X1 U6522 ( .A1(n8646), .A2(n5424), .ZN(n5015) );
  NAND2_X1 U6523 ( .A1(n4314), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5014) );
  INV_X1 U6524 ( .A(n5016), .ZN(n5018) );
  INV_X1 U6525 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6526 ( .A1(n5018), .A2(n5017), .ZN(n5021) );
  NAND2_X1 U6527 ( .A1(n5016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5019) );
  MUX2_X1 U6528 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5019), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5020) );
  XNOR2_X2 U6529 ( .A(n5022), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8501) );
  AND2_X4 U6530 ( .A1(n8503), .A2(n5023), .ZN(n5239) );
  NAND2_X1 U6531 ( .A1(n5239), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5027) );
  AND2_X2 U6532 ( .A1(n8501), .A2(n5024), .ZN(n5067) );
  NAND2_X1 U6533 ( .A1(n5067), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6534 ( .A1(n4319), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6535 ( .A1(n5239), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U6536 ( .A1(n5409), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6537 ( .A1(n4320), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5028) );
  INV_X1 U6538 ( .A(n8178), .ZN(n6563) );
  NOR2_X1 U6539 ( .A1(n6563), .A2(n7463), .ZN(n5418) );
  NAND2_X1 U6540 ( .A1(n5067), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6541 ( .A1(n4323), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6542 ( .A1(n5239), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6543 ( .A1(n4319), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5031) );
  AND4_X2 U6544 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5031), .ZN(n6915)
         );
  INV_X1 U6545 ( .A(SI_0_), .ZN(n5036) );
  INV_X1 U6546 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5035) );
  OAI21_X1 U6547 ( .B1(n4401), .B2(n5036), .A(n5035), .ZN(n5037) );
  AND2_X1 U6548 ( .A1(n5038), .A2(n5037), .ZN(n8514) );
  MUX2_X1 U6549 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8514), .S(n6700), .Z(n9951) );
  NAND2_X1 U6550 ( .A1(n5067), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6551 ( .A1(n5068), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6552 ( .A1(n5074), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6553 ( .A1(n4318), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5039) );
  XNOR2_X1 U6554 ( .A(n5044), .B(n5043), .ZN(n6554) );
  NAND2_X1 U6555 ( .A1(n4313), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5047) );
  INV_X1 U6556 ( .A(n8109), .ZN(n5045) );
  NAND2_X1 U6557 ( .A1(n5048), .A2(n6448), .ZN(n5580) );
  NAND2_X1 U6558 ( .A1(n5445), .A2(n5580), .ZN(n9919) );
  INV_X1 U6559 ( .A(n9919), .ZN(n5060) );
  NAND2_X1 U6560 ( .A1(n4324), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6561 ( .A1(n5067), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6562 ( .A1(n4319), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6563 ( .A1(n5239), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5049) );
  NAND4_X2 U6564 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5637)
         );
  INV_X1 U6565 ( .A(n5637), .ZN(n6935) );
  XNOR2_X1 U6566 ( .A(n5054), .B(n5053), .ZN(n6546) );
  NAND2_X1 U6567 ( .A1(n5204), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5058) );
  INV_X4 U6568 ( .A(n6700), .ZN(n6574) );
  OR2_X1 U6569 ( .A1(n5055), .A2(n8498), .ZN(n5056) );
  XNOR2_X1 U6570 ( .A(n5056), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U6571 ( .A1(n6574), .A2(n8120), .ZN(n5057) );
  NAND2_X1 U6572 ( .A1(n5637), .A2(n9968), .ZN(n5446) );
  NAND2_X2 U6573 ( .A1(n5447), .A2(n5446), .ZN(n9933) );
  INV_X1 U6574 ( .A(n9933), .ZN(n5059) );
  NAND2_X1 U6575 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  NAND2_X1 U6576 ( .A1(n5061), .A2(n5447), .ZN(n9905) );
  XNOR2_X1 U6577 ( .A(n5063), .B(n5062), .ZN(n6542) );
  NAND2_X1 U6578 ( .A1(n4314), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6579 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4352), .ZN(n5064) );
  XNOR2_X1 U6580 ( .A(n5064), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U6581 ( .A1(n6574), .A2(n6824), .ZN(n5065) );
  INV_X1 U6582 ( .A(n4312), .ZN(n9973) );
  NAND2_X1 U6583 ( .A1(n5067), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5072) );
  INV_X1 U6584 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U6585 ( .A1(n4323), .A2(n9911), .ZN(n5071) );
  NAND2_X1 U6586 ( .A1(n4320), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6587 ( .A1(n5239), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5069) );
  NAND4_X1 U6588 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9835)
         );
  XNOR2_X1 U6589 ( .A(n9973), .B(n9835), .ZN(n9904) );
  INV_X1 U6590 ( .A(n9904), .ZN(n5583) );
  NAND2_X1 U6591 ( .A1(n9905), .A2(n5583), .ZN(n5073) );
  INV_X1 U6592 ( .A(n9835), .ZN(n6453) );
  NAND2_X1 U6593 ( .A1(n6453), .A2(n4312), .ZN(n5436) );
  NAND2_X1 U6594 ( .A1(n5073), .A2(n5436), .ZN(n7089) );
  NAND2_X1 U6595 ( .A1(n5239), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6596 ( .A1(n5067), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6597 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5085) );
  OAI21_X1 U6598 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5085), .ZN(n9815) );
  INV_X1 U6599 ( .A(n9815), .ZN(n7086) );
  NAND2_X1 U6600 ( .A1(n4324), .A2(n7086), .ZN(n5076) );
  NAND2_X1 U6601 ( .A1(n4320), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5075) );
  INV_X1 U6602 ( .A(n8102), .ZN(n6456) );
  NAND2_X1 U6603 ( .A1(n4314), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6604 ( .A1(n5081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U6605 ( .A(n5082), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U6606 ( .A1(n6574), .A2(n6823), .ZN(n5083) );
  NAND2_X1 U6607 ( .A1(n6456), .A2(n9811), .ZN(n5437) );
  NAND2_X1 U6608 ( .A1(n5437), .A2(n9889), .ZN(n7084) );
  NAND2_X1 U6609 ( .A1(n4345), .A2(n9889), .ZN(n5100) );
  NAND2_X1 U6610 ( .A1(n5239), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6611 ( .A1(n5067), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5089) );
  NOR2_X1 U6612 ( .A1(n5085), .A2(n7021), .ZN(n5101) );
  AND2_X1 U6613 ( .A1(n5085), .A2(n7021), .ZN(n5086) );
  NOR2_X1 U6614 ( .A1(n5101), .A2(n5086), .ZN(n7015) );
  NAND2_X1 U6615 ( .A1(n4323), .A2(n7015), .ZN(n5088) );
  NAND2_X1 U6616 ( .A1(n4320), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5087) );
  NAND4_X1 U6617 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n8101)
         );
  INV_X1 U6618 ( .A(n8101), .ZN(n5099) );
  XNOR2_X1 U6619 ( .A(n5092), .B(n5091), .ZN(n6549) );
  NAND2_X1 U6620 ( .A1(n5204), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6621 ( .A1(n5093), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5094) );
  MUX2_X1 U6622 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5094), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5096) );
  NOR2_X1 U6623 ( .A1(n5093), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5119) );
  INV_X1 U6624 ( .A(n5119), .ZN(n5095) );
  NAND2_X1 U6625 ( .A1(n6574), .A2(n6821), .ZN(n5097) );
  NAND2_X1 U6626 ( .A1(n5099), .A2(n4315), .ZN(n5438) );
  NAND2_X1 U6627 ( .A1(n5239), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6628 ( .A1(n5067), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6629 ( .A1(n5101), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5123) );
  OR2_X1 U6630 ( .A1(n5101), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6631 ( .A1(n5123), .A2(n5102), .ZN(n9862) );
  INV_X1 U6632 ( .A(n9862), .ZN(n7149) );
  NAND2_X1 U6633 ( .A1(n4324), .A2(n7149), .ZN(n5104) );
  NAND2_X1 U6634 ( .A1(n4320), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5103) );
  NAND4_X1 U6635 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n8100)
         );
  INV_X1 U6636 ( .A(n8100), .ZN(n5112) );
  OR2_X1 U6637 ( .A1(n5119), .A2(n8498), .ZN(n5107) );
  XNOR2_X1 U6638 ( .A(n5107), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U6639 ( .A1(n5204), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6574), .B2(
        n6820), .ZN(n5111) );
  OR2_X1 U6640 ( .A1(n5117), .A2(n6557), .ZN(n5110) );
  NAND2_X1 U6641 ( .A1(n5112), .A2(n9858), .ZN(n7071) );
  INV_X1 U6642 ( .A(n9858), .ZN(n7152) );
  NAND2_X1 U6643 ( .A1(n7152), .A2(n8100), .ZN(n5460) );
  INV_X1 U6644 ( .A(n7113), .ZN(n5113) );
  NOR2_X1 U6645 ( .A1(n7117), .A2(n5113), .ZN(n5114) );
  XNOR2_X1 U6646 ( .A(n5116), .B(n5115), .ZN(n6561) );
  NAND2_X1 U6647 ( .A1(n5119), .A2(n5118), .ZN(n5133) );
  NAND2_X1 U6648 ( .A1(n5133), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U6649 ( .A(n5120), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U6650 ( .A1(n5204), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6574), .B2(
        n6843), .ZN(n5121) );
  NAND2_X1 U6651 ( .A1(n5239), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6652 ( .A1(n5067), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6653 ( .A1(n5123), .A2(n5122), .ZN(n5124) );
  AND2_X1 U6654 ( .A1(n5137), .A2(n5124), .ZN(n7261) );
  NAND2_X1 U6655 ( .A1(n4324), .A2(n7261), .ZN(n5126) );
  NAND2_X1 U6656 ( .A1(n4319), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5125) );
  NAND4_X1 U6657 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n8099)
         );
  INV_X1 U6658 ( .A(n8099), .ZN(n7231) );
  NAND2_X1 U6659 ( .A1(n7231), .A2(n7080), .ZN(n5462) );
  INV_X1 U6660 ( .A(n7070), .ZN(n5129) );
  INV_X1 U6661 ( .A(n7071), .ZN(n5440) );
  NOR2_X1 U6662 ( .A1(n5129), .A2(n5440), .ZN(n5130) );
  XNOR2_X1 U6663 ( .A(n5132), .B(n5131), .ZN(n6566) );
  NAND2_X1 U6664 ( .A1(n6566), .A2(n5424), .ZN(n5136) );
  NAND2_X1 U6665 ( .A1(n5146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U6666 ( .A(n5134), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6854) );
  AOI22_X1 U6667 ( .A1(n5204), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6574), .B2(
        n6854), .ZN(n5135) );
  NAND2_X1 U6668 ( .A1(n5136), .A2(n5135), .ZN(n7240) );
  NAND2_X1 U6669 ( .A1(n5239), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6670 ( .A1(n5067), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6671 ( .A1(n5137), .A2(n9471), .ZN(n5138) );
  NAND2_X1 U6672 ( .A1(n5151), .A2(n5138), .ZN(n7236) );
  INV_X1 U6673 ( .A(n7236), .ZN(n5139) );
  NAND2_X1 U6674 ( .A1(n4323), .A2(n5139), .ZN(n5141) );
  NAND2_X1 U6675 ( .A1(n4319), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5140) );
  NAND4_X1 U6676 ( .A1(n5143), .A2(n5142), .A3(n5141), .A4(n5140), .ZN(n8097)
         );
  XNOR2_X1 U6677 ( .A(n7240), .B(n8097), .ZN(n7178) );
  INV_X1 U6678 ( .A(n8097), .ZN(n7404) );
  NAND2_X1 U6679 ( .A1(n7240), .A2(n7404), .ZN(n5467) );
  XNOR2_X1 U6680 ( .A(n5145), .B(n5144), .ZN(n6578) );
  NAND2_X1 U6681 ( .A1(n6578), .A2(n5424), .ZN(n5149) );
  OR2_X1 U6682 ( .A1(n5162), .A2(n8498), .ZN(n5147) );
  XNOR2_X1 U6683 ( .A(n5147), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U6684 ( .A1(n5204), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6574), .B2(
        n6921), .ZN(n5148) );
  NAND2_X1 U6685 ( .A1(n5149), .A2(n5148), .ZN(n7475) );
  NAND2_X1 U6686 ( .A1(n5239), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6687 ( .A1(n5067), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5155) );
  AND2_X1 U6688 ( .A1(n5151), .A2(n5150), .ZN(n5152) );
  NOR2_X1 U6689 ( .A1(n5168), .A2(n5152), .ZN(n7409) );
  NAND2_X1 U6690 ( .A1(n4323), .A2(n7409), .ZN(n5154) );
  NAND2_X1 U6691 ( .A1(n4320), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5153) );
  NAND4_X1 U6692 ( .A1(n5156), .A2(n5155), .A3(n5154), .A4(n5153), .ZN(n8096)
         );
  INV_X1 U6693 ( .A(n8096), .ZN(n5157) );
  OR2_X1 U6694 ( .A1(n7475), .A2(n5157), .ZN(n5472) );
  NAND2_X1 U6695 ( .A1(n7475), .A2(n5157), .ZN(n5158) );
  NAND2_X1 U6696 ( .A1(n5472), .A2(n5158), .ZN(n7316) );
  INV_X1 U6697 ( .A(n7316), .ZN(n5586) );
  INV_X1 U6698 ( .A(n5158), .ZN(n5474) );
  XNOR2_X1 U6699 ( .A(n5160), .B(n5159), .ZN(n6598) );
  NAND2_X1 U6700 ( .A1(n6598), .A2(n5424), .ZN(n5167) );
  NAND2_X1 U6701 ( .A1(n5162), .A2(n5161), .ZN(n5188) );
  NAND2_X1 U6702 ( .A1(n5188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6703 ( .A1(n5164), .A2(n5163), .ZN(n5176) );
  OR2_X1 U6704 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  AOI22_X1 U6705 ( .A1(n5204), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6574), .B2(
        n7189), .ZN(n5166) );
  NAND2_X1 U6706 ( .A1(n5239), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6707 ( .A1(n5067), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5172) );
  OR2_X1 U6708 ( .A1(n5168), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6709 ( .A1(n5168), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5180) );
  AND2_X1 U6710 ( .A1(n5169), .A2(n5180), .ZN(n9876) );
  NAND2_X1 U6711 ( .A1(n4324), .A2(n9876), .ZN(n5171) );
  NAND2_X1 U6712 ( .A1(n4319), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5170) );
  NAND4_X1 U6713 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n8095)
         );
  INV_X1 U6714 ( .A(n8095), .ZN(n5174) );
  NAND2_X1 U6715 ( .A1(n9877), .A2(n5174), .ZN(n5478) );
  NAND2_X1 U6716 ( .A1(n5473), .A2(n5478), .ZN(n7592) );
  NAND2_X1 U6717 ( .A1(n5176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5177) );
  XNOR2_X1 U6718 ( .A(n5177), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8136) );
  AOI22_X1 U6719 ( .A1(n5204), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6574), .B2(
        n8136), .ZN(n5178) );
  NAND2_X1 U6720 ( .A1(n5067), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6721 ( .A1(n5180), .A2(n9816), .ZN(n5181) );
  NAND2_X1 U6722 ( .A1(n5193), .A2(n5181), .ZN(n9831) );
  INV_X1 U6723 ( .A(n9831), .ZN(n7438) );
  NAND2_X1 U6724 ( .A1(n4323), .A2(n7438), .ZN(n5184) );
  NAND2_X1 U6725 ( .A1(n4320), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6726 ( .A1(n5239), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5182) );
  NAND4_X1 U6727 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n8094)
         );
  INV_X1 U6728 ( .A(n8094), .ZN(n5199) );
  NAND2_X1 U6729 ( .A1(n9827), .A2(n5199), .ZN(n5577) );
  XNOR2_X1 U6730 ( .A(n5187), .B(n5186), .ZN(n6667) );
  NAND2_X1 U6731 ( .A1(n6667), .A2(n5424), .ZN(n5191) );
  NAND2_X1 U6732 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6733 ( .A(n5189), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7352) );
  AOI22_X1 U6734 ( .A1(n5204), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6574), .B2(
        n7352), .ZN(n5190) );
  NAND2_X1 U6735 ( .A1(n5191), .A2(n5190), .ZN(n7663) );
  NAND2_X1 U6736 ( .A1(n5239), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6737 ( .A1(n5067), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5197) );
  AND2_X1 U6738 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  NOR2_X1 U6739 ( .A1(n5207), .A2(n5194), .ZN(n7658) );
  NAND2_X1 U6740 ( .A1(n4324), .A2(n7658), .ZN(n5196) );
  NAND2_X1 U6741 ( .A1(n4319), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5195) );
  NAND4_X1 U6742 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n8093)
         );
  INV_X1 U6743 ( .A(n8093), .ZN(n5200) );
  OR2_X1 U6744 ( .A1(n7663), .A2(n5200), .ZN(n5576) );
  OR2_X1 U6745 ( .A1(n9827), .A2(n5199), .ZN(n7520) );
  AND2_X1 U6746 ( .A1(n5576), .A2(n7520), .ZN(n5483) );
  NAND2_X1 U6747 ( .A1(n7663), .A2(n5200), .ZN(n5575) );
  XNOR2_X1 U6748 ( .A(n5202), .B(n5201), .ZN(n6732) );
  NAND2_X1 U6749 ( .A1(n6732), .A2(n5424), .ZN(n5206) );
  OAI21_X1 U6750 ( .B1(n5203), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6751 ( .A(n5217), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7452) );
  AOI22_X1 U6752 ( .A1(n4314), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6574), .B2(
        n7452), .ZN(n5205) );
  NAND2_X1 U6753 ( .A1(n5239), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6754 ( .A1(n5409), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6755 ( .A1(n5207), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5221) );
  OR2_X1 U6756 ( .A1(n5207), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5208) );
  AND2_X1 U6757 ( .A1(n5221), .A2(n5208), .ZN(n7706) );
  NAND2_X1 U6758 ( .A1(n4323), .A2(n7706), .ZN(n5210) );
  NAND2_X1 U6759 ( .A1(n4320), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5209) );
  NAND4_X1 U6760 ( .A1(n5212), .A2(n5211), .A3(n5210), .A4(n5209), .ZN(n8092)
         );
  INV_X1 U6761 ( .A(n8092), .ZN(n6467) );
  OR2_X1 U6762 ( .A1(n7575), .A2(n6467), .ZN(n5490) );
  NAND2_X1 U6763 ( .A1(n7575), .A2(n6467), .ZN(n5489) );
  XNOR2_X1 U6764 ( .A(n5215), .B(n5214), .ZN(n6759) );
  NAND2_X1 U6765 ( .A1(n6759), .A2(n5424), .ZN(n5220) );
  NAND2_X1 U6766 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NAND2_X1 U6767 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6768 ( .A(n5231), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7644) );
  AOI22_X1 U6769 ( .A1(n6574), .A2(n7644), .B1(n4314), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6770 ( .A1(n5067), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6771 ( .A1(n5221), .A2(n9441), .ZN(n5222) );
  NAND2_X1 U6772 ( .A1(n5237), .A2(n5222), .ZN(n9642) );
  INV_X1 U6773 ( .A(n9642), .ZN(n7680) );
  NAND2_X1 U6774 ( .A1(n4324), .A2(n7680), .ZN(n5225) );
  NAND2_X1 U6775 ( .A1(n4320), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6776 ( .A1(n5239), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5223) );
  NAND4_X1 U6777 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n8091)
         );
  INV_X1 U6778 ( .A(n8091), .ZN(n5227) );
  OR2_X1 U6779 ( .A1(n9638), .A2(n5227), .ZN(n5495) );
  NAND2_X1 U6780 ( .A1(n9638), .A2(n5227), .ZN(n5494) );
  INV_X1 U6781 ( .A(n7674), .ZN(n5591) );
  NAND2_X1 U6782 ( .A1(n7673), .A2(n5495), .ZN(n7738) );
  XNOR2_X1 U6783 ( .A(n5229), .B(n5228), .ZN(n6959) );
  NAND2_X1 U6784 ( .A1(n6959), .A2(n5424), .ZN(n5235) );
  NAND2_X1 U6785 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  NAND2_X1 U6786 ( .A1(n5232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5233) );
  XNOR2_X1 U6787 ( .A(n5233), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7807) );
  AOI22_X1 U6788 ( .A1(n7807), .A2(n6574), .B1(n4314), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6789 ( .A1(n5067), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5243) );
  INV_X1 U6790 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7905) );
  NAND2_X1 U6791 ( .A1(n5237), .A2(n7905), .ZN(n5238) );
  AND2_X1 U6792 ( .A1(n5252), .A2(n5238), .ZN(n7908) );
  NAND2_X1 U6793 ( .A1(n4324), .A2(n7908), .ZN(n5242) );
  NAND2_X1 U6794 ( .A1(n4320), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6795 ( .A1(n5239), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5240) );
  NAND4_X1 U6796 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n8090)
         );
  INV_X1 U6797 ( .A(n8090), .ZN(n5244) );
  OR2_X1 U6798 ( .A1(n7744), .A2(n5244), .ZN(n5497) );
  NAND2_X1 U6799 ( .A1(n7744), .A2(n5244), .ZN(n5498) );
  NAND2_X1 U6800 ( .A1(n5497), .A2(n5498), .ZN(n7734) );
  INV_X1 U6801 ( .A(n7734), .ZN(n7737) );
  XNOR2_X1 U6802 ( .A(n5246), .B(n5245), .ZN(n7059) );
  NAND2_X1 U6803 ( .A1(n7059), .A2(n5424), .ZN(n5251) );
  NOR2_X1 U6804 ( .A1(n5247), .A2(n8498), .ZN(n5248) );
  MUX2_X1 U6805 ( .A(n8498), .B(n5248), .S(P2_IR_REG_16__SCAN_IN), .Z(n5249)
         );
  AOI22_X1 U6806 ( .A1(n4314), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6574), .B2(
        n7877), .ZN(n5250) );
  NAND2_X1 U6807 ( .A1(n5239), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6808 ( .A1(n5067), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6809 ( .A1(n5252), .A2(n9544), .ZN(n5253) );
  AND2_X1 U6810 ( .A1(n5277), .A2(n5253), .ZN(n8012) );
  NAND2_X1 U6811 ( .A1(n4324), .A2(n8012), .ZN(n5255) );
  NAND2_X1 U6812 ( .A1(n4319), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5254) );
  NAND4_X1 U6813 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n8089)
         );
  INV_X1 U6814 ( .A(n8089), .ZN(n7896) );
  OR2_X1 U6815 ( .A1(n8459), .A2(n7896), .ZN(n5502) );
  NAND2_X1 U6816 ( .A1(n8459), .A2(n7896), .ZN(n5501) );
  INV_X1 U6817 ( .A(n7827), .ZN(n7832) );
  XNOR2_X1 U6818 ( .A(n5259), .B(n5258), .ZN(n7061) );
  NAND2_X1 U6819 ( .A1(n7061), .A2(n5424), .ZN(n5265) );
  NAND2_X1 U6820 ( .A1(n5260), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5261) );
  MUX2_X1 U6821 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5261), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5263) );
  AND2_X1 U6822 ( .A1(n5263), .A2(n5262), .ZN(n8150) );
  AOI22_X1 U6823 ( .A1(n5204), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6574), .B2(
        n8150), .ZN(n5264) );
  XNOR2_X1 U6824 ( .A(n5277), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U6825 ( .A1(n8372), .A2(n4323), .ZN(n5269) );
  NAND2_X1 U6826 ( .A1(n5239), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6827 ( .A1(n5067), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6828 ( .A1(n4320), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5266) );
  NAND4_X1 U6829 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n8088)
         );
  XNOR2_X1 U6830 ( .A(n8453), .B(n8056), .ZN(n8378) );
  XNOR2_X1 U6831 ( .A(n5272), .B(n5271), .ZN(n7243) );
  NAND2_X1 U6832 ( .A1(n7243), .A2(n5424), .ZN(n5275) );
  NAND2_X1 U6833 ( .A1(n5262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6834 ( .A(n5273), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8151) );
  AOI22_X1 U6835 ( .A1(n5204), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6574), .B2(
        n8151), .ZN(n5274) );
  INV_X1 U6836 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5276) );
  OAI21_X1 U6837 ( .B1(n5277), .B2(n9419), .A(n5276), .ZN(n5280) );
  AND2_X1 U6838 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5278) );
  NAND2_X1 U6839 ( .A1(n5280), .A2(n5290), .ZN(n8358) );
  OR2_X1 U6840 ( .A1(n5408), .A2(n8358), .ZN(n5284) );
  NAND2_X1 U6841 ( .A1(n5239), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6842 ( .A1(n5409), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6843 ( .A1(n4319), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5281) );
  NAND4_X1 U6844 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n8087)
         );
  OR2_X1 U6845 ( .A1(n8357), .A2(n7970), .ZN(n5513) );
  NAND2_X1 U6846 ( .A1(n8357), .A2(n7970), .ZN(n5506) );
  NAND2_X1 U6847 ( .A1(n5513), .A2(n5506), .ZN(n8349) );
  NOR2_X1 U6848 ( .A1(n8453), .A2(n8056), .ZN(n8350) );
  NOR2_X1 U6849 ( .A1(n8349), .A2(n8350), .ZN(n5285) );
  NAND2_X1 U6850 ( .A1(n8348), .A2(n5285), .ZN(n8351) );
  NAND2_X1 U6851 ( .A1(n8351), .A2(n5506), .ZN(n8338) );
  XNOR2_X1 U6852 ( .A(n5287), .B(n5286), .ZN(n7342) );
  NAND2_X1 U6853 ( .A1(n7342), .A2(n5424), .ZN(n5289) );
  AOI22_X1 U6854 ( .A1(n5204), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6574), .B2(
        n8254), .ZN(n5288) );
  INV_X1 U6855 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6856 ( .A1(n5290), .A2(n9481), .ZN(n5291) );
  NAND2_X1 U6857 ( .A1(n5309), .A2(n5291), .ZN(n7974) );
  OR2_X1 U6858 ( .A1(n7974), .A2(n5408), .ZN(n5293) );
  AOI22_X1 U6859 ( .A1(n5239), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n5067), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5292) );
  OAI211_X1 U6860 ( .C1(n5412), .C2(n5294), .A(n5293), .B(n5292), .ZN(n8086)
         );
  INV_X1 U6861 ( .A(n8086), .ZN(n8058) );
  OR2_X1 U6862 ( .A1(n8443), .A2(n8058), .ZN(n5514) );
  NAND2_X1 U6863 ( .A1(n8443), .A2(n8058), .ZN(n5515) );
  XNOR2_X1 U6864 ( .A(n5296), .B(n5295), .ZN(n7431) );
  NAND2_X1 U6865 ( .A1(n7431), .A2(n5424), .ZN(n5298) );
  NAND2_X1 U6866 ( .A1(n5204), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6867 ( .A(n5309), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U6868 ( .A1(n8330), .A2(n4324), .ZN(n5303) );
  INV_X1 U6869 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U6870 ( .A1(n5239), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6871 ( .A1(n5409), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5299) );
  OAI211_X1 U6872 ( .C1(n8487), .C2(n5412), .A(n5300), .B(n5299), .ZN(n5301)
         );
  INV_X1 U6873 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6874 ( .A1(n5303), .A2(n5302), .ZN(n8085) );
  INV_X1 U6875 ( .A(n8085), .ZN(n7985) );
  NAND2_X1 U6876 ( .A1(n8329), .A2(n7985), .ZN(n5519) );
  NAND2_X1 U6877 ( .A1(n5522), .A2(n5519), .ZN(n8322) );
  NAND2_X1 U6878 ( .A1(n8325), .A2(n5522), .ZN(n8309) );
  XNOR2_X1 U6879 ( .A(n5305), .B(n5304), .ZN(n7461) );
  NAND2_X1 U6880 ( .A1(n7461), .A2(n5424), .ZN(n5307) );
  NAND2_X1 U6881 ( .A1(n5204), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6882 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5308) );
  INV_X1 U6883 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8031) );
  INV_X1 U6884 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7990) );
  OAI21_X1 U6885 ( .B1(n5309), .B2(n8031), .A(n7990), .ZN(n5310) );
  AND2_X1 U6886 ( .A1(n5322), .A2(n5310), .ZN(n8315) );
  NAND2_X1 U6887 ( .A1(n8315), .A2(n4323), .ZN(n5316) );
  INV_X1 U6888 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6889 ( .A1(n5239), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U6890 ( .A1(n5409), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5311) );
  OAI211_X1 U6891 ( .C1(n5313), .C2(n5412), .A(n5312), .B(n5311), .ZN(n5314)
         );
  INV_X1 U6892 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6893 ( .A1(n5316), .A2(n5315), .ZN(n8084) );
  INV_X1 U6894 ( .A(n8084), .ZN(n6471) );
  XNOR2_X1 U6895 ( .A(n8433), .B(n6471), .ZN(n8310) );
  NAND2_X1 U6896 ( .A1(n8433), .A2(n6471), .ZN(n5518) );
  XNOR2_X1 U6897 ( .A(n5318), .B(n5317), .ZN(n7609) );
  NAND2_X1 U6898 ( .A1(n7609), .A2(n5424), .ZN(n5320) );
  NAND2_X1 U6899 ( .A1(n4314), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5319) );
  INV_X1 U6900 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U6901 ( .A1(n5322), .A2(n9530), .ZN(n5323) );
  AND2_X1 U6902 ( .A1(n5335), .A2(n5323), .ZN(n8301) );
  NAND2_X1 U6903 ( .A1(n8301), .A2(n4324), .ZN(n5329) );
  INV_X1 U6904 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6905 ( .A1(n4318), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6906 ( .A1(n5409), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5324) );
  OAI211_X1 U6907 ( .C1(n5326), .C2(n5412), .A(n5325), .B(n5324), .ZN(n5327)
         );
  INV_X1 U6908 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6909 ( .A1(n5329), .A2(n5328), .ZN(n8083) );
  INV_X1 U6910 ( .A(n8083), .ZN(n7964) );
  NAND2_X1 U6911 ( .A1(n8299), .A2(n7964), .ZN(n5511) );
  XNOR2_X1 U6912 ( .A(n5331), .B(n5330), .ZN(n7666) );
  NAND2_X1 U6913 ( .A1(n7666), .A2(n5424), .ZN(n5333) );
  NAND2_X1 U6914 ( .A1(n5204), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5332) );
  INV_X1 U6915 ( .A(n5335), .ZN(n5334) );
  NAND2_X1 U6916 ( .A1(n5335), .A2(n9531), .ZN(n5336) );
  NAND2_X1 U6917 ( .A1(n5347), .A2(n5336), .ZN(n8284) );
  OR2_X1 U6918 ( .A1(n8284), .A2(n5408), .ZN(n5342) );
  INV_X1 U6919 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6920 ( .A1(n5239), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6921 ( .A1(n5409), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5337) );
  OAI211_X1 U6922 ( .C1(n5339), .C2(n5412), .A(n5338), .B(n5337), .ZN(n5340)
         );
  INV_X1 U6923 ( .A(n5340), .ZN(n5341) );
  NAND2_X1 U6924 ( .A1(n5342), .A2(n5341), .ZN(n8082) );
  XNOR2_X1 U6925 ( .A(n8421), .B(n8082), .ZN(n8281) );
  INV_X1 U6926 ( .A(n8082), .ZN(n5533) );
  NAND2_X1 U6927 ( .A1(n8421), .A2(n5533), .ZN(n5512) );
  XNOR2_X1 U6928 ( .A(n5344), .B(n5343), .ZN(n7709) );
  NAND2_X1 U6929 ( .A1(n7709), .A2(n5424), .ZN(n5346) );
  NAND2_X1 U6930 ( .A1(n4314), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5345) );
  INV_X1 U6931 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U6932 ( .A1(n5347), .A2(n9504), .ZN(n5348) );
  AND2_X1 U6933 ( .A1(n5359), .A2(n5348), .ZN(n8272) );
  NAND2_X1 U6934 ( .A1(n8272), .A2(n4323), .ZN(n5353) );
  INV_X1 U6935 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U6936 ( .A1(n4318), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6937 ( .A1(n5067), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5349) );
  OAI211_X1 U6938 ( .C1(n8481), .C2(n5412), .A(n5350), .B(n5349), .ZN(n5351)
         );
  INV_X1 U6939 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6940 ( .A1(n8271), .A2(n8020), .ZN(n5535) );
  NAND2_X1 U6941 ( .A1(n5532), .A2(n5535), .ZN(n8267) );
  INV_X1 U6942 ( .A(n8267), .ZN(n8262) );
  XNOR2_X1 U6943 ( .A(n5355), .B(n5354), .ZN(n7793) );
  NAND2_X1 U6944 ( .A1(n7793), .A2(n5424), .ZN(n5357) );
  NAND2_X1 U6945 ( .A1(n5204), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5356) );
  INV_X1 U6946 ( .A(n5359), .ZN(n5358) );
  NAND2_X1 U6947 ( .A1(n5358), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5370) );
  INV_X1 U6948 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U6949 ( .A1(n5359), .A2(n7999), .ZN(n5360) );
  NAND2_X1 U6950 ( .A1(n5370), .A2(n5360), .ZN(n7997) );
  INV_X1 U6951 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U6952 ( .A1(n5239), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6953 ( .A1(n5409), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5361) );
  OAI211_X1 U6954 ( .C1(n8477), .C2(n5412), .A(n5362), .B(n5361), .ZN(n5363)
         );
  INV_X1 U6955 ( .A(n5363), .ZN(n5364) );
  NAND2_X1 U6956 ( .A1(n5365), .A2(n5364), .ZN(n8080) );
  NAND2_X1 U6957 ( .A1(n8253), .A2(n8065), .ZN(n5433) );
  NAND2_X1 U6958 ( .A1(n7857), .A2(n5424), .ZN(n5369) );
  NAND2_X1 U6959 ( .A1(n5204), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5368) );
  INV_X1 U6960 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U6961 ( .A1(n5370), .A2(n9527), .ZN(n5371) );
  NAND2_X1 U6962 ( .A1(n8070), .A2(n4324), .ZN(n5377) );
  INV_X1 U6963 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6964 ( .A1(n5239), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6965 ( .A1(n5409), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5372) );
  OAI211_X1 U6966 ( .C1(n5374), .C2(n5412), .A(n5373), .B(n5372), .ZN(n5375)
         );
  INV_X1 U6967 ( .A(n5375), .ZN(n5376) );
  NAND2_X1 U6968 ( .A1(n5377), .A2(n5376), .ZN(n8079) );
  INV_X1 U6969 ( .A(n8079), .ZN(n7953) );
  NAND2_X1 U6970 ( .A1(n8406), .A2(n7953), .ZN(n8218) );
  INV_X1 U6971 ( .A(n8232), .ZN(n5540) );
  NOR2_X1 U6972 ( .A1(n8228), .A2(n5540), .ZN(n5378) );
  NAND2_X1 U6973 ( .A1(n8509), .A2(n5424), .ZN(n5382) );
  NAND2_X1 U6974 ( .A1(n5204), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5381) );
  XNOR2_X1 U6975 ( .A(n5395), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U6976 ( .A1(n8223), .A2(n4323), .ZN(n5388) );
  INV_X1 U6977 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6978 ( .A1(n4318), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6979 ( .A1(n5409), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5383) );
  OAI211_X1 U6980 ( .C1(n5385), .C2(n5412), .A(n5384), .B(n5383), .ZN(n5386)
         );
  INV_X1 U6981 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6982 ( .A1(n5388), .A2(n5387), .ZN(n8078) );
  INV_X1 U6983 ( .A(n8078), .ZN(n6474) );
  NAND2_X1 U6984 ( .A1(n8401), .A2(n6474), .ZN(n5546) );
  INV_X1 U6985 ( .A(n8218), .ZN(n5543) );
  NOR2_X1 U6986 ( .A1(n8216), .A2(n5543), .ZN(n5389) );
  NAND2_X1 U6987 ( .A1(n8230), .A2(n5389), .ZN(n8215) );
  NAND2_X1 U6988 ( .A1(n8215), .A2(n5545), .ZN(n8201) );
  NAND2_X1 U6989 ( .A1(n8506), .A2(n5424), .ZN(n5393) );
  NAND2_X1 U6990 ( .A1(n5204), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5392) );
  INV_X1 U6991 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5394) );
  OAI21_X1 U6992 ( .B1(n5395), .B2(n9540), .A(n5394), .ZN(n5398) );
  INV_X1 U6993 ( .A(n5395), .ZN(n5397) );
  AND2_X1 U6994 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5396) );
  NAND2_X1 U6995 ( .A1(n5397), .A2(n5396), .ZN(n8191) );
  NAND2_X1 U6996 ( .A1(n5398), .A2(n8191), .ZN(n5797) );
  INV_X1 U6997 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U6998 ( .A1(n5239), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6999 ( .A1(n5409), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5399) );
  OAI211_X1 U7000 ( .C1(n8471), .C2(n5412), .A(n5400), .B(n5399), .ZN(n5401)
         );
  INV_X1 U7001 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U7002 ( .A1(n5403), .A2(n5402), .ZN(n8077) );
  NAND2_X1 U7003 ( .A1(n8201), .A2(n8204), .ZN(n8200) );
  NAND2_X1 U7004 ( .A1(n8200), .A2(n5550), .ZN(n6480) );
  NAND2_X1 U7005 ( .A1(n8638), .A2(n5424), .ZN(n5407) );
  NAND2_X1 U7006 ( .A1(n4314), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5406) );
  OR2_X1 U7007 ( .A1(n8191), .A2(n5408), .ZN(n5415) );
  INV_X1 U7008 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7009 ( .A1(n5409), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7010 ( .A1(n4318), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5410) );
  OAI211_X1 U7011 ( .C1(n5412), .C2(n6498), .A(n5411), .B(n5410), .ZN(n5413)
         );
  INV_X1 U7012 ( .A(n5413), .ZN(n5414) );
  NAND2_X1 U7013 ( .A1(n5415), .A2(n5414), .ZN(n8076) );
  INV_X1 U7014 ( .A(n8076), .ZN(n5416) );
  INV_X1 U7015 ( .A(n5560), .ZN(n5417) );
  NAND2_X1 U7016 ( .A1(n8196), .A2(n5416), .ZN(n5561) );
  MUX2_X1 U7017 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4401), .Z(n5422) );
  XNOR2_X1 U7018 ( .A(n5422), .B(SI_31_), .ZN(n5423) );
  NAND2_X1 U7019 ( .A1(n8654), .A2(n5424), .ZN(n5427) );
  NAND2_X1 U7020 ( .A1(n5204), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5426) );
  OR2_X1 U7021 ( .A1(n8175), .A2(n8178), .ZN(n5567) );
  NAND2_X1 U7022 ( .A1(n8182), .A2(n6595), .ZN(n5428) );
  NAND2_X1 U7023 ( .A1(n8175), .A2(n8178), .ZN(n5571) );
  XNOR2_X1 U7024 ( .A(n5430), .B(n7343), .ZN(n5431) );
  AOI21_X1 U7025 ( .B1(n9898), .B2(n6482), .A(n5431), .ZN(n5611) );
  NOR2_X1 U7026 ( .A1(n7463), .A2(n7343), .ZN(n5432) );
  INV_X1 U7027 ( .A(n5547), .ZN(n5555) );
  INV_X1 U7028 ( .A(n5570), .ZN(n5559) );
  NAND2_X1 U7029 ( .A1(n5437), .A2(n5438), .ZN(n5435) );
  NAND2_X1 U7030 ( .A1(n9889), .A2(n7113), .ZN(n5434) );
  MUX2_X1 U7031 ( .A(n5435), .B(n5434), .S(n5570), .Z(n5458) );
  AOI21_X1 U7032 ( .B1(n5437), .B2(n5436), .A(n5458), .ZN(n5441) );
  INV_X1 U7033 ( .A(n5438), .ZN(n5439) );
  NOR3_X1 U7034 ( .A1(n5441), .A2(n5440), .A3(n5439), .ZN(n5455) );
  INV_X1 U7035 ( .A(n5580), .ZN(n5443) );
  INV_X1 U7036 ( .A(n9951), .ZN(n6914) );
  NAND2_X1 U7037 ( .A1(n8104), .A2(n6914), .ZN(n5578) );
  INV_X1 U7038 ( .A(n5578), .ZN(n5442) );
  OAI211_X1 U7039 ( .C1(n5443), .C2(n5442), .A(n5447), .B(n5579), .ZN(n5444)
         );
  NAND2_X1 U7040 ( .A1(n5444), .A2(n5446), .ZN(n5451) );
  AOI21_X1 U7041 ( .B1(n5630), .B2(n5578), .A(n5445), .ZN(n5449) );
  NAND2_X1 U7042 ( .A1(n5580), .A2(n5446), .ZN(n5448) );
  OAI21_X1 U7043 ( .B1(n5449), .B2(n5448), .A(n5447), .ZN(n5450) );
  MUX2_X1 U7044 ( .A(n5451), .B(n5450), .S(n5570), .Z(n5453) );
  INV_X1 U7045 ( .A(n5458), .ZN(n5452) );
  NAND3_X1 U7046 ( .A1(n5453), .A2(n5452), .A3(n5583), .ZN(n5454) );
  OAI21_X1 U7047 ( .B1(n5455), .B2(n5559), .A(n5454), .ZN(n5461) );
  INV_X1 U7048 ( .A(n9889), .ZN(n5456) );
  AOI21_X1 U7049 ( .B1(n9973), .B2(n9835), .A(n5456), .ZN(n5457) );
  OAI211_X1 U7050 ( .C1(n5458), .C2(n5457), .A(n5460), .B(n7113), .ZN(n5459)
         );
  AOI22_X1 U7051 ( .A1(n5461), .A2(n5460), .B1(n5559), .B2(n5459), .ZN(n5466)
         );
  OAI21_X1 U7052 ( .B1(n7071), .B2(n5570), .A(n7070), .ZN(n5465) );
  MUX2_X1 U7053 ( .A(n5463), .B(n5462), .S(n5570), .Z(n5464) );
  OAI211_X1 U7054 ( .C1(n5466), .C2(n5465), .A(n7178), .B(n5464), .ZN(n5471)
         );
  INV_X1 U7055 ( .A(n5467), .ZN(n5468) );
  NAND3_X1 U7056 ( .A1(n7520), .A2(n5473), .A3(n5570), .ZN(n5480) );
  OAI21_X1 U7057 ( .B1(n5474), .B2(n5468), .A(n5480), .ZN(n5470) );
  INV_X1 U7058 ( .A(n7240), .ZN(n9995) );
  NAND3_X1 U7059 ( .A1(n9995), .A2(n8097), .A3(n5570), .ZN(n5469) );
  NAND4_X1 U7060 ( .A1(n5471), .A2(n5472), .A3(n5470), .A4(n5469), .ZN(n5482)
         );
  NAND2_X1 U7061 ( .A1(n5473), .A2(n5472), .ZN(n5475) );
  MUX2_X1 U7062 ( .A(n5475), .B(n5474), .S(n5570), .Z(n5477) );
  INV_X1 U7063 ( .A(n5478), .ZN(n5476) );
  NOR2_X1 U7064 ( .A1(n5477), .A2(n5476), .ZN(n5481) );
  NAND3_X1 U7065 ( .A1(n5577), .A2(n5559), .A3(n5478), .ZN(n5479) );
  AOI22_X1 U7066 ( .A1(n5482), .A2(n5481), .B1(n5480), .B2(n5479), .ZN(n5486)
         );
  INV_X1 U7067 ( .A(n5483), .ZN(n5484) );
  OAI21_X1 U7068 ( .B1(n5486), .B2(n5484), .A(n5575), .ZN(n5488) );
  NAND2_X1 U7069 ( .A1(n5575), .A2(n5577), .ZN(n5485) );
  OAI21_X1 U7070 ( .B1(n5486), .B2(n5485), .A(n5576), .ZN(n5487) );
  MUX2_X1 U7071 ( .A(n5488), .B(n5487), .S(n5570), .Z(n5493) );
  INV_X1 U7072 ( .A(n5490), .ZN(n5491) );
  MUX2_X1 U7073 ( .A(n5213), .B(n5491), .S(n5570), .Z(n5492) );
  MUX2_X1 U7074 ( .A(n5495), .B(n5494), .S(n5570), .Z(n5496) );
  NAND2_X1 U7075 ( .A1(n7737), .A2(n5496), .ZN(n5500) );
  MUX2_X1 U7076 ( .A(n5498), .B(n5497), .S(n5570), .Z(n5499) );
  MUX2_X1 U7077 ( .A(n5502), .B(n5501), .S(n5570), .Z(n5503) );
  INV_X1 U7078 ( .A(n8453), .ZN(n8375) );
  OAI21_X1 U7079 ( .B1(n8375), .B2(n8088), .A(n5506), .ZN(n5504) );
  MUX2_X1 U7080 ( .A(n5504), .B(n8350), .S(n5570), .Z(n5505) );
  INV_X1 U7081 ( .A(n5506), .ZN(n5507) );
  OAI21_X1 U7082 ( .B1(n5517), .B2(n5507), .A(n5514), .ZN(n5508) );
  NAND3_X1 U7083 ( .A1(n5508), .A2(n5519), .A3(n5515), .ZN(n5509) );
  NAND2_X1 U7084 ( .A1(n8318), .A2(n8084), .ZN(n5524) );
  NAND3_X1 U7085 ( .A1(n5509), .A2(n5522), .A3(n5524), .ZN(n5510) );
  NOR2_X1 U7086 ( .A1(n5512), .A2(n5559), .ZN(n5530) );
  NAND2_X1 U7087 ( .A1(n5514), .A2(n5513), .ZN(n5516) );
  OAI21_X1 U7088 ( .B1(n5517), .B2(n5516), .A(n5515), .ZN(n5523) );
  INV_X1 U7089 ( .A(n5518), .ZN(n5521) );
  INV_X1 U7090 ( .A(n5519), .ZN(n5520) );
  AOI211_X1 U7091 ( .C1(n5523), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5527)
         );
  NAND3_X1 U7092 ( .A1(n5525), .A2(n5559), .A3(n5524), .ZN(n5526) );
  OAI21_X1 U7093 ( .B1(n5533), .B2(n8421), .A(n5532), .ZN(n5534) );
  NAND2_X1 U7094 ( .A1(n5534), .A2(n5559), .ZN(n5537) );
  INV_X1 U7095 ( .A(n5535), .ZN(n5536) );
  INV_X1 U7096 ( .A(n5539), .ZN(n5542) );
  NOR2_X1 U7097 ( .A1(n5542), .A2(n5540), .ZN(n5541) );
  AOI21_X1 U7098 ( .B1(n5543), .B2(n5559), .A(n8216), .ZN(n5544) );
  INV_X1 U7099 ( .A(n5545), .ZN(n5549) );
  NAND2_X1 U7100 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  MUX2_X1 U7101 ( .A(n5549), .B(n5548), .S(n5570), .Z(n5552) );
  INV_X1 U7102 ( .A(n5550), .ZN(n5551) );
  AOI211_X1 U7103 ( .C1(n8473), .C2(n5570), .A(n5555), .B(n5556), .ZN(n5564)
         );
  NAND2_X1 U7104 ( .A1(n5560), .A2(n5561), .ZN(n6475) );
  AOI21_X1 U7105 ( .B1(n5559), .B2(n5560), .A(n5558), .ZN(n5563) );
  MUX2_X1 U7106 ( .A(n5561), .B(n5560), .S(n5570), .Z(n5562) );
  XOR2_X1 U7107 ( .A(n6595), .B(n8182), .Z(n5566) );
  OR2_X1 U7108 ( .A1(n8182), .A2(n6595), .ZN(n5565) );
  NAND2_X1 U7109 ( .A1(n5571), .A2(n5565), .ZN(n5574) );
  INV_X1 U7110 ( .A(n5567), .ZN(n5568) );
  INV_X1 U7111 ( .A(n6972), .ZN(n9952) );
  INV_X1 U7112 ( .A(n5628), .ZN(n5573) );
  INV_X1 U7113 ( .A(n5574), .ZN(n5599) );
  INV_X1 U7114 ( .A(n6475), .ZN(n6481) );
  INV_X1 U7115 ( .A(n8204), .ZN(n5597) );
  INV_X1 U7116 ( .A(n8349), .ZN(n5593) );
  NAND2_X1 U7117 ( .A1(n7520), .A2(n5577), .ZN(n6466) );
  NAND2_X1 U7118 ( .A1(n6973), .A2(n5578), .ZN(n9953) );
  NOR2_X1 U7119 ( .A1(n9953), .A2(n5629), .ZN(n5582) );
  INV_X1 U7120 ( .A(n7084), .ZN(n7090) );
  INV_X1 U7121 ( .A(n6446), .ZN(n5581) );
  NAND4_X1 U7122 ( .A1(n5582), .A2(n7090), .A3(n5059), .A4(n5581), .ZN(n5585)
         );
  NAND2_X1 U7123 ( .A1(n5583), .A2(n9887), .ZN(n5584) );
  NOR3_X1 U7124 ( .A1(n5585), .A2(n5584), .A3(n7117), .ZN(n5587) );
  NAND4_X1 U7125 ( .A1(n5587), .A2(n5586), .A3(n7070), .A4(n7178), .ZN(n5588)
         );
  NOR2_X1 U7126 ( .A1(n5588), .A2(n7592), .ZN(n5589) );
  NAND4_X1 U7127 ( .A1(n7570), .A2(n7522), .A3(n4750), .A4(n5589), .ZN(n5590)
         );
  NOR4_X1 U7128 ( .A1(n7832), .A2(n7734), .A3(n5591), .A4(n5590), .ZN(n5592)
         );
  NAND4_X1 U7129 ( .A1(n8337), .A2(n5593), .A3(n5592), .A4(n5270), .ZN(n5594)
         );
  NOR4_X1 U7130 ( .A1(n8291), .A2(n8310), .A3(n8322), .A4(n5594), .ZN(n5595)
         );
  NAND4_X1 U7131 ( .A1(n8247), .A2(n8262), .A3(n5595), .A4(n8281), .ZN(n5596)
         );
  NOR4_X1 U7132 ( .A1(n5597), .A2(n8216), .A3(n8228), .A4(n5596), .ZN(n5598)
         );
  NAND4_X1 U7133 ( .A1(n5600), .A2(n5599), .A3(n6481), .A4(n5598), .ZN(n5601)
         );
  XNOR2_X1 U7134 ( .A(n5601), .B(n7343), .ZN(n5602) );
  OAI22_X1 U7135 ( .A1(n5602), .A2(n5630), .B1(n6478), .B2(n5628), .ZN(n5603)
         );
  NAND2_X1 U7136 ( .A1(n6507), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6696) );
  OAI21_X1 U7137 ( .B1(n5611), .B2(n5610), .A(n7667), .ZN(n5627) );
  NAND2_X1 U7138 ( .A1(n4396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5616) );
  MUX2_X1 U7139 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5616), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5617) );
  NAND2_X1 U7140 ( .A1(n5617), .A2(n5011), .ZN(n5786) );
  NAND2_X1 U7141 ( .A1(n5618), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5619) );
  MUX2_X1 U7142 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5619), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5620) );
  NAND2_X1 U7143 ( .A1(n5620), .A2(n4396), .ZN(n7795) );
  NOR2_X1 U7144 ( .A1(n5786), .A2(n7795), .ZN(n5621) );
  INV_X1 U7145 ( .A(n9944), .ZN(n8035) );
  AND2_X1 U7146 ( .A1(n5629), .A2(n7343), .ZN(n5798) );
  INV_X1 U7147 ( .A(n6703), .ZN(n8511) );
  NAND2_X1 U7148 ( .A1(n5625), .A2(n5630), .ZN(n5799) );
  INV_X1 U7149 ( .A(n5799), .ZN(n6699) );
  INV_X1 U7150 ( .A(n5622), .ZN(n5623) );
  AND2_X2 U7151 ( .A1(n6699), .A2(n5623), .ZN(n9832) );
  NAND4_X1 U7152 ( .A1(n8035), .A2(n5798), .A3(n8511), .A4(n9832), .ZN(n5624)
         );
  OAI211_X1 U7153 ( .C1(n5625), .C2(n6696), .A(n5624), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5626) );
  NAND2_X1 U7154 ( .A1(n5627), .A2(n5626), .ZN(P2_U3244) );
  NAND2_X1 U7155 ( .A1(n8104), .A2(n9951), .ZN(n6445) );
  INV_X1 U7156 ( .A(n6445), .ZN(n6963) );
  NAND2_X1 U7157 ( .A1(n6963), .A2(n5638), .ZN(n6916) );
  NAND2_X1 U7158 ( .A1(n6914), .A2(n5662), .ZN(n5632) );
  AND2_X1 U7159 ( .A1(n6916), .A2(n5632), .ZN(n6909) );
  NAND2_X1 U7160 ( .A1(n9833), .A2(n5638), .ZN(n5634) );
  INV_X1 U7161 ( .A(n5633), .ZN(n5635) );
  NAND2_X1 U7162 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  AND2_X1 U7163 ( .A1(n5637), .A2(n5638), .ZN(n5640) );
  XNOR2_X1 U7164 ( .A(n9930), .B(n4322), .ZN(n5639) );
  NAND2_X1 U7165 ( .A1(n5640), .A2(n5639), .ZN(n5644) );
  INV_X1 U7166 ( .A(n5639), .ZN(n6936) );
  INV_X1 U7167 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7168 ( .A1(n6936), .A2(n5641), .ZN(n5642) );
  NAND2_X1 U7169 ( .A1(n5644), .A2(n5642), .ZN(n9838) );
  NAND2_X1 U7170 ( .A1(n6937), .A2(n5644), .ZN(n5650) );
  AND2_X1 U7171 ( .A1(n9835), .A2(n9898), .ZN(n5646) );
  XNOR2_X1 U7172 ( .A(n4312), .B(n5761), .ZN(n5645) );
  NAND2_X1 U7173 ( .A1(n5646), .A2(n5645), .ZN(n5651) );
  INV_X1 U7174 ( .A(n5645), .ZN(n5648) );
  INV_X1 U7175 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7176 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  AND2_X1 U7177 ( .A1(n5651), .A2(n5649), .ZN(n6938) );
  NAND2_X1 U7178 ( .A1(n5650), .A2(n6938), .ZN(n6940) );
  XNOR2_X1 U7179 ( .A(n9811), .B(n5761), .ZN(n5652) );
  NAND2_X1 U7180 ( .A1(n8102), .A2(n9898), .ZN(n5653) );
  XNOR2_X1 U7181 ( .A(n5652), .B(n5653), .ZN(n9809) );
  INV_X1 U7182 ( .A(n5652), .ZN(n5654) );
  NAND2_X1 U7183 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  AND2_X1 U7184 ( .A1(n8101), .A2(n9898), .ZN(n5657) );
  XNOR2_X1 U7185 ( .A(n4315), .B(n5761), .ZN(n5656) );
  NAND2_X1 U7186 ( .A1(n5657), .A2(n5656), .ZN(n5661) );
  INV_X1 U7187 ( .A(n5656), .ZN(n5659) );
  INV_X1 U7188 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7189 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  AND2_X1 U7190 ( .A1(n5661), .A2(n5660), .ZN(n7017) );
  NAND2_X1 U7191 ( .A1(n7016), .A2(n5661), .ZN(n9853) );
  INV_X1 U7192 ( .A(n9853), .ZN(n5664) );
  XNOR2_X1 U7193 ( .A(n9858), .B(n5769), .ZN(n5666) );
  NAND2_X1 U7194 ( .A1(n8100), .A2(n9898), .ZN(n5665) );
  XNOR2_X1 U7195 ( .A(n5666), .B(n5665), .ZN(n9852) );
  NAND2_X1 U7196 ( .A1(n5664), .A2(n5663), .ZN(n9856) );
  NAND2_X1 U7197 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  XNOR2_X1 U7198 ( .A(n7080), .B(n5761), .ZN(n5668) );
  AND2_X1 U7199 ( .A1(n8099), .A2(n9898), .ZN(n5669) );
  NAND2_X1 U7200 ( .A1(n5668), .A2(n5669), .ZN(n5672) );
  INV_X1 U7201 ( .A(n5668), .ZN(n7232) );
  INV_X1 U7202 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U7203 ( .A1(n7232), .A2(n5670), .ZN(n5671) );
  AND2_X1 U7204 ( .A1(n5672), .A2(n5671), .ZN(n7125) );
  XNOR2_X1 U7205 ( .A(n7240), .B(n5761), .ZN(n5673) );
  AND2_X1 U7206 ( .A1(n8097), .A2(n9898), .ZN(n5674) );
  NAND2_X1 U7207 ( .A1(n5673), .A2(n5674), .ZN(n5678) );
  INV_X1 U7208 ( .A(n5673), .ZN(n7405) );
  INV_X1 U7209 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U7210 ( .A1(n7405), .A2(n5675), .ZN(n5676) );
  AND2_X1 U7211 ( .A1(n5678), .A2(n5676), .ZN(n7228) );
  XNOR2_X1 U7212 ( .A(n7475), .B(n5761), .ZN(n5680) );
  NAND2_X1 U7213 ( .A1(n8096), .A2(n9898), .ZN(n5681) );
  XNOR2_X1 U7214 ( .A(n5680), .B(n5681), .ZN(n7419) );
  AND2_X1 U7215 ( .A1(n7419), .A2(n5678), .ZN(n5679) );
  INV_X1 U7216 ( .A(n5680), .ZN(n5682) );
  NAND2_X1 U7217 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  XNOR2_X1 U7218 ( .A(n9877), .B(n5769), .ZN(n5684) );
  NAND2_X1 U7219 ( .A1(n8095), .A2(n9898), .ZN(n5685) );
  XNOR2_X1 U7220 ( .A(n5684), .B(n5685), .ZN(n7421) );
  INV_X1 U7221 ( .A(n5684), .ZN(n5687) );
  INV_X1 U7222 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7223 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  NAND2_X1 U7224 ( .A1(n7423), .A2(n5688), .ZN(n9821) );
  XNOR2_X1 U7225 ( .A(n9827), .B(n5769), .ZN(n5689) );
  NAND2_X1 U7226 ( .A1(n8094), .A2(n9898), .ZN(n5690) );
  NAND2_X1 U7227 ( .A1(n5689), .A2(n5690), .ZN(n9819) );
  INV_X1 U7228 ( .A(n5689), .ZN(n5692) );
  INV_X1 U7229 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7230 ( .A1(n5692), .A2(n5691), .ZN(n9820) );
  XNOR2_X1 U7231 ( .A(n7663), .B(n5769), .ZN(n5694) );
  NAND2_X1 U7232 ( .A1(n8093), .A2(n9898), .ZN(n5693) );
  XNOR2_X1 U7233 ( .A(n5694), .B(n5693), .ZN(n7657) );
  XNOR2_X1 U7234 ( .A(n7575), .B(n5761), .ZN(n5695) );
  AND2_X1 U7235 ( .A1(n8092), .A2(n9898), .ZN(n5696) );
  NAND2_X1 U7236 ( .A1(n5695), .A2(n5696), .ZN(n5700) );
  INV_X1 U7237 ( .A(n5695), .ZN(n5698) );
  INV_X1 U7238 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7239 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  AND2_X1 U7240 ( .A1(n5700), .A2(n5699), .ZN(n7700) );
  XNOR2_X1 U7241 ( .A(n9638), .B(n5761), .ZN(n5701) );
  NAND2_X1 U7242 ( .A1(n8091), .A2(n9898), .ZN(n5702) );
  XNOR2_X1 U7243 ( .A(n5701), .B(n5702), .ZN(n9636) );
  INV_X1 U7244 ( .A(n5701), .ZN(n5703) );
  NAND2_X1 U7245 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7246 ( .A1(n9635), .A2(n5704), .ZN(n7901) );
  XNOR2_X1 U7247 ( .A(n8459), .B(n5761), .ZN(n8007) );
  AND2_X1 U7248 ( .A1(n8089), .A2(n9898), .ZN(n5707) );
  AND2_X1 U7249 ( .A1(n8090), .A2(n9898), .ZN(n5706) );
  XNOR2_X1 U7250 ( .A(n7744), .B(n5761), .ZN(n7902) );
  AOI22_X1 U7251 ( .A1(n8007), .A2(n5707), .B1(n5706), .B2(n7902), .ZN(n5705)
         );
  NAND2_X1 U7252 ( .A1(n7901), .A2(n5705), .ZN(n5712) );
  INV_X1 U7253 ( .A(n8007), .ZN(n5710) );
  OAI21_X1 U7254 ( .B1(n7902), .B2(n5706), .A(n5707), .ZN(n5709) );
  INV_X1 U7255 ( .A(n7902), .ZN(n8003) );
  INV_X1 U7256 ( .A(n5706), .ZN(n8004) );
  INV_X1 U7257 ( .A(n5707), .ZN(n8006) );
  AND2_X1 U7258 ( .A1(n8004), .A2(n8006), .ZN(n5708) );
  AOI22_X1 U7259 ( .A1(n5710), .A2(n5709), .B1(n8003), .B2(n5708), .ZN(n5711)
         );
  XNOR2_X1 U7260 ( .A(n8453), .B(n5761), .ZN(n5713) );
  AND2_X1 U7261 ( .A1(n8088), .A2(n9898), .ZN(n5714) );
  NAND2_X1 U7262 ( .A1(n5713), .A2(n5714), .ZN(n5718) );
  INV_X1 U7263 ( .A(n5713), .ZN(n8052) );
  INV_X1 U7264 ( .A(n5714), .ZN(n5715) );
  NAND2_X1 U7265 ( .A1(n8052), .A2(n5715), .ZN(n5716) );
  NAND2_X1 U7266 ( .A1(n5718), .A2(n5716), .ZN(n7892) );
  XNOR2_X1 U7267 ( .A(n8357), .B(n5761), .ZN(n5719) );
  AND2_X1 U7268 ( .A1(n8087), .A2(n9898), .ZN(n5720) );
  NAND2_X1 U7269 ( .A1(n5719), .A2(n5720), .ZN(n5724) );
  INV_X1 U7270 ( .A(n5719), .ZN(n7971) );
  INV_X1 U7271 ( .A(n5720), .ZN(n5721) );
  NAND2_X1 U7272 ( .A1(n7971), .A2(n5721), .ZN(n5722) );
  AND2_X1 U7273 ( .A1(n5724), .A2(n5722), .ZN(n8050) );
  NAND2_X1 U7274 ( .A1(n5723), .A2(n8050), .ZN(n7969) );
  XNOR2_X1 U7275 ( .A(n8443), .B(n5761), .ZN(n5726) );
  NAND2_X1 U7276 ( .A1(n8086), .A2(n9898), .ZN(n5727) );
  XNOR2_X1 U7277 ( .A(n5726), .B(n5727), .ZN(n7980) );
  AND2_X1 U7278 ( .A1(n7980), .A2(n5724), .ZN(n5725) );
  NAND2_X1 U7279 ( .A1(n7969), .A2(n5725), .ZN(n7976) );
  INV_X1 U7280 ( .A(n5726), .ZN(n5728) );
  NAND2_X1 U7281 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  XNOR2_X1 U7282 ( .A(n8329), .B(n5761), .ZN(n5730) );
  AND2_X1 U7283 ( .A1(n8085), .A2(n9898), .ZN(n5731) );
  NAND2_X1 U7284 ( .A1(n5730), .A2(n5731), .ZN(n5735) );
  INV_X1 U7285 ( .A(n5730), .ZN(n7986) );
  INV_X1 U7286 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7287 ( .A1(n7986), .A2(n5732), .ZN(n5733) );
  NAND2_X1 U7288 ( .A1(n5735), .A2(n5733), .ZN(n8028) );
  XNOR2_X1 U7289 ( .A(n8433), .B(n5761), .ZN(n5739) );
  NAND2_X1 U7290 ( .A1(n8084), .A2(n9898), .ZN(n5737) );
  XNOR2_X1 U7291 ( .A(n5739), .B(n5737), .ZN(n7983) );
  INV_X1 U7292 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7293 ( .A1(n5739), .A2(n5738), .ZN(n5740) );
  XNOR2_X1 U7294 ( .A(n8299), .B(n5769), .ZN(n5742) );
  NAND2_X1 U7295 ( .A1(n8083), .A2(n9898), .ZN(n8038) );
  NAND2_X1 U7296 ( .A1(n8039), .A2(n8038), .ZN(n5745) );
  INV_X1 U7297 ( .A(n5741), .ZN(n5743) );
  NAND2_X1 U7298 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  XNOR2_X1 U7299 ( .A(n8421), .B(n5761), .ZN(n5747) );
  XNOR2_X1 U7300 ( .A(n8271), .B(n5769), .ZN(n8018) );
  NAND2_X1 U7301 ( .A1(n8082), .A2(n9898), .ZN(n7961) );
  AOI21_X1 U7302 ( .B1(n8018), .B2(n8020), .A(n7961), .ZN(n5746) );
  NAND2_X1 U7303 ( .A1(n8081), .A2(n9898), .ZN(n8022) );
  NAND2_X1 U7304 ( .A1(n8018), .A2(n8022), .ZN(n5748) );
  XNOR2_X1 U7305 ( .A(n8253), .B(n5761), .ZN(n5750) );
  AND2_X1 U7306 ( .A1(n8080), .A2(n9898), .ZN(n5751) );
  NAND2_X1 U7307 ( .A1(n5750), .A2(n5751), .ZN(n5754) );
  INV_X1 U7308 ( .A(n5750), .ZN(n8066) );
  INV_X1 U7309 ( .A(n5751), .ZN(n5752) );
  NAND2_X1 U7310 ( .A1(n8066), .A2(n5752), .ZN(n5753) );
  AND2_X1 U7311 ( .A1(n5754), .A2(n5753), .ZN(n7996) );
  NAND2_X1 U7312 ( .A1(n7995), .A2(n5754), .ZN(n5759) );
  XNOR2_X1 U7313 ( .A(n8406), .B(n5761), .ZN(n5755) );
  AND2_X1 U7314 ( .A1(n8079), .A2(n9898), .ZN(n5756) );
  NAND2_X1 U7315 ( .A1(n5755), .A2(n5756), .ZN(n5760) );
  INV_X1 U7316 ( .A(n5755), .ZN(n7954) );
  INV_X1 U7317 ( .A(n5756), .ZN(n5757) );
  NAND2_X1 U7318 ( .A1(n7954), .A2(n5757), .ZN(n5758) );
  AND2_X1 U7319 ( .A1(n5760), .A2(n5758), .ZN(n8062) );
  NAND2_X1 U7320 ( .A1(n7950), .A2(n5760), .ZN(n5767) );
  XNOR2_X1 U7321 ( .A(n8401), .B(n5761), .ZN(n5762) );
  AND2_X1 U7322 ( .A1(n8078), .A2(n9898), .ZN(n5763) );
  NAND2_X1 U7323 ( .A1(n5762), .A2(n5763), .ZN(n5768) );
  INV_X1 U7324 ( .A(n5762), .ZN(n5765) );
  INV_X1 U7325 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7326 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  AND2_X1 U7327 ( .A1(n5768), .A2(n5766), .ZN(n7951) );
  NAND2_X1 U7328 ( .A1(n5767), .A2(n7951), .ZN(n7955) );
  NAND2_X1 U7329 ( .A1(n7955), .A2(n5768), .ZN(n5772) );
  NAND2_X1 U7330 ( .A1(n8077), .A2(n9898), .ZN(n5770) );
  XNOR2_X1 U7331 ( .A(n5770), .B(n5769), .ZN(n5771) );
  XNOR2_X1 U7332 ( .A(n5772), .B(n5771), .ZN(n5792) );
  INV_X1 U7333 ( .A(n5792), .ZN(n5791) );
  NOR4_X1 U7334 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5776) );
  NOR4_X1 U7335 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5775) );
  NOR4_X1 U7336 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5774) );
  NOR4_X1 U7337 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5773) );
  NAND4_X1 U7338 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5784)
         );
  NOR2_X1 U7339 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n5780) );
  NOR4_X1 U7340 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5779) );
  NOR4_X1 U7341 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5778) );
  NOR4_X1 U7342 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5777) );
  NAND4_X1 U7343 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5783)
         );
  XOR2_X1 U7344 ( .A(n7710), .B(P2_B_REG_SCAN_IN), .Z(n5781) );
  NAND2_X1 U7345 ( .A1(n7795), .A2(n5781), .ZN(n5782) );
  NOR2_X1 U7346 ( .A1(n7710), .A2(n7858), .ZN(n9946) );
  INV_X1 U7347 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9945) );
  AND2_X1 U7348 ( .A1(n9943), .A2(n9945), .ZN(n5785) );
  INV_X1 U7349 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U7350 ( .A1(n9943), .A2(n9948), .ZN(n5788) );
  AND2_X1 U7351 ( .A1(n5786), .A2(n7795), .ZN(n9950) );
  INV_X1 U7352 ( .A(n9950), .ZN(n5787) );
  NAND2_X1 U7353 ( .A1(n5788), .A2(n5787), .ZN(n6964) );
  NOR2_X1 U7354 ( .A1(n6966), .A2(n6964), .ZN(n5789) );
  NAND2_X1 U7355 ( .A1(n6489), .A2(n5789), .ZN(n5793) );
  AND2_X1 U7356 ( .A1(n10002), .A2(n5799), .ZN(n5790) );
  NAND2_X1 U7357 ( .A1(n5791), .A2(n9841), .ZN(n5806) );
  NAND2_X1 U7358 ( .A1(n5793), .A2(n6969), .ZN(n8036) );
  NOR2_X1 U7359 ( .A1(n9944), .A2(n10002), .ZN(n5794) );
  AND2_X2 U7360 ( .A1(n6699), .A2(n5622), .ZN(n9834) );
  AOI22_X1 U7361 ( .A1(n8078), .A2(n9832), .B1(n8076), .B2(n9834), .ZN(n8202)
         );
  INV_X1 U7362 ( .A(n5797), .ZN(n8208) );
  NOR2_X1 U7363 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  NAND2_X1 U7364 ( .A1(n8036), .A2(n6488), .ZN(n5802) );
  AOI22_X1 U7365 ( .A1(n8208), .A2(n8046), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5803) );
  NOR2_X1 U7366 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5809) );
  NOR2_X1 U7367 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5808) );
  NAND4_X1 U7368 ( .A1(n5809), .A2(n5808), .A3(n5834), .A4(n6129), .ZN(n5813)
         );
  NAND4_X1 U7369 ( .A1(n5811), .A2(n5810), .A3(n6174), .A4(n5866), .ZN(n5812)
         );
  INV_X1 U7370 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5816) );
  INV_X1 U7371 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5817) );
  INV_X1 U7372 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5818) );
  INV_X1 U7373 ( .A(n5828), .ZN(n5826) );
  NAND2_X1 U7374 ( .A1(n5858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7375 ( .A1(n6232), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7376 ( .A1(n5827), .A2(n5828), .ZN(n5899) );
  NAND2_X1 U7377 ( .A1(n4344), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5829) );
  INV_X1 U7378 ( .A(n6151), .ZN(n5835) );
  NOR2_X1 U7379 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n5835), .ZN(n5836) );
  INV_X1 U7380 ( .A(n6173), .ZN(n5838) );
  NOR2_X1 U7381 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5837) );
  NAND2_X1 U7382 ( .A1(n5838), .A2(n5837), .ZN(n5871) );
  NAND2_X1 U7383 ( .A1(n5840), .A2(n5839), .ZN(n5873) );
  NAND2_X2 U7384 ( .A1(n6385), .A2(n8947), .ZN(n5875) );
  NAND2_X1 U7385 ( .A1(n5846), .A2(n5845), .ZN(n5848) );
  OR2_X1 U7386 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U7387 ( .A1(n4351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5850) );
  NAND2_X2 U7388 ( .A1(n6393), .A2(n5851), .ZN(n6504) );
  OR2_X4 U7389 ( .A1(n5875), .A2(n5877), .ZN(n6379) );
  NAND2_X1 U7390 ( .A1(n6744), .A2(n5893), .ZN(n5865) );
  NAND2_X1 U7391 ( .A1(n4401), .A2(SI_0_), .ZN(n5853) );
  INV_X1 U7392 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7393 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  OR2_X1 U7394 ( .A1(n5861), .A2(n5860), .ZN(n5855) );
  NAND2_X1 U7395 ( .A1(n5855), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5857) );
  INV_X1 U7396 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5860) );
  INV_X1 U7397 ( .A(n5861), .ZN(n5862) );
  NAND2_X4 U7398 ( .A1(n5875), .A2(n6504), .ZN(n6380) );
  AOI22_X1 U7399 ( .A1(n7270), .A2(n5880), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n5877), .ZN(n5864) );
  NAND2_X1 U7400 ( .A1(n5865), .A2(n5864), .ZN(n6736) );
  INV_X1 U7401 ( .A(n6736), .ZN(n5876) );
  NAND2_X1 U7402 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  NAND2_X1 U7403 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5870) );
  XNOR2_X1 U7404 ( .A(n5870), .B(n5869), .ZN(n5878) );
  NAND2_X1 U7405 ( .A1(n5871), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  MUX2_X1 U7406 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5872), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5874) );
  NAND2_X1 U7407 ( .A1(n5876), .A2(n7222), .ZN(n5883) );
  NAND2_X1 U7408 ( .A1(n5878), .A2(n6418), .ZN(n5879) );
  AND2_X2 U7409 ( .A1(n5880), .A2(n5879), .ZN(n5909) );
  AND2_X1 U7410 ( .A1(n5882), .A2(n5881), .ZN(n6738) );
  NAND2_X1 U7411 ( .A1(n6738), .A2(n6736), .ZN(n6737) );
  AND2_X1 U7412 ( .A1(n5883), .A2(n6737), .ZN(n5894) );
  NAND2_X1 U7413 ( .A1(n6232), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7414 ( .A1(n4325), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7415 ( .A1(n4344), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7416 ( .A1(n7041), .A2(n4316), .ZN(n5891) );
  INV_X1 U7417 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7418 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5888) );
  NAND2_X1 U7419 ( .A1(n5921), .A2(n6553), .ZN(n5889) );
  NAND2_X1 U7420 ( .A1(n7101), .A2(n6346), .ZN(n5890) );
  NAND2_X1 U7421 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  XNOR2_X1 U7422 ( .A(n5892), .B(n7222), .ZN(n5895) );
  NAND2_X1 U7423 ( .A1(n5894), .A2(n5895), .ZN(n6751) );
  AOI22_X1 U7424 ( .A1(n7041), .A2(n5909), .B1(n7101), .B2(n5893), .ZN(n6752)
         );
  NAND2_X1 U7425 ( .A1(n6751), .A2(n6752), .ZN(n5898) );
  INV_X1 U7426 ( .A(n5894), .ZN(n5897) );
  INV_X1 U7427 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U7428 ( .A1(n5897), .A2(n5896), .ZN(n6750) );
  NAND2_X1 U7429 ( .A1(n5898), .A2(n6750), .ZN(n7934) );
  NAND2_X1 U7430 ( .A1(n5914), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7431 ( .A1(n4344), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7432 ( .A1(n6232), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5900) );
  INV_X1 U7433 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7434 ( .A1(n4311), .A2(n6546), .ZN(n5906) );
  INV_X1 U7435 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6541) );
  OR2_X1 U7436 ( .A1(n5927), .A2(n6541), .ZN(n5905) );
  OAI211_X1 U7437 ( .C1(n6506), .C2(n6777), .A(n5906), .B(n5905), .ZN(n5907)
         );
  INV_X2 U7438 ( .A(n5907), .ZN(n7943) );
  OAI22_X1 U7439 ( .A1(n7303), .A2(n6379), .B1(n7943), .B2(n6380), .ZN(n5908)
         );
  XNOR2_X1 U7440 ( .A(n5908), .B(n7222), .ZN(n5911) );
  OAI22_X1 U7441 ( .A1(n7303), .A2(n6378), .B1(n7943), .B2(n6379), .ZN(n5910)
         );
  NAND2_X1 U7442 ( .A1(n5911), .A2(n5910), .ZN(n5912) );
  AND2_X2 U7443 ( .A1(n5913), .A2(n5912), .ZN(n7935) );
  NAND2_X1 U7444 ( .A1(n7934), .A2(n7935), .ZN(n7933) );
  NAND2_X1 U7445 ( .A1(n7933), .A2(n5913), .ZN(n6950) );
  INV_X1 U7446 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7447 ( .A1(n6298), .A2(n5915), .ZN(n5920) );
  NAND2_X1 U7448 ( .A1(n5916), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7449 ( .A1(n6232), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7450 ( .A1(n4344), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5917) );
  AND4_X2 U7451 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n7938)
         );
  NAND2_X1 U7452 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U7453 ( .A1(n5924), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  INV_X1 U7454 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7455 ( .A(n5926), .B(n5925), .ZN(n6676) );
  INV_X1 U7456 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6543) );
  OR2_X1 U7457 ( .A1(n5927), .A2(n6543), .ZN(n5929) );
  OR2_X1 U7458 ( .A1(n5943), .A2(n6542), .ZN(n5928) );
  OAI22_X1 U7459 ( .A1(n7938), .A2(n6379), .B1(n9761), .B2(n6380), .ZN(n5930)
         );
  XNOR2_X1 U7460 ( .A(n5930), .B(n6255), .ZN(n5931) );
  OAI22_X1 U7461 ( .A1(n7938), .A2(n6378), .B1(n9761), .B2(n6379), .ZN(n5932)
         );
  XNOR2_X1 U7462 ( .A(n5931), .B(n5932), .ZN(n6947) );
  INV_X1 U7463 ( .A(n5931), .ZN(n5933) );
  OR2_X1 U7464 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U7465 ( .A1(n5916), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5939) );
  INV_X1 U7466 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7467 ( .A(n5935), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U7468 ( .A1(n6298), .A2(n7291), .ZN(n5938) );
  NAND2_X1 U7469 ( .A1(n6232), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7470 ( .A1(n4344), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7471 ( .A1(n5940), .A2(n5860), .ZN(n5942) );
  XNOR2_X1 U7472 ( .A(n5942), .B(n5941), .ZN(n6804) );
  INV_X1 U7473 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6552) );
  OR2_X1 U7474 ( .A1(n5927), .A2(n6552), .ZN(n5945) );
  OR2_X1 U7475 ( .A1(n5943), .A2(n6551), .ZN(n5944) );
  OAI211_X1 U7476 ( .C1(n8655), .C2(n6804), .A(n5945), .B(n5944), .ZN(n7292)
         );
  OAI22_X1 U7477 ( .A1(n7302), .A2(n6379), .B1(n7217), .B2(n6380), .ZN(n5946)
         );
  XNOR2_X1 U7478 ( .A(n5946), .B(n6255), .ZN(n5950) );
  OR2_X1 U7479 ( .A1(n7302), .A2(n6378), .ZN(n5948) );
  NAND2_X1 U7480 ( .A1(n7292), .A2(n6356), .ZN(n5947) );
  NAND2_X1 U7481 ( .A1(n5948), .A2(n5947), .ZN(n5951) );
  INV_X1 U7482 ( .A(n5951), .ZN(n5949) );
  AND2_X1 U7483 ( .A1(n5950), .A2(n5949), .ZN(n7005) );
  INV_X1 U7484 ( .A(n5950), .ZN(n5952) );
  NAND2_X1 U7485 ( .A1(n5952), .A2(n5951), .ZN(n7006) );
  NAND2_X1 U7486 ( .A1(n5916), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7487 ( .A1(n5965), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U7488 ( .B1(n5965), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5985), .ZN(
        n7285) );
  INV_X1 U7489 ( .A(n7285), .ZN(n7374) );
  NAND2_X1 U7490 ( .A1(n6298), .A2(n7374), .ZN(n5957) );
  INV_X2 U7491 ( .A(n5954), .ZN(n8649) );
  NAND2_X1 U7492 ( .A1(n8649), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7493 ( .A1(n8650), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7494 ( .A1(n5959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5961) );
  INV_X1 U7495 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5960) );
  XNOR2_X1 U7496 ( .A(n5961), .B(n5960), .ZN(n6658) );
  OR2_X1 U7497 ( .A1(n5927), .A2(n6556), .ZN(n5963) );
  OAI211_X1 U7498 ( .C1(n8655), .C2(n6658), .A(n5963), .B(n5962), .ZN(n7287)
         );
  XNOR2_X1 U7499 ( .A(n5964), .B(n7222), .ZN(n5982) );
  OAI22_X1 U7500 ( .A1(n7392), .A2(n6378), .B1(n9773), .B2(n6379), .ZN(n5981)
         );
  OR2_X1 U7501 ( .A1(n5982), .A2(n5981), .ZN(n7366) );
  NAND2_X1 U7502 ( .A1(n5916), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5970) );
  AOI21_X1 U7503 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5966) );
  NOR2_X1 U7504 ( .A1(n5966), .A2(n5965), .ZN(n7210) );
  NAND2_X1 U7505 ( .A1(n6298), .A2(n7210), .ZN(n5969) );
  NAND2_X1 U7506 ( .A1(n8649), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7507 ( .A1(n8650), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5967) );
  NOR2_X1 U7508 ( .A1(n5971), .A2(n5860), .ZN(n5972) );
  MUX2_X1 U7509 ( .A(n5860), .B(n5972), .S(P1_IR_REG_5__SCAN_IN), .Z(n5973) );
  INV_X1 U7510 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U7511 ( .A1(n5974), .A2(n5959), .ZN(n6637) );
  INV_X1 U7512 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6550) );
  OR2_X1 U7513 ( .A1(n5927), .A2(n6550), .ZN(n5976) );
  OR2_X1 U7514 ( .A1(n5943), .A2(n6549), .ZN(n5975) );
  OAI211_X1 U7515 ( .C1(n8655), .C2(n6637), .A(n5976), .B(n5975), .ZN(n7338)
         );
  INV_X1 U7516 ( .A(n7338), .ZN(n9768) );
  OAI22_X1 U7517 ( .A1(n7369), .A2(n6379), .B1(n9768), .B2(n6380), .ZN(n5977)
         );
  XNOR2_X1 U7518 ( .A(n5977), .B(n7222), .ZN(n7364) );
  OR2_X1 U7519 ( .A1(n7369), .A2(n6378), .ZN(n5979) );
  NAND2_X1 U7520 ( .A1(n7338), .A2(n6356), .ZN(n5978) );
  NAND2_X1 U7521 ( .A1(n5979), .A2(n5978), .ZN(n7330) );
  OR2_X1 U7522 ( .A1(n7364), .A2(n7330), .ZN(n5980) );
  NAND2_X1 U7523 ( .A1(n7363), .A2(n4852), .ZN(n7159) );
  NAND3_X1 U7524 ( .A1(n7366), .A2(n7364), .A3(n7330), .ZN(n5983) );
  NAND2_X1 U7525 ( .A1(n5982), .A2(n5981), .ZN(n7365) );
  AND2_X1 U7526 ( .A1(n5983), .A2(n7365), .ZN(n7158) );
  NAND2_X1 U7527 ( .A1(n5916), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5990) );
  AND2_X1 U7528 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NOR2_X1 U7529 ( .A1(n6002), .A2(n5986), .ZN(n7398) );
  NAND2_X1 U7530 ( .A1(n6298), .A2(n7398), .ZN(n5989) );
  NAND2_X1 U7531 ( .A1(n8649), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7532 ( .A1(n8650), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5987) );
  OR2_X1 U7533 ( .A1(n5959), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7534 ( .A1(n6008), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7535 ( .A(n5992), .B(n5991), .ZN(n6619) );
  INV_X1 U7536 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6562) );
  OR2_X1 U7537 ( .A1(n5927), .A2(n6562), .ZN(n5994) );
  OR2_X1 U7538 ( .A1(n5943), .A2(n6561), .ZN(n5993) );
  OAI22_X1 U7539 ( .A1(n7504), .A2(n6379), .B1(n9780), .B2(n6380), .ZN(n5995)
         );
  XNOR2_X1 U7540 ( .A(n5995), .B(n6255), .ZN(n7161) );
  INV_X1 U7541 ( .A(n7161), .ZN(n5998) );
  OR2_X1 U7542 ( .A1(n7504), .A2(n6378), .ZN(n5997) );
  NAND2_X1 U7543 ( .A1(n7385), .A2(n6356), .ZN(n5996) );
  NAND2_X1 U7544 ( .A1(n5997), .A2(n5996), .ZN(n7160) );
  NAND2_X1 U7545 ( .A1(n5998), .A2(n7160), .ZN(n5999) );
  INV_X1 U7546 ( .A(n7160), .ZN(n6000) );
  AOI21_X2 U7547 ( .B1(n7159), .B2(n6001), .A(n4846), .ZN(n7250) );
  NAND2_X1 U7548 ( .A1(n5916), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7549 ( .A1(n6002), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7550 ( .A1(n6002), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6003) );
  AND2_X1 U7551 ( .A1(n6022), .A2(n6003), .ZN(n7581) );
  NAND2_X1 U7552 ( .A1(n6298), .A2(n7581), .ZN(n6006) );
  NAND2_X1 U7553 ( .A1(n8649), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7554 ( .A1(n8650), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7555 ( .A1(n7510), .A2(n6378), .ZN(n6012) );
  NOR2_X1 U7556 ( .A1(n6008), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6015) );
  OR2_X1 U7557 ( .A1(n6015), .A2(n5860), .ZN(n6009) );
  XNOR2_X1 U7558 ( .A(n6009), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7559 ( .A1(n8639), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5921), .B2(
        n6612), .ZN(n6010) );
  NAND2_X1 U7560 ( .A1(n7559), .A2(n6356), .ZN(n6011) );
  NAND2_X1 U7561 ( .A1(n6012), .A2(n6011), .ZN(n7248) );
  OAI22_X1 U7562 ( .A1(n7510), .A2(n6379), .B1(n7583), .B2(n6380), .ZN(n6013)
         );
  XNOR2_X1 U7563 ( .A(n6013), .B(n7222), .ZN(n7247) );
  NAND2_X1 U7564 ( .A1(n6578), .A2(n8645), .ZN(n6020) );
  NAND2_X1 U7565 ( .A1(n6015), .A2(n6014), .ZN(n6017) );
  NAND2_X1 U7566 ( .A1(n6017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  MUX2_X1 U7567 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6016), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6018) );
  AOI22_X1 U7568 ( .A1(n8639), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5921), .B2(
        n6688), .ZN(n6019) );
  NAND2_X1 U7569 ( .A1(n6020), .A2(n6019), .ZN(n7535) );
  NAND2_X1 U7570 ( .A1(n7535), .A2(n6346), .ZN(n6029) );
  NAND2_X1 U7571 ( .A1(n5916), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7572 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  AND2_X1 U7573 ( .A1(n6041), .A2(n6023), .ZN(n7513) );
  NAND2_X1 U7574 ( .A1(n6298), .A2(n7513), .ZN(n6026) );
  NAND2_X1 U7575 ( .A1(n8649), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7576 ( .A1(n8650), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6024) );
  NAND4_X1 U7577 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n8970)
         );
  NAND2_X1 U7578 ( .A1(n8970), .A2(n6356), .ZN(n6028) );
  NAND2_X1 U7579 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  XNOR2_X1 U7580 ( .A(n6030), .B(n6255), .ZN(n6031) );
  AOI22_X1 U7581 ( .A1(n7535), .A2(n6356), .B1(n8970), .B2(n5909), .ZN(n6032)
         );
  NAND2_X1 U7582 ( .A1(n6031), .A2(n6032), .ZN(n6036) );
  INV_X1 U7583 ( .A(n6031), .ZN(n6034) );
  INV_X1 U7584 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U7585 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  NAND2_X1 U7586 ( .A1(n6036), .A2(n6035), .ZN(n7467) );
  NAND2_X1 U7587 ( .A1(n7465), .A2(n6036), .ZN(n7487) );
  NAND2_X1 U7588 ( .A1(n6598), .A2(n8645), .ZN(n6039) );
  NAND2_X1 U7589 ( .A1(n6056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6037) );
  XNOR2_X1 U7590 ( .A(n6037), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7591 ( .A1(n8639), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5921), .B2(
        n6724), .ZN(n6038) );
  NAND2_X1 U7592 ( .A1(n6039), .A2(n6038), .ZN(n7613) );
  NAND2_X1 U7593 ( .A1(n7613), .A2(n6346), .ZN(n6048) );
  NAND2_X1 U7594 ( .A1(n5916), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7595 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  AND2_X1 U7596 ( .A1(n6061), .A2(n6042), .ZN(n7488) );
  NAND2_X1 U7597 ( .A1(n6298), .A2(n7488), .ZN(n6045) );
  NAND2_X1 U7598 ( .A1(n8649), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7599 ( .A1(n8650), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7600 ( .A1(n7618), .A2(n6379), .ZN(n6047) );
  NAND2_X1 U7601 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  XNOR2_X1 U7602 ( .A(n6049), .B(n7222), .ZN(n6052) );
  NAND2_X1 U7603 ( .A1(n7613), .A2(n6356), .ZN(n6051) );
  OR2_X1 U7604 ( .A1(n7618), .A2(n6378), .ZN(n6050) );
  NAND2_X1 U7605 ( .A1(n6051), .A2(n6050), .ZN(n6053) );
  NAND2_X1 U7606 ( .A1(n6052), .A2(n6053), .ZN(n7485) );
  INV_X1 U7607 ( .A(n6052), .ZN(n6055) );
  INV_X1 U7608 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7609 ( .A1(n6055), .A2(n6054), .ZN(n7484) );
  NAND2_X1 U7610 ( .A1(n6596), .A2(n8645), .ZN(n6059) );
  OAI21_X1 U7611 ( .B1(n6056), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6057) );
  XNOR2_X1 U7612 ( .A(n6057), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U7613 ( .A1(n8639), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5921), .B2(
        n6996), .ZN(n6058) );
  NAND2_X1 U7614 ( .A1(n6059), .A2(n6058), .ZN(n7697) );
  NAND2_X1 U7615 ( .A1(n7697), .A2(n6346), .ZN(n6068) );
  NAND2_X1 U7616 ( .A1(n5916), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6066) );
  AND2_X1 U7617 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  NOR2_X1 U7618 ( .A1(n6079), .A2(n6062), .ZN(n7623) );
  NAND2_X1 U7619 ( .A1(n6298), .A2(n7623), .ZN(n6065) );
  NAND2_X1 U7620 ( .A1(n8650), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7621 ( .A1(n8649), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7622 ( .A1(n9612), .A2(n6379), .ZN(n6067) );
  NAND2_X1 U7623 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  XNOR2_X1 U7624 ( .A(n6069), .B(n6255), .ZN(n6073) );
  NOR2_X1 U7625 ( .A1(n9612), .A2(n6378), .ZN(n6070) );
  AOI21_X1 U7626 ( .B1(n7697), .B2(n6356), .A(n6070), .ZN(n6072) );
  XNOR2_X1 U7627 ( .A(n6073), .B(n6072), .ZN(n7694) );
  OR2_X1 U7628 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U7629 ( .A1(n7691), .A2(n6074), .ZN(n9616) );
  NAND2_X1 U7630 ( .A1(n6667), .A2(n8645), .ZN(n6078) );
  NAND2_X1 U7631 ( .A1(n6075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6076) );
  XNOR2_X1 U7632 ( .A(n6076), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8992) );
  AOI22_X1 U7633 ( .A1(n8639), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5921), .B2(
        n8992), .ZN(n6077) );
  NAND2_X1 U7634 ( .A1(n6078), .A2(n6077), .ZN(n7637) );
  NAND2_X1 U7635 ( .A1(n7637), .A2(n6346), .ZN(n6088) );
  NAND2_X1 U7636 ( .A1(n6079), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6099) );
  INV_X1 U7637 ( .A(n6079), .ZN(n6081) );
  INV_X1 U7638 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7639 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  NAND2_X1 U7640 ( .A1(n6099), .A2(n6082), .ZN(n9624) );
  INV_X1 U7641 ( .A(n9624), .ZN(n7638) );
  NAND2_X1 U7642 ( .A1(n6298), .A2(n7638), .ZN(n6086) );
  NAND2_X1 U7643 ( .A1(n5916), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7644 ( .A1(n8650), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7645 ( .A1(n8649), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7646 ( .A1(n7782), .A2(n6379), .ZN(n6087) );
  NAND2_X1 U7647 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  XNOR2_X1 U7648 ( .A(n6089), .B(n6255), .ZN(n6093) );
  NOR2_X1 U7649 ( .A1(n7782), .A2(n6378), .ZN(n6090) );
  AOI21_X1 U7650 ( .B1(n7637), .B2(n6356), .A(n6090), .ZN(n6092) );
  XNOR2_X1 U7651 ( .A(n6093), .B(n6092), .ZN(n9617) );
  NAND2_X1 U7652 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  NAND2_X1 U7653 ( .A1(n6732), .A2(n8645), .ZN(n6097) );
  OR2_X1 U7654 ( .A1(n5833), .A2(n5860), .ZN(n6095) );
  XNOR2_X1 U7655 ( .A(n6095), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U7656 ( .A1(n8639), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5921), .B2(
        n9674), .ZN(n6096) );
  NAND2_X1 U7657 ( .A1(n8707), .A2(n6346), .ZN(n6106) );
  NAND2_X1 U7658 ( .A1(n5916), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7659 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  AND2_X1 U7660 ( .A1(n6114), .A2(n6100), .ZN(n7716) );
  NAND2_X1 U7661 ( .A1(n6298), .A2(n7716), .ZN(n6103) );
  NAND2_X1 U7662 ( .A1(n8650), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7663 ( .A1(n6232), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6101) );
  NAND4_X1 U7664 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n9607)
         );
  NAND2_X1 U7665 ( .A1(n9607), .A2(n6356), .ZN(n6105) );
  NAND2_X1 U7666 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  XNOR2_X1 U7667 ( .A(n6107), .B(n6255), .ZN(n7713) );
  AND2_X1 U7668 ( .A1(n9607), .A2(n5909), .ZN(n6108) );
  AOI21_X1 U7669 ( .B1(n8707), .B2(n6356), .A(n6108), .ZN(n7712) );
  AND2_X1 U7670 ( .A1(n7713), .A2(n7712), .ZN(n6109) );
  NAND2_X1 U7671 ( .A1(n6759), .A2(n8645), .ZN(n6112) );
  OR2_X1 U7672 ( .A1(n6110), .A2(n5860), .ZN(n6130) );
  XNOR2_X1 U7673 ( .A(n6130), .B(n6129), .ZN(n9002) );
  INV_X1 U7674 ( .A(n9002), .ZN(n9689) );
  AOI22_X1 U7675 ( .A1(n8639), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5921), .B2(
        n9689), .ZN(n6111) );
  NAND2_X1 U7676 ( .A1(n9346), .A2(n6346), .ZN(n6121) );
  NAND2_X1 U7677 ( .A1(n5916), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6119) );
  INV_X1 U7678 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U7679 ( .A1(n6114), .A2(n7770), .ZN(n6115) );
  AND2_X1 U7680 ( .A1(n6136), .A2(n6115), .ZN(n7769) );
  NAND2_X1 U7681 ( .A1(n6298), .A2(n7769), .ZN(n6118) );
  NAND2_X1 U7682 ( .A1(n6232), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7683 ( .A1(n8650), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6116) );
  NAND4_X1 U7684 ( .A1(n6119), .A2(n6118), .A3(n6117), .A4(n6116), .ZN(n8966)
         );
  NAND2_X1 U7685 ( .A1(n8966), .A2(n6356), .ZN(n6120) );
  NAND2_X1 U7686 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  XNOR2_X1 U7687 ( .A(n6122), .B(n6255), .ZN(n7767) );
  AND2_X1 U7688 ( .A1(n8966), .A2(n5909), .ZN(n6123) );
  AOI21_X1 U7689 ( .B1(n9346), .B2(n6356), .A(n6123), .ZN(n6125) );
  NAND2_X1 U7690 ( .A1(n7767), .A2(n6125), .ZN(n6124) );
  NAND2_X1 U7691 ( .A1(n7765), .A2(n6124), .ZN(n6128) );
  INV_X1 U7692 ( .A(n7767), .ZN(n6126) );
  INV_X1 U7693 ( .A(n6125), .ZN(n7766) );
  NAND2_X1 U7694 ( .A1(n6126), .A2(n7766), .ZN(n6127) );
  NAND2_X1 U7695 ( .A1(n6128), .A2(n6127), .ZN(n7848) );
  NAND2_X1 U7696 ( .A1(n6959), .A2(n8645), .ZN(n6134) );
  NAND2_X1 U7697 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  NAND2_X1 U7698 ( .A1(n6131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6132) );
  XNOR2_X1 U7699 ( .A(n6132), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9708) );
  AOI22_X1 U7700 ( .A1(n8639), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5921), .B2(
        n9708), .ZN(n6133) );
  NAND2_X1 U7701 ( .A1(n9339), .A2(n6346), .ZN(n6143) );
  NAND2_X1 U7702 ( .A1(n5916), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7703 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  AND2_X1 U7704 ( .A1(n6158), .A2(n6137), .ZN(n7869) );
  NAND2_X1 U7705 ( .A1(n6298), .A2(n7869), .ZN(n6140) );
  NAND2_X1 U7706 ( .A1(n8649), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7707 ( .A1(n8650), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6138) );
  NAND4_X1 U7708 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n8965)
         );
  NAND2_X1 U7709 ( .A1(n8965), .A2(n6356), .ZN(n6142) );
  NAND2_X1 U7710 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  XNOR2_X1 U7711 ( .A(n6144), .B(n6255), .ZN(n7850) );
  AND2_X1 U7712 ( .A1(n8965), .A2(n5909), .ZN(n6145) );
  AOI21_X1 U7713 ( .B1(n9339), .B2(n6356), .A(n6145), .ZN(n6147) );
  NAND2_X1 U7714 ( .A1(n7850), .A2(n6147), .ZN(n6146) );
  NAND2_X1 U7715 ( .A1(n7848), .A2(n6146), .ZN(n6150) );
  INV_X1 U7716 ( .A(n7850), .ZN(n6148) );
  INV_X1 U7717 ( .A(n6147), .ZN(n7849) );
  NAND2_X1 U7718 ( .A1(n6148), .A2(n7849), .ZN(n6149) );
  NAND2_X1 U7719 ( .A1(n7059), .A2(n8645), .ZN(n6155) );
  NAND2_X1 U7720 ( .A1(n6110), .A2(n6151), .ZN(n6152) );
  NAND2_X1 U7721 ( .A1(n6152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U7722 ( .A(n6153), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U7723 ( .A1(n8639), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5921), .B2(
        n9720), .ZN(n6154) );
  NAND2_X1 U7724 ( .A1(n9336), .A2(n6346), .ZN(n6165) );
  NAND2_X1 U7725 ( .A1(n5916), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6163) );
  INV_X1 U7726 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7727 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  AND2_X1 U7728 ( .A1(n6180), .A2(n6159), .ZN(n9256) );
  NAND2_X1 U7729 ( .A1(n6298), .A2(n9256), .ZN(n6162) );
  NAND2_X1 U7730 ( .A1(n8649), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7731 ( .A1(n8650), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6160) );
  OR2_X1 U7732 ( .A1(n8579), .A2(n6379), .ZN(n6164) );
  NAND2_X1 U7733 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  XNOR2_X1 U7734 ( .A(n6166), .B(n6255), .ZN(n6169) );
  NOR2_X1 U7735 ( .A1(n8579), .A2(n6378), .ZN(n6167) );
  AOI21_X1 U7736 ( .B1(n9336), .B2(n6356), .A(n6167), .ZN(n6168) );
  NAND2_X1 U7737 ( .A1(n6169), .A2(n6168), .ZN(n6172) );
  OR2_X1 U7738 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7739 ( .A1(n6172), .A2(n6170), .ZN(n8568) );
  INV_X1 U7740 ( .A(n8568), .ZN(n6171) );
  NAND2_X1 U7741 ( .A1(n7061), .A2(n8645), .ZN(n6178) );
  NAND2_X1 U7742 ( .A1(n6173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6175) );
  OR2_X1 U7743 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  NAND2_X1 U7744 ( .A1(n6175), .A2(n6174), .ZN(n6194) );
  AOI22_X1 U7745 ( .A1(n8639), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5921), .B2(
        n9731), .ZN(n6177) );
  NAND2_X1 U7746 ( .A1(n9329), .A2(n6346), .ZN(n6187) );
  NAND2_X1 U7747 ( .A1(n5916), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6185) );
  INV_X1 U7748 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7749 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  AND2_X1 U7750 ( .A1(n6200), .A2(n6181), .ZN(n9228) );
  NAND2_X1 U7751 ( .A1(n6298), .A2(n9228), .ZN(n6184) );
  NAND2_X1 U7752 ( .A1(n6232), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7753 ( .A1(n8650), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6182) );
  NAND4_X1 U7754 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n9222)
         );
  NAND2_X1 U7755 ( .A1(n9222), .A2(n6356), .ZN(n6186) );
  NAND2_X1 U7756 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  XNOR2_X1 U7757 ( .A(n6188), .B(n7222), .ZN(n6190) );
  AND2_X1 U7758 ( .A1(n9222), .A2(n5909), .ZN(n6189) );
  AOI21_X1 U7759 ( .B1(n9329), .B2(n6356), .A(n6189), .ZN(n6191) );
  XNOR2_X1 U7760 ( .A(n6190), .B(n6191), .ZN(n8576) );
  NAND2_X1 U7761 ( .A1(n8575), .A2(n8576), .ZN(n8574) );
  INV_X1 U7762 ( .A(n6190), .ZN(n6192) );
  NAND2_X1 U7763 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  AND2_X2 U7764 ( .A1(n8574), .A2(n6193), .ZN(n6210) );
  NAND2_X1 U7765 ( .A1(n7243), .A2(n8645), .ZN(n6197) );
  NAND2_X1 U7766 ( .A1(n6194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6195) );
  XNOR2_X1 U7767 ( .A(n6195), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U7768 ( .A1(n8639), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5921), .B2(
        n9747), .ZN(n6196) );
  NAND2_X1 U7769 ( .A1(n9324), .A2(n6346), .ZN(n6207) );
  NAND2_X1 U7770 ( .A1(n5916), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6205) );
  INV_X1 U7771 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7772 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  AND2_X1 U7773 ( .A1(n6216), .A2(n6201), .ZN(n9214) );
  NAND2_X1 U7774 ( .A1(n6298), .A2(n9214), .ZN(n6204) );
  NAND2_X1 U7775 ( .A1(n8649), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7776 ( .A1(n8650), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6202) );
  OR2_X1 U7777 ( .A1(n9197), .A2(n6379), .ZN(n6206) );
  NAND2_X1 U7778 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  XNOR2_X1 U7779 ( .A(n6208), .B(n7222), .ZN(n6211) );
  NOR2_X1 U7780 ( .A1(n9197), .A2(n6378), .ZN(n6209) );
  AOI21_X1 U7781 ( .B1(n9324), .B2(n6356), .A(n6209), .ZN(n8616) );
  NAND2_X1 U7782 ( .A1(n7342), .A2(n8645), .ZN(n6213) );
  AOI22_X1 U7783 ( .A1(n8639), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9018), .B2(
        n5921), .ZN(n6212) );
  INV_X1 U7784 ( .A(n6216), .ZN(n6214) );
  NAND2_X1 U7785 ( .A1(n6214), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6228) );
  INV_X1 U7786 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7787 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  AND2_X1 U7788 ( .A1(n6228), .A2(n6217), .ZN(n9204) );
  NAND2_X1 U7789 ( .A1(n6298), .A2(n9204), .ZN(n6221) );
  NAND2_X1 U7790 ( .A1(n8649), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7791 ( .A1(n5916), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7792 ( .A1(n8650), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6218) );
  OAI22_X1 U7793 ( .A1(n9208), .A2(n6380), .B1(n9182), .B2(n6379), .ZN(n6222)
         );
  XNOR2_X1 U7794 ( .A(n6222), .B(n7222), .ZN(n6224) );
  OAI22_X1 U7795 ( .A1(n9208), .A2(n6379), .B1(n9182), .B2(n6378), .ZN(n6223)
         );
  NAND2_X1 U7796 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AND2_X1 U7797 ( .A1(n8592), .A2(n6225), .ZN(n8538) );
  NAND2_X1 U7798 ( .A1(n7431), .A2(n8645), .ZN(n6227) );
  NAND2_X1 U7799 ( .A1(n8639), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7800 ( .A1(n9316), .A2(n6346), .ZN(n6236) );
  INV_X1 U7801 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U7802 ( .A1(n6228), .A2(n8596), .ZN(n6229) );
  NAND2_X1 U7803 ( .A1(n6248), .A2(n6229), .ZN(n9185) );
  NAND2_X1 U7804 ( .A1(n5916), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7805 ( .A1(n8650), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6230) );
  AND2_X1 U7806 ( .A1(n6231), .A2(n6230), .ZN(n6234) );
  NAND2_X1 U7807 ( .A1(n6232), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U7808 ( .C1(n9185), .C2(n6425), .A(n6234), .B(n6233), .ZN(n9162)
         );
  NAND2_X1 U7809 ( .A1(n9162), .A2(n6356), .ZN(n6235) );
  NAND2_X1 U7810 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  XNOR2_X1 U7811 ( .A(n6237), .B(n6255), .ZN(n6239) );
  AND2_X1 U7812 ( .A1(n9162), .A2(n5909), .ZN(n6238) );
  AOI21_X1 U7813 ( .B1(n9316), .B2(n6356), .A(n6238), .ZN(n6240) );
  NAND2_X1 U7814 ( .A1(n6239), .A2(n6240), .ZN(n6244) );
  INV_X1 U7815 ( .A(n6239), .ZN(n6242) );
  INV_X1 U7816 ( .A(n6240), .ZN(n6241) );
  NAND2_X1 U7817 ( .A1(n6242), .A2(n6241), .ZN(n6243) );
  NAND2_X1 U7818 ( .A1(n6244), .A2(n6243), .ZN(n8591) );
  INV_X1 U7819 ( .A(n6244), .ZN(n8549) );
  NAND2_X1 U7820 ( .A1(n7461), .A2(n8645), .ZN(n6246) );
  NAND2_X1 U7821 ( .A1(n8639), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7822 ( .A1(n9310), .A2(n6346), .ZN(n6254) );
  INV_X1 U7823 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7824 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  AND2_X1 U7825 ( .A1(n6267), .A2(n6249), .ZN(n9167) );
  NAND2_X1 U7826 ( .A1(n9167), .A2(n6298), .ZN(n6252) );
  AOI22_X1 U7827 ( .A1(n5916), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n8649), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7828 ( .A1(n8650), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6250) );
  INV_X1 U7829 ( .A(n9183), .ZN(n8964) );
  NAND2_X1 U7830 ( .A1(n8964), .A2(n6356), .ZN(n6253) );
  NAND2_X1 U7831 ( .A1(n6254), .A2(n6253), .ZN(n6256) );
  XNOR2_X1 U7832 ( .A(n6256), .B(n6255), .ZN(n6258) );
  NOR2_X1 U7833 ( .A1(n9183), .A2(n6378), .ZN(n6257) );
  AOI21_X1 U7834 ( .B1(n9310), .B2(n6356), .A(n6257), .ZN(n6259) );
  NAND2_X1 U7835 ( .A1(n6258), .A2(n6259), .ZN(n6263) );
  INV_X1 U7836 ( .A(n6258), .ZN(n6261) );
  INV_X1 U7837 ( .A(n6259), .ZN(n6260) );
  NAND2_X1 U7838 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  AND2_X1 U7839 ( .A1(n6263), .A2(n6262), .ZN(n8548) );
  NAND2_X1 U7840 ( .A1(n8547), .A2(n6263), .ZN(n6276) );
  NAND2_X1 U7841 ( .A1(n7609), .A2(n8645), .ZN(n6265) );
  NAND2_X1 U7842 ( .A1(n8639), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6264) );
  INV_X1 U7843 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U7844 ( .A1(n6267), .A2(n8607), .ZN(n6268) );
  NAND2_X1 U7845 ( .A1(n6281), .A2(n6268), .ZN(n9146) );
  OR2_X1 U7846 ( .A1(n9146), .A2(n6425), .ZN(n6273) );
  INV_X1 U7847 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U7848 ( .A1(n5916), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7849 ( .A1(n8650), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7850 ( .C1(n5954), .C2(n9147), .A(n6270), .B(n6269), .ZN(n6271)
         );
  INV_X1 U7851 ( .A(n6271), .ZN(n6272) );
  AOI22_X1 U7852 ( .A1(n9305), .A2(n6356), .B1(n5909), .B2(n9161), .ZN(n6275)
         );
  NAND2_X1 U7853 ( .A1(n6276), .A2(n6275), .ZN(n8602) );
  OAI22_X1 U7854 ( .A1(n9144), .A2(n6380), .B1(n8553), .B2(n6379), .ZN(n6274)
         );
  XNOR2_X1 U7855 ( .A(n6274), .B(n7222), .ZN(n8605) );
  NAND2_X1 U7856 ( .A1(n7666), .A2(n8645), .ZN(n6278) );
  NAND2_X1 U7857 ( .A1(n8639), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6277) );
  INV_X1 U7858 ( .A(n6281), .ZN(n6279) );
  INV_X1 U7859 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7860 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U7861 ( .A1(n6296), .A2(n6282), .ZN(n9129) );
  OR2_X1 U7862 ( .A1(n9129), .A2(n6425), .ZN(n6288) );
  INV_X1 U7863 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7864 ( .A1(n5916), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7865 ( .A1(n8650), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6283) );
  OAI211_X1 U7866 ( .C1(n5954), .C2(n6285), .A(n6284), .B(n6283), .ZN(n6286)
         );
  INV_X1 U7867 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U7868 ( .A1(n6288), .A2(n6287), .ZN(n8963) );
  OAI22_X1 U7869 ( .A1(n9132), .A2(n6380), .B1(n9153), .B2(n6379), .ZN(n6289)
         );
  XOR2_X1 U7870 ( .A(n7222), .B(n6289), .Z(n6290) );
  NAND2_X1 U7871 ( .A1(n8531), .A2(n6290), .ZN(n6292) );
  OAI22_X1 U7872 ( .A1(n9132), .A2(n6379), .B1(n9153), .B2(n6378), .ZN(n8528)
         );
  INV_X1 U7873 ( .A(n8531), .ZN(n6291) );
  INV_X1 U7874 ( .A(n6290), .ZN(n8529) );
  NAND2_X1 U7875 ( .A1(n7709), .A2(n8645), .ZN(n6294) );
  NAND2_X1 U7876 ( .A1(n8639), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6293) );
  INV_X1 U7877 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7878 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  AND2_X1 U7879 ( .A1(n6316), .A2(n6297), .ZN(n9119) );
  NAND2_X1 U7880 ( .A1(n9119), .A2(n6298), .ZN(n6304) );
  INV_X1 U7881 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7882 ( .A1(n5916), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7883 ( .A1(n8650), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6299) );
  OAI211_X1 U7884 ( .C1(n5954), .C2(n6301), .A(n6300), .B(n6299), .ZN(n6302)
         );
  INV_X1 U7885 ( .A(n6302), .ZN(n6303) );
  OAI22_X1 U7886 ( .A1(n9122), .A2(n6380), .B1(n9107), .B2(n6379), .ZN(n6305)
         );
  XNOR2_X1 U7887 ( .A(n6305), .B(n7222), .ZN(n6309) );
  OR2_X1 U7888 ( .A1(n9122), .A2(n6379), .ZN(n6307) );
  NAND2_X1 U7889 ( .A1(n9136), .A2(n5909), .ZN(n6306) );
  NAND2_X1 U7890 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  NOR2_X1 U7891 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  AOI21_X1 U7892 ( .B1(n6309), .B2(n6308), .A(n6310), .ZN(n8584) );
  NAND2_X1 U7893 ( .A1(n8585), .A2(n8584), .ZN(n8583) );
  INV_X1 U7894 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U7895 ( .A1(n8583), .A2(n6311), .ZN(n8558) );
  NAND2_X1 U7896 ( .A1(n7793), .A2(n8645), .ZN(n6313) );
  NAND2_X1 U7897 ( .A1(n8639), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7898 ( .A1(n9290), .A2(n6346), .ZN(n6324) );
  INV_X1 U7899 ( .A(n6316), .ZN(n6314) );
  NAND2_X1 U7900 ( .A1(n6314), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6328) );
  INV_X1 U7901 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7902 ( .A1(n6316), .A2(n6315), .ZN(n6317) );
  NAND2_X1 U7903 ( .A1(n6328), .A2(n6317), .ZN(n9101) );
  INV_X1 U7904 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U7905 ( .A1(n5916), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7906 ( .A1(n8650), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6318) );
  OAI211_X1 U7907 ( .C1(n5954), .C2(n9100), .A(n6319), .B(n6318), .ZN(n6320)
         );
  INV_X1 U7908 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U7909 ( .A1(n9090), .A2(n6356), .ZN(n6323) );
  NAND2_X1 U7910 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  XNOR2_X1 U7911 ( .A(n6325), .B(n7222), .ZN(n6340) );
  AOI22_X1 U7912 ( .A1(n9290), .A2(n6356), .B1(n5909), .B2(n9090), .ZN(n6341)
         );
  XNOR2_X1 U7913 ( .A(n6340), .B(n6341), .ZN(n8559) );
  NAND2_X1 U7914 ( .A1(n7857), .A2(n8645), .ZN(n6327) );
  NAND2_X1 U7915 ( .A1(n8639), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7916 ( .A1(n9283), .A2(n6346), .ZN(n6337) );
  INV_X1 U7917 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U7918 ( .A1(n6328), .A2(n8629), .ZN(n6329) );
  NAND2_X1 U7919 ( .A1(n9083), .A2(n6298), .ZN(n6335) );
  INV_X1 U7920 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7921 ( .A1(n5916), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7922 ( .A1(n8650), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6330) );
  OAI211_X1 U7923 ( .C1(n5954), .C2(n6332), .A(n6331), .B(n6330), .ZN(n6333)
         );
  INV_X1 U7924 ( .A(n6333), .ZN(n6334) );
  NAND2_X1 U7925 ( .A1(n8962), .A2(n6356), .ZN(n6336) );
  NAND2_X1 U7926 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  XNOR2_X1 U7927 ( .A(n6338), .B(n7222), .ZN(n6363) );
  AND2_X1 U7928 ( .A1(n8962), .A2(n5909), .ZN(n6339) );
  AOI21_X1 U7929 ( .B1(n9283), .B2(n6356), .A(n6339), .ZN(n6361) );
  XNOR2_X1 U7930 ( .A(n6363), .B(n6361), .ZN(n8627) );
  INV_X1 U7931 ( .A(n6340), .ZN(n6342) );
  NAND2_X1 U7932 ( .A1(n6342), .A2(n6341), .ZN(n8624) );
  NAND2_X1 U7933 ( .A1(n8509), .A2(n8645), .ZN(n6345) );
  NAND2_X1 U7934 ( .A1(n8639), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U7935 ( .A1(n9280), .A2(n6346), .ZN(n6354) );
  XNOR2_X1 U7936 ( .A(n6368), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U7937 ( .A1(n8524), .A2(n6298), .ZN(n6352) );
  INV_X1 U7938 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7939 ( .A1(n5916), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7940 ( .A1(n8650), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6347) );
  OAI211_X1 U7941 ( .C1(n6349), .C2(n5954), .A(n6348), .B(n6347), .ZN(n6350)
         );
  INV_X1 U7942 ( .A(n6350), .ZN(n6351) );
  NAND2_X1 U7943 ( .A1(n9091), .A2(n6356), .ZN(n6353) );
  NAND2_X1 U7944 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  XNOR2_X1 U7945 ( .A(n6355), .B(n7222), .ZN(n6360) );
  NAND2_X1 U7946 ( .A1(n9280), .A2(n6356), .ZN(n6358) );
  NAND2_X1 U7947 ( .A1(n9091), .A2(n5909), .ZN(n6357) );
  NAND2_X1 U7948 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NOR2_X1 U7949 ( .A1(n6360), .A2(n6359), .ZN(n6365) );
  AOI21_X1 U7950 ( .B1(n6360), .B2(n6359), .A(n6365), .ZN(n8517) );
  INV_X1 U7951 ( .A(n6361), .ZN(n6362) );
  NAND2_X1 U7952 ( .A1(n6363), .A2(n6362), .ZN(n8518) );
  NAND2_X1 U7953 ( .A1(n8516), .A2(n6364), .ZN(n8515) );
  NAND2_X1 U7954 ( .A1(n8506), .A2(n8645), .ZN(n6367) );
  NAND2_X1 U7955 ( .A1(n8639), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6366) );
  INV_X1 U7956 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8521) );
  INV_X1 U7957 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6438) );
  OAI21_X1 U7958 ( .B1(n6368), .B2(n8521), .A(n6438), .ZN(n6371) );
  INV_X1 U7959 ( .A(n6368), .ZN(n6370) );
  AND2_X1 U7960 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6369) );
  NAND2_X1 U7961 ( .A1(n6370), .A2(n6369), .ZN(n9051) );
  NAND2_X1 U7962 ( .A1(n6371), .A2(n9051), .ZN(n9064) );
  INV_X1 U7963 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7964 ( .A1(n5916), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7965 ( .A1(n8650), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U7966 ( .C1(n5954), .C2(n6374), .A(n6373), .B(n6372), .ZN(n6375)
         );
  INV_X1 U7967 ( .A(n6375), .ZN(n6376) );
  OAI22_X1 U7968 ( .A1(n9067), .A2(n6379), .B1(n9049), .B2(n6378), .ZN(n6383)
         );
  OAI22_X1 U7969 ( .A1(n9067), .A2(n6380), .B1(n9049), .B2(n6379), .ZN(n6381)
         );
  XNOR2_X1 U7970 ( .A(n6381), .B(n7222), .ZN(n6382) );
  XOR2_X1 U7971 ( .A(n6383), .B(n6382), .Z(n6384) );
  NAND2_X1 U7972 ( .A1(n5878), .A2(n6386), .ZN(n7033) );
  INV_X1 U7973 ( .A(n7033), .ZN(n6387) );
  NAND3_X1 U7974 ( .A1(n6388), .A2(P1_B_REG_SCAN_IN), .A3(n7752), .ZN(n6392)
         );
  INV_X1 U7975 ( .A(n7752), .ZN(n6390) );
  INV_X1 U7976 ( .A(P1_B_REG_SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7977 ( .A1(n6390), .A2(n6389), .ZN(n6391) );
  AND2_X1 U7978 ( .A1(n6392), .A2(n6391), .ZN(n6394) );
  NOR4_X1 U7979 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6398) );
  NOR4_X1 U7980 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6397) );
  NOR4_X1 U7981 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6396) );
  NOR4_X1 U7982 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6395) );
  NAND4_X1 U7983 ( .A1(n6398), .A2(n6397), .A3(n6396), .A4(n6395), .ZN(n6404)
         );
  NOR2_X1 U7984 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6402) );
  NOR4_X1 U7985 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6401) );
  NOR4_X1 U7986 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6400) );
  NOR4_X1 U7987 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6399) );
  NAND4_X1 U7988 ( .A1(n6402), .A2(n6401), .A3(n6400), .A4(n6399), .ZN(n6403)
         );
  NOR2_X1 U7989 ( .A1(n6404), .A2(n6403), .ZN(n6766) );
  NAND2_X1 U7990 ( .A1(n6766), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7991 ( .A1(n6768), .A2(n6405), .ZN(n6406) );
  INV_X1 U7992 ( .A(n6393), .ZN(n7862) );
  NAND2_X1 U7993 ( .A1(n7862), .A2(n7752), .ZN(n6764) );
  NAND2_X1 U7994 ( .A1(n6406), .A2(n6764), .ZN(n6742) );
  INV_X1 U7995 ( .A(n6742), .ZN(n6410) );
  INV_X1 U7996 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7997 ( .A1(n6768), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U7998 ( .A1(n7862), .A2(n6388), .ZN(n6408) );
  INV_X1 U7999 ( .A(n6433), .ZN(n6416) );
  NAND2_X1 U8000 ( .A1(n6411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6412) );
  MUX2_X1 U8001 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6412), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n6413) );
  NAND2_X1 U8002 ( .A1(n6413), .A2(n4351), .ZN(n7669) );
  AND2_X1 U8003 ( .A1(n7669), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6414) );
  INV_X1 U8004 ( .A(n7098), .ZN(n8952) );
  OR2_X1 U8005 ( .A1(n6416), .A2(n8952), .ZN(n6420) );
  INV_X1 U8006 ( .A(n7030), .ZN(n6745) );
  NOR2_X1 U8007 ( .A1(n6420), .A2(n6745), .ZN(n6415) );
  NOR2_X1 U8008 ( .A1(n7033), .A2(n8947), .ZN(n7224) );
  AND2_X1 U8009 ( .A1(n6416), .A2(n7098), .ZN(n6417) );
  NAND2_X1 U8010 ( .A1(n7224), .A2(n6417), .ZN(n6436) );
  INV_X1 U8011 ( .A(n6772), .ZN(n6419) );
  INV_X1 U8012 ( .A(n6420), .ZN(n6422) );
  OR2_X1 U8013 ( .A1(n7026), .A2(n7025), .ZN(n8953) );
  INV_X1 U8014 ( .A(n8953), .ZN(n6421) );
  NAND2_X1 U8015 ( .A1(n6422), .A2(n6421), .ZN(n6439) );
  INV_X1 U8016 ( .A(n6439), .ZN(n6424) );
  OR2_X1 U8017 ( .A1(n9051), .A2(n6425), .ZN(n6431) );
  INV_X1 U8018 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8019 ( .A1(n8649), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8020 ( .A1(n8650), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6426) );
  OAI211_X1 U8021 ( .C1(n6428), .C2(n5899), .A(n6427), .B(n6426), .ZN(n6429)
         );
  INV_X1 U8022 ( .A(n6429), .ZN(n6430) );
  AND3_X1 U8023 ( .A1(n6432), .A2(n6504), .A3(n7669), .ZN(n6434) );
  OR2_X1 U8024 ( .A1(n9347), .A2(n6433), .ZN(n6739) );
  NAND2_X1 U8025 ( .A1(n6434), .A2(n6739), .ZN(n6435) );
  NAND2_X1 U8026 ( .A1(n6435), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6437) );
  OAI22_X1 U8027 ( .A1(n9064), .A2(n9625), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6438), .ZN(n6441) );
  NOR2_X1 U8028 ( .A1(n8631), .A2(n9611), .ZN(n6440) );
  AOI211_X1 U8029 ( .C1(n9608), .C2(n9072), .A(n6441), .B(n6440), .ZN(n6442)
         );
  INV_X1 U8030 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8031 ( .A1(n6446), .A2(n6445), .ZN(n6450) );
  NAND2_X1 U8032 ( .A1(n6447), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U8033 ( .A1(n6450), .A2(n6449), .ZN(n9932) );
  NAND2_X1 U8034 ( .A1(n9932), .A2(n9933), .ZN(n6452) );
  NAND2_X1 U8035 ( .A1(n6935), .A2(n9968), .ZN(n6451) );
  NAND2_X1 U8036 ( .A1(n6452), .A2(n6451), .ZN(n9903) );
  NAND2_X1 U8037 ( .A1(n9903), .A2(n9904), .ZN(n6455) );
  NAND2_X1 U8038 ( .A1(n6453), .A2(n9973), .ZN(n6454) );
  NAND2_X1 U8039 ( .A1(n6455), .A2(n6454), .ZN(n7083) );
  NAND2_X1 U8040 ( .A1(n6456), .A2(n9979), .ZN(n6457) );
  NAND2_X1 U8041 ( .A1(n8101), .A2(n4315), .ZN(n6458) );
  NAND2_X1 U8042 ( .A1(n8100), .A2(n9858), .ZN(n6459) );
  NAND2_X1 U8043 ( .A1(n6460), .A2(n6459), .ZN(n7068) );
  INV_X1 U8044 ( .A(n7068), .ZN(n6461) );
  NAND2_X1 U8045 ( .A1(n7264), .A2(n7231), .ZN(n6462) );
  OR2_X1 U8046 ( .A1(n7475), .A2(n8096), .ZN(n6464) );
  AND2_X2 U8047 ( .A1(n7312), .A2(n6464), .ZN(n7593) );
  NAND2_X1 U8048 ( .A1(n9877), .A2(n8095), .ZN(n6465) );
  OAI22_X2 U8049 ( .A1(n7672), .A2(n7674), .B1(n8091), .B2(n9638), .ZN(n7735)
         );
  NAND2_X1 U8050 ( .A1(n8357), .A2(n8087), .ZN(n6469) );
  NAND2_X1 U8051 ( .A1(n8433), .A2(n8084), .ZN(n6472) );
  OAI22_X2 U8052 ( .A1(n8229), .A2(n8231), .B1(n8406), .B2(n8079), .ZN(n8214)
         );
  AOI22_X2 U8053 ( .A1(n8214), .A2(n8216), .B1(n4485), .B2(n6474), .ZN(n8205)
         );
  OAI22_X1 U8054 ( .A1(n8205), .A2(n8204), .B1(n8077), .B2(n8207), .ZN(n6476)
         );
  XNOR2_X1 U8055 ( .A(n6476), .B(n6475), .ZN(n8189) );
  XNOR2_X1 U8056 ( .A(n7944), .B(n6970), .ZN(n6477) );
  NOR2_X1 U8057 ( .A1(n6478), .A2(n7343), .ZN(n6479) );
  NAND2_X1 U8058 ( .A1(n6479), .A2(n7944), .ZN(n7594) );
  XOR2_X1 U8059 ( .A(n6481), .B(n6480), .Z(n6486) );
  INV_X1 U8060 ( .A(n9832), .ZN(n8055) );
  NAND2_X1 U8061 ( .A1(n8511), .A2(P2_B_REG_SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8062 ( .A1(n9834), .A2(n6483), .ZN(n8177) );
  OAI22_X1 U8063 ( .A1(n6484), .A2(n8055), .B1(n6595), .B2(n8177), .ZN(n6485)
         );
  AOI21_X1 U8064 ( .B1(n6486), .B2(n9922), .A(n6485), .ZN(n8199) );
  NAND2_X1 U8065 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  INV_X1 U8066 ( .A(n7475), .ZN(n7327) );
  INV_X1 U8067 ( .A(n7663), .ZN(n10003) );
  NAND2_X1 U8068 ( .A1(n8328), .A2(n8318), .ZN(n8298) );
  INV_X1 U8069 ( .A(n6487), .ZN(n8206) );
  INV_X1 U8070 ( .A(n10004), .ZN(n9926) );
  OAI211_X1 U8071 ( .C1(n6499), .C2(n8206), .A(n9926), .B(n8181), .ZN(n8193)
         );
  NAND2_X1 U8072 ( .A1(n6969), .A2(n6964), .ZN(n6494) );
  NOR2_X1 U8073 ( .A1(n6966), .A2(n6494), .ZN(n6490) );
  NAND2_X1 U8074 ( .A1(n8196), .A2(n6492), .ZN(n6493) );
  INV_X1 U8075 ( .A(n6494), .ZN(n6495) );
  AND2_X1 U8076 ( .A1(n6966), .A2(n6495), .ZN(n6496) );
  MUX2_X1 U8077 ( .A(n6498), .B(n6497), .S(n10012), .Z(n6502) );
  NAND2_X1 U8078 ( .A1(n8196), .A2(n6500), .ZN(n6501) );
  NAND2_X1 U8079 ( .A1(n6502), .A2(n6501), .ZN(P2_U3517) );
  INV_X1 U8080 ( .A(n7669), .ZN(n6503) );
  NAND2_X1 U8081 ( .A1(n7030), .A2(n6504), .ZN(n6505) );
  NAND2_X1 U8082 ( .A1(n6505), .A2(n7669), .ZN(n6518) );
  NAND2_X1 U8083 ( .A1(n6518), .A2(n6506), .ZN(n6586) );
  NAND2_X1 U8084 ( .A1(n6586), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8085 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U8086 ( .A1(n6688), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6508) );
  OAI21_X1 U8087 ( .B1(n6688), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6508), .ZN(
        n6516) );
  INV_X1 U8088 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6514) );
  INV_X1 U8089 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6513) );
  INV_X1 U8090 ( .A(n6804), .ZN(n6511) );
  INV_X1 U8091 ( .A(n6676), .ZN(n6525) );
  INV_X1 U8092 ( .A(n6777), .ZN(n6790) );
  INV_X1 U8093 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7109) );
  MUX2_X1 U8094 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7109), .S(n6553), .Z(n6645)
         );
  NAND2_X1 U8095 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6792) );
  INV_X1 U8096 ( .A(n6792), .ZN(n6644) );
  AND2_X1 U8097 ( .A1(n6645), .A2(n6644), .ZN(n6642) );
  AOI21_X1 U8098 ( .B1(n6553), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6642), .ZN(
        n6787) );
  XOR2_X1 U8099 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6777), .Z(n6786) );
  NOR2_X1 U8100 ( .A1(n6787), .A2(n6786), .ZN(n6785) );
  AOI21_X1 U8101 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6790), .A(n6785), .ZN(
        n6679) );
  INV_X1 U8102 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7308) );
  XNOR2_X1 U8103 ( .A(n6676), .B(n7308), .ZN(n6678) );
  INV_X1 U8104 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6509) );
  MUX2_X1 U8105 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6509), .S(n6804), .Z(n6510)
         );
  INV_X1 U8106 ( .A(n6510), .ZN(n6797) );
  XNOR2_X1 U8107 ( .A(n6637), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6630) );
  INV_X1 U8108 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6512) );
  AOI22_X1 U8109 ( .A1(n6631), .A2(n6630), .B1(n6637), .B2(n6512), .ZN(n6662)
         );
  MUX2_X1 U8110 ( .A(n6513), .B(P1_REG2_REG_6__SCAN_IN), .S(n6658), .Z(n6663)
         );
  NAND2_X1 U8111 ( .A1(n6662), .A2(n6663), .ZN(n6661) );
  XOR2_X1 U8112 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6619), .Z(n6618) );
  XNOR2_X1 U8113 ( .A(n6612), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U8114 ( .A1(n8951), .A2(n4309), .ZN(n9375) );
  NAND2_X1 U8115 ( .A1(n6518), .A2(n9375), .ZN(n9014) );
  INV_X1 U8116 ( .A(n9014), .ZN(n6534) );
  INV_X1 U8117 ( .A(n6423), .ZN(n6582) );
  NOR2_X1 U8118 ( .A1(n6515), .A2(n6516), .ZN(n6687) );
  AOI211_X1 U8119 ( .C1(n6516), .C2(n6515), .A(n9715), .B(n6687), .ZN(n6538)
         );
  NOR2_X1 U8120 ( .A1(n6423), .A2(P1_U3084), .ZN(n9372) );
  AND2_X1 U8121 ( .A1(n9372), .A2(n8951), .ZN(n6517) );
  INV_X1 U8122 ( .A(n6612), .ZN(n6567) );
  MUX2_X1 U8123 ( .A(n7058), .B(P1_REG1_REG_2__SCAN_IN), .S(n6777), .Z(n6521)
         );
  INV_X1 U8124 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6519) );
  MUX2_X1 U8125 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6519), .S(n6553), .Z(n6648)
         );
  AND2_X1 U8126 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6649) );
  NAND2_X1 U8127 ( .A1(n6648), .A2(n6649), .ZN(n6779) );
  NAND2_X1 U8128 ( .A1(n6553), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8129 ( .A1(n6779), .A2(n6778), .ZN(n6520) );
  NAND2_X1 U8130 ( .A1(n6521), .A2(n6520), .ZN(n6782) );
  NAND2_X1 U8131 ( .A1(n6790), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8132 ( .A1(n6782), .A2(n6671), .ZN(n6524) );
  INV_X1 U8133 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6522) );
  MUX2_X1 U8134 ( .A(n6522), .B(P1_REG1_REG_3__SCAN_IN), .S(n6676), .Z(n6523)
         );
  NAND2_X1 U8135 ( .A1(n6524), .A2(n6523), .ZN(n6674) );
  NAND2_X1 U8136 ( .A1(n6525), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6526) );
  AND2_X1 U8137 ( .A1(n6674), .A2(n6526), .ZN(n6801) );
  INV_X1 U8138 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7148) );
  MUX2_X1 U8139 ( .A(n7148), .B(P1_REG1_REG_4__SCAN_IN), .S(n6804), .Z(n6800)
         );
  NAND2_X1 U8140 ( .A1(n6801), .A2(n6800), .ZN(n6799) );
  NAND2_X1 U8141 ( .A1(n6804), .A2(n7148), .ZN(n6527) );
  NAND2_X1 U8142 ( .A1(n6799), .A2(n6527), .ZN(n6633) );
  INV_X1 U8143 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9796) );
  MUX2_X1 U8144 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9796), .S(n6637), .Z(n6632)
         );
  OR2_X1 U8145 ( .A1(n6633), .A2(n6632), .ZN(n6635) );
  OR2_X1 U8146 ( .A1(n6637), .A2(n9796), .ZN(n6528) );
  AND2_X1 U8147 ( .A1(n6635), .A2(n6528), .ZN(n6657) );
  INV_X1 U8148 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9798) );
  MUX2_X1 U8149 ( .A(n9798), .B(P1_REG1_REG_6__SCAN_IN), .S(n6658), .Z(n6656)
         );
  NAND2_X1 U8150 ( .A1(n6657), .A2(n6656), .ZN(n6655) );
  NAND2_X1 U8151 ( .A1(n6658), .A2(n9798), .ZN(n6621) );
  NAND2_X1 U8152 ( .A1(n6655), .A2(n6621), .ZN(n6529) );
  INV_X1 U8153 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9800) );
  MUX2_X1 U8154 ( .A(n9800), .B(P1_REG1_REG_7__SCAN_IN), .S(n6619), .Z(n6620)
         );
  NAND2_X1 U8155 ( .A1(n6529), .A2(n6620), .ZN(n6624) );
  NAND2_X1 U8156 ( .A1(n6619), .A2(n9800), .ZN(n6530) );
  NAND2_X1 U8157 ( .A1(n6624), .A2(n6530), .ZN(n6607) );
  INV_X1 U8158 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7565) );
  MUX2_X1 U8159 ( .A(n7565), .B(P1_REG1_REG_8__SCAN_IN), .S(n6612), .Z(n6606)
         );
  OR2_X1 U8160 ( .A1(n6607), .A2(n6606), .ZN(n6609) );
  OAI21_X1 U8161 ( .B1(n6567), .B2(n7565), .A(n6609), .ZN(n6532) );
  INV_X1 U8162 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9804) );
  INV_X1 U8163 ( .A(n6688), .ZN(n6591) );
  AOI22_X1 U8164 ( .A1(n6688), .A2(n9804), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6591), .ZN(n6531) );
  NOR2_X1 U8165 ( .A1(n6532), .A2(n6531), .ZN(n6683) );
  AOI21_X1 U8166 ( .B1(n6532), .B2(n6531), .A(n6683), .ZN(n6533) );
  NOR2_X1 U8167 ( .A1(n9756), .A2(n6533), .ZN(n6537) );
  OR2_X1 U8168 ( .A1(P1_U3083), .A2(n6535), .ZN(n9759) );
  INV_X1 U8169 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10057) );
  OAI22_X1 U8170 ( .A1(n6994), .A2(n6591), .B1(n9759), .B2(n10057), .ZN(n6536)
         );
  OR4_X1 U8171 ( .A1(n7468), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(P1_U3250)
         );
  XNOR2_X1 U8172 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U8173 ( .A(n8510), .ZN(n7947) );
  INV_X1 U8174 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6540) );
  OR2_X2 U8175 ( .A1(n4401), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8513) );
  INV_X1 U8176 ( .A(n6824), .ZN(n6717) );
  OAI222_X1 U8177 ( .A1(n7947), .A2(n6540), .B1(n8513), .B2(n6542), .C1(
        P2_U3152), .C2(n6717), .ZN(P2_U3355) );
  OR2_X2 U8178 ( .A1(n4401), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9369) );
  OAI222_X1 U8179 ( .A1(n9369), .A2(n6541), .B1(n9378), .B2(n6546), .C1(n4309), 
        .C2(n6777), .ZN(P1_U3351) );
  OAI222_X1 U8180 ( .A1(n9369), .A2(n6543), .B1(n9378), .B2(n6542), .C1(
        P1_U3084), .C2(n6676), .ZN(P1_U3350) );
  INV_X1 U8181 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6544) );
  OAI222_X1 U8182 ( .A1(n7947), .A2(n6544), .B1(n8513), .B2(n6554), .C1(
        P2_U3152), .C2(n5045), .ZN(P2_U3357) );
  INV_X1 U8183 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6545) );
  INV_X1 U8184 ( .A(n6823), .ZN(n6889) );
  OAI222_X1 U8185 ( .A1(n7947), .A2(n6545), .B1(n8513), .B2(n6551), .C1(
        P2_U3152), .C2(n6889), .ZN(P2_U3354) );
  INV_X1 U8186 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6547) );
  INV_X1 U8187 ( .A(n8120), .ZN(n6711) );
  OAI222_X1 U8188 ( .A1(n7947), .A2(n6547), .B1(n8513), .B2(n6546), .C1(
        P2_U3152), .C2(n6711), .ZN(P2_U3356) );
  INV_X1 U8189 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6548) );
  INV_X1 U8190 ( .A(n6821), .ZN(n6901) );
  OAI222_X1 U8191 ( .A1(n7947), .A2(n6548), .B1(n8513), .B2(n6549), .C1(
        P2_U3152), .C2(n6901), .ZN(P2_U3353) );
  OAI222_X1 U8192 ( .A1(n9369), .A2(n6550), .B1(n9378), .B2(n6549), .C1(n4309), 
        .C2(n6637), .ZN(P1_U3348) );
  OAI222_X1 U8193 ( .A1(n9369), .A2(n6552), .B1(n9378), .B2(n6551), .C1(
        P1_U3084), .C2(n6804), .ZN(P1_U3349) );
  INV_X1 U8194 ( .A(n6553), .ZN(n6647) );
  OAI222_X1 U8195 ( .A1(n9369), .A2(n6555), .B1(n9378), .B2(n6554), .C1(n4309), 
        .C2(n6647), .ZN(P1_U3352) );
  OAI222_X1 U8196 ( .A1(n9369), .A2(n6556), .B1(n9378), .B2(n6557), .C1(
        P1_U3084), .C2(n6658), .ZN(P1_U3347) );
  INV_X1 U8197 ( .A(n6820), .ZN(n6876) );
  OAI222_X1 U8198 ( .A1(n7947), .A2(n6558), .B1(n8513), .B2(n6557), .C1(
        P2_U3152), .C2(n6876), .ZN(P2_U3352) );
  NAND2_X1 U8199 ( .A1(n7096), .A2(n7098), .ZN(n6559) );
  OAI21_X1 U8200 ( .B1(n7098), .B2(n6407), .A(n6559), .ZN(P1_U3441) );
  INV_X1 U8201 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6560) );
  INV_X1 U8202 ( .A(n6843), .ZN(n6835) );
  OAI222_X1 U8203 ( .A1(n7947), .A2(n6560), .B1(n8513), .B2(n6561), .C1(
        P2_U3152), .C2(n6835), .ZN(P2_U3351) );
  OAI222_X1 U8204 ( .A1(n9369), .A2(n6562), .B1(n9378), .B2(n6561), .C1(n4309), 
        .C2(n6619), .ZN(P1_U3346) );
  INV_X1 U8205 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8206 ( .A1(P2_U3966), .A2(n6563), .ZN(n6564) );
  OAI21_X1 U8207 ( .B1(P2_U3966), .B2(n6565), .A(n6564), .ZN(P2_U3583) );
  INV_X1 U8208 ( .A(n6566), .ZN(n6569) );
  OAI222_X1 U8209 ( .A1(n9369), .A2(n6568), .B1(n9378), .B2(n6569), .C1(
        P1_U3084), .C2(n6567), .ZN(P1_U3345) );
  INV_X1 U8210 ( .A(n6854), .ZN(n6859) );
  OAI222_X1 U8211 ( .A1(n7947), .A2(n6570), .B1(n8513), .B2(n6569), .C1(
        P2_U3152), .C2(n6859), .ZN(P2_U3350) );
  INV_X1 U8212 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6763) );
  INV_X1 U8213 ( .A(n6768), .ZN(n6571) );
  INV_X1 U8214 ( .A(n9760), .ZN(n6572) );
  OAI21_X1 U8215 ( .B1(n6572), .B2(P1_D_REG_0__SCAN_IN), .A(n6764), .ZN(n6573)
         );
  OAI21_X1 U8216 ( .B1(n6763), .B2(n7098), .A(n6573), .ZN(P1_U3440) );
  NAND2_X1 U8217 ( .A1(n8035), .A2(n6699), .ZN(n6577) );
  NAND2_X1 U8218 ( .A1(n9944), .A2(n6696), .ZN(n6575) );
  NAND2_X1 U8219 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  NOR2_X1 U8220 ( .A1(n9866), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8221 ( .A(n6578), .ZN(n6592) );
  INV_X1 U8222 ( .A(n6921), .ZN(n6927) );
  OAI222_X1 U8223 ( .A1(n8513), .A2(n6592), .B1(n6927), .B2(P2_U3152), .C1(
        n6579), .C2(n7947), .ZN(P2_U3349) );
  INV_X1 U8224 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6590) );
  NOR2_X1 U8225 ( .A1(n8951), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U8226 ( .B1(n6423), .B2(n6580), .A(n4465), .ZN(n6793) );
  INV_X1 U8227 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6749) );
  INV_X1 U8228 ( .A(n8951), .ZN(n9025) );
  NAND2_X1 U8229 ( .A1(n9025), .A2(n6792), .ZN(n6581) );
  OAI211_X1 U8230 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6749), .A(n6582), .B(n6581), .ZN(n6583) );
  NAND3_X1 U8231 ( .A1(n6793), .A2(P1_STATE_REG_SCAN_IN), .A3(n6583), .ZN(
        n6585) );
  INV_X1 U8232 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6584) );
  OAI22_X1 U8233 ( .A1(n6586), .A2(n6585), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6584), .ZN(n6587) );
  INV_X1 U8234 ( .A(n6587), .ZN(n6589) );
  NAND3_X1 U8235 ( .A1(n9736), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6749), .ZN(
        n6588) );
  OAI211_X1 U8236 ( .C1(n9759), .C2(n6590), .A(n6589), .B(n6588), .ZN(P1_U3241) );
  OAI222_X1 U8237 ( .A1(n9369), .A2(n6593), .B1(n9378), .B2(n6592), .C1(n6591), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  NAND2_X1 U8238 ( .A1(n8103), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6594) );
  OAI21_X1 U8239 ( .B1(n8103), .B2(n6595), .A(n6594), .ZN(P2_U3582) );
  INV_X1 U8240 ( .A(n6596), .ZN(n6602) );
  AOI22_X1 U8241 ( .A1(n8136), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8510), .ZN(n6597) );
  OAI21_X1 U8242 ( .B1(n6602), .B2(n8513), .A(n6597), .ZN(P2_U3347) );
  INV_X1 U8243 ( .A(n6598), .ZN(n6600) );
  INV_X1 U8244 ( .A(n6724), .ZN(n6719) );
  OAI222_X1 U8245 ( .A1(n9369), .A2(n6599), .B1(n9378), .B2(n6600), .C1(n6719), 
        .C2(n4309), .ZN(P1_U3343) );
  INV_X1 U8246 ( .A(n7189), .ZN(n7198) );
  OAI222_X1 U8247 ( .A1(n7947), .A2(n6601), .B1(n7198), .B2(P2_U3152), .C1(
        n8513), .C2(n6600), .ZN(P2_U3348) );
  INV_X1 U8248 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6603) );
  OAI222_X1 U8249 ( .A1(n9369), .A2(n6603), .B1(n9378), .B2(n6602), .C1(n6990), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  XOR2_X1 U8250 ( .A(n6605), .B(n6604), .Z(n6615) );
  NAND2_X1 U8251 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  NAND3_X1 U8252 ( .A1(n9736), .A2(n6609), .A3(n6608), .ZN(n6610) );
  NAND2_X1 U8253 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7251) );
  NAND2_X1 U8254 ( .A1(n6610), .A2(n7251), .ZN(n6611) );
  AOI21_X1 U8255 ( .B1(n6612), .B2(n9748), .A(n6611), .ZN(n6614) );
  INV_X1 U8256 ( .A(n9759), .ZN(n7002) );
  NAND2_X1 U8257 ( .A1(n7002), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6613) );
  OAI211_X1 U8258 ( .C1(n6615), .C2(n9715), .A(n6614), .B(n6613), .ZN(P1_U3249) );
  AOI21_X1 U8259 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n6629) );
  INV_X1 U8260 ( .A(n6619), .ZN(n6626) );
  AND2_X1 U8261 ( .A1(n4309), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7165) );
  INV_X1 U8262 ( .A(n6620), .ZN(n6622) );
  NAND3_X1 U8263 ( .A1(n6655), .A2(n6622), .A3(n6621), .ZN(n6623) );
  AOI21_X1 U8264 ( .B1(n6624), .B2(n6623), .A(n9756), .ZN(n6625) );
  AOI211_X1 U8265 ( .C1(n9748), .C2(n6626), .A(n7165), .B(n6625), .ZN(n6628)
         );
  INV_X1 U8266 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9398) );
  OR2_X1 U8267 ( .A1(n9759), .A2(n9398), .ZN(n6627) );
  OAI211_X1 U8268 ( .C1(n6629), .C2(n9715), .A(n6628), .B(n6627), .ZN(P1_U3248) );
  INV_X1 U8269 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6641) );
  XNOR2_X1 U8270 ( .A(n6631), .B(n6630), .ZN(n6639) );
  NAND2_X1 U8271 ( .A1(n4309), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U8272 ( .A1(n6633), .A2(n6632), .ZN(n6634) );
  NAND3_X1 U8273 ( .A1(n9736), .A2(n6635), .A3(n6634), .ZN(n6636) );
  OAI211_X1 U8274 ( .C1(n6994), .C2(n6637), .A(n7334), .B(n6636), .ZN(n6638)
         );
  AOI21_X1 U8275 ( .B1(n9746), .B2(n6639), .A(n6638), .ZN(n6640) );
  OAI21_X1 U8276 ( .B1(n9759), .B2(n6641), .A(n6640), .ZN(P1_U3246) );
  INV_X1 U8277 ( .A(n6642), .ZN(n6643) );
  OAI211_X1 U8278 ( .C1(n6645), .C2(n6644), .A(n9746), .B(n6643), .ZN(n6646)
         );
  OAI21_X1 U8279 ( .B1(n6994), .B2(n6647), .A(n6646), .ZN(n6653) );
  INV_X1 U8280 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6651) );
  OAI211_X1 U8281 ( .C1(n6649), .C2(n6648), .A(n9736), .B(n6779), .ZN(n6650)
         );
  OAI21_X1 U8282 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6651), .A(n6650), .ZN(n6652) );
  AOI211_X1 U8283 ( .C1(n7002), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6653), .B(
        n6652), .ZN(n6654) );
  INV_X1 U8284 ( .A(n6654), .ZN(P1_U3242) );
  INV_X1 U8285 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6666) );
  OAI21_X1 U8286 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(n6660) );
  AND2_X1 U8287 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7371) );
  NOR2_X1 U8288 ( .A1(n6994), .A2(n6658), .ZN(n6659) );
  AOI211_X1 U8289 ( .C1(n9736), .C2(n6660), .A(n7371), .B(n6659), .ZN(n6665)
         );
  OAI211_X1 U8290 ( .C1(n6663), .C2(n6662), .A(n9746), .B(n6661), .ZN(n6664)
         );
  OAI211_X1 U8291 ( .C1(n6666), .C2(n9759), .A(n6665), .B(n6664), .ZN(P1_U3247) );
  INV_X1 U8292 ( .A(n6667), .ZN(n6669) );
  INV_X1 U8293 ( .A(n8992), .ZN(n6993) );
  OAI222_X1 U8294 ( .A1(n9369), .A2(n6668), .B1(n9378), .B2(n6669), .C1(n4309), 
        .C2(n6993), .ZN(P1_U3341) );
  INV_X1 U8295 ( .A(n7352), .ZN(n7348) );
  OAI222_X1 U8296 ( .A1(n7947), .A2(n6670), .B1(n8513), .B2(n6669), .C1(
        P2_U3152), .C2(n7348), .ZN(P2_U3346) );
  NAND2_X1 U8297 ( .A1(n4309), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6953) );
  MUX2_X1 U8298 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6522), .S(n6676), .Z(n6672)
         );
  NAND3_X1 U8299 ( .A1(n6672), .A2(n6782), .A3(n6671), .ZN(n6673) );
  NAND3_X1 U8300 ( .A1(n9736), .A2(n6674), .A3(n6673), .ZN(n6675) );
  OAI211_X1 U8301 ( .C1(n6994), .C2(n6676), .A(n6953), .B(n6675), .ZN(n6681)
         );
  AOI211_X1 U8302 ( .C1(n6679), .C2(n6678), .A(n6677), .B(n9715), .ZN(n6680)
         );
  AOI211_X1 U8303 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n7002), .A(n6681), .B(
        n6680), .ZN(n6682) );
  INV_X1 U8304 ( .A(n6682), .ZN(P1_U3244) );
  NOR2_X1 U8305 ( .A1(n6688), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6684) );
  NOR2_X1 U8306 ( .A1(n6684), .A2(n6683), .ZN(n6686) );
  INV_X1 U8307 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9605) );
  AOI22_X1 U8308 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6719), .B1(n6724), .B2(
        n9605), .ZN(n6685) );
  NOR2_X1 U8309 ( .A1(n6686), .A2(n6685), .ZN(n6718) );
  AOI21_X1 U8310 ( .B1(n6686), .B2(n6685), .A(n6718), .ZN(n6695) );
  NAND2_X1 U8311 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7489) );
  OAI21_X1 U8312 ( .B1(n6994), .B2(n6719), .A(n7489), .ZN(n6693) );
  INV_X1 U8313 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6689) );
  MUX2_X1 U8314 ( .A(n6689), .B(P1_REG2_REG_10__SCAN_IN), .S(n6724), .Z(n6690)
         );
  AOI211_X1 U8315 ( .C1(n6691), .C2(n6690), .A(n6723), .B(n9715), .ZN(n6692)
         );
  AOI211_X1 U8316 ( .C1(n7002), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n6693), .B(
        n6692), .ZN(n6694) );
  OAI21_X1 U8317 ( .B1(n6695), .B2(n9756), .A(n6694), .ZN(P1_U3251) );
  NOR2_X1 U8318 ( .A1(n5622), .A2(P2_U3152), .ZN(n8507) );
  INV_X1 U8319 ( .A(n6696), .ZN(n7667) );
  AOI21_X1 U8320 ( .B1(n6697), .B2(n8507), .A(n7667), .ZN(n6698) );
  OAI21_X1 U8321 ( .B1(n9944), .B2(n6699), .A(n6698), .ZN(n6701) );
  NAND2_X1 U8322 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  NAND2_X1 U8323 ( .A1(n6702), .A2(n8103), .ZN(n6712) );
  NOR2_X1 U8324 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9911), .ZN(n6944) );
  INV_X1 U8325 ( .A(n6702), .ZN(n6704) );
  INV_X1 U8326 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8327 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6705), .S(n8109), .Z(n8111)
         );
  NAND3_X1 U8328 ( .A1(n8111), .A2(P2_REG1_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U8329 ( .A1(n8109), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8122) );
  INV_X1 U8330 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U8331 ( .A(n10016), .B(P2_REG1_REG_2__SCAN_IN), .S(n8120), .Z(n8124)
         );
  AOI21_X1 U8332 ( .B1(n8123), .B2(n8122), .A(n8124), .ZN(n8121) );
  AOI21_X1 U8333 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n8120), .A(n8121), .ZN(
        n6826) );
  INV_X1 U8334 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10018) );
  MUX2_X1 U8335 ( .A(n10018), .B(P2_REG1_REG_3__SCAN_IN), .S(n6824), .Z(n6825)
         );
  XNOR2_X1 U8336 ( .A(n6826), .B(n6825), .ZN(n6706) );
  NOR2_X1 U8337 ( .A1(n9868), .A2(n6706), .ZN(n6707) );
  AOI211_X1 U8338 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9866), .A(n6944), .B(
        n6707), .ZN(n6716) );
  NAND2_X1 U8339 ( .A1(n6824), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6708) );
  OAI21_X1 U8340 ( .B1(n6824), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6708), .ZN(
        n6709) );
  INV_X1 U8341 ( .A(n6709), .ZN(n6714) );
  INV_X1 U8342 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9937) );
  XOR2_X1 U8343 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8120), .Z(n8119) );
  INV_X1 U8344 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6710) );
  AND2_X1 U8345 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8106) );
  OAI21_X1 U8346 ( .B1(n6710), .B2(n5045), .A(n8105), .ZN(n8118) );
  NAND2_X1 U8347 ( .A1(n8119), .A2(n8118), .ZN(n8117) );
  OAI21_X1 U8348 ( .B1(n9937), .B2(n6711), .A(n8117), .ZN(n6713) );
  NAND2_X1 U8349 ( .A1(n6712), .A2(n8511), .ZN(n9869) );
  OAI211_X1 U8350 ( .C1(n6714), .C2(n6713), .A(n9865), .B(n6810), .ZN(n6715)
         );
  OAI211_X1 U8351 ( .C1(n9867), .C2(n6717), .A(n6716), .B(n6715), .ZN(P2_U3248) );
  AOI21_X1 U8352 ( .B1(n9605), .B2(n6719), .A(n6718), .ZN(n6721) );
  INV_X1 U8353 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9664) );
  AOI22_X1 U8354 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6990), .B1(n6996), .B2(
        n9664), .ZN(n6720) );
  NOR2_X1 U8355 ( .A1(n6721), .A2(n6720), .ZN(n6989) );
  AOI21_X1 U8356 ( .B1(n6721), .B2(n6720), .A(n6989), .ZN(n6731) );
  INV_X1 U8357 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U8358 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6996), .B1(n6990), .B2(
        n6722), .ZN(n6726) );
  OAI21_X1 U8359 ( .B1(n6726), .B2(n6725), .A(n6995), .ZN(n6729) );
  NAND2_X1 U8360 ( .A1(n7002), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U8361 ( .A1(n4309), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7686) );
  OAI211_X1 U8362 ( .C1(n6994), .C2(n6990), .A(n6727), .B(n7686), .ZN(n6728)
         );
  AOI21_X1 U8363 ( .B1(n6729), .B2(n9746), .A(n6728), .ZN(n6730) );
  OAI21_X1 U8364 ( .B1(n6731), .B2(n9756), .A(n6730), .ZN(P1_U3252) );
  INV_X1 U8365 ( .A(n6732), .ZN(n6735) );
  INV_X1 U8366 ( .A(n9369), .ZN(n9376) );
  AOI22_X1 U8367 ( .A1(n9674), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9376), .ZN(n6733) );
  OAI21_X1 U8368 ( .B1(n6735), .B2(n9378), .A(n6733), .ZN(P1_U3340) );
  INV_X1 U8369 ( .A(n7452), .ZN(n7447) );
  OAI222_X1 U8370 ( .A1(n8513), .A2(n6735), .B1(n7447), .B2(P2_U3152), .C1(
        n6734), .C2(n7947), .ZN(P2_U3345) );
  OAI21_X1 U8371 ( .B1(n6738), .B2(n6736), .A(n6737), .ZN(n6791) );
  AOI22_X1 U8372 ( .A1(n8626), .A2(n6791), .B1(n8611), .B2(n7270), .ZN(n6741)
         );
  NAND2_X1 U8373 ( .A1(n9621), .A2(n6739), .ZN(n7940) );
  AOI22_X1 U8374 ( .A1(n7940), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9608), .B2(
        n7041), .ZN(n6740) );
  NAND2_X1 U8375 ( .A1(n6741), .A2(n6740), .ZN(P1_U3230) );
  AND2_X1 U8376 ( .A1(n8781), .A2(n8947), .ZN(n7100) );
  AND2_X1 U8377 ( .A1(n6744), .A2(n7034), .ZN(n8915) );
  NOR2_X1 U8378 ( .A1(n7046), .A2(n8915), .ZN(n8799) );
  NAND2_X1 U8379 ( .A1(n8953), .A2(n7033), .ZN(n6746) );
  INV_X1 U8380 ( .A(n7041), .ZN(n7937) );
  OAI22_X1 U8381 ( .A1(n8799), .A2(n6746), .B1(n7937), .B2(n9250), .ZN(n7269)
         );
  INV_X1 U8382 ( .A(n7269), .ZN(n6747) );
  OAI21_X1 U8383 ( .B1(n7034), .B2(n7033), .A(n6747), .ZN(n6774) );
  NAND2_X1 U8384 ( .A1(n6774), .A2(n9802), .ZN(n6748) );
  OAI21_X1 U8385 ( .B1(n9802), .B2(n6749), .A(n6748), .ZN(P1_U3523) );
  NAND2_X1 U8386 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  XNOR2_X1 U8387 ( .A(n6753), .B(n6752), .ZN(n6758) );
  INV_X1 U8388 ( .A(n9608), .ZN(n8630) );
  INV_X1 U8389 ( .A(n6744), .ZN(n6754) );
  OAI22_X1 U8390 ( .A1(n8630), .A2(n7303), .B1(n6754), .B2(n9611), .ZN(n6756)
         );
  NOR2_X1 U8391 ( .A1(n8637), .A2(n7032), .ZN(n6755) );
  AOI211_X1 U8392 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7940), .A(n6756), .B(
        n6755), .ZN(n6757) );
  OAI21_X1 U8393 ( .B1(n6758), .B2(n9618), .A(n6757), .ZN(P1_U3220) );
  INV_X1 U8394 ( .A(n6759), .ZN(n6762) );
  INV_X1 U8395 ( .A(n7644), .ZN(n7648) );
  INV_X1 U8396 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6760) );
  OAI222_X1 U8397 ( .A1(n8513), .A2(n6762), .B1(n7648), .B2(P2_U3152), .C1(
        n6760), .C2(n7947), .ZN(P2_U3344) );
  INV_X1 U8398 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6761) );
  OAI222_X1 U8399 ( .A1(n4309), .A2(n9002), .B1(n9378), .B2(n6762), .C1(n6761), 
        .C2(n9369), .ZN(P1_U3339) );
  NAND2_X1 U8400 ( .A1(n6768), .A2(n6763), .ZN(n6765) );
  NAND2_X1 U8401 ( .A1(n6765), .A2(n6764), .ZN(n6770) );
  INV_X1 U8402 ( .A(n6766), .ZN(n6767) );
  NAND2_X1 U8403 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  NAND2_X1 U8404 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  INV_X2 U8405 ( .A(n9792), .ZN(n9794) );
  INV_X1 U8406 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8407 ( .A1(n6774), .A2(n9794), .ZN(n6775) );
  OAI21_X1 U8408 ( .B1(n9794), .B2(n6776), .A(n6775), .ZN(P1_U3454) );
  INV_X1 U8409 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9386) );
  INV_X1 U8410 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6784) );
  INV_X1 U8411 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7058) );
  MUX2_X1 U8412 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7058), .S(n6777), .Z(n6780)
         );
  NAND3_X1 U8413 ( .A1(n6780), .A2(n6779), .A3(n6778), .ZN(n6781) );
  NAND3_X1 U8414 ( .A1(n9736), .A2(n6782), .A3(n6781), .ZN(n6783) );
  OAI21_X1 U8415 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6784), .A(n6783), .ZN(n6789) );
  AOI211_X1 U8416 ( .C1(n6787), .C2(n6786), .A(n6785), .B(n9715), .ZN(n6788)
         );
  AOI211_X1 U8417 ( .C1(n9748), .C2(n6790), .A(n6789), .B(n6788), .ZN(n6795)
         );
  MUX2_X1 U8418 ( .A(n6792), .B(n6791), .S(n8951), .Z(n6794) );
  OAI211_X1 U8419 ( .C1(n6794), .C2(n6423), .A(P1_U4006), .B(n6793), .ZN(n6808) );
  OAI211_X1 U8420 ( .C1(n9386), .C2(n9759), .A(n6795), .B(n6808), .ZN(P1_U3243) );
  INV_X1 U8421 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6809) );
  OAI21_X1 U8422 ( .B1(n6798), .B2(n6797), .A(n6796), .ZN(n6806) );
  OAI21_X1 U8423 ( .B1(n6801), .B2(n6800), .A(n6799), .ZN(n6802) );
  AND2_X1 U8424 ( .A1(n4309), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7010) );
  AOI21_X1 U8425 ( .B1(n9736), .B2(n6802), .A(n7010), .ZN(n6803) );
  OAI21_X1 U8426 ( .B1(n6994), .B2(n6804), .A(n6803), .ZN(n6805) );
  AOI21_X1 U8427 ( .B1(n9746), .B2(n6806), .A(n6805), .ZN(n6807) );
  OAI211_X1 U8428 ( .C1(n9759), .C2(n6809), .A(n6808), .B(n6807), .ZN(P1_U3245) );
  INV_X1 U8429 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8430 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6811), .S(n6823), .Z(n6812)
         );
  INV_X1 U8431 ( .A(n6812), .ZN(n6880) );
  AOI21_X1 U8432 ( .B1(n6823), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6879), .ZN(
        n6894) );
  NAND2_X1 U8433 ( .A1(n6821), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6813) );
  OAI21_X1 U8434 ( .B1(n6821), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6813), .ZN(
        n6893) );
  NOR2_X1 U8435 ( .A1(n6894), .A2(n6893), .ZN(n6892) );
  AOI21_X1 U8436 ( .B1(n6821), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6892), .ZN(
        n6869) );
  INV_X1 U8437 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6814) );
  MUX2_X1 U8438 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6814), .S(n6820), .Z(n6815)
         );
  INV_X1 U8439 ( .A(n6815), .ZN(n6868) );
  NOR2_X1 U8440 ( .A1(n6869), .A2(n6868), .ZN(n6867) );
  AOI21_X1 U8441 ( .B1(n6820), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6867), .ZN(
        n6818) );
  NAND2_X1 U8442 ( .A1(n6843), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6816) );
  OAI21_X1 U8443 ( .B1(n6843), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6816), .ZN(
        n6817) );
  AOI211_X1 U8444 ( .C1(n6818), .C2(n6817), .A(n6838), .B(n7879), .ZN(n6837)
         );
  NOR2_X1 U8445 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5122), .ZN(n7127) );
  AOI21_X1 U8446 ( .B1(n9866), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7127), .ZN(
        n6834) );
  INV_X1 U8447 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8448 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6819), .S(n6843), .Z(n6832)
         );
  INV_X1 U8449 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6830) );
  MUX2_X1 U8450 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6830), .S(n6820), .Z(n6872)
         );
  NAND2_X1 U8451 ( .A1(n6821), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6829) );
  INV_X1 U8452 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6822) );
  MUX2_X1 U8453 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6822), .S(n6821), .Z(n6898)
         );
  INV_X1 U8454 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10020) );
  MUX2_X1 U8455 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10020), .S(n6823), .Z(n6885)
         );
  NAND2_X1 U8456 ( .A1(n6824), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6828) );
  OR2_X1 U8457 ( .A1(n6826), .A2(n6825), .ZN(n6827) );
  NAND2_X1 U8458 ( .A1(n6828), .A2(n6827), .ZN(n6886) );
  NAND2_X1 U8459 ( .A1(n6885), .A2(n6886), .ZN(n6884) );
  OAI21_X1 U8460 ( .B1(n6889), .B2(n10020), .A(n6884), .ZN(n6897) );
  NAND2_X1 U8461 ( .A1(n6898), .A2(n6897), .ZN(n6896) );
  NAND2_X1 U8462 ( .A1(n6829), .A2(n6896), .ZN(n6873) );
  NAND2_X1 U8463 ( .A1(n6872), .A2(n6873), .ZN(n6871) );
  OAI21_X1 U8464 ( .B1(n6876), .B2(n6830), .A(n6871), .ZN(n6831) );
  NAND2_X1 U8465 ( .A1(n6832), .A2(n6831), .ZN(n6844) );
  OAI211_X1 U8466 ( .C1(n6832), .C2(n6831), .A(n9864), .B(n6844), .ZN(n6833)
         );
  OAI211_X1 U8467 ( .C1(n9867), .C2(n6835), .A(n6834), .B(n6833), .ZN(n6836)
         );
  OR2_X1 U8468 ( .A1(n6837), .A2(n6836), .ZN(P2_U3252) );
  NAND2_X1 U8469 ( .A1(n6854), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6839) );
  OAI21_X1 U8470 ( .B1(n6854), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6839), .ZN(
        n6840) );
  AOI211_X1 U8471 ( .C1(n6841), .C2(n6840), .A(n6853), .B(n7879), .ZN(n6852)
         );
  NOR2_X1 U8472 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9471), .ZN(n6842) );
  AOI21_X1 U8473 ( .B1(n9866), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6842), .ZN(
        n6850) );
  NAND2_X1 U8474 ( .A1(n6843), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8475 ( .A1(n6845), .A2(n6844), .ZN(n6848) );
  INV_X1 U8476 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6846) );
  MUX2_X1 U8477 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6846), .S(n6854), .Z(n6847)
         );
  NAND2_X1 U8478 ( .A1(n6847), .A2(n6848), .ZN(n6858) );
  OAI211_X1 U8479 ( .C1(n6848), .C2(n6847), .A(n9864), .B(n6858), .ZN(n6849)
         );
  OAI211_X1 U8480 ( .C1(n9867), .C2(n6859), .A(n6850), .B(n6849), .ZN(n6851)
         );
  OR2_X1 U8481 ( .A1(n6852), .A2(n6851), .ZN(P2_U3253) );
  NAND2_X1 U8482 ( .A1(n6921), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6855) );
  OAI21_X1 U8483 ( .B1(n6921), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6855), .ZN(
        n6856) );
  NOR2_X1 U8484 ( .A1(n6857), .A2(n6856), .ZN(n6920) );
  AOI211_X1 U8485 ( .C1(n6857), .C2(n6856), .A(n6920), .B(n7879), .ZN(n6866)
         );
  NOR2_X1 U8486 ( .A1(n5150), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7411) );
  AOI21_X1 U8487 ( .B1(n9866), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7411), .ZN(
        n6864) );
  OAI21_X1 U8488 ( .B1(n6859), .B2(n6846), .A(n6858), .ZN(n6862) );
  INV_X1 U8489 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6860) );
  MUX2_X1 U8490 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6860), .S(n6921), .Z(n6861)
         );
  NAND2_X1 U8491 ( .A1(n6861), .A2(n6862), .ZN(n6926) );
  OAI211_X1 U8492 ( .C1(n6862), .C2(n6861), .A(n9864), .B(n6926), .ZN(n6863)
         );
  OAI211_X1 U8493 ( .C1(n9867), .C2(n6927), .A(n6864), .B(n6863), .ZN(n6865)
         );
  OR2_X1 U8494 ( .A1(n6866), .A2(n6865), .ZN(P2_U3254) );
  AOI211_X1 U8495 ( .C1(n6869), .C2(n6868), .A(n6867), .B(n7879), .ZN(n6878)
         );
  INV_X1 U8496 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9501) );
  NOR2_X1 U8497 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9501), .ZN(n6870) );
  AOI21_X1 U8498 ( .B1(n9866), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6870), .ZN(
        n6875) );
  OAI211_X1 U8499 ( .C1(n6873), .C2(n6872), .A(n9864), .B(n6871), .ZN(n6874)
         );
  OAI211_X1 U8500 ( .C1(n9867), .C2(n6876), .A(n6875), .B(n6874), .ZN(n6877)
         );
  OR2_X1 U8501 ( .A1(n6878), .A2(n6877), .ZN(P2_U3251) );
  AOI211_X1 U8502 ( .C1(n6881), .C2(n6880), .A(n6879), .B(n7879), .ZN(n6891)
         );
  INV_X1 U8503 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6882) );
  NOR2_X1 U8504 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6882), .ZN(n6883) );
  AOI21_X1 U8505 ( .B1(n9866), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6883), .ZN(
        n6888) );
  OAI211_X1 U8506 ( .C1(n6886), .C2(n6885), .A(n9864), .B(n6884), .ZN(n6887)
         );
  OAI211_X1 U8507 ( .C1(n9867), .C2(n6889), .A(n6888), .B(n6887), .ZN(n6890)
         );
  OR2_X1 U8508 ( .A1(n6891), .A2(n6890), .ZN(P2_U3249) );
  AOI211_X1 U8509 ( .C1(n6894), .C2(n6893), .A(n6892), .B(n7879), .ZN(n6903)
         );
  AND2_X1 U8510 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6895) );
  AOI21_X1 U8511 ( .B1(n9866), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6895), .ZN(
        n6900) );
  OAI211_X1 U8512 ( .C1(n6898), .C2(n6897), .A(n9864), .B(n6896), .ZN(n6899)
         );
  OAI211_X1 U8513 ( .C1(n9867), .C2(n6901), .A(n6900), .B(n6899), .ZN(n6902)
         );
  OR2_X1 U8514 ( .A1(n6903), .A2(n6902), .ZN(P2_U3250) );
  AND2_X1 U8515 ( .A1(n8036), .A2(n6904), .ZN(n9848) );
  INV_X1 U8516 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6913) );
  INV_X1 U8517 ( .A(n9844), .ZN(n9851) );
  NAND2_X1 U8518 ( .A1(n8104), .A2(n9832), .ZN(n6906) );
  NAND2_X1 U8519 ( .A1(n5637), .A2(n9834), .ZN(n6905) );
  NAND2_X1 U8520 ( .A1(n6906), .A2(n6905), .ZN(n6974) );
  AOI22_X1 U8521 ( .A1(n9851), .A2(n6974), .B1(n9859), .B2(n9958), .ZN(n6912)
         );
  OAI21_X1 U8522 ( .B1(n6909), .B2(n6908), .A(n6907), .ZN(n6910) );
  NAND2_X1 U8523 ( .A1(n9841), .A2(n6910), .ZN(n6911) );
  OAI211_X1 U8524 ( .C1(n9848), .C2(n6913), .A(n6912), .B(n6911), .ZN(P2_U3224) );
  INV_X1 U8525 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U8526 ( .A1(n9841), .A2(n9898), .ZN(n8064) );
  OAI22_X1 U8527 ( .A1(n6915), .A2(n8064), .B1(n9854), .B2(n6914), .ZN(n6917)
         );
  NAND2_X1 U8528 ( .A1(n6917), .A2(n6916), .ZN(n6919) );
  NOR2_X1 U8529 ( .A1(n6447), .A2(n8057), .ZN(n6980) );
  AOI22_X1 U8530 ( .A1(n9851), .A2(n6980), .B1(n9859), .B2(n9951), .ZN(n6918)
         );
  OAI211_X1 U8531 ( .C1(n9479), .C2(n9848), .A(n6919), .B(n6918), .ZN(P2_U3234) );
  NAND2_X1 U8532 ( .A1(n7189), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6922) );
  OAI21_X1 U8533 ( .B1(n7189), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6922), .ZN(
        n6923) );
  AOI211_X1 U8534 ( .C1(n6924), .C2(n6923), .A(n7188), .B(n7879), .ZN(n6934)
         );
  INV_X1 U8535 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U8536 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9542), .ZN(n6925) );
  AOI21_X1 U8537 ( .B1(n9866), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6925), .ZN(
        n6932) );
  OAI21_X1 U8538 ( .B1(n6927), .B2(n6860), .A(n6926), .ZN(n6930) );
  INV_X1 U8539 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6928) );
  MUX2_X1 U8540 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6928), .S(n7189), .Z(n6929)
         );
  NAND2_X1 U8541 ( .A1(n6929), .A2(n6930), .ZN(n7197) );
  OAI211_X1 U8542 ( .C1(n6930), .C2(n6929), .A(n9864), .B(n7197), .ZN(n6931)
         );
  OAI211_X1 U8543 ( .C1(n9867), .C2(n7198), .A(n6932), .B(n6931), .ZN(n6933)
         );
  OR2_X1 U8544 ( .A1(n6934), .A2(n6933), .ZN(P2_U3255) );
  NOR3_X1 U8545 ( .A1(n8064), .A2(n6936), .A3(n6935), .ZN(n6942) );
  INV_X1 U8546 ( .A(n6938), .ZN(n6939) );
  AOI21_X1 U8547 ( .B1(n6937), .B2(n6939), .A(n9854), .ZN(n6941) );
  OAI21_X1 U8548 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(n6946) );
  AOI22_X1 U8549 ( .A1(n9832), .A2(n5637), .B1(n8102), .B2(n9834), .ZN(n9906)
         );
  NOR2_X1 U8550 ( .A1(n9844), .A2(n9906), .ZN(n6943) );
  AOI211_X1 U8551 ( .C1(n9859), .C2(n4312), .A(n6944), .B(n6943), .ZN(n6945)
         );
  OAI211_X1 U8552 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9863), .A(n6946), .B(
        n6945), .ZN(P2_U3220) );
  OAI21_X1 U8553 ( .B1(n6947), .B2(n6950), .A(n6948), .ZN(n6951) );
  NAND2_X1 U8554 ( .A1(n6951), .A2(n8626), .ZN(n6958) );
  INV_X1 U8555 ( .A(n9611), .ZN(n8599) );
  INV_X1 U8556 ( .A(n6953), .ZN(n6954) );
  AOI21_X1 U8557 ( .B1(n8599), .B2(n8977), .A(n6954), .ZN(n6955) );
  OAI21_X1 U8558 ( .B1(n7302), .B2(n8630), .A(n6955), .ZN(n6956) );
  AOI21_X1 U8559 ( .B1(n8611), .B2(n6952), .A(n6956), .ZN(n6957) );
  OAI211_X1 U8560 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9625), .A(n6958), .B(
        n6957), .ZN(P1_U3216) );
  INV_X1 U8561 ( .A(n6959), .ZN(n6961) );
  INV_X1 U8562 ( .A(n7807), .ZN(n7815) );
  OAI222_X1 U8563 ( .A1(n7947), .A2(n6960), .B1(n8513), .B2(n6961), .C1(
        P2_U3152), .C2(n7815), .ZN(P2_U3343) );
  INV_X1 U8564 ( .A(n9708), .ZN(n9004) );
  OAI222_X1 U8565 ( .A1(n9369), .A2(n6962), .B1(n9378), .B2(n6961), .C1(
        P1_U3084), .C2(n9004), .ZN(P1_U3338) );
  XNOR2_X1 U8566 ( .A(n6446), .B(n6963), .ZN(n9961) );
  INV_X1 U8567 ( .A(n6964), .ZN(n6965) );
  AND2_X1 U8568 ( .A1(n6966), .A2(n6965), .ZN(n6967) );
  NAND2_X1 U8569 ( .A1(n6968), .A2(n6967), .ZN(n6971) );
  OR2_X1 U8570 ( .A1(n6970), .A2(n7343), .ZN(n7173) );
  NAND2_X1 U8571 ( .A1(n7602), .A2(n7173), .ZN(n9900) );
  AOI211_X1 U8572 ( .C1(n9951), .C2(n9958), .A(n10004), .B(n9924), .ZN(n9957)
         );
  INV_X1 U8573 ( .A(n6971), .ZN(n6985) );
  NAND2_X1 U8574 ( .A1(n6985), .A2(n7343), .ZN(n8192) );
  NOR2_X1 U8575 ( .A1(n6972), .A2(n5629), .ZN(n9896) );
  AOI22_X1 U8576 ( .A1(n9957), .A2(n9929), .B1(n9931), .B2(n9958), .ZN(n6979)
         );
  XNOR2_X1 U8577 ( .A(n6973), .B(n6446), .ZN(n6975) );
  AOI21_X1 U8578 ( .B1(n6975), .B2(n9922), .A(n6974), .ZN(n9959) );
  OAI21_X1 U8579 ( .B1(n6913), .B2(n9894), .A(n9959), .ZN(n6976) );
  MUX2_X1 U8580 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6976), .S(n9938), .Z(n6977)
         );
  INV_X1 U8581 ( .A(n6977), .ZN(n6978) );
  OAI211_X1 U8582 ( .C1(n9961), .C2(n8385), .A(n6979), .B(n6978), .ZN(P2_U3295) );
  INV_X1 U8583 ( .A(n9953), .ZN(n6988) );
  AOI21_X1 U8584 ( .B1(n9922), .B2(n9953), .A(n6980), .ZN(n9955) );
  OAI21_X1 U8585 ( .B1(n9894), .B2(n9479), .A(n9955), .ZN(n6983) );
  INV_X1 U8586 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6981) );
  NOR2_X1 U8587 ( .A1(n9938), .A2(n6981), .ZN(n6982) );
  AOI21_X1 U8588 ( .B1(n9938), .B2(n6983), .A(n6982), .ZN(n6987) );
  NAND2_X1 U8589 ( .A1(n6985), .A2(n6984), .ZN(n7531) );
  INV_X1 U8590 ( .A(n7531), .ZN(n7324) );
  OAI21_X1 U8591 ( .B1(n7324), .B2(n9931), .A(n9951), .ZN(n6986) );
  OAI211_X1 U8592 ( .C1(n6988), .C2(n8385), .A(n6987), .B(n6986), .ZN(P2_U3296) );
  AOI21_X1 U8593 ( .B1(n9664), .B2(n6990), .A(n6989), .ZN(n6992) );
  INV_X1 U8594 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U8595 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6993), .B1(n8992), .B2(
        n9659), .ZN(n6991) );
  NOR2_X1 U8596 ( .A1(n6992), .A2(n6991), .ZN(n8994) );
  AOI21_X1 U8597 ( .B1(n6992), .B2(n6991), .A(n8994), .ZN(n7004) );
  NAND2_X1 U8598 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9609) );
  OAI21_X1 U8599 ( .B1(n6994), .B2(n6993), .A(n9609), .ZN(n7001) );
  OAI21_X1 U8600 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6996), .A(n6995), .ZN(
        n6999) );
  NAND2_X1 U8601 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n8992), .ZN(n6997) );
  OAI21_X1 U8602 ( .B1(n8992), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6997), .ZN(
        n6998) );
  NOR2_X1 U8603 ( .A1(n6998), .A2(n6999), .ZN(n8979) );
  AOI211_X1 U8604 ( .C1(n6999), .C2(n6998), .A(n8979), .B(n9715), .ZN(n7000)
         );
  AOI211_X1 U8605 ( .C1(n7002), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7001), .B(
        n7000), .ZN(n7003) );
  OAI21_X1 U8606 ( .B1(n7004), .B2(n9756), .A(n7003), .ZN(P1_U3253) );
  INV_X1 U8607 ( .A(n7005), .ZN(n7007) );
  NAND2_X1 U8608 ( .A1(n7007), .A2(n7006), .ZN(n7008) );
  INV_X1 U8609 ( .A(n7369), .ZN(n8974) );
  NOR2_X1 U8610 ( .A1(n9611), .A2(n7938), .ZN(n7009) );
  AOI211_X1 U8611 ( .C1(n9608), .C2(n8974), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OAI21_X1 U8612 ( .B1(n7217), .B2(n8637), .A(n7011), .ZN(n7012) );
  AOI21_X1 U8613 ( .B1(n7291), .B2(n8634), .A(n7012), .ZN(n7013) );
  OAI21_X1 U8614 ( .B1(n7014), .B2(n9618), .A(n7013), .ZN(P1_U3228) );
  INV_X1 U8615 ( .A(n7015), .ZN(n9893) );
  OAI211_X1 U8616 ( .C1(n7018), .C2(n7017), .A(n7016), .B(n9841), .ZN(n7024)
         );
  NAND2_X1 U8617 ( .A1(n8102), .A2(n9832), .ZN(n7020) );
  NAND2_X1 U8618 ( .A1(n8100), .A2(n9834), .ZN(n7019) );
  AND2_X1 U8619 ( .A1(n7020), .A2(n7019), .ZN(n9892) );
  OAI22_X1 U8620 ( .A1(n9844), .A2(n9892), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7021), .ZN(n7022) );
  AOI21_X1 U8621 ( .B1(n9859), .B2(n4315), .A(n7022), .ZN(n7023) );
  OAI211_X1 U8622 ( .C1(n9863), .C2(n9893), .A(n7024), .B(n7023), .ZN(P2_U3229) );
  MUX2_X1 U8623 ( .A(n8956), .B(n7026), .S(n7025), .Z(n7786) );
  INV_X1 U8624 ( .A(n7100), .ZN(n7027) );
  NAND2_X1 U8625 ( .A1(n7029), .A2(n7028), .ZN(n7043) );
  OAI21_X1 U8626 ( .B1(n7028), .B2(n7029), .A(n7043), .ZN(n7104) );
  NAND2_X1 U8627 ( .A1(n8956), .A2(n9018), .ZN(n8787) );
  INV_X1 U8628 ( .A(n8947), .ZN(n8911) );
  NAND2_X1 U8629 ( .A1(n6385), .A2(n8911), .ZN(n8906) );
  XNOR2_X1 U8630 ( .A(n4408), .B(n7046), .ZN(n7031) );
  AOI222_X1 U8631 ( .A1(n9237), .A2(n7031), .B1(n8977), .B2(n9234), .C1(n6744), 
        .C2(n9232), .ZN(n7103) );
  NAND2_X1 U8632 ( .A1(n7032), .A2(n7034), .ZN(n7052) );
  OAI211_X1 U8633 ( .C1(n7034), .C2(n7032), .A(n9646), .B(n7052), .ZN(n7035)
         );
  INV_X1 U8634 ( .A(n7035), .ZN(n7106) );
  AOI21_X1 U8635 ( .B1(n9347), .B2(n7101), .A(n7106), .ZN(n7036) );
  OAI211_X1 U8636 ( .C1(n9653), .C2(n7104), .A(n7103), .B(n7036), .ZN(n7038)
         );
  NAND2_X1 U8637 ( .A1(n7038), .A2(n9802), .ZN(n7037) );
  OAI21_X1 U8638 ( .B1(n9802), .B2(n6519), .A(n7037), .ZN(P1_U3524) );
  INV_X1 U8639 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U8640 ( .A1(n7038), .A2(n9794), .ZN(n7039) );
  OAI21_X1 U8641 ( .B1(n9794), .B2(n7040), .A(n7039), .ZN(P1_U3457) );
  INV_X1 U8642 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7055) );
  INV_X1 U8643 ( .A(n7786), .ZN(n7543) );
  NAND2_X1 U8644 ( .A1(n7041), .A2(n7101), .ZN(n7042) );
  NAND2_X1 U8645 ( .A1(n7303), .A2(n5907), .ZN(n8919) );
  NAND2_X1 U8646 ( .A1(n8977), .A2(n7943), .ZN(n8920) );
  AND2_X1 U8647 ( .A1(n8919), .A2(n8920), .ZN(n8800) );
  NAND2_X1 U8648 ( .A1(n8919), .A2(n8920), .ZN(n7044) );
  OAI21_X1 U8649 ( .B1(n7045), .B2(n7044), .A(n7134), .ZN(n7051) );
  OAI22_X1 U8650 ( .A1(n7937), .A2(n9248), .B1(n7938), .B2(n9250), .ZN(n7050)
         );
  NAND2_X1 U8651 ( .A1(n7937), .A2(n7101), .ZN(n7047) );
  XNOR2_X1 U8652 ( .A(n8922), .B(n7044), .ZN(n7048) );
  NOR2_X1 U8653 ( .A1(n7048), .A2(n9246), .ZN(n7049) );
  AOI211_X1 U8654 ( .C1(n7543), .C2(n7051), .A(n7050), .B(n7049), .ZN(n7381)
         );
  AOI21_X1 U8655 ( .B1(n5907), .B2(n7052), .A(n7296), .ZN(n7379) );
  AOI22_X1 U8656 ( .A1(n7379), .A2(n9646), .B1(n9347), .B2(n5907), .ZN(n7053)
         );
  NAND2_X1 U8657 ( .A1(n7381), .A2(n7053), .ZN(n7056) );
  NAND2_X1 U8658 ( .A1(n7056), .A2(n9794), .ZN(n7054) );
  OAI21_X1 U8659 ( .B1(n9794), .B2(n7055), .A(n7054), .ZN(P1_U3460) );
  NAND2_X1 U8660 ( .A1(n7056), .A2(n9802), .ZN(n7057) );
  OAI21_X1 U8661 ( .B1(n9802), .B2(n7058), .A(n7057), .ZN(P1_U3525) );
  INV_X1 U8662 ( .A(n7059), .ZN(n7066) );
  AOI22_X1 U8663 ( .A1(n9720), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9376), .ZN(n7060) );
  OAI21_X1 U8664 ( .B1(n7066), .B2(n9378), .A(n7060), .ZN(P1_U3337) );
  INV_X1 U8665 ( .A(n7061), .ZN(n7065) );
  AOI22_X1 U8666 ( .A1(n9731), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9376), .ZN(n7062) );
  OAI21_X1 U8667 ( .B1(n7065), .B2(n9378), .A(n7062), .ZN(P1_U3336) );
  INV_X2 U8668 ( .A(P1_U4006), .ZN(n8978) );
  NAND2_X1 U8669 ( .A1(n8978), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7063) );
  OAI21_X1 U8670 ( .B1(n9049), .B2(n8978), .A(n7063), .ZN(P1_U3583) );
  INV_X1 U8671 ( .A(n8150), .ZN(n8145) );
  INV_X1 U8672 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7064) );
  OAI222_X1 U8673 ( .A1(n8513), .A2(n7065), .B1(n8145), .B2(P2_U3152), .C1(
        n7064), .C2(n7947), .ZN(P2_U3341) );
  OAI222_X1 U8674 ( .A1(n7947), .A2(n7067), .B1(n7885), .B2(P2_U3152), .C1(
        n8513), .C2(n7066), .ZN(P2_U3342) );
  XNOR2_X1 U8675 ( .A(n7068), .B(n7070), .ZN(n7259) );
  AOI211_X1 U8676 ( .C1(n7080), .C2(n7111), .A(n10004), .B(n7182), .ZN(n7260)
         );
  NAND2_X1 U8677 ( .A1(n7069), .A2(n9922), .ZN(n7076) );
  AOI21_X1 U8678 ( .B1(n7114), .B2(n7071), .A(n7070), .ZN(n7075) );
  NAND2_X1 U8679 ( .A1(n8100), .A2(n9832), .ZN(n7073) );
  NAND2_X1 U8680 ( .A1(n8097), .A2(n9834), .ZN(n7072) );
  NAND2_X1 U8681 ( .A1(n7073), .A2(n7072), .ZN(n7128) );
  INV_X1 U8682 ( .A(n7128), .ZN(n7074) );
  OAI21_X1 U8683 ( .B1(n7076), .B2(n7075), .A(n7074), .ZN(n7266) );
  AOI211_X1 U8684 ( .C1(n7259), .C2(n10008), .A(n7260), .B(n7266), .ZN(n7082)
         );
  INV_X1 U8685 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7077) );
  OAI22_X1 U8686 ( .A1(n8494), .A2(n7264), .B1(n10012), .B2(n7077), .ZN(n7078)
         );
  INV_X1 U8687 ( .A(n7078), .ZN(n7079) );
  OAI21_X1 U8688 ( .B1(n7082), .B2(n10010), .A(n7079), .ZN(P2_U3472) );
  AOI22_X1 U8689 ( .A1(n6492), .A2(n7080), .B1(n10024), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7081) );
  OAI21_X1 U8690 ( .B1(n7082), .B2(n10024), .A(n7081), .ZN(P2_U3527) );
  XNOR2_X1 U8691 ( .A(n7084), .B(n7083), .ZN(n9983) );
  AND2_X1 U8692 ( .A1(n9912), .A2(n9811), .ZN(n7085) );
  OR2_X1 U8693 ( .A1(n7085), .A2(n9886), .ZN(n9980) );
  NAND2_X1 U8694 ( .A1(n9931), .A2(n9811), .ZN(n7088) );
  NAND2_X1 U8695 ( .A1(n9928), .A2(n7086), .ZN(n7087) );
  OAI211_X1 U8696 ( .C1(n7531), .C2(n9980), .A(n7088), .B(n7087), .ZN(n7094)
         );
  INV_X1 U8697 ( .A(n7089), .ZN(n7091) );
  OAI211_X1 U8698 ( .C1(n7091), .C2(n7090), .A(n4345), .B(n9922), .ZN(n7092)
         );
  AOI22_X1 U8699 ( .A1(n9832), .A2(n9835), .B1(n8101), .B2(n9834), .ZN(n9806)
         );
  NAND2_X1 U8700 ( .A1(n7092), .A2(n9806), .ZN(n9981) );
  MUX2_X1 U8701 ( .A(n9981), .B(P2_REG2_REG_4__SCAN_IN), .S(n9942), .Z(n7093)
         );
  AOI211_X1 U8702 ( .C1(n9934), .C2(n9983), .A(n7094), .B(n7093), .ZN(n7095)
         );
  INV_X1 U8703 ( .A(n7095), .ZN(P2_U3292) );
  NAND2_X1 U8704 ( .A1(n7097), .A2(n7096), .ZN(n7397) );
  AND2_X1 U8705 ( .A1(n7098), .A2(n6386), .ZN(n7099) );
  AOI22_X1 U8706 ( .A1(n9255), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7224), .B2(
        n7101), .ZN(n7102) );
  OAI211_X1 U8707 ( .C1(n7786), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7105)
         );
  NAND2_X1 U8708 ( .A1(n7105), .A2(n9263), .ZN(n7108) );
  NAND2_X1 U8709 ( .A1(n9203), .A2(n7106), .ZN(n7107) );
  OAI211_X1 U8710 ( .C1(n7109), .C2(n9263), .A(n7108), .B(n7107), .ZN(P1_U3290) );
  XOR2_X1 U8711 ( .A(n7110), .B(n7117), .Z(n7156) );
  AOI21_X1 U8712 ( .B1(n9884), .B2(n9858), .A(n10004), .ZN(n7112) );
  AND2_X1 U8713 ( .A1(n7112), .A2(n7111), .ZN(n7150) );
  NAND2_X1 U8714 ( .A1(n9891), .A2(n7113), .ZN(n7116) );
  INV_X1 U8715 ( .A(n7114), .ZN(n7115) );
  AOI21_X1 U8716 ( .B1(n7117), .B2(n7116), .A(n7115), .ZN(n7118) );
  AOI22_X1 U8717 ( .A1(n9832), .A2(n8101), .B1(n8099), .B2(n9834), .ZN(n9849)
         );
  OAI21_X1 U8718 ( .B1(n7118), .B2(n9907), .A(n9849), .ZN(n7153) );
  AOI211_X1 U8719 ( .C1(n7156), .C2(n10008), .A(n7150), .B(n7153), .ZN(n7123)
         );
  AOI22_X1 U8720 ( .A1(n6492), .A2(n9858), .B1(n10024), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7119) );
  OAI21_X1 U8721 ( .B1(n7123), .B2(n10024), .A(n7119), .ZN(P2_U3526) );
  INV_X1 U8722 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7120) );
  OAI22_X1 U8723 ( .A1(n8494), .A2(n7152), .B1(n10012), .B2(n7120), .ZN(n7121)
         );
  INV_X1 U8724 ( .A(n7121), .ZN(n7122) );
  OAI21_X1 U8725 ( .B1(n7123), .B2(n10010), .A(n7122), .ZN(P2_U3469) );
  INV_X1 U8726 ( .A(n7261), .ZN(n7131) );
  OAI211_X1 U8727 ( .C1(n4398), .C2(n7125), .A(n7230), .B(n9841), .ZN(n7130)
         );
  NOR2_X1 U8728 ( .A1(n5795), .A2(n7264), .ZN(n7126) );
  AOI211_X1 U8729 ( .C1(n9851), .C2(n7128), .A(n7127), .B(n7126), .ZN(n7129)
         );
  OAI211_X1 U8730 ( .C1(n9863), .C2(n7131), .A(n7130), .B(n7129), .ZN(P2_U3215) );
  INV_X1 U8731 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7145) );
  INV_X1 U8732 ( .A(n7298), .ZN(n7132) );
  OAI21_X1 U8733 ( .B1(n7132), .B2(n7217), .A(n7208), .ZN(n7295) );
  NAND2_X1 U8734 ( .A1(n7303), .A2(n7943), .ZN(n7133) );
  NAND2_X1 U8735 ( .A1(n7134), .A2(n7133), .ZN(n7301) );
  INV_X1 U8736 ( .A(n7938), .ZN(n8976) );
  NAND2_X1 U8737 ( .A1(n8976), .A2(n9761), .ZN(n8848) );
  NAND2_X1 U8738 ( .A1(n7938), .A2(n6952), .ZN(n8924) );
  NAND2_X1 U8739 ( .A1(n7301), .A2(n8798), .ZN(n7300) );
  NAND2_X1 U8740 ( .A1(n7938), .A2(n9761), .ZN(n7135) );
  NAND2_X1 U8741 ( .A1(n7300), .A2(n7135), .ZN(n7136) );
  NAND2_X1 U8742 ( .A1(n7302), .A2(n7292), .ZN(n8663) );
  INV_X1 U8743 ( .A(n7302), .ZN(n8975) );
  NAND2_X1 U8744 ( .A1(n8975), .A2(n7217), .ZN(n8854) );
  OAI21_X1 U8745 ( .B1(n7136), .B2(n8797), .A(n7219), .ZN(n7142) );
  OAI22_X1 U8746 ( .A1(n7938), .A2(n9248), .B1(n7369), .B2(n9250), .ZN(n7141)
         );
  NAND2_X1 U8747 ( .A1(n7137), .A2(n8919), .ZN(n7299) );
  INV_X1 U8748 ( .A(n8798), .ZN(n7138) );
  XNOR2_X1 U8749 ( .A(n8665), .B(n8797), .ZN(n7139) );
  NOR2_X1 U8750 ( .A1(n7139), .A2(n9246), .ZN(n7140) );
  AOI211_X1 U8751 ( .C1(n7543), .C2(n7142), .A(n7141), .B(n7140), .ZN(n7290)
         );
  NAND2_X1 U8752 ( .A1(n9347), .A2(n7292), .ZN(n7143) );
  OAI211_X1 U8753 ( .C1(n9786), .C2(n7295), .A(n7290), .B(n7143), .ZN(n7146)
         );
  NAND2_X1 U8754 ( .A1(n7146), .A2(n9794), .ZN(n7144) );
  OAI21_X1 U8755 ( .B1(n9794), .B2(n7145), .A(n7144), .ZN(P1_U3466) );
  NAND2_X1 U8756 ( .A1(n7146), .A2(n9802), .ZN(n7147) );
  OAI21_X1 U8757 ( .B1(n9802), .B2(n7148), .A(n7147), .ZN(P1_U3527) );
  AOI22_X1 U8758 ( .A1(n9929), .A2(n7150), .B1(n7149), .B2(n9928), .ZN(n7151)
         );
  OAI21_X1 U8759 ( .B1(n7152), .B2(n8374), .A(n7151), .ZN(n7155) );
  MUX2_X1 U8760 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7153), .S(n9938), .Z(n7154)
         );
  AOI211_X1 U8761 ( .C1(n7156), .C2(n9934), .A(n7155), .B(n7154), .ZN(n7157)
         );
  INV_X1 U8762 ( .A(n7157), .ZN(P2_U3290) );
  NAND2_X1 U8763 ( .A1(n7159), .A2(n7158), .ZN(n7163) );
  XNOR2_X1 U8764 ( .A(n7161), .B(n7160), .ZN(n7162) );
  XNOR2_X1 U8765 ( .A(n7163), .B(n7162), .ZN(n7169) );
  NOR2_X1 U8766 ( .A1(n9611), .A2(n7392), .ZN(n7164) );
  AOI211_X1 U8767 ( .C1(n9608), .C2(n8971), .A(n7165), .B(n7164), .ZN(n7166)
         );
  OAI21_X1 U8768 ( .B1(n9780), .B2(n8637), .A(n7166), .ZN(n7167) );
  AOI21_X1 U8769 ( .B1(n7398), .B2(n8634), .A(n7167), .ZN(n7168) );
  OAI21_X1 U8770 ( .B1(n7169), .B2(n9618), .A(n7168), .ZN(P1_U3211) );
  NAND2_X1 U8771 ( .A1(n7171), .A2(n7178), .ZN(n7172) );
  NAND2_X1 U8772 ( .A1(n4758), .A2(n7172), .ZN(n9994) );
  INV_X1 U8773 ( .A(n7173), .ZN(n7174) );
  NAND2_X1 U8774 ( .A1(n9938), .A2(n7174), .ZN(n7320) );
  NAND2_X1 U8775 ( .A1(n8099), .A2(n9832), .ZN(n7176) );
  NAND2_X1 U8776 ( .A1(n8096), .A2(n9834), .ZN(n7175) );
  AND2_X1 U8777 ( .A1(n7176), .A2(n7175), .ZN(n7237) );
  OAI21_X1 U8778 ( .B1(n4844), .B2(n7178), .A(n7177), .ZN(n7179) );
  NAND2_X1 U8779 ( .A1(n7179), .A2(n9922), .ZN(n7180) );
  OAI211_X1 U8780 ( .C1(n9994), .C2(n7602), .A(n7237), .B(n7180), .ZN(n9997)
         );
  NAND2_X1 U8781 ( .A1(n9997), .A2(n9938), .ZN(n7187) );
  INV_X1 U8782 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7181) );
  OAI22_X1 U8783 ( .A1(n9938), .A2(n7181), .B1(n7236), .B2(n9894), .ZN(n7185)
         );
  NOR2_X1 U8784 ( .A1(n7182), .A2(n9995), .ZN(n7183) );
  OR2_X1 U8785 ( .A1(n7321), .A2(n7183), .ZN(n9996) );
  NOR2_X1 U8786 ( .A1(n9996), .A2(n7531), .ZN(n7184) );
  AOI211_X1 U8787 ( .C1(n9931), .C2(n7240), .A(n7185), .B(n7184), .ZN(n7186)
         );
  OAI211_X1 U8788 ( .C1(n9994), .C2(n7320), .A(n7187), .B(n7186), .ZN(P2_U3288) );
  INV_X1 U8789 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7190) );
  MUX2_X1 U8790 ( .A(n7190), .B(P2_REG2_REG_11__SCAN_IN), .S(n8136), .Z(n7191)
         );
  INV_X1 U8791 ( .A(n7191), .ZN(n8133) );
  OAI21_X1 U8792 ( .B1(n8136), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8131), .ZN(
        n7194) );
  NAND2_X1 U8793 ( .A1(n7352), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7192) );
  OAI21_X1 U8794 ( .B1(n7352), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7192), .ZN(
        n7193) );
  NOR2_X1 U8795 ( .A1(n7193), .A2(n7194), .ZN(n7351) );
  AOI211_X1 U8796 ( .C1(n7194), .C2(n7193), .A(n7351), .B(n7879), .ZN(n7207)
         );
  INV_X1 U8797 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7195) );
  MUX2_X1 U8798 ( .A(n7195), .B(P2_REG1_REG_12__SCAN_IN), .S(n7352), .Z(n7201)
         );
  INV_X1 U8799 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8800 ( .A1(n8136), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7199) );
  MUX2_X1 U8801 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7196), .S(n8136), .Z(n8138)
         );
  OAI21_X1 U8802 ( .B1(n7198), .B2(n6928), .A(n7197), .ZN(n8139) );
  NAND2_X1 U8803 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
  NAND2_X1 U8804 ( .A1(n7199), .A2(n8137), .ZN(n7200) );
  NOR2_X1 U8805 ( .A1(n7200), .A2(n7201), .ZN(n7347) );
  AOI21_X1 U8806 ( .B1(n7201), .B2(n7200), .A(n7347), .ZN(n7205) );
  NAND2_X1 U8807 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7659) );
  INV_X1 U8808 ( .A(n7659), .ZN(n7202) );
  AOI21_X1 U8809 ( .B1(n9866), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7202), .ZN(
        n7204) );
  NAND2_X1 U8810 ( .A1(n8169), .A2(n7352), .ZN(n7203) );
  OAI211_X1 U8811 ( .C1(n9868), .C2(n7205), .A(n7204), .B(n7203), .ZN(n7206)
         );
  OR2_X1 U8812 ( .A1(n7207), .A2(n7206), .ZN(P2_U3257) );
  AOI21_X1 U8813 ( .B1(n7208), .B2(n7338), .A(n9786), .ZN(n7209) );
  NAND2_X1 U8814 ( .A1(n7209), .A2(n7274), .ZN(n9767) );
  INV_X1 U8815 ( .A(n9767), .ZN(n7216) );
  INV_X1 U8816 ( .A(n7210), .ZN(n7341) );
  OR2_X1 U8817 ( .A1(n7392), .A2(n9250), .ZN(n9766) );
  OAI21_X1 U8818 ( .B1(n9145), .B2(n7341), .A(n9766), .ZN(n7215) );
  INV_X1 U8819 ( .A(n8663), .ZN(n7211) );
  NAND2_X1 U8820 ( .A1(n7369), .A2(n7338), .ZN(n8664) );
  NAND2_X1 U8821 ( .A1(n8974), .A2(n9768), .ZN(n8853) );
  INV_X1 U8822 ( .A(n8801), .ZN(n7279) );
  XNOR2_X1 U8823 ( .A(n7382), .B(n7279), .ZN(n7212) );
  NAND2_X1 U8824 ( .A1(n7212), .A2(n9237), .ZN(n7214) );
  OR2_X1 U8825 ( .A1(n7302), .A2(n9248), .ZN(n7213) );
  NAND2_X1 U8826 ( .A1(n7214), .A2(n7213), .ZN(n9770) );
  AOI211_X1 U8827 ( .C1(n7216), .C2(n9168), .A(n7215), .B(n9770), .ZN(n7227)
         );
  NAND2_X1 U8828 ( .A1(n7302), .A2(n7217), .ZN(n7218) );
  INV_X1 U8829 ( .A(n7278), .ZN(n7220) );
  AOI21_X1 U8830 ( .B1(n8801), .B2(n7221), .A(n7220), .ZN(n9771) );
  AND2_X1 U8831 ( .A1(n8953), .A2(n7222), .ZN(n7223) );
  INV_X1 U8832 ( .A(n9265), .ZN(n9173) );
  OAI22_X1 U8833 ( .A1(n9260), .A2(n9768), .B1(n6512), .B2(n9263), .ZN(n7225)
         );
  AOI21_X1 U8834 ( .B1(n9771), .B2(n9173), .A(n7225), .ZN(n7226) );
  OAI21_X1 U8835 ( .B1(n7227), .B2(n9205), .A(n7226), .ZN(P1_U3286) );
  INV_X1 U8836 ( .A(n7228), .ZN(n7229) );
  AOI21_X1 U8837 ( .B1(n7230), .B2(n7229), .A(n9854), .ZN(n7235) );
  NOR3_X1 U8838 ( .A1(n8064), .A2(n7232), .A3(n7231), .ZN(n7234) );
  OAI21_X1 U8839 ( .B1(n7235), .B2(n7234), .A(n7233), .ZN(n7242) );
  NOR2_X1 U8840 ( .A1(n9863), .A2(n7236), .ZN(n7239) );
  OAI22_X1 U8841 ( .A1(n9844), .A2(n7237), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9471), .ZN(n7238) );
  AOI211_X1 U8842 ( .C1(n9859), .C2(n7240), .A(n7239), .B(n7238), .ZN(n7241)
         );
  NAND2_X1 U8843 ( .A1(n7242), .A2(n7241), .ZN(P2_U3223) );
  INV_X1 U8844 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7244) );
  INV_X1 U8845 ( .A(n7243), .ZN(n7245) );
  INV_X1 U8846 ( .A(n9747), .ZN(n9010) );
  OAI222_X1 U8847 ( .A1(n9369), .A2(n7244), .B1(n9378), .B2(n7245), .C1(n4309), 
        .C2(n9010), .ZN(P1_U3335) );
  INV_X1 U8848 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7246) );
  INV_X1 U8849 ( .A(n8151), .ZN(n8165) );
  OAI222_X1 U8850 ( .A1(n7947), .A2(n7246), .B1(n8513), .B2(n7245), .C1(
        P2_U3152), .C2(n8165), .ZN(P2_U3340) );
  XOR2_X1 U8851 ( .A(n7248), .B(n7247), .Z(n7249) );
  XNOR2_X1 U8852 ( .A(n7250), .B(n7249), .ZN(n7258) );
  INV_X1 U8853 ( .A(n7581), .ZN(n7255) );
  INV_X1 U8854 ( .A(n7251), .ZN(n7252) );
  AOI21_X1 U8855 ( .B1(n8599), .B2(n8972), .A(n7252), .ZN(n7254) );
  NAND2_X1 U8856 ( .A1(n9608), .A2(n8970), .ZN(n7253) );
  OAI211_X1 U8857 ( .C1(n9625), .C2(n7255), .A(n7254), .B(n7253), .ZN(n7256)
         );
  AOI21_X1 U8858 ( .B1(n8611), .B2(n7559), .A(n7256), .ZN(n7257) );
  OAI21_X1 U8859 ( .B1(n7258), .B2(n9618), .A(n7257), .ZN(P1_U3219) );
  INV_X1 U8860 ( .A(n7259), .ZN(n7268) );
  NAND2_X1 U8861 ( .A1(n7260), .A2(n9929), .ZN(n7263) );
  AOI22_X1 U8862 ( .A1(n9942), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7261), .B2(
        n9928), .ZN(n7262) );
  OAI211_X1 U8863 ( .C1(n7264), .C2(n8374), .A(n7263), .B(n7262), .ZN(n7265)
         );
  AOI21_X1 U8864 ( .B1(n9938), .B2(n7266), .A(n7265), .ZN(n7267) );
  OAI21_X1 U8865 ( .B1(n8385), .B2(n7268), .A(n7267), .ZN(P2_U3289) );
  INV_X1 U8866 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7273) );
  AOI22_X1 U8867 ( .A1(n7269), .A2(n9263), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9255), .ZN(n7272) );
  INV_X1 U8868 ( .A(n9260), .ZN(n9174) );
  OAI21_X1 U8869 ( .B1(n9240), .B2(n9174), .A(n7270), .ZN(n7271) );
  OAI211_X1 U8870 ( .C1(n9263), .C2(n7273), .A(n7272), .B(n7271), .ZN(P1_U3291) );
  INV_X1 U8871 ( .A(n9240), .ZN(n7792) );
  INV_X1 U8872 ( .A(n7396), .ZN(n7276) );
  NAND2_X1 U8873 ( .A1(n7274), .A2(n7287), .ZN(n7275) );
  NAND2_X1 U8874 ( .A1(n7276), .A2(n7275), .ZN(n9774) );
  NAND2_X1 U8875 ( .A1(n8974), .A2(n7338), .ZN(n7277) );
  NAND2_X1 U8876 ( .A1(n7278), .A2(n7277), .ZN(n7394) );
  NAND2_X1 U8877 ( .A1(n7392), .A2(n7287), .ZN(n8850) );
  INV_X1 U8878 ( .A(n7392), .ZN(n8973) );
  NAND2_X1 U8879 ( .A1(n8973), .A2(n9773), .ZN(n8659) );
  INV_X1 U8880 ( .A(n8803), .ZN(n8660) );
  XNOR2_X1 U8881 ( .A(n7394), .B(n8660), .ZN(n7284) );
  OR2_X1 U8882 ( .A1(n7382), .A2(n7279), .ZN(n7280) );
  NAND2_X1 U8883 ( .A1(n7280), .A2(n8664), .ZN(n8661) );
  XNOR2_X1 U8884 ( .A(n8661), .B(n8803), .ZN(n7282) );
  OAI22_X1 U8885 ( .A1(n7369), .A2(n9248), .B1(n7504), .B2(n9250), .ZN(n7281)
         );
  AOI21_X1 U8886 ( .B1(n7282), .B2(n9237), .A(n7281), .ZN(n7283) );
  OAI21_X1 U8887 ( .B1(n7284), .B2(n7786), .A(n7283), .ZN(n9775) );
  NAND2_X1 U8888 ( .A1(n9775), .A2(n9263), .ZN(n7289) );
  OAI22_X1 U8889 ( .A1(n9263), .A2(n6513), .B1(n7285), .B2(n9145), .ZN(n7286)
         );
  AOI21_X1 U8890 ( .B1(n9174), .B2(n7287), .A(n7286), .ZN(n7288) );
  OAI211_X1 U8891 ( .C1(n7792), .C2(n9774), .A(n7289), .B(n7288), .ZN(P1_U3285) );
  MUX2_X1 U8892 ( .A(n6509), .B(n7290), .S(n9263), .Z(n7294) );
  AOI22_X1 U8893 ( .A1(n9174), .A2(n7292), .B1(n7291), .B2(n9255), .ZN(n7293)
         );
  OAI211_X1 U8894 ( .C1(n7792), .C2(n7295), .A(n7294), .B(n7293), .ZN(P1_U3287) );
  OR2_X1 U8895 ( .A1(n7296), .A2(n9761), .ZN(n7297) );
  NAND2_X1 U8896 ( .A1(n7298), .A2(n7297), .ZN(n9762) );
  XNOR2_X1 U8897 ( .A(n7299), .B(n8798), .ZN(n7307) );
  OAI21_X1 U8898 ( .B1(n7301), .B2(n8798), .A(n7300), .ZN(n7305) );
  OAI22_X1 U8899 ( .A1(n7303), .A2(n9248), .B1(n7302), .B2(n9250), .ZN(n7304)
         );
  AOI21_X1 U8900 ( .B1(n7305), .B2(n7543), .A(n7304), .ZN(n7306) );
  OAI21_X1 U8901 ( .B1(n9246), .B2(n7307), .A(n7306), .ZN(n9763) );
  NAND2_X1 U8902 ( .A1(n9763), .A2(n9263), .ZN(n7311) );
  OAI22_X1 U8903 ( .A1(n9263), .A2(n7308), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9145), .ZN(n7309) );
  AOI21_X1 U8904 ( .B1(n9174), .B2(n6952), .A(n7309), .ZN(n7310) );
  OAI211_X1 U8905 ( .C1(n7792), .C2(n9762), .A(n7311), .B(n7310), .ZN(P1_U3288) );
  OAI21_X1 U8906 ( .B1(n7313), .B2(n7316), .A(n7312), .ZN(n7474) );
  INV_X1 U8907 ( .A(n7602), .ZN(n9910) );
  NAND2_X1 U8908 ( .A1(n8097), .A2(n9832), .ZN(n7315) );
  NAND2_X1 U8909 ( .A1(n8095), .A2(n9834), .ZN(n7314) );
  NAND2_X1 U8910 ( .A1(n7315), .A2(n7314), .ZN(n7408) );
  XNOR2_X1 U8911 ( .A(n7317), .B(n7316), .ZN(n7318) );
  NOR2_X1 U8912 ( .A1(n7318), .A2(n9907), .ZN(n7319) );
  AOI211_X1 U8913 ( .C1(n7474), .C2(n9910), .A(n7408), .B(n7319), .ZN(n7478)
         );
  INV_X1 U8914 ( .A(n7320), .ZN(n9914) );
  INV_X1 U8915 ( .A(n7321), .ZN(n7323) );
  INV_X1 U8916 ( .A(n7595), .ZN(n7322) );
  AOI21_X1 U8917 ( .B1(n7475), .B2(n7323), .A(n7322), .ZN(n7476) );
  NAND2_X1 U8918 ( .A1(n7476), .A2(n7324), .ZN(n7326) );
  AOI22_X1 U8919 ( .A1(n9942), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7409), .B2(
        n9928), .ZN(n7325) );
  OAI211_X1 U8920 ( .C1(n7327), .C2(n8374), .A(n7326), .B(n7325), .ZN(n7328)
         );
  AOI21_X1 U8921 ( .B1(n7474), .B2(n9914), .A(n7328), .ZN(n7329) );
  OAI21_X1 U8922 ( .B1(n7478), .B2(n9942), .A(n7329), .ZN(P2_U3287) );
  XOR2_X1 U8923 ( .A(n7363), .B(n7364), .Z(n7332) );
  INV_X1 U8924 ( .A(n7330), .ZN(n7331) );
  NAND2_X1 U8925 ( .A1(n7332), .A2(n7331), .ZN(n7362) );
  OAI21_X1 U8926 ( .B1(n7332), .B2(n7331), .A(n7362), .ZN(n7333) );
  NAND2_X1 U8927 ( .A1(n7333), .A2(n8626), .ZN(n7340) );
  INV_X1 U8928 ( .A(n7334), .ZN(n7335) );
  AOI21_X1 U8929 ( .B1(n8599), .B2(n8975), .A(n7335), .ZN(n7336) );
  OAI21_X1 U8930 ( .B1(n7392), .B2(n8630), .A(n7336), .ZN(n7337) );
  AOI21_X1 U8931 ( .B1(n8611), .B2(n7338), .A(n7337), .ZN(n7339) );
  OAI211_X1 U8932 ( .C1(n9625), .C2(n7341), .A(n7340), .B(n7339), .ZN(P1_U3225) );
  INV_X1 U8933 ( .A(n7342), .ZN(n7345) );
  OAI222_X1 U8934 ( .A1(n7947), .A2(n7344), .B1(n8513), .B2(n7345), .C1(n7343), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8935 ( .A1(n9369), .A2(n7346), .B1(n9378), .B2(n7345), .C1(
        P1_U3084), .C2(n9168), .ZN(P1_U3334) );
  AOI21_X1 U8936 ( .B1(n7348), .B2(n7195), .A(n7347), .ZN(n7350) );
  INV_X1 U8937 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7727) );
  AOI22_X1 U8938 ( .A1(n7452), .A2(n7727), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7447), .ZN(n7349) );
  NOR2_X1 U8939 ( .A1(n7350), .A2(n7349), .ZN(n7446) );
  AOI21_X1 U8940 ( .B1(n7350), .B2(n7349), .A(n7446), .ZN(n7361) );
  NOR2_X1 U8941 ( .A1(n7452), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7353) );
  AOI21_X1 U8942 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7452), .A(n7353), .ZN(
        n7354) );
  OAI21_X1 U8943 ( .B1(n7355), .B2(n7354), .A(n7451), .ZN(n7356) );
  NAND2_X1 U8944 ( .A1(n7356), .A2(n9865), .ZN(n7360) );
  INV_X1 U8945 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8946 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7703) );
  OAI21_X1 U8947 ( .B1(n8174), .B2(n7357), .A(n7703), .ZN(n7358) );
  AOI21_X1 U8948 ( .B1(n7452), .B2(n8169), .A(n7358), .ZN(n7359) );
  OAI211_X1 U8949 ( .C1(n7361), .C2(n9868), .A(n7360), .B(n7359), .ZN(P2_U3258) );
  OAI21_X1 U8950 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(n7368) );
  NAND2_X1 U8951 ( .A1(n7366), .A2(n7365), .ZN(n7367) );
  XNOR2_X1 U8952 ( .A(n7368), .B(n7367), .ZN(n7376) );
  NOR2_X1 U8953 ( .A1(n9611), .A2(n7369), .ZN(n7370) );
  AOI211_X1 U8954 ( .C1(n9608), .C2(n8972), .A(n7371), .B(n7370), .ZN(n7372)
         );
  OAI21_X1 U8955 ( .B1(n9773), .B2(n8637), .A(n7372), .ZN(n7373) );
  AOI21_X1 U8956 ( .B1(n7374), .B2(n8634), .A(n7373), .ZN(n7375) );
  OAI21_X1 U8957 ( .B1(n7376), .B2(n9618), .A(n7375), .ZN(P1_U3237) );
  AOI22_X1 U8958 ( .A1(n9257), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9255), .ZN(n7377) );
  OAI21_X1 U8959 ( .B1(n7943), .B2(n9260), .A(n7377), .ZN(n7378) );
  AOI21_X1 U8960 ( .B1(n9240), .B2(n7379), .A(n7378), .ZN(n7380) );
  OAI21_X1 U8961 ( .B1(n7381), .B2(n9205), .A(n7380), .ZN(P1_U3289) );
  AND2_X1 U8962 ( .A1(n8850), .A2(n8664), .ZN(n8855) );
  NAND2_X1 U8963 ( .A1(n7382), .A2(n8855), .ZN(n7384) );
  NAND2_X1 U8964 ( .A1(n8853), .A2(n8659), .ZN(n7383) );
  NAND2_X1 U8965 ( .A1(n8850), .A2(n7383), .ZN(n8927) );
  NAND2_X1 U8966 ( .A1(n7384), .A2(n8927), .ZN(n7388) );
  NAND2_X1 U8967 ( .A1(n7504), .A2(n7385), .ZN(n8839) );
  NAND2_X1 U8968 ( .A1(n8972), .A2(n9780), .ZN(n8928) );
  NAND2_X1 U8969 ( .A1(n8839), .A2(n8928), .ZN(n8805) );
  INV_X1 U8970 ( .A(n8805), .ZN(n7386) );
  NAND2_X1 U8971 ( .A1(n7388), .A2(n8805), .ZN(n7389) );
  NAND2_X1 U8972 ( .A1(n4406), .A2(n7389), .ZN(n7391) );
  OAI22_X1 U8973 ( .A1(n7392), .A2(n9248), .B1(n7510), .B2(n9250), .ZN(n7390)
         );
  AOI21_X1 U8974 ( .B1(n7391), .B2(n9237), .A(n7390), .ZN(n9779) );
  NAND2_X1 U8975 ( .A1(n7392), .A2(n9773), .ZN(n7393) );
  OAI21_X1 U8976 ( .B1(n7395), .B2(n8805), .A(n7506), .ZN(n9782) );
  NAND2_X1 U8977 ( .A1(n9782), .A2(n9173), .ZN(n7403) );
  NAND2_X1 U8978 ( .A1(n7396), .A2(n9780), .ZN(n7558) );
  OAI211_X1 U8979 ( .C1(n7396), .C2(n9780), .A(n7558), .B(n9646), .ZN(n9778)
         );
  INV_X1 U8980 ( .A(n9778), .ZN(n7401) );
  NOR2_X1 U8981 ( .A1(n7397), .A2(n9018), .ZN(n9254) );
  AOI22_X1 U8982 ( .A1(n9257), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7398), .B2(
        n9255), .ZN(n7399) );
  OAI21_X1 U8983 ( .B1(n9780), .B2(n9260), .A(n7399), .ZN(n7400) );
  AOI21_X1 U8984 ( .B1(n7401), .B2(n9254), .A(n7400), .ZN(n7402) );
  OAI211_X1 U8985 ( .C1(n9257), .C2(n9779), .A(n7403), .B(n7402), .ZN(P1_U3284) );
  INV_X1 U8986 ( .A(n7233), .ZN(n7407) );
  NOR3_X1 U8987 ( .A1(n8064), .A2(n7405), .A3(n7404), .ZN(n7406) );
  AOI21_X1 U8988 ( .B1(n7407), .B2(n9841), .A(n7406), .ZN(n7420) );
  INV_X1 U8989 ( .A(n7408), .ZN(n7414) );
  INV_X1 U8990 ( .A(n7409), .ZN(n7410) );
  OR2_X1 U8991 ( .A1(n9863), .A2(n7410), .ZN(n7413) );
  INV_X1 U8992 ( .A(n7411), .ZN(n7412) );
  OAI211_X1 U8993 ( .C1(n9844), .C2(n7414), .A(n7413), .B(n7412), .ZN(n7417)
         );
  NOR2_X1 U8994 ( .A1(n7415), .A2(n9854), .ZN(n7416) );
  AOI211_X1 U8995 ( .C1(n9859), .C2(n7475), .A(n7417), .B(n7416), .ZN(n7418)
         );
  OAI21_X1 U8996 ( .B1(n7420), .B2(n7419), .A(n7418), .ZN(P2_U3233) );
  INV_X1 U8997 ( .A(n9877), .ZN(n7430) );
  AOI21_X1 U8998 ( .B1(n7422), .B2(n7421), .A(n9854), .ZN(n7424) );
  NAND2_X1 U8999 ( .A1(n7424), .A2(n7423), .ZN(n7429) );
  NAND2_X1 U9000 ( .A1(n8096), .A2(n9832), .ZN(n7426) );
  NAND2_X1 U9001 ( .A1(n8094), .A2(n9834), .ZN(n7425) );
  AND2_X1 U9002 ( .A1(n7426), .A2(n7425), .ZN(n7601) );
  OAI22_X1 U9003 ( .A1(n9844), .A2(n7601), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9542), .ZN(n7427) );
  AOI21_X1 U9004 ( .B1(n9876), .B2(n8046), .A(n7427), .ZN(n7428) );
  OAI211_X1 U9005 ( .C1(n7430), .C2(n5795), .A(n7429), .B(n7428), .ZN(P2_U3219) );
  INV_X1 U9006 ( .A(n7431), .ZN(n7444) );
  OAI222_X1 U9007 ( .A1(n8513), .A2(n7444), .B1(P2_U3152), .B2(n5629), .C1(
        n7432), .C2(n7947), .ZN(P2_U3338) );
  XNOR2_X1 U9008 ( .A(n7433), .B(n4750), .ZN(n7498) );
  INV_X1 U9009 ( .A(n7498), .ZN(n7443) );
  XNOR2_X1 U9010 ( .A(n7434), .B(n4750), .ZN(n7437) );
  NAND2_X1 U9011 ( .A1(n8095), .A2(n9832), .ZN(n7436) );
  NAND2_X1 U9012 ( .A1(n8093), .A2(n9834), .ZN(n7435) );
  AND2_X1 U9013 ( .A1(n7436), .A2(n7435), .ZN(n9817) );
  OAI21_X1 U9014 ( .B1(n7437), .B2(n9907), .A(n9817), .ZN(n7496) );
  AOI211_X1 U9015 ( .C1(n9827), .C2(n7596), .A(n10004), .B(n7528), .ZN(n7497)
         );
  NAND2_X1 U9016 ( .A1(n7497), .A2(n9929), .ZN(n7440) );
  AOI22_X1 U9017 ( .A1(n9942), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7438), .B2(
        n9928), .ZN(n7439) );
  OAI211_X1 U9018 ( .C1(n4480), .C2(n8374), .A(n7440), .B(n7439), .ZN(n7441)
         );
  AOI21_X1 U9019 ( .B1(n7496), .B2(n9938), .A(n7441), .ZN(n7442) );
  OAI21_X1 U9020 ( .B1(n7443), .B2(n8385), .A(n7442), .ZN(P2_U3285) );
  OAI222_X1 U9021 ( .A1(n9369), .A2(n7445), .B1(n9378), .B2(n7444), .C1(n8947), 
        .C2(n4309), .ZN(P1_U3333) );
  AOI21_X1 U9022 ( .B1(n7447), .B2(n7727), .A(n7446), .ZN(n7449) );
  INV_X1 U9023 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7804) );
  AOI22_X1 U9024 ( .A1(n7644), .A2(n7804), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7648), .ZN(n7448) );
  NOR2_X1 U9025 ( .A1(n7449), .A2(n7448), .ZN(n7647) );
  AOI21_X1 U9026 ( .B1(n7449), .B2(n7448), .A(n7647), .ZN(n7460) );
  INV_X1 U9027 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7450) );
  AOI22_X1 U9028 ( .A1(n7644), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7450), .B2(
        n7648), .ZN(n7454) );
  OAI21_X1 U9029 ( .B1(n7454), .B2(n7453), .A(n7643), .ZN(n7455) );
  NAND2_X1 U9030 ( .A1(n7455), .A2(n9865), .ZN(n7459) );
  INV_X1 U9031 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9032 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9632) );
  OAI21_X1 U9033 ( .B1(n8174), .B2(n7456), .A(n9632), .ZN(n7457) );
  AOI21_X1 U9034 ( .B1(n7644), .B2(n8169), .A(n7457), .ZN(n7458) );
  OAI211_X1 U9035 ( .C1(n7460), .C2(n9868), .A(n7459), .B(n7458), .ZN(P2_U3259) );
  INV_X1 U9036 ( .A(n7461), .ZN(n7948) );
  INV_X1 U9037 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7462) );
  OAI222_X1 U9038 ( .A1(n8513), .A2(n7948), .B1(P2_U3152), .B2(n7463), .C1(
        n7462), .C2(n7947), .ZN(P2_U3337) );
  INV_X1 U9039 ( .A(n7465), .ZN(n7466) );
  AOI21_X1 U9040 ( .B1(n7467), .B2(n7464), .A(n7466), .ZN(n7473) );
  NAND2_X1 U9041 ( .A1(n8634), .A2(n7513), .ZN(n7470) );
  AOI21_X1 U9042 ( .B1(n8599), .B2(n8971), .A(n7468), .ZN(n7469) );
  OAI211_X1 U9043 ( .C1(n7618), .C2(n8630), .A(n7470), .B(n7469), .ZN(n7471)
         );
  AOI21_X1 U9044 ( .B1(n8611), .B2(n7535), .A(n7471), .ZN(n7472) );
  OAI21_X1 U9045 ( .B1(n7473), .B2(n9618), .A(n7472), .ZN(P1_U3229) );
  INV_X1 U9046 ( .A(n7474), .ZN(n7479) );
  AOI22_X1 U9047 ( .A1(n7476), .A2(n9926), .B1(n9987), .B2(n7475), .ZN(n7477)
         );
  OAI211_X1 U9048 ( .C1(n7479), .C2(n7594), .A(n7478), .B(n7477), .ZN(n7481)
         );
  NAND2_X1 U9049 ( .A1(n7481), .A2(n10026), .ZN(n7480) );
  OAI21_X1 U9050 ( .B1(n10026), .B2(n6860), .A(n7480), .ZN(P2_U3529) );
  INV_X1 U9051 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9052 ( .A1(n7481), .A2(n10012), .ZN(n7482) );
  OAI21_X1 U9053 ( .B1(n10012), .B2(n7483), .A(n7482), .ZN(P2_U3478) );
  NAND2_X1 U9054 ( .A1(n7485), .A2(n7484), .ZN(n7486) );
  XNOR2_X1 U9055 ( .A(n7487), .B(n7486), .ZN(n7495) );
  INV_X1 U9056 ( .A(n7488), .ZN(n7545) );
  INV_X1 U9057 ( .A(n7489), .ZN(n7490) );
  AOI21_X1 U9058 ( .B1(n8599), .B2(n8970), .A(n7490), .ZN(n7492) );
  INV_X1 U9059 ( .A(n9612), .ZN(n8968) );
  NAND2_X1 U9060 ( .A1(n8968), .A2(n9608), .ZN(n7491) );
  OAI211_X1 U9061 ( .C1(n9625), .C2(n7545), .A(n7492), .B(n7491), .ZN(n7493)
         );
  AOI21_X1 U9062 ( .B1(n8611), .B2(n7613), .A(n7493), .ZN(n7494) );
  OAI21_X1 U9063 ( .B1(n7495), .B2(n9618), .A(n7494), .ZN(P1_U3215) );
  AOI211_X1 U9064 ( .C1(n7498), .C2(n10008), .A(n7497), .B(n7496), .ZN(n7503)
         );
  INV_X1 U9065 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7499) );
  NOR2_X1 U9066 ( .A1(n10012), .A2(n7499), .ZN(n7500) );
  AOI21_X1 U9067 ( .B1(n6500), .B2(n9827), .A(n7500), .ZN(n7501) );
  OAI21_X1 U9068 ( .B1(n7503), .B2(n10010), .A(n7501), .ZN(P2_U3484) );
  AOI22_X1 U9069 ( .A1(n6492), .A2(n9827), .B1(n10024), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n7502) );
  OAI21_X1 U9070 ( .B1(n7503), .B2(n10024), .A(n7502), .ZN(P2_U3531) );
  NAND2_X1 U9071 ( .A1(n7504), .A2(n9780), .ZN(n7505) );
  NAND2_X1 U9072 ( .A1(n7510), .A2(n7559), .ZN(n8679) );
  INV_X1 U9073 ( .A(n7535), .ZN(n9785) );
  NAND2_X1 U9074 ( .A1(n9785), .A2(n8970), .ZN(n8680) );
  INV_X1 U9075 ( .A(n8970), .ZN(n7507) );
  NAND2_X1 U9076 ( .A1(n7507), .A2(n7535), .ZN(n8671) );
  XNOR2_X1 U9077 ( .A(n7537), .B(n8808), .ZN(n9791) );
  INV_X1 U9078 ( .A(n9791), .ZN(n7518) );
  NAND2_X1 U9079 ( .A1(n9263), .A2(n7543), .ZN(n7590) );
  XNOR2_X1 U9080 ( .A(n7617), .B(n8808), .ZN(n7509) );
  OAI222_X1 U9081 ( .A1(n9250), .A2(n7618), .B1(n9248), .B2(n7510), .C1(n9246), 
        .C2(n7509), .ZN(n9788) );
  INV_X1 U9082 ( .A(n7511), .ZN(n7557) );
  INV_X1 U9083 ( .A(n7546), .ZN(n7512) );
  OAI21_X1 U9084 ( .B1(n9785), .B2(n7557), .A(n7512), .ZN(n9787) );
  AOI22_X1 U9085 ( .A1(n9205), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7513), .B2(
        n9255), .ZN(n7515) );
  NAND2_X1 U9086 ( .A1(n9174), .A2(n7535), .ZN(n7514) );
  OAI211_X1 U9087 ( .C1(n9787), .C2(n7792), .A(n7515), .B(n7514), .ZN(n7516)
         );
  AOI21_X1 U9088 ( .B1(n9788), .B2(n9263), .A(n7516), .ZN(n7517) );
  OAI21_X1 U9089 ( .B1(n7518), .B2(n7590), .A(n7517), .ZN(P1_U3282) );
  XNOR2_X1 U9090 ( .A(n7519), .B(n7522), .ZN(n10009) );
  INV_X1 U9091 ( .A(n10009), .ZN(n7534) );
  NAND2_X1 U9092 ( .A1(n7521), .A2(n7520), .ZN(n7523) );
  XNOR2_X1 U9093 ( .A(n7523), .B(n7522), .ZN(n7526) );
  NAND2_X1 U9094 ( .A1(n8094), .A2(n9832), .ZN(n7525) );
  NAND2_X1 U9095 ( .A1(n8092), .A2(n9834), .ZN(n7524) );
  AND2_X1 U9096 ( .A1(n7525), .A2(n7524), .ZN(n7661) );
  OAI21_X1 U9097 ( .B1(n7526), .B2(n9907), .A(n7661), .ZN(n10006) );
  INV_X1 U9098 ( .A(n7574), .ZN(n7527) );
  OAI21_X1 U9099 ( .B1(n10003), .B2(n7528), .A(n7527), .ZN(n10005) );
  AOI22_X1 U9100 ( .A1(n9942), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7658), .B2(
        n9928), .ZN(n7530) );
  NAND2_X1 U9101 ( .A1(n9931), .A2(n7663), .ZN(n7529) );
  OAI211_X1 U9102 ( .C1(n10005), .C2(n7531), .A(n7530), .B(n7529), .ZN(n7532)
         );
  AOI21_X1 U9103 ( .B1(n10006), .B2(n9938), .A(n7532), .ZN(n7533) );
  OAI21_X1 U9104 ( .B1(n7534), .B2(n8385), .A(n7533), .ZN(P2_U3284) );
  AND2_X1 U9105 ( .A1(n7535), .A2(n8970), .ZN(n7536) );
  OR2_X1 U9106 ( .A1(n7613), .A2(n7618), .ZN(n8676) );
  NAND2_X1 U9107 ( .A1(n7613), .A2(n7618), .ZN(n8672) );
  NAND2_X1 U9108 ( .A1(n8676), .A2(n8672), .ZN(n8807) );
  XNOR2_X1 U9109 ( .A(n7614), .B(n8807), .ZN(n7544) );
  INV_X1 U9110 ( .A(n8680), .ZN(n7538) );
  OAI21_X1 U9111 ( .B1(n7617), .B2(n7538), .A(n8671), .ZN(n7539) );
  XNOR2_X1 U9112 ( .A(n7539), .B(n8807), .ZN(n7541) );
  AOI22_X1 U9113 ( .A1(n8968), .A2(n9234), .B1(n9232), .B2(n8970), .ZN(n7540)
         );
  OAI21_X1 U9114 ( .B1(n7541), .B2(n9246), .A(n7540), .ZN(n7542) );
  AOI21_X1 U9115 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n9603) );
  OAI22_X1 U9116 ( .A1(n9263), .A2(n6689), .B1(n7545), .B2(n9145), .ZN(n7550)
         );
  INV_X1 U9117 ( .A(n7613), .ZN(n9600) );
  OAI21_X1 U9118 ( .B1(n7546), .B2(n9600), .A(n9646), .ZN(n7547) );
  OR2_X1 U9119 ( .A1(n7611), .A2(n7547), .ZN(n9599) );
  INV_X1 U9120 ( .A(n9254), .ZN(n7548) );
  NOR2_X1 U9121 ( .A1(n9599), .A2(n7548), .ZN(n7549) );
  AOI211_X1 U9122 ( .C1(n9174), .C2(n7613), .A(n7550), .B(n7549), .ZN(n7551)
         );
  OAI21_X1 U9123 ( .B1(n9603), .B2(n9205), .A(n7551), .ZN(P1_U3281) );
  INV_X1 U9124 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7562) );
  OAI21_X1 U9125 ( .B1(n7552), .B2(n7554), .A(n7553), .ZN(n7589) );
  XNOR2_X1 U9126 ( .A(n7555), .B(n8809), .ZN(n7556) );
  AOI222_X1 U9127 ( .A1(n9237), .A2(n7556), .B1(n8970), .B2(n9234), .C1(n8972), 
        .C2(n9232), .ZN(n7584) );
  AOI21_X1 U9128 ( .B1(n7559), .B2(n7558), .A(n7557), .ZN(n7587) );
  AOI22_X1 U9129 ( .A1(n7587), .A2(n9646), .B1(n9347), .B2(n7559), .ZN(n7560)
         );
  OAI211_X1 U9130 ( .C1(n7589), .C2(n9653), .A(n7584), .B(n7560), .ZN(n7563)
         );
  NAND2_X1 U9131 ( .A1(n7563), .A2(n9794), .ZN(n7561) );
  OAI21_X1 U9132 ( .B1(n9794), .B2(n7562), .A(n7561), .ZN(P1_U3478) );
  NAND2_X1 U9133 ( .A1(n7563), .A2(n9802), .ZN(n7564) );
  OAI21_X1 U9134 ( .B1(n9802), .B2(n7565), .A(n7564), .ZN(P1_U3531) );
  NAND2_X1 U9135 ( .A1(n7566), .A2(n7570), .ZN(n7567) );
  NAND2_X1 U9136 ( .A1(n7568), .A2(n7567), .ZN(n7722) );
  XNOR2_X1 U9137 ( .A(n7569), .B(n7570), .ZN(n7573) );
  NAND2_X1 U9138 ( .A1(n8091), .A2(n9834), .ZN(n7572) );
  NAND2_X1 U9139 ( .A1(n8093), .A2(n9832), .ZN(n7571) );
  NAND2_X1 U9140 ( .A1(n7572), .A2(n7571), .ZN(n7702) );
  AOI21_X1 U9141 ( .B1(n7573), .B2(n9922), .A(n7702), .ZN(n7724) );
  INV_X1 U9142 ( .A(n7724), .ZN(n7579) );
  OAI211_X1 U9143 ( .C1(n7574), .C2(n7732), .A(n9926), .B(n4395), .ZN(n7723)
         );
  AOI22_X1 U9144 ( .A1(n9942), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7706), .B2(
        n9928), .ZN(n7577) );
  NAND2_X1 U9145 ( .A1(n7575), .A2(n9931), .ZN(n7576) );
  OAI211_X1 U9146 ( .C1(n7723), .C2(n8192), .A(n7577), .B(n7576), .ZN(n7578)
         );
  AOI21_X1 U9147 ( .B1(n7579), .B2(n9938), .A(n7578), .ZN(n7580) );
  OAI21_X1 U9148 ( .B1(n7722), .B2(n8385), .A(n7580), .ZN(P2_U3283) );
  AOI22_X1 U9149 ( .A1(n9205), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7581), .B2(
        n9255), .ZN(n7582) );
  OAI21_X1 U9150 ( .B1(n7583), .B2(n9260), .A(n7582), .ZN(n7586) );
  NOR2_X1 U9151 ( .A1(n7584), .A2(n9257), .ZN(n7585) );
  AOI211_X1 U9152 ( .C1(n7587), .C2(n9240), .A(n7586), .B(n7585), .ZN(n7588)
         );
  OAI21_X1 U9153 ( .B1(n7590), .B2(n7589), .A(n7588), .ZN(P1_U3283) );
  OAI21_X1 U9154 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(n7603) );
  INV_X1 U9155 ( .A(n7603), .ZN(n9879) );
  INV_X1 U9156 ( .A(n7594), .ZN(n10000) );
  AOI21_X1 U9157 ( .B1(n7595), .B2(n9877), .A(n10004), .ZN(n7597) );
  AND2_X1 U9158 ( .A1(n7597), .A2(n7596), .ZN(n9878) );
  OAI211_X1 U9159 ( .C1(n7599), .C2(n4747), .A(n7598), .B(n9922), .ZN(n7600)
         );
  OAI211_X1 U9160 ( .C1(n7603), .C2(n7602), .A(n7601), .B(n7600), .ZN(n9875)
         );
  AOI211_X1 U9161 ( .C1(n9879), .C2(n10000), .A(n9878), .B(n9875), .ZN(n7608)
         );
  INV_X1 U9162 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7604) );
  NOR2_X1 U9163 ( .A1(n10012), .A2(n7604), .ZN(n7605) );
  AOI21_X1 U9164 ( .B1(n6500), .B2(n9877), .A(n7605), .ZN(n7606) );
  OAI21_X1 U9165 ( .B1(n7608), .B2(n10010), .A(n7606), .ZN(P2_U3481) );
  AOI22_X1 U9166 ( .A1(n6492), .A2(n9877), .B1(n10024), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7607) );
  OAI21_X1 U9167 ( .B1(n7608), .B2(n10024), .A(n7607), .ZN(P2_U3530) );
  INV_X1 U9168 ( .A(n7609), .ZN(n7945) );
  OAI222_X1 U9169 ( .A1(n9369), .A2(n7610), .B1(n9378), .B2(n7945), .C1(n4309), 
        .C2(n5878), .ZN(P1_U3331) );
  INV_X1 U9170 ( .A(n7697), .ZN(n9660) );
  OR2_X1 U9171 ( .A1(n7611), .A2(n9660), .ZN(n7612) );
  NAND2_X1 U9172 ( .A1(n7636), .A2(n7612), .ZN(n9661) );
  INV_X1 U9173 ( .A(n7618), .ZN(n8969) );
  OR2_X1 U9174 ( .A1(n7697), .A2(n9612), .ZN(n8687) );
  NAND2_X1 U9175 ( .A1(n7697), .A2(n9612), .ZN(n8841) );
  INV_X1 U9176 ( .A(n8813), .ZN(n7615) );
  OAI21_X1 U9177 ( .B1(n7616), .B2(n7615), .A(n7628), .ZN(n7622) );
  NAND2_X1 U9178 ( .A1(n8676), .A2(n8680), .ZN(n8875) );
  NAND2_X1 U9179 ( .A1(n8672), .A2(n8671), .ZN(n8683) );
  NAND2_X1 U9180 ( .A1(n8683), .A2(n8676), .ZN(n8840) );
  XNOR2_X1 U9181 ( .A(n7632), .B(n8813), .ZN(n7620) );
  OAI22_X1 U9182 ( .A1(n7618), .A2(n9248), .B1(n7782), .B2(n9250), .ZN(n7619)
         );
  AOI21_X1 U9183 ( .B1(n7620), .B2(n9237), .A(n7619), .ZN(n7621) );
  OAI21_X1 U9184 ( .B1(n7622), .B2(n7786), .A(n7621), .ZN(n9662) );
  NAND2_X1 U9185 ( .A1(n9662), .A2(n9263), .ZN(n7626) );
  INV_X1 U9186 ( .A(n7623), .ZN(n7690) );
  OAI22_X1 U9187 ( .A1(n9263), .A2(n6722), .B1(n7690), .B2(n9145), .ZN(n7624)
         );
  AOI21_X1 U9188 ( .B1(n9174), .B2(n7697), .A(n7624), .ZN(n7625) );
  OAI211_X1 U9189 ( .C1(n7792), .C2(n9661), .A(n7626), .B(n7625), .ZN(P1_U3280) );
  NAND2_X1 U9190 ( .A1(n7697), .A2(n8968), .ZN(n7627) );
  OR2_X1 U9191 ( .A1(n7637), .A2(n7782), .ZN(n8691) );
  NAND2_X1 U9192 ( .A1(n7637), .A2(n7782), .ZN(n8842) );
  NAND2_X1 U9193 ( .A1(n8691), .A2(n8842), .ZN(n7633) );
  OR2_X1 U9194 ( .A1(n7629), .A2(n7633), .ZN(n7630) );
  NAND2_X1 U9195 ( .A1(n7755), .A2(n7630), .ZN(n9654) );
  INV_X1 U9196 ( .A(n8841), .ZN(n7631) );
  INV_X1 U9197 ( .A(n7633), .ZN(n8814) );
  XNOR2_X1 U9198 ( .A(n7758), .B(n8814), .ZN(n7634) );
  OAI222_X1 U9199 ( .A1(n9248), .A2(n9612), .B1(n9250), .B2(n8699), .C1(n9246), 
        .C2(n7634), .ZN(n9656) );
  INV_X1 U9200 ( .A(n7637), .ZN(n9614) );
  INV_X1 U9201 ( .A(n7776), .ZN(n7635) );
  AOI211_X1 U9202 ( .C1(n7637), .C2(n7636), .A(n9786), .B(n7635), .ZN(n9657)
         );
  NAND2_X1 U9203 ( .A1(n9657), .A2(n9254), .ZN(n7640) );
  AOI22_X1 U9204 ( .A1(n9257), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7638), .B2(
        n9255), .ZN(n7639) );
  OAI211_X1 U9205 ( .C1(n9614), .C2(n9260), .A(n7640), .B(n7639), .ZN(n7641)
         );
  AOI21_X1 U9206 ( .B1(n9656), .B2(n9263), .A(n7641), .ZN(n7642) );
  OAI21_X1 U9207 ( .B1(n9654), .B2(n9265), .A(n7642), .ZN(P1_U3279) );
  OAI21_X1 U9208 ( .B1(n7644), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7643), .ZN(
        n7814) );
  XNOR2_X1 U9209 ( .A(n7814), .B(n7807), .ZN(n7646) );
  INV_X1 U9210 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U9211 ( .A1(n7646), .A2(n7645), .ZN(n7816) );
  OAI21_X1 U9212 ( .B1(n7646), .B2(n7645), .A(n7816), .ZN(n7654) );
  AOI21_X1 U9213 ( .B1(n7648), .B2(n7804), .A(n7647), .ZN(n7806) );
  XNOR2_X1 U9214 ( .A(n7806), .B(n7815), .ZN(n7649) );
  NAND2_X1 U9215 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7649), .ZN(n7808) );
  OAI211_X1 U9216 ( .C1(n7649), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9864), .B(
        n7808), .ZN(n7652) );
  AND2_X1 U9217 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7650) );
  AOI21_X1 U9218 ( .B1(n9866), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7650), .ZN(
        n7651) );
  OAI211_X1 U9219 ( .C1(n9867), .C2(n7815), .A(n7652), .B(n7651), .ZN(n7653)
         );
  AOI21_X1 U9220 ( .B1(n9865), .B2(n7654), .A(n7653), .ZN(n7655) );
  INV_X1 U9221 ( .A(n7655), .ZN(P2_U3260) );
  AOI21_X1 U9222 ( .B1(n7657), .B2(n9826), .A(n7656), .ZN(n7665) );
  NAND2_X1 U9223 ( .A1(n8046), .A2(n7658), .ZN(n7660) );
  OAI211_X1 U9224 ( .C1(n7661), .C2(n9844), .A(n7660), .B(n7659), .ZN(n7662)
         );
  AOI21_X1 U9225 ( .B1(n9859), .B2(n7663), .A(n7662), .ZN(n7664) );
  OAI21_X1 U9226 ( .B1(n7665), .B2(n9854), .A(n7664), .ZN(P2_U3226) );
  INV_X1 U9227 ( .A(n7666), .ZN(n7671) );
  AOI21_X1 U9228 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8510), .A(n7667), .ZN(
        n7668) );
  OAI21_X1 U9229 ( .B1(n7671), .B2(n8513), .A(n7668), .ZN(P2_U3335) );
  NOR2_X1 U9230 ( .A1(n7669), .A2(n4309), .ZN(n8954) );
  AOI21_X1 U9231 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9376), .A(n8954), .ZN(
        n7670) );
  OAI21_X1 U9232 ( .B1(n7671), .B2(n9378), .A(n7670), .ZN(P1_U3330) );
  XNOR2_X1 U9233 ( .A(n7672), .B(n7674), .ZN(n7800) );
  INV_X1 U9234 ( .A(n7800), .ZN(n7685) );
  OAI211_X1 U9235 ( .C1(n7675), .C2(n7674), .A(n7673), .B(n9922), .ZN(n7678)
         );
  NAND2_X1 U9236 ( .A1(n8092), .A2(n9832), .ZN(n7677) );
  NAND2_X1 U9237 ( .A1(n8090), .A2(n9834), .ZN(n7676) );
  AND2_X1 U9238 ( .A1(n7677), .A2(n7676), .ZN(n9633) );
  NAND2_X1 U9239 ( .A1(n7678), .A2(n9633), .ZN(n7798) );
  INV_X1 U9240 ( .A(n7743), .ZN(n7679) );
  AOI211_X1 U9241 ( .C1(n9638), .C2(n4395), .A(n10004), .B(n7679), .ZN(n7799)
         );
  NAND2_X1 U9242 ( .A1(n7799), .A2(n9929), .ZN(n7682) );
  AOI22_X1 U9243 ( .A1(n9942), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7680), .B2(
        n9928), .ZN(n7681) );
  OAI211_X1 U9244 ( .C1(n4481), .C2(n8374), .A(n7682), .B(n7681), .ZN(n7683)
         );
  AOI21_X1 U9245 ( .B1(n7798), .B2(n9938), .A(n7683), .ZN(n7684) );
  OAI21_X1 U9246 ( .B1(n7685), .B2(n8385), .A(n7684), .ZN(P2_U3282) );
  INV_X1 U9247 ( .A(n7686), .ZN(n7687) );
  AOI21_X1 U9248 ( .B1(n8599), .B2(n8969), .A(n7687), .ZN(n7689) );
  INV_X1 U9249 ( .A(n7782), .ZN(n8967) );
  NAND2_X1 U9250 ( .A1(n8967), .A2(n9608), .ZN(n7688) );
  OAI211_X1 U9251 ( .C1(n9625), .C2(n7690), .A(n7689), .B(n7688), .ZN(n7696)
         );
  INV_X1 U9252 ( .A(n7691), .ZN(n7692) );
  AOI211_X1 U9253 ( .C1(n7694), .C2(n7693), .A(n9618), .B(n7692), .ZN(n7695)
         );
  AOI211_X1 U9254 ( .C1(n8611), .C2(n7697), .A(n7696), .B(n7695), .ZN(n7698)
         );
  INV_X1 U9255 ( .A(n7698), .ZN(P1_U3234) );
  OAI211_X1 U9256 ( .C1(n7701), .C2(n7700), .A(n7699), .B(n9841), .ZN(n7708)
         );
  INV_X1 U9257 ( .A(n7702), .ZN(n7704) );
  OAI21_X1 U9258 ( .B1(n9844), .B2(n7704), .A(n7703), .ZN(n7705) );
  AOI21_X1 U9259 ( .B1(n7706), .B2(n8046), .A(n7705), .ZN(n7707) );
  OAI211_X1 U9260 ( .C1(n7732), .C2(n5795), .A(n7708), .B(n7707), .ZN(P2_U3236) );
  INV_X1 U9261 ( .A(n7709), .ZN(n7751) );
  AOI22_X1 U9262 ( .A1(n7710), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n8510), .ZN(n7711) );
  OAI21_X1 U9263 ( .B1(n7751), .B2(n8513), .A(n7711), .ZN(P2_U3334) );
  XNOR2_X1 U9264 ( .A(n7713), .B(n7712), .ZN(n7714) );
  XNOR2_X1 U9265 ( .A(n7715), .B(n7714), .ZN(n7721) );
  INV_X1 U9266 ( .A(n7716), .ZN(n7788) );
  AND2_X1 U9267 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9673) );
  NOR2_X1 U9268 ( .A1(n9611), .A2(n7782), .ZN(n7717) );
  AOI211_X1 U9269 ( .C1(n9608), .C2(n8966), .A(n9673), .B(n7717), .ZN(n7718)
         );
  OAI21_X1 U9270 ( .B1(n9625), .B2(n7788), .A(n7718), .ZN(n7719) );
  AOI21_X1 U9271 ( .B1(n8611), .B2(n8707), .A(n7719), .ZN(n7720) );
  OAI21_X1 U9272 ( .B1(n7721), .B2(n9618), .A(n7720), .ZN(P1_U3232) );
  OR2_X1 U9273 ( .A1(n7722), .A2(n9962), .ZN(n7726) );
  AND2_X1 U9274 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  AND2_X1 U9275 ( .A1(n7726), .A2(n7725), .ZN(n7730) );
  MUX2_X1 U9276 ( .A(n7730), .B(n7727), .S(n10024), .Z(n7728) );
  OAI21_X1 U9277 ( .B1(n7732), .B2(n8451), .A(n7728), .ZN(P2_U3533) );
  INV_X1 U9278 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7729) );
  MUX2_X1 U9279 ( .A(n7730), .B(n7729), .S(n10010), .Z(n7731) );
  OAI21_X1 U9280 ( .B1(n7732), .B2(n8494), .A(n7731), .ZN(P2_U3490) );
  OAI21_X1 U9281 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7842) );
  INV_X1 U9282 ( .A(n7842), .ZN(n7749) );
  OAI211_X1 U9283 ( .C1(n7738), .C2(n7737), .A(n7736), .B(n9922), .ZN(n7741)
         );
  NAND2_X1 U9284 ( .A1(n8089), .A2(n9834), .ZN(n7740) );
  NAND2_X1 U9285 ( .A1(n8091), .A2(n9832), .ZN(n7739) );
  AND2_X1 U9286 ( .A1(n7740), .A2(n7739), .ZN(n7906) );
  NAND2_X1 U9287 ( .A1(n7741), .A2(n7906), .ZN(n7840) );
  INV_X1 U9288 ( .A(n7744), .ZN(n7911) );
  INV_X1 U9289 ( .A(n7834), .ZN(n7742) );
  AOI211_X1 U9290 ( .C1(n7744), .C2(n7743), .A(n10004), .B(n7742), .ZN(n7841)
         );
  NAND2_X1 U9291 ( .A1(n7841), .A2(n9929), .ZN(n7746) );
  AOI22_X1 U9292 ( .A1(n9942), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7908), .B2(
        n9928), .ZN(n7745) );
  OAI211_X1 U9293 ( .C1(n7911), .C2(n8374), .A(n7746), .B(n7745), .ZN(n7747)
         );
  AOI21_X1 U9294 ( .B1(n7840), .B2(n9938), .A(n7747), .ZN(n7748) );
  OAI21_X1 U9295 ( .B1(n7749), .B2(n8385), .A(n7748), .ZN(P2_U3281) );
  INV_X1 U9296 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7750) );
  OAI222_X1 U9297 ( .A1(P1_U3084), .A2(n7752), .B1(n9378), .B2(n7751), .C1(
        n7750), .C2(n9369), .ZN(P1_U3329) );
  INV_X1 U9298 ( .A(n7753), .ZN(n7754) );
  INV_X1 U9299 ( .A(n8707), .ZN(n9649) );
  XNOR2_X1 U9300 ( .A(n9346), .B(n8703), .ZN(n8817) );
  XNOR2_X1 U9301 ( .A(n7864), .B(n8817), .ZN(n9349) );
  INV_X1 U9302 ( .A(n8691), .ZN(n7757) );
  OR2_X1 U9303 ( .A1(n8707), .A2(n8699), .ZN(n8690) );
  NAND2_X1 U9304 ( .A1(n8707), .A2(n8699), .ZN(n8876) );
  NAND2_X1 U9305 ( .A1(n7781), .A2(n8815), .ZN(n7780) );
  NAND2_X1 U9306 ( .A1(n7780), .A2(n8876), .ZN(n7871) );
  XNOR2_X1 U9307 ( .A(n7871), .B(n8817), .ZN(n7759) );
  OAI222_X1 U9308 ( .A1(n9250), .A2(n9247), .B1(n9248), .B2(n8699), .C1(n9246), 
        .C2(n7759), .ZN(n9344) );
  INV_X1 U9309 ( .A(n7777), .ZN(n7760) );
  AOI211_X1 U9310 ( .C1(n9346), .C2(n7760), .A(n9786), .B(n7866), .ZN(n9345)
         );
  NAND2_X1 U9311 ( .A1(n9345), .A2(n9254), .ZN(n7762) );
  AOI22_X1 U9312 ( .A1(n9205), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7769), .B2(
        n9255), .ZN(n7761) );
  OAI211_X1 U9313 ( .C1(n8712), .C2(n9260), .A(n7762), .B(n7761), .ZN(n7763)
         );
  AOI21_X1 U9314 ( .B1(n9344), .B2(n9263), .A(n7763), .ZN(n7764) );
  OAI21_X1 U9315 ( .B1(n9349), .B2(n9265), .A(n7764), .ZN(P1_U3277) );
  XNOR2_X1 U9316 ( .A(n7767), .B(n7766), .ZN(n7768) );
  XNOR2_X1 U9317 ( .A(n7765), .B(n7768), .ZN(n7775) );
  NAND2_X1 U9318 ( .A1(n8634), .A2(n7769), .ZN(n7772) );
  NOR2_X1 U9319 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7770), .ZN(n9688) );
  AOI21_X1 U9320 ( .B1(n8599), .B2(n9607), .A(n9688), .ZN(n7771) );
  OAI211_X1 U9321 ( .C1(n9247), .C2(n8630), .A(n7772), .B(n7771), .ZN(n7773)
         );
  AOI21_X1 U9322 ( .B1(n9346), .B2(n8611), .A(n7773), .ZN(n7774) );
  OAI21_X1 U9323 ( .B1(n7775), .B2(n9618), .A(n7774), .ZN(P1_U3213) );
  AND2_X1 U9324 ( .A1(n7776), .A2(n8707), .ZN(n7778) );
  OR2_X1 U9325 ( .A1(n7778), .A2(n7777), .ZN(n9650) );
  XOR2_X1 U9326 ( .A(n7779), .B(n8815), .Z(n7787) );
  OAI21_X1 U9327 ( .B1(n8815), .B2(n7781), .A(n7780), .ZN(n7784) );
  OAI22_X1 U9328 ( .A1(n8703), .A2(n9250), .B1(n7782), .B2(n9248), .ZN(n7783)
         );
  AOI21_X1 U9329 ( .B1(n7784), .B2(n9237), .A(n7783), .ZN(n7785) );
  OAI21_X1 U9330 ( .B1(n7787), .B2(n7786), .A(n7785), .ZN(n9651) );
  NAND2_X1 U9331 ( .A1(n9651), .A2(n9263), .ZN(n7791) );
  OAI22_X1 U9332 ( .A1(n9263), .A2(n4509), .B1(n7788), .B2(n9145), .ZN(n7789)
         );
  AOI21_X1 U9333 ( .B1(n8707), .B2(n9174), .A(n7789), .ZN(n7790) );
  OAI211_X1 U9334 ( .C1(n7792), .C2(n9650), .A(n7791), .B(n7790), .ZN(P1_U3278) );
  INV_X1 U9335 ( .A(n7793), .ZN(n7796) );
  OAI222_X1 U9336 ( .A1(n9369), .A2(n7794), .B1(n9378), .B2(n7796), .C1(
        P1_U3084), .C2(n6388), .ZN(P1_U3328) );
  OAI222_X1 U9337 ( .A1(n7947), .A2(n7797), .B1(n8513), .B2(n7796), .C1(n7795), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  INV_X1 U9338 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7801) );
  AOI211_X1 U9339 ( .C1(n7800), .C2(n10008), .A(n7799), .B(n7798), .ZN(n7803)
         );
  MUX2_X1 U9340 ( .A(n7801), .B(n7803), .S(n10012), .Z(n7802) );
  OAI21_X1 U9341 ( .B1(n4481), .B2(n8494), .A(n7802), .ZN(P2_U3493) );
  MUX2_X1 U9342 ( .A(n7804), .B(n7803), .S(n10026), .Z(n7805) );
  OAI21_X1 U9343 ( .B1(n4481), .B2(n8451), .A(n7805), .ZN(P2_U3534) );
  NAND2_X1 U9344 ( .A1(n7807), .A2(n7806), .ZN(n7809) );
  NAND2_X1 U9345 ( .A1(n7809), .A2(n7808), .ZN(n7811) );
  XNOR2_X1 U9346 ( .A(n7877), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7810) );
  NOR2_X1 U9347 ( .A1(n7810), .A2(n7811), .ZN(n7883) );
  AOI21_X1 U9348 ( .B1(n7811), .B2(n7810), .A(n7883), .ZN(n7824) );
  INV_X1 U9349 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7813) );
  OR2_X1 U9350 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9544), .ZN(n7812) );
  OAI21_X1 U9351 ( .B1(n8174), .B2(n7813), .A(n7812), .ZN(n7822) );
  NAND2_X1 U9352 ( .A1(n7815), .A2(n7814), .ZN(n7817) );
  NAND2_X1 U9353 ( .A1(n7817), .A2(n7816), .ZN(n7820) );
  NAND2_X1 U9354 ( .A1(n7877), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7818) );
  OAI21_X1 U9355 ( .B1(n7877), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7818), .ZN(
        n7819) );
  NOR2_X1 U9356 ( .A1(n7819), .A2(n7820), .ZN(n7876) );
  AOI211_X1 U9357 ( .C1(n7820), .C2(n7819), .A(n7876), .B(n7879), .ZN(n7821)
         );
  AOI211_X1 U9358 ( .C1(n8169), .C2(n7877), .A(n7822), .B(n7821), .ZN(n7823)
         );
  OAI21_X1 U9359 ( .B1(n7824), .B2(n9868), .A(n7823), .ZN(P2_U3261) );
  AOI21_X1 U9360 ( .B1(n7827), .B2(n7826), .A(n7825), .ZN(n7828) );
  INV_X1 U9361 ( .A(n7828), .ZN(n8461) );
  INV_X1 U9362 ( .A(n7829), .ZN(n7830) );
  AOI21_X1 U9363 ( .B1(n7832), .B2(n7831), .A(n7830), .ZN(n7833) );
  AOI22_X1 U9364 ( .A1(n9834), .A2(n8088), .B1(n8090), .B2(n9832), .ZN(n8010)
         );
  OAI21_X1 U9365 ( .B1(n7833), .B2(n9907), .A(n8010), .ZN(n8457) );
  INV_X1 U9366 ( .A(n8459), .ZN(n7837) );
  AOI211_X1 U9367 ( .C1(n8459), .C2(n7834), .A(n10004), .B(n8368), .ZN(n8458)
         );
  NAND2_X1 U9368 ( .A1(n8458), .A2(n9929), .ZN(n7836) );
  AOI22_X1 U9369 ( .A1(n9942), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8012), .B2(
        n9928), .ZN(n7835) );
  OAI211_X1 U9370 ( .C1(n7837), .C2(n8374), .A(n7836), .B(n7835), .ZN(n7838)
         );
  AOI21_X1 U9371 ( .B1(n8457), .B2(n9938), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9372 ( .B1(n8461), .B2(n8385), .A(n7839), .ZN(P2_U3280) );
  INV_X1 U9373 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7843) );
  AOI211_X1 U9374 ( .C1(n7842), .C2(n10008), .A(n7841), .B(n7840), .ZN(n7845)
         );
  MUX2_X1 U9375 ( .A(n7843), .B(n7845), .S(n10012), .Z(n7844) );
  OAI21_X1 U9376 ( .B1(n7911), .B2(n8494), .A(n7844), .ZN(P2_U3496) );
  INV_X1 U9377 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7846) );
  MUX2_X1 U9378 ( .A(n7846), .B(n7845), .S(n10026), .Z(n7847) );
  OAI21_X1 U9379 ( .B1(n7911), .B2(n8451), .A(n7847), .ZN(P2_U3535) );
  XNOR2_X1 U9380 ( .A(n7850), .B(n7849), .ZN(n7851) );
  XNOR2_X1 U9381 ( .A(n7848), .B(n7851), .ZN(n7856) );
  NAND2_X1 U9382 ( .A1(n8634), .A2(n7869), .ZN(n7853) );
  AND2_X1 U9383 ( .A1(n4309), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9707) );
  AOI21_X1 U9384 ( .B1(n9233), .B2(n9608), .A(n9707), .ZN(n7852) );
  OAI211_X1 U9385 ( .C1(n8703), .C2(n9611), .A(n7853), .B(n7852), .ZN(n7854)
         );
  AOI21_X1 U9386 ( .B1(n9339), .B2(n8611), .A(n7854), .ZN(n7855) );
  OAI21_X1 U9387 ( .B1(n7856), .B2(n9618), .A(n7855), .ZN(P1_U3239) );
  INV_X1 U9388 ( .A(n7857), .ZN(n7861) );
  AOI22_X1 U9389 ( .A1(n7858), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n8510), .ZN(n7859) );
  OAI21_X1 U9390 ( .B1(n7861), .B2(n8513), .A(n7859), .ZN(P2_U3332) );
  OAI222_X1 U9391 ( .A1(n4309), .A2(n7862), .B1(n9378), .B2(n7861), .C1(n7860), 
        .C2(n9369), .ZN(P1_U3327) );
  NOR2_X1 U9392 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NOR2_X1 U9393 ( .A1(n7865), .A2(n4848), .ZN(n7915) );
  AND2_X1 U9394 ( .A1(n7916), .A2(n8965), .ZN(n8883) );
  NAND2_X1 U9395 ( .A1(n9339), .A2(n9247), .ZN(n8838) );
  INV_X1 U9396 ( .A(n8838), .ZN(n8714) );
  XNOR2_X1 U9397 ( .A(n7915), .B(n8818), .ZN(n9343) );
  INV_X1 U9398 ( .A(n7866), .ZN(n7868) );
  INV_X1 U9399 ( .A(n9253), .ZN(n7867) );
  AOI21_X1 U9400 ( .B1(n9339), .B2(n7868), .A(n7867), .ZN(n9340) );
  AOI22_X1 U9401 ( .A1(n9205), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7869), .B2(
        n9255), .ZN(n7870) );
  OAI21_X1 U9402 ( .B1(n7916), .B2(n9260), .A(n7870), .ZN(n7874) );
  OR2_X1 U9403 ( .A1(n9346), .A2(n8703), .ZN(n8879) );
  XNOR2_X1 U9404 ( .A(n7921), .B(n8818), .ZN(n7872) );
  AOI222_X1 U9405 ( .A1(n9237), .A2(n7872), .B1(n9233), .B2(n9234), .C1(n8966), 
        .C2(n9232), .ZN(n9342) );
  NOR2_X1 U9406 ( .A1(n9342), .A2(n9205), .ZN(n7873) );
  AOI211_X1 U9407 ( .C1(n9340), .C2(n9240), .A(n7874), .B(n7873), .ZN(n7875)
         );
  OAI21_X1 U9408 ( .B1(n9343), .B2(n9265), .A(n7875), .ZN(P1_U3276) );
  NAND2_X1 U9409 ( .A1(n8150), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7878) );
  OAI21_X1 U9410 ( .B1(n8150), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7878), .ZN(
        n7880) );
  AOI211_X1 U9411 ( .C1(n7881), .C2(n7880), .A(n8149), .B(n7879), .ZN(n7891)
         );
  INV_X1 U9412 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9419) );
  NOR2_X1 U9413 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9419), .ZN(n7882) );
  AOI21_X1 U9414 ( .B1(n9866), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7882), .ZN(
        n7889) );
  XNOR2_X1 U9415 ( .A(n8145), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7887) );
  INV_X1 U9416 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7884) );
  AOI21_X1 U9417 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7886) );
  NAND2_X1 U9418 ( .A1(n7887), .A2(n7886), .ZN(n8144) );
  OAI211_X1 U9419 ( .C1(n7887), .C2(n7886), .A(n9864), .B(n8144), .ZN(n7888)
         );
  OAI211_X1 U9420 ( .C1(n9867), .C2(n8145), .A(n7889), .B(n7888), .ZN(n7890)
         );
  OR2_X1 U9421 ( .A1(n7891), .A2(n7890), .ZN(P2_U3262) );
  AOI21_X1 U9422 ( .B1(n7893), .B2(n7892), .A(n9854), .ZN(n7895) );
  NAND2_X1 U9423 ( .A1(n7895), .A2(n7894), .ZN(n7900) );
  OAI22_X1 U9424 ( .A1(n7970), .A2(n8057), .B1(n7896), .B2(n8055), .ZN(n8379)
         );
  INV_X1 U9425 ( .A(n8379), .ZN(n7897) );
  OAI22_X1 U9426 ( .A1(n9844), .A2(n7897), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9419), .ZN(n7898) );
  AOI21_X1 U9427 ( .B1(n8372), .B2(n8046), .A(n7898), .ZN(n7899) );
  OAI211_X1 U9428 ( .C1(n8375), .C2(n5795), .A(n7900), .B(n7899), .ZN(P2_U3230) );
  INV_X1 U9429 ( .A(n8064), .ZN(n8037) );
  NAND2_X1 U9430 ( .A1(n8037), .A2(n8090), .ZN(n7904) );
  NAND2_X1 U9431 ( .A1(n9841), .A2(n8004), .ZN(n7903) );
  XNOR2_X1 U9432 ( .A(n7901), .B(n7902), .ZN(n8005) );
  MUX2_X1 U9433 ( .A(n7904), .B(n7903), .S(n8005), .Z(n7910) );
  OAI22_X1 U9434 ( .A1(n9844), .A2(n7906), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7905), .ZN(n7907) );
  AOI21_X1 U9435 ( .B1(n7908), .B2(n8046), .A(n7907), .ZN(n7909) );
  OAI211_X1 U9436 ( .C1(n7911), .C2(n5795), .A(n7910), .B(n7909), .ZN(P2_U3243) );
  INV_X1 U9437 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7913) );
  INV_X1 U9438 ( .A(n8638), .ZN(n8505) );
  OAI222_X1 U9439 ( .A1(n9369), .A2(n7913), .B1(n4309), .B2(n7912), .C1(n9378), 
        .C2(n8505), .ZN(P1_U3324) );
  OR2_X1 U9440 ( .A1(n9336), .A2(n8579), .ZN(n8885) );
  NAND2_X1 U9441 ( .A1(n9336), .A2(n8579), .ZN(n8834) );
  NAND2_X1 U9442 ( .A1(n8885), .A2(n8834), .ZN(n9243) );
  OR2_X1 U9443 ( .A1(n9324), .A2(n9197), .ZN(n8724) );
  NAND2_X1 U9444 ( .A1(n9324), .A2(n9197), .ZN(n8869) );
  NAND2_X1 U9445 ( .A1(n8724), .A2(n8869), .ZN(n9219) );
  NAND2_X1 U9446 ( .A1(n9208), .A2(n9182), .ZN(n7917) );
  NAND2_X1 U9447 ( .A1(n9316), .A2(n9162), .ZN(n7918) );
  INV_X1 U9448 ( .A(n9316), .ZN(n9189) );
  INV_X1 U9449 ( .A(n9162), .ZN(n9198) );
  OR2_X1 U9450 ( .A1(n9310), .A2(n9183), .ZN(n8737) );
  NAND2_X1 U9451 ( .A1(n9310), .A2(n9183), .ZN(n8734) );
  NAND2_X1 U9452 ( .A1(n8737), .A2(n8734), .ZN(n9170) );
  INV_X1 U9453 ( .A(n9310), .ZN(n8557) );
  NAND2_X1 U9454 ( .A1(n9144), .A2(n8553), .ZN(n7919) );
  NAND2_X1 U9455 ( .A1(n9290), .A2(n9116), .ZN(n8758) );
  NAND2_X1 U9456 ( .A1(n9086), .A2(n8758), .ZN(n9105) );
  NAND2_X1 U9457 ( .A1(n9096), .A2(n9105), .ZN(n9097) );
  NAND2_X1 U9458 ( .A1(n9097), .A2(n7920), .ZN(n9080) );
  NAND2_X1 U9459 ( .A1(n9280), .A2(n8631), .ZN(n8898) );
  XNOR2_X1 U9460 ( .A(n9036), .B(n8827), .ZN(n9282) );
  INV_X1 U9461 ( .A(n8834), .ZN(n7922) );
  NAND2_X1 U9462 ( .A1(n9329), .A2(n9249), .ZN(n8835) );
  NAND2_X1 U9463 ( .A1(n9231), .A2(n8835), .ZN(n9218) );
  OR2_X1 U9464 ( .A1(n9329), .A2(n9249), .ZN(n9217) );
  AND2_X1 U9465 ( .A1(n8724), .A2(n9217), .ZN(n8867) );
  INV_X1 U9466 ( .A(n8869), .ZN(n7923) );
  OR2_X1 U9467 ( .A1(n9202), .A2(n9182), .ZN(n8728) );
  NAND2_X1 U9468 ( .A1(n9202), .A2(n9182), .ZN(n8726) );
  NAND2_X1 U9469 ( .A1(n8728), .A2(n8726), .ZN(n9194) );
  INV_X1 U9470 ( .A(n8726), .ZN(n8865) );
  NAND2_X1 U9471 ( .A1(n9316), .A2(n9198), .ZN(n8796) );
  INV_X1 U9472 ( .A(n9170), .ZN(n9159) );
  OR2_X1 U9473 ( .A1(n9316), .A2(n9198), .ZN(n9156) );
  NAND3_X1 U9474 ( .A1(n9157), .A2(n9159), .A3(n9156), .ZN(n9158) );
  NAND2_X1 U9475 ( .A1(n9158), .A2(n8734), .ZN(n9150) );
  NAND2_X1 U9476 ( .A1(n9298), .A2(n9153), .ZN(n8746) );
  NAND2_X1 U9477 ( .A1(n9135), .A2(n9134), .ZN(n9133) );
  NAND2_X1 U9478 ( .A1(n9133), .A2(n8862), .ZN(n9113) );
  XNOR2_X1 U9479 ( .A(n9295), .B(n9107), .ZN(n9114) );
  AND2_X1 U9480 ( .A1(n9295), .A2(n9107), .ZN(n8744) );
  OR2_X1 U9481 ( .A1(n9283), .A2(n9108), .ZN(n8792) );
  AND2_X1 U9482 ( .A1(n8792), .A2(n9086), .ZN(n8935) );
  AND2_X1 U9483 ( .A1(n9283), .A2(n9108), .ZN(n8896) );
  NAND2_X1 U9484 ( .A1(n7924), .A2(n8827), .ZN(n9041) );
  OAI211_X1 U9485 ( .C1(n7924), .C2(n8827), .A(n9041), .B(n9237), .ZN(n7926)
         );
  NAND2_X1 U9486 ( .A1(n8962), .A2(n9232), .ZN(n7925) );
  OAI211_X1 U9487 ( .C1(n9049), .C2(n9250), .A(n7926), .B(n7925), .ZN(n9278)
         );
  INV_X1 U9488 ( .A(n9280), .ZN(n8527) );
  NAND2_X1 U9489 ( .A1(n9213), .A2(n9208), .ZN(n9199) );
  NOR2_X1 U9490 ( .A1(n9165), .A2(n9305), .ZN(n9143) );
  NAND2_X1 U9491 ( .A1(n9143), .A2(n9132), .ZN(n9126) );
  INV_X1 U9492 ( .A(n9283), .ZN(n9085) );
  INV_X1 U9493 ( .A(n9081), .ZN(n7928) );
  INV_X1 U9494 ( .A(n9063), .ZN(n7927) );
  AOI211_X1 U9495 ( .C1(n9280), .C2(n7928), .A(n9786), .B(n7927), .ZN(n9279)
         );
  NAND2_X1 U9496 ( .A1(n9279), .A2(n9203), .ZN(n7930) );
  AOI22_X1 U9497 ( .A1(n8524), .A2(n9255), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9205), .ZN(n7929) );
  OAI211_X1 U9498 ( .C1(n8527), .C2(n9260), .A(n7930), .B(n7929), .ZN(n7931)
         );
  AOI21_X1 U9499 ( .B1(n9278), .B2(n9263), .A(n7931), .ZN(n7932) );
  OAI21_X1 U9500 ( .B1(n9282), .B2(n9265), .A(n7932), .ZN(P1_U3264) );
  OAI21_X1 U9501 ( .B1(n7935), .B2(n7934), .A(n7933), .ZN(n7936) );
  NAND2_X1 U9502 ( .A1(n7936), .A2(n8626), .ZN(n7942) );
  OAI22_X1 U9503 ( .A1(n8630), .A2(n7938), .B1(n7937), .B2(n9611), .ZN(n7939)
         );
  AOI21_X1 U9504 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7940), .A(n7939), .ZN(
        n7941) );
  OAI211_X1 U9505 ( .C1(n7943), .C2(n8637), .A(n7942), .B(n7941), .ZN(P1_U3235) );
  OAI222_X1 U9506 ( .A1(n7947), .A2(n7946), .B1(n8513), .B2(n7945), .C1(n7944), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9507 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7949) );
  OAI222_X1 U9508 ( .A1(n9369), .A2(n7949), .B1(n9378), .B2(n7948), .C1(n6386), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  INV_X1 U9509 ( .A(n7951), .ZN(n7952) );
  AOI21_X1 U9510 ( .B1(n7950), .B2(n7952), .A(n9854), .ZN(n7957) );
  NOR3_X1 U9511 ( .A1(n7954), .A2(n7953), .A3(n8064), .ZN(n7956) );
  OAI21_X1 U9512 ( .B1(n7957), .B2(n7956), .A(n7955), .ZN(n7960) );
  AOI22_X1 U9513 ( .A1(n8077), .A2(n9834), .B1(n9832), .B2(n8079), .ZN(n8219)
         );
  OAI22_X1 U9514 ( .A1(n8219), .A2(n9844), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9540), .ZN(n7958) );
  AOI21_X1 U9515 ( .B1(n8223), .B2(n8046), .A(n7958), .ZN(n7959) );
  OAI211_X1 U9516 ( .C1(n4485), .C2(n5795), .A(n7960), .B(n7959), .ZN(P2_U3216) );
  AOI22_X1 U9517 ( .A1(n7963), .A2(n9841), .B1(n8037), .B2(n8082), .ZN(n7968)
         );
  OAI22_X1 U9518 ( .A1(n8020), .A2(n8057), .B1(n7964), .B2(n8055), .ZN(n8279)
         );
  AOI22_X1 U9519 ( .A1(n8279), .A2(n9851), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7965) );
  OAI21_X1 U9520 ( .B1(n8284), .B2(n9863), .A(n7965), .ZN(n7966) );
  AOI21_X1 U9521 ( .B1(n8421), .B2(n9859), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9522 ( .B1(n8017), .B2(n7968), .A(n7967), .ZN(P2_U3218) );
  INV_X1 U9523 ( .A(n7969), .ZN(n7973) );
  NOR3_X1 U9524 ( .A1(n7971), .A2(n7970), .A3(n8064), .ZN(n7972) );
  AOI21_X1 U9525 ( .B1(n7973), .B2(n9841), .A(n7972), .ZN(n7981) );
  AOI22_X1 U9526 ( .A1(n8085), .A2(n9834), .B1(n9832), .B2(n8087), .ZN(n8339)
         );
  INV_X1 U9527 ( .A(n7974), .ZN(n8342) );
  NAND2_X1 U9528 ( .A1(n8046), .A2(n8342), .ZN(n7975) );
  NAND2_X1 U9529 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8172) );
  OAI211_X1 U9530 ( .C1(n8339), .C2(n9844), .A(n7975), .B(n8172), .ZN(n7978)
         );
  NOR2_X1 U9531 ( .A1(n7976), .A2(n9854), .ZN(n7977) );
  AOI211_X1 U9532 ( .C1(n9859), .C2(n8443), .A(n7978), .B(n7977), .ZN(n7979)
         );
  OAI21_X1 U9533 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(P2_U3221) );
  INV_X1 U9534 ( .A(n7983), .ZN(n7984) );
  AOI21_X1 U9535 ( .B1(n7982), .B2(n7984), .A(n9854), .ZN(n7989) );
  NOR3_X1 U9536 ( .A1(n7986), .A2(n7985), .A3(n8064), .ZN(n7988) );
  OAI21_X1 U9537 ( .B1(n7989), .B2(n7988), .A(n7987), .ZN(n7993) );
  AOI22_X1 U9538 ( .A1(n8083), .A2(n9834), .B1(n9832), .B2(n8085), .ZN(n8311)
         );
  OAI22_X1 U9539 ( .A1(n9844), .A2(n8311), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7990), .ZN(n7991) );
  AOI21_X1 U9540 ( .B1(n8315), .B2(n8046), .A(n7991), .ZN(n7992) );
  OAI211_X1 U9541 ( .C1(n8318), .C2(n5795), .A(n7993), .B(n7992), .ZN(P2_U3225) );
  OAI211_X1 U9542 ( .C1(n7994), .C2(n7996), .A(n7995), .B(n9841), .ZN(n8002)
         );
  INV_X1 U9543 ( .A(n7997), .ZN(n8255) );
  NOR2_X1 U9544 ( .A1(n8020), .A2(n8055), .ZN(n7998) );
  AOI21_X1 U9545 ( .B1(n8079), .B2(n9834), .A(n7998), .ZN(n8248) );
  OAI22_X1 U9546 ( .A1(n8248), .A2(n9844), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7999), .ZN(n8000) );
  AOI21_X1 U9547 ( .B1(n8255), .B2(n8046), .A(n8000), .ZN(n8001) );
  OAI211_X1 U9548 ( .C1(n8479), .C2(n5795), .A(n8002), .B(n8001), .ZN(P2_U3227) );
  AOI22_X1 U9549 ( .A1(n8005), .A2(n8004), .B1(n8003), .B2(n7901), .ZN(n8009)
         );
  XNOR2_X1 U9550 ( .A(n8007), .B(n8006), .ZN(n8008) );
  XNOR2_X1 U9551 ( .A(n8009), .B(n8008), .ZN(n8015) );
  OAI22_X1 U9552 ( .A1(n9844), .A2(n8010), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9544), .ZN(n8011) );
  AOI21_X1 U9553 ( .B1(n8012), .B2(n8046), .A(n8011), .ZN(n8014) );
  NAND2_X1 U9554 ( .A1(n8459), .A2(n9859), .ZN(n8013) );
  OAI211_X1 U9555 ( .C1(n8015), .C2(n9854), .A(n8014), .B(n8013), .ZN(P2_U3228) );
  NOR2_X1 U9556 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  XNOR2_X1 U9557 ( .A(n8019), .B(n8018), .ZN(n8023) );
  OAI22_X1 U9558 ( .A1(n8023), .A2(n9854), .B1(n8020), .B2(n8064), .ZN(n8021)
         );
  OAI21_X1 U9559 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8027) );
  AND2_X1 U9560 ( .A1(n8082), .A2(n9832), .ZN(n8024) );
  AOI21_X1 U9561 ( .B1(n8080), .B2(n9834), .A(n8024), .ZN(n8264) );
  OAI22_X1 U9562 ( .A1(n8264), .A2(n9844), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9504), .ZN(n8025) );
  AOI21_X1 U9563 ( .B1(n8272), .B2(n8046), .A(n8025), .ZN(n8026) );
  OAI211_X1 U9564 ( .C1(n4756), .C2(n5795), .A(n8027), .B(n8026), .ZN(P2_U3231) );
  AOI21_X1 U9565 ( .B1(n8029), .B2(n8028), .A(n9854), .ZN(n8030) );
  NAND2_X1 U9566 ( .A1(n8030), .A2(n7982), .ZN(n8034) );
  AOI22_X1 U9567 ( .A1(n8084), .A2(n9834), .B1(n9832), .B2(n8086), .ZN(n8326)
         );
  OAI22_X1 U9568 ( .A1(n9844), .A2(n8326), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8031), .ZN(n8032) );
  AOI21_X1 U9569 ( .B1(n8330), .B2(n8046), .A(n8032), .ZN(n8033) );
  OAI211_X1 U9570 ( .C1(n8489), .C2(n5795), .A(n8034), .B(n8033), .ZN(P2_U3235) );
  NAND2_X1 U9571 ( .A1(n8299), .A2(n9987), .ZN(n8428) );
  NAND2_X1 U9572 ( .A1(n8036), .A2(n8035), .ZN(n8049) );
  NAND2_X1 U9573 ( .A1(n8037), .A2(n8083), .ZN(n8041) );
  NAND2_X1 U9574 ( .A1(n9841), .A2(n8038), .ZN(n8040) );
  MUX2_X1 U9575 ( .A(n8041), .B(n8040), .S(n8039), .Z(n8048) );
  NAND2_X1 U9576 ( .A1(n8082), .A2(n9834), .ZN(n8043) );
  NAND2_X1 U9577 ( .A1(n8084), .A2(n9832), .ZN(n8042) );
  NAND2_X1 U9578 ( .A1(n8043), .A2(n8042), .ZN(n8293) );
  INV_X1 U9579 ( .A(n8293), .ZN(n8044) );
  OAI22_X1 U9580 ( .A1(n9844), .A2(n8044), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9530), .ZN(n8045) );
  AOI21_X1 U9581 ( .B1(n8301), .B2(n8046), .A(n8045), .ZN(n8047) );
  OAI211_X1 U9582 ( .C1(n8428), .C2(n8049), .A(n8048), .B(n8047), .ZN(P2_U3237) );
  INV_X1 U9583 ( .A(n8050), .ZN(n8051) );
  AOI21_X1 U9584 ( .B1(n7894), .B2(n8051), .A(n9854), .ZN(n8054) );
  NOR3_X1 U9585 ( .A1(n8052), .A2(n8056), .A3(n8064), .ZN(n8053) );
  OAI21_X1 U9586 ( .B1(n8054), .B2(n8053), .A(n7969), .ZN(n8061) );
  OAI22_X1 U9587 ( .A1(n8058), .A2(n8057), .B1(n8056), .B2(n8055), .ZN(n8353)
         );
  AND2_X1 U9588 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8156) );
  NOR2_X1 U9589 ( .A1(n9863), .A2(n8358), .ZN(n8059) );
  AOI211_X1 U9590 ( .C1(n9851), .C2(n8353), .A(n8156), .B(n8059), .ZN(n8060)
         );
  OAI211_X1 U9591 ( .C1(n8495), .C2(n5795), .A(n8061), .B(n8060), .ZN(P2_U3240) );
  INV_X1 U9592 ( .A(n8406), .ZN(n8075) );
  INV_X1 U9593 ( .A(n8062), .ZN(n8063) );
  AOI21_X1 U9594 ( .B1(n7995), .B2(n8063), .A(n9854), .ZN(n8068) );
  NOR3_X1 U9595 ( .A1(n8066), .A2(n8065), .A3(n8064), .ZN(n8067) );
  OAI21_X1 U9596 ( .B1(n8068), .B2(n8067), .A(n7950), .ZN(n8074) );
  AND2_X1 U9597 ( .A1(n8080), .A2(n9832), .ZN(n8069) );
  AOI21_X1 U9598 ( .B1(n8078), .B2(n9834), .A(n8069), .ZN(n8235) );
  INV_X1 U9599 ( .A(n8235), .ZN(n8072) );
  INV_X1 U9600 ( .A(n8070), .ZN(n8239) );
  OAI22_X1 U9601 ( .A1(n8239), .A2(n9863), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9527), .ZN(n8071) );
  AOI21_X1 U9602 ( .B1(n8072), .B2(n9851), .A(n8071), .ZN(n8073) );
  OAI211_X1 U9603 ( .C1(n8075), .C2(n5795), .A(n8074), .B(n8073), .ZN(P2_U3242) );
  MUX2_X1 U9604 ( .A(n8076), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8103), .Z(
        P2_U3581) );
  MUX2_X1 U9605 ( .A(n8077), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8103), .Z(
        P2_U3580) );
  MUX2_X1 U9606 ( .A(n8078), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8103), .Z(
        P2_U3579) );
  MUX2_X1 U9607 ( .A(n8079), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8103), .Z(
        P2_U3578) );
  MUX2_X1 U9608 ( .A(n8080), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8103), .Z(
        P2_U3577) );
  MUX2_X1 U9609 ( .A(n8081), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8103), .Z(
        P2_U3576) );
  MUX2_X1 U9610 ( .A(n8082), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8103), .Z(
        P2_U3575) );
  MUX2_X1 U9611 ( .A(n8083), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8103), .Z(
        P2_U3574) );
  MUX2_X1 U9612 ( .A(n8084), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8103), .Z(
        P2_U3573) );
  MUX2_X1 U9613 ( .A(n8085), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8103), .Z(
        P2_U3572) );
  MUX2_X1 U9614 ( .A(n8086), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8103), .Z(
        P2_U3571) );
  MUX2_X1 U9615 ( .A(n8087), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8103), .Z(
        P2_U3570) );
  MUX2_X1 U9616 ( .A(n8088), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8103), .Z(
        P2_U3569) );
  MUX2_X1 U9617 ( .A(n8089), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8098), .Z(
        P2_U3568) );
  MUX2_X1 U9618 ( .A(n8090), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8098), .Z(
        P2_U3567) );
  MUX2_X1 U9619 ( .A(n8091), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8098), .Z(
        P2_U3566) );
  MUX2_X1 U9620 ( .A(n8092), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8098), .Z(
        P2_U3565) );
  MUX2_X1 U9621 ( .A(n8093), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8098), .Z(
        P2_U3564) );
  MUX2_X1 U9622 ( .A(n8094), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8098), .Z(
        P2_U3563) );
  MUX2_X1 U9623 ( .A(n8095), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8098), .Z(
        P2_U3562) );
  MUX2_X1 U9624 ( .A(n8096), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8098), .Z(
        P2_U3561) );
  MUX2_X1 U9625 ( .A(n8097), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8098), .Z(
        P2_U3560) );
  MUX2_X1 U9626 ( .A(n8099), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8098), .Z(
        P2_U3559) );
  MUX2_X1 U9627 ( .A(n8100), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8103), .Z(
        P2_U3558) );
  MUX2_X1 U9628 ( .A(n8101), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8103), .Z(
        P2_U3557) );
  MUX2_X1 U9629 ( .A(n8102), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8103), .Z(
        P2_U3556) );
  MUX2_X1 U9630 ( .A(n9835), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8103), .Z(
        P2_U3555) );
  MUX2_X1 U9631 ( .A(n5637), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8103), .Z(
        P2_U3554) );
  MUX2_X1 U9632 ( .A(n9833), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8103), .Z(
        P2_U3553) );
  MUX2_X1 U9633 ( .A(n8104), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8103), .Z(
        P2_U3552) );
  OAI211_X1 U9634 ( .C1(n8107), .C2(n8106), .A(n9865), .B(n8105), .ZN(n8116)
         );
  AOI22_X1 U9635 ( .A1(n9866), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8115) );
  NAND2_X1 U9636 ( .A1(n8169), .A2(n8109), .ZN(n8114) );
  INV_X1 U9637 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n8110) );
  INV_X1 U9638 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U9639 ( .A1(n8110), .A2(n10013), .ZN(n8112) );
  OAI211_X1 U9640 ( .C1(n8112), .C2(n8111), .A(n9864), .B(n8123), .ZN(n8113)
         );
  NAND4_X1 U9641 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(
        P2_U3246) );
  OAI211_X1 U9642 ( .C1(n8119), .C2(n8118), .A(n9865), .B(n8117), .ZN(n8130)
         );
  AOI22_X1 U9643 ( .A1(n9866), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8129) );
  NAND2_X1 U9644 ( .A1(n8169), .A2(n8120), .ZN(n8128) );
  INV_X1 U9645 ( .A(n8121), .ZN(n8126) );
  NAND3_X1 U9646 ( .A1(n8124), .A2(n8123), .A3(n8122), .ZN(n8125) );
  NAND3_X1 U9647 ( .A1(n9864), .A2(n8126), .A3(n8125), .ZN(n8127) );
  NAND4_X1 U9648 ( .A1(n8130), .A2(n8129), .A3(n8128), .A4(n8127), .ZN(
        P2_U3247) );
  OAI21_X1 U9649 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8134) );
  NAND2_X1 U9650 ( .A1(n9865), .A2(n8134), .ZN(n8143) );
  NOR2_X1 U9651 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9816), .ZN(n8135) );
  AOI21_X1 U9652 ( .B1(n9866), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8135), .ZN(
        n8142) );
  NAND2_X1 U9653 ( .A1(n8169), .A2(n8136), .ZN(n8141) );
  OAI211_X1 U9654 ( .C1(n8139), .C2(n8138), .A(n9864), .B(n8137), .ZN(n8140)
         );
  NAND4_X1 U9655 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(
        P2_U3256) );
  INV_X1 U9656 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8146) );
  OAI21_X1 U9657 ( .B1(n8146), .B2(n8145), .A(n8144), .ZN(n8148) );
  INV_X1 U9658 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8449) );
  AOI22_X1 U9659 ( .A1(n8151), .A2(n8449), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8165), .ZN(n8147) );
  NOR2_X1 U9660 ( .A1(n8148), .A2(n8147), .ZN(n8164) );
  AOI21_X1 U9661 ( .B1(n8148), .B2(n8147), .A(n8164), .ZN(n8159) );
  INV_X1 U9662 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U9663 ( .A1(n8153), .A2(n8152), .ZN(n8162) );
  OAI21_X1 U9664 ( .B1(n8153), .B2(n8152), .A(n8162), .ZN(n8154) );
  NAND2_X1 U9665 ( .A1(n8154), .A2(n9865), .ZN(n8158) );
  NOR2_X1 U9666 ( .A1(n9867), .A2(n8165), .ZN(n8155) );
  AOI211_X1 U9667 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n9866), .A(n8156), .B(
        n8155), .ZN(n8157) );
  OAI211_X1 U9668 ( .C1(n8159), .C2(n9868), .A(n8158), .B(n8157), .ZN(P2_U3263) );
  INV_X1 U9669 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U9670 ( .A1(n8160), .A2(n8165), .ZN(n8161) );
  NAND2_X1 U9671 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  XNOR2_X1 U9672 ( .A(n8163), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8168) );
  AOI21_X1 U9673 ( .B1(n8449), .B2(n8165), .A(n8164), .ZN(n8166) );
  XOR2_X1 U9674 ( .A(n8166), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8167) );
  AOI22_X1 U9675 ( .A1(n8168), .A2(n9865), .B1(n9864), .B2(n8167), .ZN(n8171)
         );
  INV_X1 U9676 ( .A(n8167), .ZN(n8170) );
  XOR2_X1 U9677 ( .A(n8185), .B(n8175), .Z(n8176) );
  NOR2_X1 U9678 ( .A1(n8176), .A2(n10004), .ZN(n8387) );
  NAND2_X1 U9679 ( .A1(n8387), .A2(n9929), .ZN(n8180) );
  NOR2_X1 U9680 ( .A1(n8178), .A2(n8177), .ZN(n8386) );
  INV_X1 U9681 ( .A(n8386), .ZN(n8390) );
  NOR2_X1 U9682 ( .A1(n9942), .A2(n8390), .ZN(n8187) );
  AOI21_X1 U9683 ( .B1(n9942), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8187), .ZN(
        n8179) );
  OAI211_X1 U9684 ( .C1(n8465), .C2(n8374), .A(n8180), .B(n8179), .ZN(P2_U3265) );
  NAND2_X1 U9685 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  NAND2_X1 U9686 ( .A1(n8183), .A2(n9926), .ZN(n8184) );
  OR2_X1 U9687 ( .A1(n8185), .A2(n8184), .ZN(n8391) );
  NOR2_X1 U9688 ( .A1(n8469), .A2(n8374), .ZN(n8186) );
  AOI211_X1 U9689 ( .C1(n9942), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8187), .B(
        n8186), .ZN(n8188) );
  OAI21_X1 U9690 ( .B1(n8192), .B2(n8391), .A(n8188), .ZN(P2_U3266) );
  NAND2_X1 U9691 ( .A1(n8189), .A2(n9934), .ZN(n8198) );
  INV_X1 U9692 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8190) );
  OAI22_X1 U9693 ( .A1(n8191), .A2(n9894), .B1(n9938), .B2(n8190), .ZN(n8195)
         );
  NOR2_X1 U9694 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  AOI211_X1 U9695 ( .C1(n9931), .C2(n8196), .A(n8195), .B(n8194), .ZN(n8197)
         );
  OAI211_X1 U9696 ( .C1(n8199), .C2(n9942), .A(n8198), .B(n8197), .ZN(P2_U3267) );
  OAI211_X1 U9697 ( .C1(n8201), .C2(n8204), .A(n8200), .B(n9922), .ZN(n8203)
         );
  NAND2_X1 U9698 ( .A1(n8203), .A2(n8202), .ZN(n8394) );
  INV_X1 U9699 ( .A(n8394), .ZN(n8213) );
  XNOR2_X1 U9700 ( .A(n8205), .B(n8204), .ZN(n8396) );
  NAND2_X1 U9701 ( .A1(n8396), .A2(n9934), .ZN(n8212) );
  AOI211_X1 U9702 ( .C1(n8207), .C2(n4487), .A(n10004), .B(n8206), .ZN(n8395)
         );
  AOI22_X1 U9703 ( .A1(n8208), .A2(n9928), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9942), .ZN(n8209) );
  OAI21_X1 U9704 ( .B1(n8473), .B2(n8374), .A(n8209), .ZN(n8210) );
  AOI21_X1 U9705 ( .B1(n8395), .B2(n9929), .A(n8210), .ZN(n8211) );
  OAI211_X1 U9706 ( .C1(n8213), .C2(n9942), .A(n8212), .B(n8211), .ZN(P2_U3268) );
  XOR2_X1 U9707 ( .A(n8214), .B(n8216), .Z(n8403) );
  NAND2_X1 U9708 ( .A1(n8215), .A2(n9922), .ZN(n8221) );
  INV_X1 U9709 ( .A(n8216), .ZN(n8217) );
  AOI21_X1 U9710 ( .B1(n8230), .B2(n8218), .A(n8217), .ZN(n8220) );
  OAI21_X1 U9711 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8399) );
  AOI211_X1 U9712 ( .C1(n8401), .C2(n8237), .A(n10004), .B(n8222), .ZN(n8400)
         );
  NAND2_X1 U9713 ( .A1(n8400), .A2(n9929), .ZN(n8225) );
  AOI22_X1 U9714 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n9942), .B1(n8223), .B2(
        n9928), .ZN(n8224) );
  OAI211_X1 U9715 ( .C1(n4485), .C2(n8374), .A(n8225), .B(n8224), .ZN(n8226)
         );
  AOI21_X1 U9716 ( .B1(n8399), .B2(n9938), .A(n8226), .ZN(n8227) );
  OAI21_X1 U9717 ( .B1(n8403), .B2(n8385), .A(n8227), .ZN(P2_U3269) );
  XNOR2_X1 U9718 ( .A(n8229), .B(n8228), .ZN(n8408) );
  AOI22_X1 U9719 ( .A1(n8406), .A2(n9931), .B1(n9942), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8243) );
  INV_X1 U9720 ( .A(n8230), .ZN(n8234) );
  OAI21_X1 U9721 ( .B1(n8234), .B2(n8233), .A(n9922), .ZN(n8236) );
  NAND2_X1 U9722 ( .A1(n8236), .A2(n8235), .ZN(n8404) );
  INV_X1 U9723 ( .A(n8237), .ZN(n8238) );
  AOI211_X1 U9724 ( .C1(n8406), .C2(n8250), .A(n10004), .B(n8238), .ZN(n8405)
         );
  INV_X1 U9725 ( .A(n8405), .ZN(n8240) );
  OAI22_X1 U9726 ( .A1(n8240), .A2(n8254), .B1(n9894), .B2(n8239), .ZN(n8241)
         );
  OAI21_X1 U9727 ( .B1(n8404), .B2(n8241), .A(n9938), .ZN(n8242) );
  OAI211_X1 U9728 ( .C1(n8408), .C2(n8385), .A(n8243), .B(n8242), .ZN(P2_U3270) );
  XNOR2_X1 U9729 ( .A(n8245), .B(n8244), .ZN(n8411) );
  INV_X1 U9730 ( .A(n8411), .ZN(n8260) );
  NAND2_X1 U9731 ( .A1(n8249), .A2(n8248), .ZN(n8409) );
  INV_X1 U9732 ( .A(n8269), .ZN(n8252) );
  INV_X1 U9733 ( .A(n8250), .ZN(n8251) );
  AOI211_X1 U9734 ( .C1(n8253), .C2(n8252), .A(n10004), .B(n8251), .ZN(n8410)
         );
  NOR2_X1 U9735 ( .A1(n9942), .A2(n8254), .ZN(n8383) );
  NAND2_X1 U9736 ( .A1(n8410), .A2(n8383), .ZN(n8257) );
  AOI22_X1 U9737 ( .A1(n9942), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8255), .B2(
        n9928), .ZN(n8256) );
  OAI211_X1 U9738 ( .C1(n8479), .C2(n8374), .A(n8257), .B(n8256), .ZN(n8258)
         );
  AOI21_X1 U9739 ( .B1(n8409), .B2(n9938), .A(n8258), .ZN(n8259) );
  OAI21_X1 U9740 ( .B1(n8260), .B2(n8385), .A(n8259), .ZN(P2_U3271) );
  OAI211_X1 U9741 ( .C1(n8263), .C2(n8262), .A(n8261), .B(n9922), .ZN(n8265)
         );
  NAND2_X1 U9742 ( .A1(n8265), .A2(n8264), .ZN(n8414) );
  INV_X1 U9743 ( .A(n8414), .ZN(n8277) );
  OAI21_X1 U9744 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8416) );
  NAND2_X1 U9745 ( .A1(n8416), .A2(n9934), .ZN(n8276) );
  INV_X1 U9746 ( .A(n8283), .ZN(n8270) );
  AOI211_X1 U9747 ( .C1(n8271), .C2(n8270), .A(n10004), .B(n8269), .ZN(n8415)
         );
  AOI22_X1 U9748 ( .A1(n9942), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8272), .B2(
        n9928), .ZN(n8273) );
  OAI21_X1 U9749 ( .B1(n4756), .B2(n8374), .A(n8273), .ZN(n8274) );
  AOI21_X1 U9750 ( .B1(n8415), .B2(n9929), .A(n8274), .ZN(n8275) );
  OAI211_X1 U9751 ( .C1(n9942), .C2(n8277), .A(n8276), .B(n8275), .ZN(P2_U3272) );
  XNOR2_X1 U9752 ( .A(n8278), .B(n4558), .ZN(n8280) );
  AOI21_X1 U9753 ( .B1(n8280), .B2(n9922), .A(n8279), .ZN(n8423) );
  NAND2_X1 U9754 ( .A1(n8282), .A2(n8281), .ZN(n8419) );
  NAND3_X1 U9755 ( .A1(n4755), .A2(n9934), .A3(n8419), .ZN(n8290) );
  AOI211_X1 U9756 ( .C1(n8421), .C2(n8300), .A(n10004), .B(n8283), .ZN(n8420)
         );
  INV_X1 U9757 ( .A(n8421), .ZN(n8287) );
  INV_X1 U9758 ( .A(n8284), .ZN(n8285) );
  AOI22_X1 U9759 ( .A1(n9942), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8285), .B2(
        n9928), .ZN(n8286) );
  OAI21_X1 U9760 ( .B1(n8287), .B2(n8374), .A(n8286), .ZN(n8288) );
  AOI21_X1 U9761 ( .B1(n8420), .B2(n9929), .A(n8288), .ZN(n8289) );
  OAI211_X1 U9762 ( .C1(n9942), .C2(n8423), .A(n8290), .B(n8289), .ZN(P2_U3273) );
  AOI21_X1 U9763 ( .B1(n8292), .B2(n8291), .A(n9907), .ZN(n8295) );
  AOI21_X1 U9764 ( .B1(n8295), .B2(n8294), .A(n8293), .ZN(n8429) );
  XNOR2_X1 U9765 ( .A(n8296), .B(n8297), .ZN(n8426) );
  NAND2_X1 U9766 ( .A1(n8426), .A2(n9934), .ZN(n8307) );
  INV_X1 U9767 ( .A(n8298), .ZN(n8313) );
  INV_X1 U9768 ( .A(n8299), .ZN(n8303) );
  OAI211_X1 U9769 ( .C1(n8313), .C2(n8303), .A(n9926), .B(n8300), .ZN(n8427)
         );
  INV_X1 U9770 ( .A(n8427), .ZN(n8305) );
  AOI22_X1 U9771 ( .A1(n9942), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8301), .B2(
        n9928), .ZN(n8302) );
  OAI21_X1 U9772 ( .B1(n8303), .B2(n8374), .A(n8302), .ZN(n8304) );
  AOI21_X1 U9773 ( .B1(n8305), .B2(n9929), .A(n8304), .ZN(n8306) );
  OAI211_X1 U9774 ( .C1(n9942), .C2(n8429), .A(n8307), .B(n8306), .ZN(P2_U3274) );
  XOR2_X1 U9775 ( .A(n8308), .B(n8310), .Z(n8435) );
  XOR2_X1 U9776 ( .A(n8310), .B(n8309), .Z(n8312) );
  OAI21_X1 U9777 ( .B1(n8312), .B2(n9907), .A(n8311), .ZN(n8431) );
  INV_X1 U9778 ( .A(n8328), .ZN(n8314) );
  AOI211_X1 U9779 ( .C1(n8433), .C2(n8314), .A(n10004), .B(n8313), .ZN(n8432)
         );
  NAND2_X1 U9780 ( .A1(n8432), .A2(n9929), .ZN(n8317) );
  AOI22_X1 U9781 ( .A1(n9942), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8315), .B2(
        n9928), .ZN(n8316) );
  OAI211_X1 U9782 ( .C1(n8318), .C2(n8374), .A(n8317), .B(n8316), .ZN(n8319)
         );
  AOI21_X1 U9783 ( .B1(n8431), .B2(n9938), .A(n8319), .ZN(n8320) );
  OAI21_X1 U9784 ( .B1(n8435), .B2(n8385), .A(n8320), .ZN(P2_U3275) );
  XOR2_X1 U9785 ( .A(n8321), .B(n8322), .Z(n8438) );
  INV_X1 U9786 ( .A(n8438), .ZN(n8335) );
  NAND2_X1 U9787 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND3_X1 U9788 ( .A1(n8325), .A2(n9922), .A3(n8324), .ZN(n8327) );
  NAND2_X1 U9789 ( .A1(n8327), .A2(n8326), .ZN(n8436) );
  AOI211_X1 U9790 ( .C1(n8329), .C2(n4475), .A(n10004), .B(n8328), .ZN(n8437)
         );
  NAND2_X1 U9791 ( .A1(n8437), .A2(n9929), .ZN(n8332) );
  AOI22_X1 U9792 ( .A1(n9942), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8330), .B2(
        n9928), .ZN(n8331) );
  OAI211_X1 U9793 ( .C1(n8489), .C2(n8374), .A(n8332), .B(n8331), .ZN(n8333)
         );
  AOI21_X1 U9794 ( .B1(n8436), .B2(n9938), .A(n8333), .ZN(n8334) );
  OAI21_X1 U9795 ( .B1(n8335), .B2(n8385), .A(n8334), .ZN(P2_U3276) );
  XOR2_X1 U9796 ( .A(n8336), .B(n8337), .Z(n8445) );
  XOR2_X1 U9797 ( .A(n8338), .B(n8337), .Z(n8340) );
  OAI21_X1 U9798 ( .B1(n8340), .B2(n9907), .A(n8339), .ZN(n8441) );
  AOI211_X1 U9799 ( .C1(n8443), .C2(n8355), .A(n10004), .B(n8341), .ZN(n8442)
         );
  NAND2_X1 U9800 ( .A1(n8442), .A2(n8383), .ZN(n8344) );
  AOI22_X1 U9801 ( .A1(n9942), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8342), .B2(
        n9928), .ZN(n8343) );
  OAI211_X1 U9802 ( .C1(n4473), .C2(n8374), .A(n8344), .B(n8343), .ZN(n8345)
         );
  AOI21_X1 U9803 ( .B1(n8441), .B2(n9938), .A(n8345), .ZN(n8346) );
  OAI21_X1 U9804 ( .B1(n8445), .B2(n8385), .A(n8346), .ZN(P2_U3277) );
  XNOR2_X1 U9805 ( .A(n8347), .B(n8349), .ZN(n8448) );
  INV_X1 U9806 ( .A(n8448), .ZN(n8364) );
  INV_X1 U9807 ( .A(n8348), .ZN(n8376) );
  OAI21_X1 U9808 ( .B1(n8376), .B2(n8350), .A(n8349), .ZN(n8352) );
  AOI21_X1 U9809 ( .B1(n8352), .B2(n8351), .A(n9907), .ZN(n8354) );
  OR2_X1 U9810 ( .A1(n8354), .A2(n8353), .ZN(n8446) );
  INV_X1 U9811 ( .A(n8355), .ZN(n8356) );
  AOI211_X1 U9812 ( .C1(n8357), .C2(n8369), .A(n10004), .B(n8356), .ZN(n8447)
         );
  NAND2_X1 U9813 ( .A1(n8447), .A2(n9929), .ZN(n8361) );
  INV_X1 U9814 ( .A(n8358), .ZN(n8359) );
  AOI22_X1 U9815 ( .A1(n9942), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8359), .B2(
        n9928), .ZN(n8360) );
  OAI211_X1 U9816 ( .C1(n8495), .C2(n8374), .A(n8361), .B(n8360), .ZN(n8362)
         );
  AOI21_X1 U9817 ( .B1(n8446), .B2(n9938), .A(n8362), .ZN(n8363) );
  OAI21_X1 U9818 ( .B1(n8364), .B2(n8385), .A(n8363), .ZN(P2_U3278) );
  OAI21_X1 U9819 ( .B1(n8366), .B2(n8378), .A(n8365), .ZN(n8367) );
  INV_X1 U9820 ( .A(n8367), .ZN(n8456) );
  INV_X1 U9821 ( .A(n8368), .ZN(n8371) );
  INV_X1 U9822 ( .A(n8369), .ZN(n8370) );
  AOI211_X1 U9823 ( .C1(n8453), .C2(n8371), .A(n10004), .B(n8370), .ZN(n8452)
         );
  AOI22_X1 U9824 ( .A1(n9942), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8372), .B2(
        n9928), .ZN(n8373) );
  OAI21_X1 U9825 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n8382) );
  AOI211_X1 U9826 ( .C1(n8378), .C2(n8377), .A(n9907), .B(n8376), .ZN(n8380)
         );
  NOR2_X1 U9827 ( .A1(n8380), .A2(n8379), .ZN(n8455) );
  NOR2_X1 U9828 ( .A1(n8455), .A2(n9942), .ZN(n8381) );
  AOI211_X1 U9829 ( .C1(n8452), .C2(n8383), .A(n8382), .B(n8381), .ZN(n8384)
         );
  OAI21_X1 U9830 ( .B1(n8456), .B2(n8385), .A(n8384), .ZN(P2_U3279) );
  INV_X1 U9831 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8388) );
  NOR2_X1 U9832 ( .A1(n8387), .A2(n8386), .ZN(n8462) );
  MUX2_X1 U9833 ( .A(n8388), .B(n8462), .S(n10026), .Z(n8389) );
  OAI21_X1 U9834 ( .B1(n8465), .B2(n8451), .A(n8389), .ZN(P2_U3551) );
  NAND2_X1 U9835 ( .A1(n8391), .A2(n8390), .ZN(n8466) );
  MUX2_X1 U9836 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8466), .S(n10026), .Z(n8392) );
  INV_X1 U9837 ( .A(n8392), .ZN(n8393) );
  OAI21_X1 U9838 ( .B1(n8469), .B2(n8451), .A(n8393), .ZN(P2_U3550) );
  INV_X1 U9839 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8397) );
  AOI211_X1 U9840 ( .C1(n8396), .C2(n10008), .A(n8395), .B(n8394), .ZN(n8470)
         );
  MUX2_X1 U9841 ( .A(n8397), .B(n8470), .S(n10026), .Z(n8398) );
  OAI21_X1 U9842 ( .B1(n8473), .B2(n8451), .A(n8398), .ZN(P2_U3548) );
  AOI211_X1 U9843 ( .C1(n9987), .C2(n8401), .A(n8400), .B(n8399), .ZN(n8402)
         );
  OAI21_X1 U9844 ( .B1(n8403), .B2(n9962), .A(n8402), .ZN(n8474) );
  MUX2_X1 U9845 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8474), .S(n10026), .Z(
        P2_U3547) );
  AOI211_X1 U9846 ( .C1(n9987), .C2(n8406), .A(n8405), .B(n8404), .ZN(n8407)
         );
  OAI21_X1 U9847 ( .B1(n8408), .B2(n9962), .A(n8407), .ZN(n8475) );
  MUX2_X1 U9848 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8475), .S(n10026), .Z(
        P2_U3546) );
  INV_X1 U9849 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8412) );
  AOI211_X1 U9850 ( .C1(n8411), .C2(n10008), .A(n8410), .B(n8409), .ZN(n8476)
         );
  MUX2_X1 U9851 ( .A(n8412), .B(n8476), .S(n10026), .Z(n8413) );
  OAI21_X1 U9852 ( .B1(n8479), .B2(n8451), .A(n8413), .ZN(P2_U3545) );
  INV_X1 U9853 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8417) );
  AOI211_X1 U9854 ( .C1(n8416), .C2(n10008), .A(n8415), .B(n8414), .ZN(n8480)
         );
  MUX2_X1 U9855 ( .A(n8417), .B(n8480), .S(n10026), .Z(n8418) );
  OAI21_X1 U9856 ( .B1(n4756), .B2(n8451), .A(n8418), .ZN(P2_U3544) );
  NAND2_X1 U9857 ( .A1(n8419), .A2(n10008), .ZN(n8424) );
  AOI21_X1 U9858 ( .B1(n9987), .B2(n8421), .A(n8420), .ZN(n8422) );
  OAI211_X1 U9859 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8422), .ZN(n8483)
         );
  MUX2_X1 U9860 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8483), .S(n10026), .Z(
        P2_U3543) );
  NAND2_X1 U9861 ( .A1(n8426), .A2(n10008), .ZN(n8430) );
  NAND4_X1 U9862 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n8484)
         );
  MUX2_X1 U9863 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8484), .S(n10026), .Z(
        P2_U3542) );
  AOI211_X1 U9864 ( .C1(n9987), .C2(n8433), .A(n8432), .B(n8431), .ZN(n8434)
         );
  OAI21_X1 U9865 ( .B1(n8435), .B2(n9962), .A(n8434), .ZN(n8485) );
  MUX2_X1 U9866 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8485), .S(n10026), .Z(
        P2_U3541) );
  INV_X1 U9867 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8439) );
  AOI211_X1 U9868 ( .C1(n8438), .C2(n10008), .A(n8437), .B(n8436), .ZN(n8486)
         );
  MUX2_X1 U9869 ( .A(n8439), .B(n8486), .S(n10026), .Z(n8440) );
  OAI21_X1 U9870 ( .B1(n8489), .B2(n8451), .A(n8440), .ZN(P2_U3540) );
  AOI211_X1 U9871 ( .C1(n9987), .C2(n8443), .A(n8442), .B(n8441), .ZN(n8444)
         );
  OAI21_X1 U9872 ( .B1(n8445), .B2(n9962), .A(n8444), .ZN(n8490) );
  MUX2_X1 U9873 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8490), .S(n10026), .Z(
        P2_U3539) );
  AOI211_X1 U9874 ( .C1(n8448), .C2(n10008), .A(n8447), .B(n8446), .ZN(n8491)
         );
  MUX2_X1 U9875 ( .A(n8449), .B(n8491), .S(n10026), .Z(n8450) );
  OAI21_X1 U9876 ( .B1(n8495), .B2(n8451), .A(n8450), .ZN(P2_U3538) );
  AOI21_X1 U9877 ( .B1(n9987), .B2(n8453), .A(n8452), .ZN(n8454) );
  OAI211_X1 U9878 ( .C1(n8456), .C2(n9962), .A(n8455), .B(n8454), .ZN(n8496)
         );
  MUX2_X1 U9879 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8496), .S(n10026), .Z(
        P2_U3537) );
  AOI211_X1 U9880 ( .C1(n9987), .C2(n8459), .A(n8458), .B(n8457), .ZN(n8460)
         );
  OAI21_X1 U9881 ( .B1(n8461), .B2(n9962), .A(n8460), .ZN(n8497) );
  MUX2_X1 U9882 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8497), .S(n10026), .Z(
        P2_U3536) );
  INV_X1 U9883 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8463) );
  MUX2_X1 U9884 ( .A(n8463), .B(n8462), .S(n10012), .Z(n8464) );
  OAI21_X1 U9885 ( .B1(n8465), .B2(n8494), .A(n8464), .ZN(P2_U3519) );
  MUX2_X1 U9886 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8466), .S(n10012), .Z(n8467) );
  INV_X1 U9887 ( .A(n8467), .ZN(n8468) );
  OAI21_X1 U9888 ( .B1(n8469), .B2(n8494), .A(n8468), .ZN(P2_U3518) );
  MUX2_X1 U9889 ( .A(n8471), .B(n8470), .S(n10012), .Z(n8472) );
  OAI21_X1 U9890 ( .B1(n8473), .B2(n8494), .A(n8472), .ZN(P2_U3516) );
  MUX2_X1 U9891 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8474), .S(n10012), .Z(
        P2_U3515) );
  MUX2_X1 U9892 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8475), .S(n10012), .Z(
        P2_U3514) );
  MUX2_X1 U9893 ( .A(n8477), .B(n8476), .S(n10012), .Z(n8478) );
  OAI21_X1 U9894 ( .B1(n8479), .B2(n8494), .A(n8478), .ZN(P2_U3513) );
  MUX2_X1 U9895 ( .A(n8481), .B(n8480), .S(n10012), .Z(n8482) );
  OAI21_X1 U9896 ( .B1(n4756), .B2(n8494), .A(n8482), .ZN(P2_U3512) );
  MUX2_X1 U9897 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8483), .S(n10012), .Z(
        P2_U3511) );
  MUX2_X1 U9898 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8484), .S(n10012), .Z(
        P2_U3510) );
  MUX2_X1 U9899 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8485), .S(n10012), .Z(
        P2_U3509) );
  MUX2_X1 U9900 ( .A(n8487), .B(n8486), .S(n10012), .Z(n8488) );
  OAI21_X1 U9901 ( .B1(n8489), .B2(n8494), .A(n8488), .ZN(P2_U3508) );
  MUX2_X1 U9902 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8490), .S(n10012), .Z(
        P2_U3507) );
  INV_X1 U9903 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8492) );
  MUX2_X1 U9904 ( .A(n8492), .B(n8491), .S(n10012), .Z(n8493) );
  OAI21_X1 U9905 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(P2_U3505) );
  MUX2_X1 U9906 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8496), .S(n10012), .Z(
        P2_U3502) );
  MUX2_X1 U9907 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8497), .S(n10012), .Z(
        P2_U3499) );
  INV_X1 U9908 ( .A(n8654), .ZN(n9368) );
  NOR4_X1 U9909 ( .A1(n5021), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n8498), .ZN(n8499) );
  AOI21_X1 U9910 ( .B1(n8510), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8499), .ZN(
        n8500) );
  OAI21_X1 U9911 ( .B1(n9368), .B2(n8513), .A(n8500), .ZN(P2_U3327) );
  INV_X1 U9912 ( .A(n8646), .ZN(n9371) );
  AOI22_X1 U9913 ( .A1(n8501), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8510), .ZN(n8502) );
  OAI21_X1 U9914 ( .B1(n9371), .B2(n8513), .A(n8502), .ZN(P2_U3328) );
  AOI22_X1 U9915 ( .A1(n8503), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8510), .ZN(n8504) );
  OAI21_X1 U9916 ( .B1(n8505), .B2(n8513), .A(n8504), .ZN(P2_U3329) );
  INV_X1 U9917 ( .A(n8506), .ZN(n9374) );
  AOI21_X1 U9918 ( .B1(n8510), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8507), .ZN(
        n8508) );
  OAI21_X1 U9919 ( .B1(n9374), .B2(n8513), .A(n8508), .ZN(P2_U3330) );
  INV_X1 U9920 ( .A(n8509), .ZN(n9379) );
  AOI22_X1 U9921 ( .A1(n8511), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8510), .ZN(n8512) );
  OAI21_X1 U9922 ( .B1(n9379), .B2(n8513), .A(n8512), .ZN(P2_U3331) );
  MUX2_X1 U9923 ( .A(n8514), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U9924 ( .A(n8515), .ZN(n8520) );
  AOI21_X1 U9925 ( .B1(n8516), .B2(n8518), .A(n8517), .ZN(n8519) );
  OAI21_X1 U9926 ( .B1(n8520), .B2(n8519), .A(n8626), .ZN(n8526) );
  OAI22_X1 U9927 ( .A1(n9108), .A2(n9611), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8521), .ZN(n8523) );
  NOR2_X1 U9928 ( .A1(n9049), .A2(n8630), .ZN(n8522) );
  AOI211_X1 U9929 ( .C1(n8524), .C2(n8634), .A(n8523), .B(n8522), .ZN(n8525)
         );
  OAI211_X1 U9930 ( .C1(n8527), .C2(n8637), .A(n8526), .B(n8525), .ZN(P1_U3212) );
  XNOR2_X1 U9931 ( .A(n8529), .B(n8528), .ZN(n8530) );
  XNOR2_X1 U9932 ( .A(n8531), .B(n8530), .ZN(n8536) );
  NAND2_X1 U9933 ( .A1(n9136), .A2(n9608), .ZN(n8533) );
  AOI22_X1 U9934 ( .A1(n9161), .A2(n8599), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8532) );
  OAI211_X1 U9935 ( .C1(n9625), .C2(n9129), .A(n8533), .B(n8532), .ZN(n8534)
         );
  AOI21_X1 U9936 ( .B1(n9298), .B2(n8611), .A(n8534), .ZN(n8535) );
  OAI21_X1 U9937 ( .B1(n8536), .B2(n9618), .A(n8535), .ZN(P1_U3214) );
  NOR2_X1 U9938 ( .A1(n9208), .A2(n9784), .ZN(n9320) );
  INV_X1 U9939 ( .A(n9320), .ZN(n8546) );
  INV_X1 U9940 ( .A(n9621), .ZN(n8545) );
  INV_X1 U9941 ( .A(n8593), .ZN(n8540) );
  NOR3_X1 U9942 ( .A1(n8537), .A2(n8614), .A3(n8538), .ZN(n8539) );
  OAI21_X1 U9943 ( .B1(n8540), .B2(n8539), .A(n8626), .ZN(n8544) );
  NAND2_X1 U9944 ( .A1(n9608), .A2(n9162), .ZN(n8541) );
  NAND2_X1 U9945 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9021) );
  OAI211_X1 U9946 ( .C1(n9197), .C2(n9611), .A(n8541), .B(n9021), .ZN(n8542)
         );
  AOI21_X1 U9947 ( .B1(n8634), .B2(n9204), .A(n8542), .ZN(n8543) );
  OAI211_X1 U9948 ( .C1(n8546), .C2(n8545), .A(n8544), .B(n8543), .ZN(P1_U3217) );
  INV_X1 U9949 ( .A(n8547), .ZN(n8551) );
  NOR3_X1 U9950 ( .A1(n8595), .A2(n8549), .A3(n8548), .ZN(n8550) );
  OAI21_X1 U9951 ( .B1(n8551), .B2(n8550), .A(n8626), .ZN(n8556) );
  AOI22_X1 U9952 ( .A1(n8599), .A2(n9162), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8552) );
  OAI21_X1 U9953 ( .B1(n8553), .B2(n8630), .A(n8552), .ZN(n8554) );
  AOI21_X1 U9954 ( .B1(n9167), .B2(n8634), .A(n8554), .ZN(n8555) );
  OAI211_X1 U9955 ( .C1(n8557), .C2(n8637), .A(n8556), .B(n8555), .ZN(P1_U3221) );
  OAI21_X1 U9956 ( .B1(n8559), .B2(n8558), .A(n8625), .ZN(n8560) );
  NAND2_X1 U9957 ( .A1(n8560), .A2(n8626), .ZN(n8564) );
  AOI22_X1 U9958 ( .A1(n9136), .A2(n8599), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        n4309), .ZN(n8561) );
  OAI21_X1 U9959 ( .B1(n9625), .B2(n9101), .A(n8561), .ZN(n8562) );
  AOI21_X1 U9960 ( .B1(n9608), .B2(n8962), .A(n8562), .ZN(n8563) );
  OAI211_X1 U9961 ( .C1(n4462), .C2(n8637), .A(n8564), .B(n8563), .ZN(P1_U3223) );
  INV_X1 U9962 ( .A(n8566), .ZN(n8567) );
  AOI21_X1 U9963 ( .B1(n8565), .B2(n8568), .A(n8567), .ZN(n8573) );
  NAND2_X1 U9964 ( .A1(n9608), .A2(n9222), .ZN(n8569) );
  NAND2_X1 U9965 ( .A1(n4309), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9714) );
  OAI211_X1 U9966 ( .C1(n9247), .C2(n9611), .A(n8569), .B(n9714), .ZN(n8570)
         );
  AOI21_X1 U9967 ( .B1(n8634), .B2(n9256), .A(n8570), .ZN(n8572) );
  NAND2_X1 U9968 ( .A1(n9336), .A2(n8611), .ZN(n8571) );
  OAI211_X1 U9969 ( .C1(n8573), .C2(n9618), .A(n8572), .B(n8571), .ZN(P1_U3224) );
  OAI21_X1 U9970 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n8577) );
  NAND2_X1 U9971 ( .A1(n8577), .A2(n8626), .ZN(n8582) );
  INV_X1 U9972 ( .A(n9197), .ZN(n9235) );
  NAND2_X1 U9973 ( .A1(n9235), .A2(n9608), .ZN(n8578) );
  NAND2_X1 U9974 ( .A1(n4309), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9732) );
  OAI211_X1 U9975 ( .C1(n8579), .C2(n9611), .A(n8578), .B(n9732), .ZN(n8580)
         );
  AOI21_X1 U9976 ( .B1(n8634), .B2(n9228), .A(n8580), .ZN(n8581) );
  OAI211_X1 U9977 ( .C1(n4455), .C2(n8637), .A(n8582), .B(n8581), .ZN(P1_U3226) );
  OAI21_X1 U9978 ( .B1(n8585), .B2(n8584), .A(n8583), .ZN(n8586) );
  NAND2_X1 U9979 ( .A1(n8586), .A2(n8626), .ZN(n8590) );
  AOI22_X1 U9980 ( .A1(n8963), .A2(n8599), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        n4309), .ZN(n8587) );
  OAI21_X1 U9981 ( .B1(n9116), .B2(n8630), .A(n8587), .ZN(n8588) );
  AOI21_X1 U9982 ( .B1(n9119), .B2(n8634), .A(n8588), .ZN(n8589) );
  OAI211_X1 U9983 ( .C1(n9122), .C2(n8637), .A(n8590), .B(n8589), .ZN(P1_U3227) );
  AND3_X1 U9984 ( .A1(n8593), .A2(n8592), .A3(n8591), .ZN(n8594) );
  OAI21_X1 U9985 ( .B1(n8595), .B2(n8594), .A(n8626), .ZN(n8601) );
  OAI22_X1 U9986 ( .A1(n8630), .A2(n9183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8596), .ZN(n8598) );
  NOR2_X1 U9987 ( .A1(n9625), .A2(n9185), .ZN(n8597) );
  AOI211_X1 U9988 ( .C1(n8599), .C2(n9221), .A(n8598), .B(n8597), .ZN(n8600)
         );
  OAI211_X1 U9989 ( .C1(n9189), .C2(n8637), .A(n8601), .B(n8600), .ZN(P1_U3231) );
  INV_X1 U9990 ( .A(n8602), .ZN(n8603) );
  NOR2_X1 U9991 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  XNOR2_X1 U9992 ( .A(n8606), .B(n8605), .ZN(n8613) );
  OAI22_X1 U9993 ( .A1(n9183), .A2(n9611), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8607), .ZN(n8608) );
  AOI21_X1 U9994 ( .B1(n9608), .B2(n8963), .A(n8608), .ZN(n8609) );
  OAI21_X1 U9995 ( .B1(n9625), .B2(n9146), .A(n8609), .ZN(n8610) );
  AOI21_X1 U9996 ( .B1(n9305), .B2(n8611), .A(n8610), .ZN(n8612) );
  OAI21_X1 U9997 ( .B1(n8613), .B2(n9618), .A(n8612), .ZN(P1_U3233) );
  INV_X1 U9998 ( .A(n8614), .ZN(n8618) );
  AOI21_X1 U9999 ( .B1(n8618), .B2(n8615), .A(n8616), .ZN(n8617) );
  AOI21_X1 U10000 ( .B1(n8537), .B2(n8618), .A(n8617), .ZN(n8623) );
  NAND2_X1 U10001 ( .A1(n9221), .A2(n9608), .ZN(n8619) );
  NAND2_X1 U10002 ( .A1(n4309), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9749) );
  OAI211_X1 U10003 ( .C1(n9249), .C2(n9611), .A(n8619), .B(n9749), .ZN(n8621)
         );
  NOR2_X1 U10004 ( .A1(n9216), .A2(n8637), .ZN(n8620) );
  AOI211_X1 U10005 ( .C1(n9214), .C2(n8634), .A(n8621), .B(n8620), .ZN(n8622)
         );
  OAI21_X1 U10006 ( .B1(n8623), .B2(n9618), .A(n8622), .ZN(P1_U3236) );
  AND2_X1 U10007 ( .A1(n8625), .A2(n8624), .ZN(n8628) );
  OAI211_X1 U10008 ( .C1(n8628), .C2(n8627), .A(n8626), .B(n8516), .ZN(n8636)
         );
  OAI22_X1 U10009 ( .A1(n9116), .A2(n9611), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8629), .ZN(n8633) );
  NOR2_X1 U10010 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  AOI211_X1 U10011 ( .C1(n9083), .C2(n8634), .A(n8633), .B(n8632), .ZN(n8635)
         );
  OAI211_X1 U10012 ( .C1(n9085), .C2(n8637), .A(n8636), .B(n8635), .ZN(
        P1_U3238) );
  NAND2_X1 U10013 ( .A1(n8638), .A2(n8645), .ZN(n8641) );
  NAND2_X1 U10014 ( .A1(n8639), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8640) );
  NOR2_X1 U10015 ( .A1(n9267), .A2(n9072), .ZN(n8658) );
  NAND2_X1 U10016 ( .A1(n5916), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10017 ( .A1(n8649), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U10018 ( .A1(n8650), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8642) );
  NAND3_X1 U10019 ( .A1(n8644), .A2(n8643), .A3(n8642), .ZN(n9027) );
  NAND2_X1 U10020 ( .A1(n8646), .A2(n8645), .ZN(n8648) );
  INV_X1 U10021 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9370) );
  OR2_X1 U10022 ( .A1(n5927), .A2(n9370), .ZN(n8647) );
  NAND2_X1 U10023 ( .A1(n5916), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U10024 ( .A1(n8649), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10025 ( .A1(n8650), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8651) );
  AND3_X1 U10026 ( .A1(n8653), .A2(n8652), .A3(n8651), .ZN(n9047) );
  OR2_X1 U10027 ( .A1(n9031), .A2(n9047), .ZN(n8790) );
  INV_X1 U10028 ( .A(n8782), .ZN(n8908) );
  INV_X1 U10029 ( .A(n9267), .ZN(n9055) );
  AND2_X1 U10030 ( .A1(n8928), .A2(n8659), .ZN(n8859) );
  OAI21_X1 U10031 ( .B1(n8661), .B2(n8660), .A(n8859), .ZN(n8662) );
  NAND2_X1 U10032 ( .A1(n8662), .A2(n8839), .ZN(n8670) );
  NAND2_X1 U10033 ( .A1(n8664), .A2(n8663), .ZN(n8849) );
  AOI21_X1 U10034 ( .B1(n8665), .B2(n8854), .A(n8849), .ZN(n8667) );
  NAND2_X1 U10035 ( .A1(n8803), .A2(n8853), .ZN(n8666) );
  OAI211_X1 U10036 ( .C1(n8667), .C2(n8666), .A(n8839), .B(n8850), .ZN(n8668)
         );
  NAND2_X1 U10037 ( .A1(n8668), .A2(n8928), .ZN(n8669) );
  INV_X1 U10038 ( .A(n8781), .ZN(n8775) );
  MUX2_X1 U10039 ( .A(n8670), .B(n8669), .S(n8775), .Z(n8682) );
  OAI211_X1 U10040 ( .C1(n8682), .C2(n4591), .A(n8671), .B(n8679), .ZN(n8675)
         );
  INV_X1 U10041 ( .A(n8875), .ZN(n8674) );
  INV_X1 U10042 ( .A(n8672), .ZN(n8673) );
  AOI21_X1 U10043 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8678) );
  AND2_X1 U10044 ( .A1(n8691), .A2(n8676), .ZN(n8677) );
  MUX2_X1 U10045 ( .A(n8678), .B(n8677), .S(n8781), .Z(n8698) );
  INV_X1 U10046 ( .A(n8679), .ZN(n8845) );
  OAI211_X1 U10047 ( .C1(n8682), .C2(n8845), .A(n8681), .B(n8680), .ZN(n8686)
         );
  NOR2_X1 U10048 ( .A1(n8683), .A2(n8775), .ZN(n8685) );
  NAND2_X1 U10049 ( .A1(n8842), .A2(n8813), .ZN(n8684) );
  AOI21_X1 U10050 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n8697) );
  NAND2_X1 U10051 ( .A1(n8691), .A2(n8687), .ZN(n8688) );
  NAND2_X1 U10052 ( .A1(n8688), .A2(n8842), .ZN(n8689) );
  NAND2_X1 U10053 ( .A1(n8690), .A2(n8689), .ZN(n8877) );
  NAND2_X1 U10054 ( .A1(n8877), .A2(n8775), .ZN(n8695) );
  NAND2_X1 U10055 ( .A1(n9346), .A2(n8703), .ZN(n8837) );
  NAND2_X1 U10056 ( .A1(n8842), .A2(n8841), .ZN(n8692) );
  NAND3_X1 U10057 ( .A1(n8692), .A2(n8781), .A3(n8691), .ZN(n8693) );
  AND2_X1 U10058 ( .A1(n8876), .A2(n8693), .ZN(n8694) );
  NAND4_X1 U10059 ( .A1(n8879), .A2(n8695), .A3(n8837), .A4(n8694), .ZN(n8696)
         );
  AOI21_X1 U10060 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n8718) );
  NAND2_X1 U10061 ( .A1(n8699), .A2(n8775), .ZN(n8705) );
  INV_X1 U10062 ( .A(n8705), .ZN(n8701) );
  NOR2_X1 U10063 ( .A1(n8966), .A2(n8781), .ZN(n8700) );
  AOI21_X1 U10064 ( .B1(n8707), .B2(n8701), .A(n8700), .ZN(n8711) );
  NAND2_X1 U10065 ( .A1(n9607), .A2(n8781), .ZN(n8704) );
  OAI22_X1 U10066 ( .A1(n8707), .A2(n8704), .B1(n8703), .B2(n8775), .ZN(n8702)
         );
  NAND2_X1 U10067 ( .A1(n8712), .A2(n8702), .ZN(n8710) );
  NOR2_X1 U10068 ( .A1(n8704), .A2(n8703), .ZN(n8708) );
  OAI21_X1 U10069 ( .B1(n8966), .B2(n8705), .A(n8707), .ZN(n8706) );
  OAI21_X1 U10070 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8709) );
  OAI211_X1 U10071 ( .C1(n8712), .C2(n8711), .A(n8710), .B(n8709), .ZN(n8713)
         );
  OR2_X1 U10072 ( .A1(n8818), .A2(n8713), .ZN(n8717) );
  MUX2_X1 U10073 ( .A(n8714), .B(n8883), .S(n8775), .Z(n8715) );
  NOR2_X1 U10074 ( .A1(n9243), .A2(n8715), .ZN(n8716) );
  OAI21_X1 U10075 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8720) );
  MUX2_X1 U10076 ( .A(n8834), .B(n8885), .S(n8781), .Z(n8719) );
  NAND3_X1 U10077 ( .A1(n8720), .A2(n9230), .A3(n8719), .ZN(n8723) );
  AND2_X1 U10078 ( .A1(n8869), .A2(n8835), .ZN(n8721) );
  MUX2_X1 U10079 ( .A(n8867), .B(n8721), .S(n8781), .Z(n8722) );
  NAND2_X1 U10080 ( .A1(n8723), .A2(n8722), .ZN(n8727) );
  NAND3_X1 U10081 ( .A1(n8727), .A2(n8724), .A3(n8728), .ZN(n8725) );
  NAND3_X1 U10082 ( .A1(n8725), .A2(n8796), .A3(n8726), .ZN(n8731) );
  NAND3_X1 U10083 ( .A1(n8727), .A2(n8869), .A3(n8726), .ZN(n8729) );
  AND2_X1 U10084 ( .A1(n9156), .A2(n8728), .ZN(n8863) );
  NAND2_X1 U10085 ( .A1(n8729), .A2(n8863), .ZN(n8730) );
  MUX2_X1 U10086 ( .A(n8731), .B(n8730), .S(n8775), .Z(n8739) );
  NAND3_X1 U10087 ( .A1(n8739), .A2(n8737), .A3(n9156), .ZN(n8732) );
  NAND2_X1 U10088 ( .A1(n8732), .A2(n8734), .ZN(n8733) );
  AOI21_X1 U10089 ( .B1(n8733), .B2(n8794), .A(n8793), .ZN(n8741) );
  AND2_X1 U10090 ( .A1(n8737), .A2(n4580), .ZN(n8736) );
  INV_X1 U10091 ( .A(n8734), .ZN(n8735) );
  OR3_X1 U10092 ( .A1(n8793), .A2(n8736), .A3(n8735), .ZN(n8866) );
  INV_X1 U10093 ( .A(n8866), .ZN(n8738) );
  OAI21_X1 U10094 ( .B1(n8866), .B2(n8737), .A(n8794), .ZN(n8861) );
  AOI21_X1 U10095 ( .B1(n8739), .B2(n8738), .A(n8861), .ZN(n8740) );
  MUX2_X1 U10096 ( .A(n8741), .B(n8740), .S(n8775), .Z(n8752) );
  AND2_X1 U10097 ( .A1(n9122), .A2(n9136), .ZN(n8747) );
  OR2_X1 U10098 ( .A1(n8747), .A2(n8744), .ZN(n8743) );
  INV_X1 U10099 ( .A(n8743), .ZN(n8742) );
  NAND2_X1 U10100 ( .A1(n8742), .A2(n9134), .ZN(n8751) );
  INV_X1 U10101 ( .A(n8747), .ZN(n8870) );
  OAI211_X1 U10102 ( .C1(n8743), .C2(n8862), .A(n9086), .B(n8870), .ZN(n8748)
         );
  INV_X1 U10103 ( .A(n8744), .ZN(n8745) );
  OAI211_X1 U10104 ( .C1(n8747), .C2(n8746), .A(n8758), .B(n8745), .ZN(n8893)
         );
  MUX2_X1 U10105 ( .A(n8748), .B(n8893), .S(n8781), .Z(n8749) );
  INV_X1 U10106 ( .A(n8749), .ZN(n8750) );
  OAI21_X1 U10107 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8764) );
  NOR2_X1 U10108 ( .A1(n8758), .A2(n8962), .ZN(n8753) );
  NOR2_X1 U10109 ( .A1(n8753), .A2(n9283), .ZN(n8755) );
  OR2_X1 U10110 ( .A1(n9283), .A2(n9086), .ZN(n8754) );
  MUX2_X1 U10111 ( .A(n8755), .B(n8754), .S(n8781), .Z(n8757) );
  NAND2_X1 U10112 ( .A1(n8962), .A2(n8781), .ZN(n8756) );
  OAI211_X1 U10113 ( .C1(n8764), .C2(n4850), .A(n8757), .B(n8756), .ZN(n8766)
         );
  NAND2_X1 U10114 ( .A1(n8758), .A2(n8962), .ZN(n8759) );
  NAND2_X1 U10115 ( .A1(n9040), .A2(n8759), .ZN(n8762) );
  NAND2_X1 U10116 ( .A1(n9283), .A2(n9086), .ZN(n8760) );
  NAND2_X1 U10117 ( .A1(n8898), .A2(n8760), .ZN(n8761) );
  MUX2_X1 U10118 ( .A(n8762), .B(n8761), .S(n8781), .Z(n8763) );
  OAI21_X1 U10119 ( .B1(n8764), .B2(n9035), .A(n8763), .ZN(n8765) );
  NAND2_X1 U10120 ( .A1(n8766), .A2(n8765), .ZN(n8769) );
  NAND2_X1 U10121 ( .A1(n9271), .A2(n9049), .ZN(n9042) );
  INV_X1 U10122 ( .A(n9070), .ZN(n8768) );
  MUX2_X1 U10123 ( .A(n8898), .B(n9040), .S(n8781), .Z(n8767) );
  NAND3_X1 U10124 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(n8772) );
  INV_X1 U10125 ( .A(n9047), .ZN(n8961) );
  NAND2_X1 U10126 ( .A1(n8961), .A2(n9027), .ZN(n8770) );
  AND2_X1 U10127 ( .A1(n9031), .A2(n8770), .ZN(n8776) );
  INV_X1 U10128 ( .A(n8776), .ZN(n8903) );
  MUX2_X1 U10129 ( .A(n9042), .B(n8832), .S(n8775), .Z(n8771) );
  NAND3_X1 U10130 ( .A1(n8772), .A2(n8903), .A3(n8771), .ZN(n8784) );
  INV_X1 U10131 ( .A(n9626), .ZN(n8774) );
  INV_X1 U10132 ( .A(n9027), .ZN(n8773) );
  AND2_X1 U10133 ( .A1(n8774), .A2(n8773), .ZN(n8789) );
  NOR3_X1 U10134 ( .A1(n8789), .A2(n8781), .A3(n8903), .ZN(n8780) );
  INV_X1 U10135 ( .A(n9072), .ZN(n8899) );
  NAND3_X1 U10136 ( .A1(n9267), .A2(n8899), .A3(n8775), .ZN(n8778) );
  NAND3_X1 U10137 ( .A1(n9055), .A2(n8781), .A3(n9072), .ZN(n8777) );
  AOI211_X1 U10138 ( .C1(n8778), .C2(n8777), .A(n8776), .B(n8782), .ZN(n8779)
         );
  AOI211_X1 U10139 ( .C1(n8782), .C2(n8781), .A(n8780), .B(n8779), .ZN(n8783)
         );
  OAI21_X1 U10140 ( .B1(n8785), .B2(n8784), .A(n8783), .ZN(n8786) );
  MUX2_X1 U10141 ( .A(n8787), .B(n8956), .S(n8786), .Z(n8788) );
  INV_X1 U10142 ( .A(n8789), .ZN(n8791) );
  NAND2_X1 U10143 ( .A1(n8791), .A2(n8790), .ZN(n8914) );
  INV_X1 U10144 ( .A(n8905), .ZN(n8945) );
  INV_X1 U10145 ( .A(n9134), .ZN(n8825) );
  INV_X1 U10146 ( .A(n8793), .ZN(n8795) );
  INV_X1 U10147 ( .A(n9219), .ZN(n8821) );
  INV_X1 U10148 ( .A(n9243), .ZN(n8820) );
  NOR2_X1 U10149 ( .A1(n8798), .A2(n8797), .ZN(n8802) );
  NAND4_X1 U10150 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n8806)
         );
  NAND2_X1 U10151 ( .A1(n8803), .A2(n4408), .ZN(n8804) );
  NOR3_X1 U10152 ( .A1(n8806), .A2(n8805), .A3(n8804), .ZN(n8811) );
  INV_X1 U10153 ( .A(n8807), .ZN(n8810) );
  AND4_X1 U10154 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(n8812)
         );
  NAND4_X1 U10155 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(n8816)
         );
  NOR3_X1 U10156 ( .A1(n8818), .A2(n8817), .A3(n8816), .ZN(n8819) );
  NAND4_X1 U10157 ( .A1(n8821), .A2(n8820), .A3(n9230), .A4(n8819), .ZN(n8822)
         );
  NOR2_X1 U10158 ( .A1(n8822), .A2(n9194), .ZN(n8823) );
  NAND4_X1 U10159 ( .A1(n9151), .A2(n9159), .A3(n9179), .A4(n8823), .ZN(n8824)
         );
  NOR4_X1 U10160 ( .A1(n9105), .A2(n9114), .A3(n8825), .A4(n8824), .ZN(n8826)
         );
  NAND3_X1 U10161 ( .A1(n8827), .A2(n9089), .A3(n8826), .ZN(n8828) );
  NOR2_X1 U10162 ( .A1(n8828), .A2(n9070), .ZN(n8829) );
  XNOR2_X1 U10163 ( .A(n9267), .B(n9072), .ZN(n9044) );
  NAND2_X1 U10164 ( .A1(n9031), .A2(n9047), .ZN(n8941) );
  NAND4_X1 U10165 ( .A1(n8945), .A2(n8829), .A3(n9044), .A4(n8941), .ZN(n8830)
         );
  OAI21_X1 U10166 ( .B1(n8914), .B2(n8830), .A(n6386), .ZN(n8831) );
  XNOR2_X1 U10167 ( .A(n8831), .B(n9018), .ZN(n8910) );
  OR2_X1 U10168 ( .A1(n9267), .A2(n8899), .ZN(n8833) );
  AND2_X1 U10169 ( .A1(n8833), .A2(n8832), .ZN(n8902) );
  INV_X1 U10170 ( .A(n8902), .ZN(n8939) );
  AND2_X1 U10171 ( .A1(n8835), .A2(n8834), .ZN(n8836) );
  NAND2_X1 U10172 ( .A1(n8869), .A2(n8836), .ZN(n8888) );
  AND2_X1 U10173 ( .A1(n8838), .A2(n8837), .ZN(n8882) );
  INV_X1 U10174 ( .A(n8882), .ZN(n8846) );
  AND3_X1 U10175 ( .A1(n8842), .A2(n8841), .A3(n8840), .ZN(n8843) );
  AND2_X1 U10176 ( .A1(n8876), .A2(n8843), .ZN(n8874) );
  INV_X1 U10177 ( .A(n8874), .ZN(n8844) );
  OR4_X1 U10178 ( .A1(n8846), .A2(n8845), .A3(n4594), .A4(n8844), .ZN(n8847)
         );
  NOR2_X1 U10179 ( .A1(n8888), .A2(n8847), .ZN(n8932) );
  INV_X1 U10180 ( .A(n7299), .ZN(n8852) );
  NAND2_X1 U10181 ( .A1(n8854), .A2(n8848), .ZN(n8923) );
  INV_X1 U10182 ( .A(n8849), .ZN(n8851) );
  AND2_X1 U10183 ( .A1(n8851), .A2(n8850), .ZN(n8926) );
  OAI211_X1 U10184 ( .C1(n8852), .C2(n8923), .A(n8926), .B(n8924), .ZN(n8860)
         );
  INV_X1 U10185 ( .A(n8853), .ZN(n8857) );
  INV_X1 U10186 ( .A(n8854), .ZN(n8856) );
  OAI21_X1 U10187 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8858) );
  NAND3_X1 U10188 ( .A1(n8860), .A2(n8859), .A3(n8858), .ZN(n8890) );
  INV_X1 U10189 ( .A(n8861), .ZN(n8873) );
  OAI21_X1 U10190 ( .B1(n8866), .B2(n8863), .A(n8862), .ZN(n8864) );
  INV_X1 U10191 ( .A(n8864), .ZN(n8872) );
  NOR2_X1 U10192 ( .A1(n8866), .A2(n8865), .ZN(n8891) );
  INV_X1 U10193 ( .A(n8867), .ZN(n8868) );
  NAND3_X1 U10194 ( .A1(n8891), .A2(n8869), .A3(n8868), .ZN(n8871) );
  NAND4_X1 U10195 ( .A1(n8873), .A2(n8872), .A3(n8871), .A4(n8870), .ZN(n8892)
         );
  OAI21_X1 U10196 ( .B1(n4591), .B2(n8875), .A(n8874), .ZN(n8880) );
  NAND2_X1 U10197 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND3_X1 U10198 ( .A1(n8880), .A2(n8879), .A3(n8878), .ZN(n8881) );
  NAND2_X1 U10199 ( .A1(n8882), .A2(n8881), .ZN(n8886) );
  INV_X1 U10200 ( .A(n8883), .ZN(n8884) );
  AND3_X1 U10201 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n8887) );
  NOR2_X1 U10202 ( .A1(n8888), .A2(n8887), .ZN(n8889) );
  OR2_X1 U10203 ( .A1(n8892), .A2(n8889), .ZN(n8934) );
  AOI21_X1 U10204 ( .B1(n8932), .B2(n8890), .A(n8934), .ZN(n8895) );
  NOR2_X1 U10205 ( .A1(n8892), .A2(n8891), .ZN(n8894) );
  OR2_X1 U10206 ( .A1(n8894), .A2(n8893), .ZN(n8936) );
  OAI211_X1 U10207 ( .C1(n8895), .C2(n8936), .A(n8935), .B(n9040), .ZN(n8904)
         );
  NAND2_X1 U10208 ( .A1(n9040), .A2(n8896), .ZN(n8897) );
  NAND3_X1 U10209 ( .A1(n9042), .A2(n8898), .A3(n8897), .ZN(n8901) );
  AND2_X1 U10210 ( .A1(n9267), .A2(n8899), .ZN(n8900) );
  AOI21_X1 U10211 ( .B1(n8902), .B2(n8901), .A(n8900), .ZN(n8942) );
  OAI211_X1 U10212 ( .C1(n8939), .C2(n8904), .A(n8942), .B(n8903), .ZN(n8907)
         );
  AOI211_X1 U10213 ( .C1(n8908), .C2(n8907), .A(n8906), .B(n8905), .ZN(n8909)
         );
  AOI21_X1 U10214 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(n8912) );
  NOR2_X1 U10215 ( .A1(n8913), .A2(n8912), .ZN(n8960) );
  INV_X1 U10216 ( .A(n8914), .ZN(n8944) );
  INV_X1 U10217 ( .A(n8915), .ZN(n8917) );
  NAND2_X1 U10218 ( .A1(n7041), .A2(n7032), .ZN(n8916) );
  NAND3_X1 U10219 ( .A1(n8917), .A2(n6385), .A3(n8916), .ZN(n8918) );
  NAND2_X1 U10220 ( .A1(n8919), .A2(n8918), .ZN(n8921) );
  OAI21_X1 U10221 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n8925) );
  AOI21_X1 U10222 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8930) );
  INV_X1 U10223 ( .A(n8926), .ZN(n8929) );
  OAI211_X1 U10224 ( .C1(n8930), .C2(n8929), .A(n8928), .B(n8927), .ZN(n8931)
         );
  AND2_X1 U10225 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NOR2_X1 U10226 ( .A1(n8934), .A2(n8933), .ZN(n8937) );
  OAI21_X1 U10227 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8938) );
  OR3_X1 U10228 ( .A1(n8939), .A2(n9035), .A3(n8938), .ZN(n8940) );
  NAND3_X1 U10229 ( .A1(n8942), .A2(n8941), .A3(n8940), .ZN(n8943) );
  NAND2_X1 U10230 ( .A1(n8944), .A2(n8943), .ZN(n8946) );
  NAND2_X1 U10231 ( .A1(n8946), .A2(n8945), .ZN(n8950) );
  NAND3_X1 U10232 ( .A1(n8950), .A2(n9018), .A3(n8947), .ZN(n8948) );
  OAI211_X1 U10233 ( .C1(n8950), .C2(n8949), .A(n8948), .B(n8954), .ZN(n8959)
         );
  NOR4_X1 U10234 ( .A1(n8953), .A2(n6423), .A3(n8952), .A4(n8951), .ZN(n8958)
         );
  INV_X1 U10235 ( .A(n8954), .ZN(n8955) );
  OAI21_X1 U10236 ( .B1(n8956), .B2(n8955), .A(P1_B_REG_SCAN_IN), .ZN(n8957)
         );
  OAI22_X1 U10237 ( .A1(n8960), .A2(n8959), .B1(n8958), .B2(n8957), .ZN(
        P1_U3240) );
  MUX2_X1 U10238 ( .A(n9027), .B(P1_DATAO_REG_31__SCAN_IN), .S(n8978), .Z(
        P1_U3586) );
  MUX2_X1 U10239 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8961), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10240 ( .A(n9072), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8978), .Z(
        P1_U3584) );
  MUX2_X1 U10241 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9091), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10242 ( .A(n8962), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8978), .Z(
        P1_U3581) );
  MUX2_X1 U10243 ( .A(n9090), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8978), .Z(
        P1_U3580) );
  MUX2_X1 U10244 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9136), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10245 ( .A(n8963), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8978), .Z(
        P1_U3578) );
  MUX2_X1 U10246 ( .A(n9161), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8978), .Z(
        P1_U3577) );
  MUX2_X1 U10247 ( .A(n8964), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8978), .Z(
        P1_U3576) );
  MUX2_X1 U10248 ( .A(n9162), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8978), .Z(
        P1_U3575) );
  MUX2_X1 U10249 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9221), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10250 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9235), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10251 ( .A(n9222), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8978), .Z(
        P1_U3572) );
  MUX2_X1 U10252 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9233), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10253 ( .A(n8965), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8978), .Z(
        P1_U3570) );
  MUX2_X1 U10254 ( .A(n8966), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8978), .Z(
        P1_U3569) );
  MUX2_X1 U10255 ( .A(n9607), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8978), .Z(
        P1_U3568) );
  MUX2_X1 U10256 ( .A(n8967), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8978), .Z(
        P1_U3567) );
  MUX2_X1 U10257 ( .A(n8968), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8978), .Z(
        P1_U3566) );
  MUX2_X1 U10258 ( .A(n8969), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8978), .Z(
        P1_U3565) );
  MUX2_X1 U10259 ( .A(n8970), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8978), .Z(
        P1_U3564) );
  MUX2_X1 U10260 ( .A(n8971), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8978), .Z(
        P1_U3563) );
  MUX2_X1 U10261 ( .A(n8972), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8978), .Z(
        P1_U3562) );
  MUX2_X1 U10262 ( .A(n8973), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8978), .Z(
        P1_U3561) );
  MUX2_X1 U10263 ( .A(n8974), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8978), .Z(
        P1_U3560) );
  MUX2_X1 U10264 ( .A(n8975), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8978), .Z(
        P1_U3559) );
  MUX2_X1 U10265 ( .A(n8976), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8978), .Z(
        P1_U3558) );
  MUX2_X1 U10266 ( .A(n8977), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8978), .Z(
        P1_U3557) );
  MUX2_X1 U10267 ( .A(n7041), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8978), .Z(
        P1_U3556) );
  MUX2_X1 U10268 ( .A(n6744), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8978), .Z(
        P1_U3555) );
  INV_X1 U10269 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9023) );
  INV_X1 U10270 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8991) );
  OR2_X1 U10271 ( .A1(n9674), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U10272 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9674), .ZN(n8980) );
  NAND2_X1 U10273 ( .A1(n8981), .A2(n8980), .ZN(n9677) );
  NOR2_X1 U10274 ( .A1(n8982), .A2(n9002), .ZN(n8983) );
  INV_X1 U10275 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9691) );
  NOR2_X1 U10276 ( .A1(n9691), .A2(n9692), .ZN(n9690) );
  NOR2_X1 U10277 ( .A1(n8983), .A2(n9690), .ZN(n8984) );
  NOR2_X1 U10278 ( .A1(n8984), .A2(n9004), .ZN(n8985) );
  INV_X1 U10279 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U10280 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9720), .ZN(n8986) );
  OAI21_X1 U10281 ( .B1(n9720), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8986), .ZN(
        n9717) );
  AOI21_X1 U10282 ( .B1(n9720), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9716), .ZN(
        n9728) );
  NAND2_X1 U10283 ( .A1(n9731), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8987) );
  OAI21_X1 U10284 ( .B1(n9731), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8987), .ZN(
        n9729) );
  NOR2_X1 U10285 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  OR2_X1 U10286 ( .A1(n9747), .A2(n8988), .ZN(n8990) );
  INV_X1 U10287 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U10288 ( .A1(n9747), .A2(n8988), .ZN(n8989) );
  AND2_X1 U10289 ( .A1(n8990), .A2(n8989), .ZN(n9744) );
  INV_X1 U10290 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9011) );
  XNOR2_X1 U10291 ( .A(n9747), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9754) );
  INV_X1 U10292 ( .A(n9731), .ZN(n9009) );
  INV_X1 U10293 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9008) );
  XOR2_X1 U10294 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9731), .Z(n9738) );
  INV_X1 U10295 ( .A(n9720), .ZN(n9007) );
  INV_X1 U10296 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9006) );
  XOR2_X1 U10297 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9720), .Z(n9722) );
  INV_X1 U10298 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9001) );
  OR2_X1 U10299 ( .A1(n9674), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8999) );
  NOR2_X1 U10300 ( .A1(n8992), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8993) );
  NOR2_X1 U10301 ( .A1(n8994), .A2(n8993), .ZN(n9682) );
  INV_X1 U10302 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8995) );
  OR2_X1 U10303 ( .A1(n9674), .A2(n8995), .ZN(n8997) );
  NAND2_X1 U10304 ( .A1(n9674), .A2(n8995), .ZN(n8996) );
  AND2_X1 U10305 ( .A1(n8997), .A2(n8996), .ZN(n9681) );
  NOR2_X1 U10306 ( .A1(n9682), .A2(n9681), .ZN(n9683) );
  INV_X1 U10307 ( .A(n9683), .ZN(n8998) );
  NOR2_X1 U10308 ( .A1(n9002), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9000) );
  AOI21_X1 U10309 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9002), .A(n9000), .ZN(
        n9698) );
  NOR2_X1 U10310 ( .A1(n9697), .A2(n9698), .ZN(n9696) );
  AOI21_X1 U10311 ( .B1(n9002), .B2(n9001), .A(n9696), .ZN(n9003) );
  NAND2_X1 U10312 ( .A1(n9708), .A2(n9003), .ZN(n9005) );
  XNOR2_X1 U10313 ( .A(n9004), .B(n9003), .ZN(n9710) );
  NAND2_X1 U10314 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9710), .ZN(n9709) );
  NAND2_X1 U10315 ( .A1(n9005), .A2(n9709), .ZN(n9723) );
  NAND2_X1 U10316 ( .A1(n9722), .A2(n9723), .ZN(n9721) );
  OAI21_X1 U10317 ( .B1(n9007), .B2(n9006), .A(n9721), .ZN(n9737) );
  NAND2_X1 U10318 ( .A1(n9738), .A2(n9737), .ZN(n9735) );
  OAI21_X1 U10319 ( .B1(n9009), .B2(n9008), .A(n9735), .ZN(n9753) );
  NOR2_X1 U10320 ( .A1(n9754), .A2(n9753), .ZN(n9752) );
  AOI21_X1 U10321 ( .B1(n9011), .B2(n9010), .A(n9752), .ZN(n9012) );
  XOR2_X1 U10322 ( .A(n9012), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9013) );
  AOI22_X1 U10323 ( .A1(n9015), .A2(n9746), .B1(n9736), .B2(n9013), .ZN(n9020)
         );
  INV_X1 U10324 ( .A(n9013), .ZN(n9017) );
  NOR2_X1 U10325 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  AOI211_X1 U10326 ( .C1(n9736), .C2(n9017), .A(n9748), .B(n9016), .ZN(n9019)
         );
  MUX2_X1 U10327 ( .A(n9020), .B(n9019), .S(n9018), .Z(n9022) );
  OAI211_X1 U10328 ( .C1(n9023), .C2(n9759), .A(n9022), .B(n9021), .ZN(
        P1_U3260) );
  NAND2_X1 U10329 ( .A1(n9050), .A2(n9644), .ZN(n9024) );
  XNOR2_X1 U10330 ( .A(n9626), .B(n9024), .ZN(n9628) );
  NAND2_X1 U10331 ( .A1(n9628), .A2(n9240), .ZN(n9030) );
  NAND2_X1 U10332 ( .A1(n9025), .A2(P1_B_REG_SCAN_IN), .ZN(n9026) );
  NAND2_X1 U10333 ( .A1(n9234), .A2(n9026), .ZN(n9048) );
  INV_X1 U10334 ( .A(n9048), .ZN(n9028) );
  NAND2_X1 U10335 ( .A1(n9028), .A2(n9027), .ZN(n9643) );
  NOR2_X1 U10336 ( .A1(n9257), .A2(n9643), .ZN(n9032) );
  AOI21_X1 U10337 ( .B1(n9257), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9032), .ZN(
        n9029) );
  OAI211_X1 U10338 ( .C1(n9260), .C2(n9626), .A(n9030), .B(n9029), .ZN(
        P1_U3261) );
  XNOR2_X1 U10339 ( .A(n9050), .B(n9031), .ZN(n9647) );
  NAND2_X1 U10340 ( .A1(n9647), .A2(n9240), .ZN(n9034) );
  AOI21_X1 U10341 ( .B1(n9257), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9032), .ZN(
        n9033) );
  OAI211_X1 U10342 ( .C1(n9644), .C2(n9260), .A(n9034), .B(n9033), .ZN(
        P1_U3262) );
  NAND2_X1 U10343 ( .A1(n9059), .A2(n9038), .ZN(n9039) );
  XNOR2_X1 U10344 ( .A(n9039), .B(n9044), .ZN(n9266) );
  INV_X1 U10345 ( .A(n9266), .ZN(n9058) );
  NAND2_X1 U10346 ( .A1(n9041), .A2(n9040), .ZN(n9069) );
  INV_X1 U10347 ( .A(n9042), .ZN(n9043) );
  NOR2_X1 U10348 ( .A1(n9068), .A2(n9043), .ZN(n9045) );
  XNOR2_X1 U10349 ( .A(n9045), .B(n9044), .ZN(n9046) );
  AOI211_X1 U10350 ( .C1(n9267), .C2(n9062), .A(n9786), .B(n9050), .ZN(n9268)
         );
  NAND2_X1 U10351 ( .A1(n9268), .A2(n9203), .ZN(n9054) );
  INV_X1 U10352 ( .A(n9051), .ZN(n9052) );
  AOI22_X1 U10353 ( .A1(n9052), .A2(n9255), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9205), .ZN(n9053) );
  OAI211_X1 U10354 ( .C1(n9055), .C2(n9260), .A(n9054), .B(n9053), .ZN(n9056)
         );
  AOI21_X1 U10355 ( .B1(n9269), .B2(n9263), .A(n9056), .ZN(n9057) );
  OAI21_X1 U10356 ( .B1(n9058), .B2(n9265), .A(n9057), .ZN(P1_U3355) );
  OR2_X1 U10357 ( .A1(n9060), .A2(n9070), .ZN(n9061) );
  AOI21_X1 U10358 ( .B1(n9271), .B2(n9063), .A(n4463), .ZN(n9272) );
  INV_X1 U10359 ( .A(n9064), .ZN(n9065) );
  AOI22_X1 U10360 ( .A1(n9065), .A2(n9255), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9205), .ZN(n9066) );
  OAI21_X1 U10361 ( .B1(n9067), .B2(n9260), .A(n9066), .ZN(n9078) );
  AOI21_X1 U10362 ( .B1(n9070), .B2(n9069), .A(n9068), .ZN(n9071) );
  INV_X1 U10363 ( .A(n9071), .ZN(n9076) );
  NAND2_X1 U10364 ( .A1(n9072), .A2(n9234), .ZN(n9073) );
  OAI21_X1 U10365 ( .B1(n9265), .B2(n9277), .A(n9079), .ZN(P1_U3263) );
  XNOR2_X1 U10366 ( .A(n9080), .B(n9089), .ZN(n9287) );
  INV_X1 U10367 ( .A(n9099), .ZN(n9082) );
  AOI21_X1 U10368 ( .B1(n9283), .B2(n9082), .A(n9081), .ZN(n9284) );
  AOI22_X1 U10369 ( .A1(n9083), .A2(n9255), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9205), .ZN(n9084) );
  OAI21_X1 U10370 ( .B1(n9085), .B2(n9260), .A(n9084), .ZN(n9094) );
  NAND2_X1 U10371 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  XOR2_X1 U10372 ( .A(n9089), .B(n9088), .Z(n9092) );
  AOI211_X1 U10373 ( .C1(n9240), .C2(n9284), .A(n9094), .B(n9093), .ZN(n9095)
         );
  OAI21_X1 U10374 ( .B1(n9287), .B2(n9265), .A(n9095), .ZN(P1_U3265) );
  OAI21_X1 U10375 ( .B1(n9096), .B2(n9105), .A(n9097), .ZN(n9098) );
  INV_X1 U10376 ( .A(n9098), .ZN(n9292) );
  AOI211_X1 U10377 ( .C1(n9290), .C2(n9117), .A(n9786), .B(n9099), .ZN(n9289)
         );
  NOR2_X1 U10378 ( .A1(n4462), .A2(n9260), .ZN(n9103) );
  OAI22_X1 U10379 ( .A1(n9101), .A2(n9145), .B1(n9100), .B2(n9263), .ZN(n9102)
         );
  AOI211_X1 U10380 ( .C1(n9289), .C2(n9203), .A(n9103), .B(n9102), .ZN(n9110)
         );
  OAI222_X1 U10381 ( .A1(n9250), .A2(n9108), .B1(n9248), .B2(n9107), .C1(n9106), .C2(n9246), .ZN(n9288) );
  NAND2_X1 U10382 ( .A1(n9288), .A2(n9263), .ZN(n9109) );
  OAI211_X1 U10383 ( .C1(n9292), .C2(n9265), .A(n9110), .B(n9109), .ZN(
        P1_U3266) );
  XNOR2_X1 U10384 ( .A(n9111), .B(n9114), .ZN(n9297) );
  AOI21_X1 U10385 ( .B1(n9114), .B2(n9113), .A(n9112), .ZN(n9115) );
  OAI222_X1 U10386 ( .A1(n9250), .A2(n9116), .B1(n9248), .B2(n9153), .C1(n9246), .C2(n9115), .ZN(n9293) );
  INV_X1 U10387 ( .A(n9117), .ZN(n9118) );
  AOI211_X1 U10388 ( .C1(n9295), .C2(n9126), .A(n9786), .B(n9118), .ZN(n9294)
         );
  NAND2_X1 U10389 ( .A1(n9294), .A2(n9203), .ZN(n9121) );
  AOI22_X1 U10390 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(n9257), .B1(n9119), .B2(
        n9255), .ZN(n9120) );
  OAI211_X1 U10391 ( .C1(n9122), .C2(n9260), .A(n9121), .B(n9120), .ZN(n9123)
         );
  AOI21_X1 U10392 ( .B1(n9293), .B2(n9263), .A(n9123), .ZN(n9124) );
  OAI21_X1 U10393 ( .B1(n9297), .B2(n9265), .A(n9124), .ZN(P1_U3267) );
  XNOR2_X1 U10394 ( .A(n9125), .B(n9134), .ZN(n9302) );
  INV_X1 U10395 ( .A(n9143), .ZN(n9128) );
  INV_X1 U10396 ( .A(n9126), .ZN(n9127) );
  AOI21_X1 U10397 ( .B1(n9298), .B2(n9128), .A(n9127), .ZN(n9299) );
  INV_X1 U10398 ( .A(n9129), .ZN(n9130) );
  AOI22_X1 U10399 ( .A1(n9257), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9130), .B2(
        n9255), .ZN(n9131) );
  OAI21_X1 U10400 ( .B1(n9132), .B2(n9260), .A(n9131), .ZN(n9140) );
  OAI211_X1 U10401 ( .C1(n9135), .C2(n9134), .A(n9133), .B(n9237), .ZN(n9138)
         );
  AOI22_X1 U10402 ( .A1(n9136), .A2(n9234), .B1(n9232), .B2(n9161), .ZN(n9137)
         );
  AND2_X1 U10403 ( .A1(n9138), .A2(n9137), .ZN(n9301) );
  NOR2_X1 U10404 ( .A1(n9301), .A2(n9257), .ZN(n9139) );
  AOI211_X1 U10405 ( .C1(n9299), .C2(n9240), .A(n9140), .B(n9139), .ZN(n9141)
         );
  OAI21_X1 U10406 ( .B1(n9302), .B2(n9265), .A(n9141), .ZN(P1_U3268) );
  XOR2_X1 U10407 ( .A(n9151), .B(n9142), .Z(n9307) );
  AOI211_X1 U10408 ( .C1(n9305), .C2(n9165), .A(n9786), .B(n9143), .ZN(n9304)
         );
  NOR2_X1 U10409 ( .A1(n9144), .A2(n9260), .ZN(n9149) );
  OAI22_X1 U10410 ( .A1(n9263), .A2(n9147), .B1(n9146), .B2(n9145), .ZN(n9148)
         );
  AOI211_X1 U10411 ( .C1(n9304), .C2(n9203), .A(n9149), .B(n9148), .ZN(n9155)
         );
  XOR2_X1 U10412 ( .A(n9151), .B(n9150), .Z(n9152) );
  OAI222_X1 U10413 ( .A1(n9250), .A2(n9153), .B1(n9248), .B2(n9183), .C1(n9152), .C2(n9246), .ZN(n9303) );
  NAND2_X1 U10414 ( .A1(n9303), .A2(n9263), .ZN(n9154) );
  OAI211_X1 U10415 ( .C1(n9307), .C2(n9265), .A(n9155), .B(n9154), .ZN(
        P1_U3269) );
  AND2_X1 U10416 ( .A1(n9157), .A2(n9156), .ZN(n9160) );
  OAI21_X1 U10417 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9163) );
  AOI222_X1 U10418 ( .A1(n9237), .A2(n9163), .B1(n9162), .B2(n9232), .C1(n9161), .C2(n9234), .ZN(n9312) );
  INV_X1 U10419 ( .A(n9165), .ZN(n9166) );
  AOI211_X1 U10420 ( .C1(n9310), .C2(n9184), .A(n9786), .B(n9166), .ZN(n9309)
         );
  AOI22_X1 U10421 ( .A1(n9309), .A2(n9168), .B1(n9255), .B2(n9167), .ZN(n9169)
         );
  AND2_X1 U10422 ( .A1(n9312), .A2(n9169), .ZN(n9177) );
  OR2_X1 U10423 ( .A1(n9171), .A2(n9170), .ZN(n9308) );
  NAND3_X1 U10424 ( .A1(n9308), .A2(n9172), .A3(n9173), .ZN(n9176) );
  AOI22_X1 U10425 ( .A1(n9310), .A2(n9174), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9205), .ZN(n9175) );
  OAI211_X1 U10426 ( .C1(n9257), .C2(n9177), .A(n9176), .B(n9175), .ZN(
        P1_U3270) );
  XNOR2_X1 U10427 ( .A(n9178), .B(n9179), .ZN(n9318) );
  XNOR2_X1 U10428 ( .A(n9180), .B(n9179), .ZN(n9181) );
  OAI222_X1 U10429 ( .A1(n9250), .A2(n9183), .B1(n9248), .B2(n9182), .C1(n9181), .C2(n9246), .ZN(n9314) );
  AOI211_X1 U10430 ( .C1(n9316), .C2(n9199), .A(n9786), .B(n9164), .ZN(n9315)
         );
  NAND2_X1 U10431 ( .A1(n9315), .A2(n9203), .ZN(n9188) );
  INV_X1 U10432 ( .A(n9185), .ZN(n9186) );
  AOI22_X1 U10433 ( .A1(n9257), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9186), .B2(
        n9255), .ZN(n9187) );
  OAI211_X1 U10434 ( .C1(n9189), .C2(n9260), .A(n9188), .B(n9187), .ZN(n9190)
         );
  AOI21_X1 U10435 ( .B1(n9314), .B2(n9263), .A(n9190), .ZN(n9191) );
  OAI21_X1 U10436 ( .B1(n9318), .B2(n9265), .A(n9191), .ZN(P1_U3271) );
  XNOR2_X1 U10437 ( .A(n9192), .B(n9194), .ZN(n9323) );
  AOI21_X1 U10438 ( .B1(n9195), .B2(n9194), .A(n9193), .ZN(n9196) );
  OAI222_X1 U10439 ( .A1(n9250), .A2(n9198), .B1(n9248), .B2(n9197), .C1(n9246), .C2(n9196), .ZN(n9321) );
  INV_X1 U10440 ( .A(n9213), .ZN(n9201) );
  INV_X1 U10441 ( .A(n9199), .ZN(n9200) );
  AOI211_X1 U10442 ( .C1(n9202), .C2(n9201), .A(n9786), .B(n9200), .ZN(n9319)
         );
  NAND2_X1 U10443 ( .A1(n9319), .A2(n9203), .ZN(n9207) );
  AOI22_X1 U10444 ( .A1(n9205), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9204), .B2(
        n9255), .ZN(n9206) );
  OAI211_X1 U10445 ( .C1(n9208), .C2(n9260), .A(n9207), .B(n9206), .ZN(n9209)
         );
  AOI21_X1 U10446 ( .B1(n9321), .B2(n9263), .A(n9209), .ZN(n9210) );
  OAI21_X1 U10447 ( .B1(n9323), .B2(n9265), .A(n9210), .ZN(P1_U3272) );
  OAI21_X1 U10448 ( .B1(n9212), .B2(n9219), .A(n9211), .ZN(n9328) );
  AOI21_X1 U10449 ( .B1(n9324), .B2(n4457), .A(n9213), .ZN(n9325) );
  AOI22_X1 U10450 ( .A1(n9257), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9214), .B2(
        n9255), .ZN(n9215) );
  OAI21_X1 U10451 ( .B1(n9216), .B2(n9260), .A(n9215), .ZN(n9225) );
  NAND2_X1 U10452 ( .A1(n9218), .A2(n9217), .ZN(n9220) );
  XNOR2_X1 U10453 ( .A(n9220), .B(n9219), .ZN(n9223) );
  AOI222_X1 U10454 ( .A1(n9237), .A2(n9223), .B1(n9222), .B2(n9232), .C1(n9221), .C2(n9234), .ZN(n9327) );
  NOR2_X1 U10455 ( .A1(n9327), .A2(n9257), .ZN(n9224) );
  AOI211_X1 U10456 ( .C1(n9325), .C2(n9240), .A(n9225), .B(n9224), .ZN(n9226)
         );
  OAI21_X1 U10457 ( .B1(n9328), .B2(n9265), .A(n9226), .ZN(P1_U3273) );
  XNOR2_X1 U10458 ( .A(n4389), .B(n9230), .ZN(n9333) );
  AOI21_X1 U10459 ( .B1(n9329), .B2(n9251), .A(n9227), .ZN(n9330) );
  AOI22_X1 U10460 ( .A1(n9257), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9228), .B2(
        n9255), .ZN(n9229) );
  OAI21_X1 U10461 ( .B1(n4455), .B2(n9260), .A(n9229), .ZN(n9239) );
  XOR2_X1 U10462 ( .A(n9231), .B(n9230), .Z(n9236) );
  AOI222_X1 U10463 ( .A1(n9237), .A2(n9236), .B1(n9235), .B2(n9234), .C1(n9233), .C2(n9232), .ZN(n9332) );
  NOR2_X1 U10464 ( .A1(n9332), .A2(n9257), .ZN(n9238) );
  AOI211_X1 U10465 ( .C1(n9330), .C2(n9240), .A(n9239), .B(n9238), .ZN(n9241)
         );
  OAI21_X1 U10466 ( .B1(n9265), .B2(n9333), .A(n9241), .ZN(P1_U3274) );
  XNOR2_X1 U10467 ( .A(n9242), .B(n9243), .ZN(n9338) );
  XNOR2_X1 U10468 ( .A(n9244), .B(n9243), .ZN(n9245) );
  OAI222_X1 U10469 ( .A1(n9250), .A2(n9249), .B1(n9248), .B2(n9247), .C1(n9246), .C2(n9245), .ZN(n9334) );
  INV_X1 U10470 ( .A(n9336), .ZN(n9261) );
  INV_X1 U10471 ( .A(n9251), .ZN(n9252) );
  AOI211_X1 U10472 ( .C1(n9336), .C2(n9253), .A(n9786), .B(n9252), .ZN(n9335)
         );
  NAND2_X1 U10473 ( .A1(n9335), .A2(n9254), .ZN(n9259) );
  AOI22_X1 U10474 ( .A1(n9257), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9256), .B2(
        n9255), .ZN(n9258) );
  OAI211_X1 U10475 ( .C1(n9261), .C2(n9260), .A(n9259), .B(n9258), .ZN(n9262)
         );
  AOI21_X1 U10476 ( .B1(n9334), .B2(n9263), .A(n9262), .ZN(n9264) );
  OAI21_X1 U10477 ( .B1(n9338), .B2(n9265), .A(n9264), .ZN(P1_U3275) );
  MUX2_X1 U10478 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9350), .S(n9802), .Z(
        P1_U3552) );
  AOI22_X1 U10479 ( .A1(n9272), .A2(n9646), .B1(n9347), .B2(n9271), .ZN(n9273)
         );
  OAI21_X1 U10480 ( .B1(n9277), .B2(n9653), .A(n9276), .ZN(n9351) );
  MUX2_X1 U10481 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9351), .S(n9802), .Z(
        P1_U3551) );
  AOI211_X1 U10482 ( .C1(n9347), .C2(n9280), .A(n9279), .B(n9278), .ZN(n9281)
         );
  OAI21_X1 U10483 ( .B1(n9282), .B2(n9653), .A(n9281), .ZN(n9352) );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9352), .S(n9802), .Z(
        P1_U3550) );
  AOI22_X1 U10485 ( .A1(n9284), .A2(n9646), .B1(n9347), .B2(n9283), .ZN(n9285)
         );
  OAI211_X1 U10486 ( .C1(n9287), .C2(n9653), .A(n9286), .B(n9285), .ZN(n9353)
         );
  MUX2_X1 U10487 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9353), .S(n9802), .Z(
        P1_U3549) );
  OAI21_X1 U10488 ( .B1(n9292), .B2(n9653), .A(n9291), .ZN(n9354) );
  MUX2_X1 U10489 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9354), .S(n9802), .Z(
        P1_U3548) );
  AOI211_X1 U10490 ( .C1(n9347), .C2(n9295), .A(n9294), .B(n9293), .ZN(n9296)
         );
  OAI21_X1 U10491 ( .B1(n9297), .B2(n9653), .A(n9296), .ZN(n9355) );
  MUX2_X1 U10492 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9355), .S(n9802), .Z(
        P1_U3547) );
  AOI22_X1 U10493 ( .A1(n9299), .A2(n9646), .B1(n9347), .B2(n9298), .ZN(n9300)
         );
  OAI211_X1 U10494 ( .C1(n9302), .C2(n9653), .A(n9301), .B(n9300), .ZN(n9356)
         );
  MUX2_X1 U10495 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9356), .S(n9802), .Z(
        P1_U3546) );
  AOI211_X1 U10496 ( .C1(n9347), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9306)
         );
  OAI21_X1 U10497 ( .B1(n9307), .B2(n9653), .A(n9306), .ZN(n9357) );
  MUX2_X1 U10498 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9357), .S(n9802), .Z(
        P1_U3545) );
  NAND3_X1 U10499 ( .A1(n9308), .A2(n9172), .A3(n9790), .ZN(n9313) );
  AOI21_X1 U10500 ( .B1(n9347), .B2(n9310), .A(n9309), .ZN(n9311) );
  NAND3_X1 U10501 ( .A1(n9313), .A2(n9312), .A3(n9311), .ZN(n9358) );
  MUX2_X1 U10502 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9358), .S(n9802), .Z(
        P1_U3544) );
  AOI211_X1 U10503 ( .C1(n9347), .C2(n9316), .A(n9315), .B(n9314), .ZN(n9317)
         );
  OAI21_X1 U10504 ( .B1(n9318), .B2(n9653), .A(n9317), .ZN(n9359) );
  MUX2_X1 U10505 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9359), .S(n9802), .Z(
        P1_U3543) );
  NOR3_X1 U10506 ( .A1(n9321), .A2(n9320), .A3(n9319), .ZN(n9322) );
  OAI21_X1 U10507 ( .B1(n9323), .B2(n9653), .A(n9322), .ZN(n9360) );
  MUX2_X1 U10508 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9360), .S(n9802), .Z(
        P1_U3542) );
  AOI22_X1 U10509 ( .A1(n9325), .A2(n9646), .B1(n9347), .B2(n9324), .ZN(n9326)
         );
  OAI211_X1 U10510 ( .C1(n9328), .C2(n9653), .A(n9327), .B(n9326), .ZN(n9361)
         );
  MUX2_X1 U10511 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9361), .S(n9802), .Z(
        P1_U3541) );
  AOI22_X1 U10512 ( .A1(n9330), .A2(n9646), .B1(n9347), .B2(n9329), .ZN(n9331)
         );
  OAI211_X1 U10513 ( .C1(n9333), .C2(n9653), .A(n9332), .B(n9331), .ZN(n9362)
         );
  MUX2_X1 U10514 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9362), .S(n9802), .Z(
        P1_U3540) );
  AOI211_X1 U10515 ( .C1(n9347), .C2(n9336), .A(n9335), .B(n9334), .ZN(n9337)
         );
  OAI21_X1 U10516 ( .B1(n9338), .B2(n9653), .A(n9337), .ZN(n9363) );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9363), .S(n9802), .Z(
        P1_U3539) );
  AOI22_X1 U10518 ( .A1(n9340), .A2(n9646), .B1(n9347), .B2(n9339), .ZN(n9341)
         );
  OAI211_X1 U10519 ( .C1(n9343), .C2(n9653), .A(n9342), .B(n9341), .ZN(n9364)
         );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9364), .S(n9802), .Z(
        P1_U3538) );
  AOI211_X1 U10521 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9348)
         );
  OAI21_X1 U10522 ( .B1(n9653), .B2(n9349), .A(n9348), .ZN(n9365) );
  MUX2_X1 U10523 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9365), .S(n9802), .Z(
        P1_U3537) );
  MUX2_X1 U10524 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9351), .S(n9794), .Z(
        P1_U3519) );
  MUX2_X1 U10525 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9352), .S(n9794), .Z(
        P1_U3518) );
  MUX2_X1 U10526 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9353), .S(n9794), .Z(
        P1_U3517) );
  MUX2_X1 U10527 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9354), .S(n9794), .Z(
        P1_U3516) );
  MUX2_X1 U10528 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9355), .S(n9794), .Z(
        P1_U3515) );
  MUX2_X1 U10529 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9356), .S(n9794), .Z(
        P1_U3514) );
  MUX2_X1 U10530 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9357), .S(n9794), .Z(
        P1_U3513) );
  MUX2_X1 U10531 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9358), .S(n9794), .Z(
        P1_U3512) );
  MUX2_X1 U10532 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9359), .S(n9794), .Z(
        P1_U3511) );
  MUX2_X1 U10533 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9360), .S(n9794), .Z(
        P1_U3510) );
  MUX2_X1 U10534 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9361), .S(n9794), .Z(
        P1_U3508) );
  MUX2_X1 U10535 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9362), .S(n9794), .Z(
        P1_U3505) );
  MUX2_X1 U10536 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9363), .S(n9794), .Z(
        P1_U3502) );
  MUX2_X1 U10537 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9364), .S(n9794), .Z(
        P1_U3499) );
  MUX2_X1 U10538 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9365), .S(n9794), .Z(
        P1_U3496) );
  NOR4_X1 U10539 ( .A1(n5824), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5860), .A4(
        P1_U3084), .ZN(n9366) );
  AOI21_X1 U10540 ( .B1(n9376), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9366), .ZN(
        n9367) );
  OAI21_X1 U10541 ( .B1(n9368), .B2(n9378), .A(n9367), .ZN(P1_U3322) );
  AOI21_X1 U10542 ( .B1(n9376), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9372), .ZN(
        n9373) );
  OAI21_X1 U10543 ( .B1(n9374), .B2(n9378), .A(n9373), .ZN(P1_U3325) );
  AOI21_X1 U10544 ( .B1(n9376), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9375), .ZN(
        n9377) );
  OAI21_X1 U10545 ( .B1(n9379), .B2(n9378), .A(n9377), .ZN(P1_U3326) );
  MUX2_X1 U10546 ( .A(n9380), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10547 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U10548 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9381) );
  AOI21_X1 U10549 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9381), .ZN(n10034) );
  NOR2_X1 U10550 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9382) );
  AOI21_X1 U10551 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9382), .ZN(n10037) );
  NOR2_X1 U10552 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9383) );
  AOI21_X1 U10553 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9383), .ZN(n10040) );
  NOR2_X1 U10554 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9384) );
  AOI21_X1 U10555 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9384), .ZN(n10043) );
  NOR2_X1 U10556 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9385) );
  AOI21_X1 U10557 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9385), .ZN(n10046) );
  NOR2_X1 U10558 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9392) );
  XNOR2_X1 U10559 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10074) );
  NAND2_X1 U10560 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9390) );
  XOR2_X1 U10561 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10072) );
  NAND2_X1 U10562 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9388) );
  XNOR2_X1 U10563 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9386), .ZN(n10060) );
  AOI21_X1 U10564 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10027) );
  INV_X1 U10565 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10031) );
  NAND3_X1 U10566 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10029) );
  OAI21_X1 U10567 ( .B1(n10027), .B2(n10031), .A(n10029), .ZN(n10059) );
  NAND2_X1 U10568 ( .A1(n10060), .A2(n10059), .ZN(n9387) );
  NAND2_X1 U10569 ( .A1(n9388), .A2(n9387), .ZN(n10071) );
  NAND2_X1 U10570 ( .A1(n10072), .A2(n10071), .ZN(n9389) );
  NAND2_X1 U10571 ( .A1(n9390), .A2(n9389), .ZN(n10073) );
  NOR2_X1 U10572 ( .A1(n10074), .A2(n10073), .ZN(n9391) );
  NAND2_X1 U10573 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10069), .ZN(n9393) );
  NOR2_X1 U10574 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10069), .ZN(n10068) );
  AOI21_X1 U10575 ( .B1(n6641), .B2(n9393), .A(n10068), .ZN(n9394) );
  NAND2_X1 U10576 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9394), .ZN(n9396) );
  XOR2_X1 U10577 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9394), .Z(n10067) );
  NAND2_X1 U10578 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10067), .ZN(n9395) );
  NAND2_X1 U10579 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U10580 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9397), .ZN(n9400) );
  XNOR2_X1 U10581 ( .A(n9398), .B(n9397), .ZN(n10066) );
  NAND2_X1 U10582 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10066), .ZN(n9399) );
  NAND2_X1 U10583 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U10584 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9401), .ZN(n9403) );
  XOR2_X1 U10585 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9401), .Z(n10061) );
  NAND2_X1 U10586 ( .A1(n10061), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U10587 ( .A1(n9403), .A2(n9402), .ZN(n9404) );
  AND2_X1 U10588 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9404), .ZN(n9405) );
  XNOR2_X1 U10589 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9404), .ZN(n10058) );
  NOR2_X1 U10590 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  NAND2_X1 U10591 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9406) );
  OAI21_X1 U10592 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9406), .ZN(n10054) );
  NAND2_X1 U10593 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9407) );
  OAI21_X1 U10594 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9407), .ZN(n10051) );
  NOR2_X1 U10595 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9408) );
  AOI21_X1 U10596 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9408), .ZN(n10048) );
  NAND2_X1 U10597 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  NAND2_X1 U10598 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  OAI21_X1 U10599 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10044), .ZN(n10042) );
  NAND2_X1 U10600 ( .A1(n10043), .A2(n10042), .ZN(n10041) );
  OAI21_X1 U10601 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10041), .ZN(n10039) );
  NAND2_X1 U10602 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U10603 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10038), .ZN(n10036) );
  NAND2_X1 U10604 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  OAI21_X1 U10605 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10035), .ZN(n10033) );
  NAND2_X1 U10606 ( .A1(n10034), .A2(n10033), .ZN(n10032) );
  OAI21_X1 U10607 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10032), .ZN(n10063) );
  NOR2_X1 U10608 ( .A1(n10064), .A2(n10063), .ZN(n9409) );
  NAND2_X1 U10609 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  OAI21_X1 U10610 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9409), .A(n10062), .ZN(
        n9594) );
  INV_X1 U10611 ( .A(SI_6_), .ZN(n9592) );
  AOI22_X1 U10612 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        SI_28_), .B2(keyinput_f4), .ZN(n9410) );
  OAI221_X1 U10613 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_28_), .C2(keyinput_f4), .A(n9410), .ZN(n9417) );
  AOI22_X1 U10614 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n9411) );
  OAI221_X1 U10615 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n9411), .ZN(n9416) );
  AOI22_X1 U10616 ( .A1(SI_14_), .A2(keyinput_f18), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n9412) );
  OAI221_X1 U10617 ( .B1(SI_14_), .B2(keyinput_f18), .C1(SI_21_), .C2(
        keyinput_f11), .A(n9412), .ZN(n9415) );
  AOI22_X1 U10618 ( .A1(SI_2_), .A2(keyinput_f30), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n9413) );
  OAI221_X1 U10619 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_17_), .C2(
        keyinput_f15), .A(n9413), .ZN(n9414) );
  NOR4_X1 U10620 ( .A1(n9417), .A2(n9416), .A3(n9415), .A4(n9414), .ZN(n9449)
         );
  XOR2_X1 U10621 ( .A(n9499), .B(keyinput_f6), .Z(n9425) );
  AOI22_X1 U10622 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(n9419), .B2(keyinput_f50), .ZN(n9418) );
  OAI221_X1 U10623 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        n9419), .C2(keyinput_f50), .A(n9418), .ZN(n9424) );
  AOI22_X1 U10624 ( .A1(SI_7_), .A2(keyinput_f25), .B1(SI_10_), .B2(
        keyinput_f22), .ZN(n9420) );
  OAI221_X1 U10625 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_10_), .C2(
        keyinput_f22), .A(n9420), .ZN(n9423) );
  AOI22_X1 U10626 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9421) );
  OAI221_X1 U10627 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9421), .ZN(n9422) );
  NOR4_X1 U10628 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9448)
         );
  INV_X1 U10629 ( .A(SI_15_), .ZN(n9523) );
  AOI22_X1 U10630 ( .A1(n9523), .A2(keyinput_f17), .B1(keyinput_f35), .B2(
        n5122), .ZN(n9426) );
  OAI221_X1 U10631 ( .B1(n9523), .B2(keyinput_f17), .C1(n5122), .C2(
        keyinput_f35), .A(n9426), .ZN(n9435) );
  INV_X1 U10632 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U10633 ( .A1(n9847), .A2(keyinput_f59), .B1(n5394), .B2(
        keyinput_f42), .ZN(n9427) );
  OAI221_X1 U10634 ( .B1(n9847), .B2(keyinput_f59), .C1(n5394), .C2(
        keyinput_f42), .A(n9427), .ZN(n9434) );
  AOI22_X1 U10635 ( .A1(n9429), .A2(keyinput_f21), .B1(keyinput_f34), .B2(
        P2_U3152), .ZN(n9428) );
  OAI221_X1 U10636 ( .B1(n9429), .B2(keyinput_f21), .C1(P2_U3152), .C2(
        keyinput_f34), .A(n9428), .ZN(n9433) );
  XNOR2_X1 U10637 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9431) );
  XNOR2_X1 U10638 ( .A(SI_24_), .B(keyinput_f8), .ZN(n9430) );
  NAND2_X1 U10639 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  NOR4_X1 U10640 ( .A1(n9435), .A2(n9434), .A3(n9433), .A4(n9432), .ZN(n9447)
         );
  AOI22_X1 U10641 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n9436) );
  OAI221_X1 U10642 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n9436), .ZN(n9445) );
  AOI22_X1 U10643 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n9437) );
  OAI221_X1 U10644 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9437), .ZN(n9444) );
  INV_X1 U10645 ( .A(SI_12_), .ZN(n9439) );
  AOI22_X1 U10646 ( .A1(n9439), .A2(keyinput_f20), .B1(n9525), .B2(
        keyinput_f16), .ZN(n9438) );
  OAI221_X1 U10647 ( .B1(n9439), .B2(keyinput_f20), .C1(n9525), .C2(
        keyinput_f16), .A(n9438), .ZN(n9443) );
  AOI22_X1 U10648 ( .A1(n9441), .A2(keyinput_f37), .B1(n9544), .B2(
        keyinput_f48), .ZN(n9440) );
  OAI221_X1 U10649 ( .B1(n9441), .B2(keyinput_f37), .C1(n9544), .C2(
        keyinput_f48), .A(n9440), .ZN(n9442) );
  NOR4_X1 U10650 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9446)
         );
  NAND4_X1 U10651 ( .A1(n9449), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(n9496)
         );
  AOI22_X1 U10652 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(SI_19_), .B2(keyinput_f13), .ZN(n9450) );
  OAI221_X1 U10653 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        SI_19_), .C2(keyinput_f13), .A(n9450), .ZN(n9457) );
  AOI22_X1 U10654 ( .A1(SI_29_), .A2(keyinput_f3), .B1(SI_5_), .B2(
        keyinput_f27), .ZN(n9451) );
  OAI221_X1 U10655 ( .B1(SI_29_), .B2(keyinput_f3), .C1(SI_5_), .C2(
        keyinput_f27), .A(n9451), .ZN(n9456) );
  AOI22_X1 U10656 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n9452) );
  OAI221_X1 U10657 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n9452), .ZN(n9455) );
  AOI22_X1 U10658 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n9453) );
  OAI221_X1 U10659 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n9453), .ZN(n9454) );
  NOR4_X1 U10660 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .ZN(n9494)
         );
  AOI22_X1 U10661 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n9458) );
  OAI221_X1 U10662 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9458), .ZN(n9465) );
  AOI22_X1 U10663 ( .A1(SI_8_), .A2(keyinput_f24), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n9459) );
  OAI221_X1 U10664 ( .B1(SI_8_), .B2(keyinput_f24), .C1(SI_25_), .C2(
        keyinput_f7), .A(n9459), .ZN(n9464) );
  AOI22_X1 U10665 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n9460) );
  OAI221_X1 U10666 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n9460), .ZN(n9463) );
  AOI22_X1 U10667 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(SI_0_), 
        .B2(keyinput_f32), .ZN(n9461) );
  OAI221_X1 U10668 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(SI_0_), .C2(keyinput_f32), .A(n9461), .ZN(n9462) );
  NOR4_X1 U10669 ( .A1(n9465), .A2(n9464), .A3(n9463), .A4(n9462), .ZN(n9493)
         );
  AOI22_X1 U10670 ( .A1(n9527), .A2(keyinput_f62), .B1(keyinput_f61), .B2(
        n9501), .ZN(n9466) );
  OAI221_X1 U10671 ( .B1(n9527), .B2(keyinput_f62), .C1(n9501), .C2(
        keyinput_f61), .A(n9466), .ZN(n9477) );
  AOI22_X1 U10672 ( .A1(n9469), .A2(keyinput_f19), .B1(n9468), .B2(keyinput_f5), .ZN(n9467) );
  OAI221_X1 U10673 ( .B1(n9469), .B2(keyinput_f19), .C1(n9468), .C2(
        keyinput_f5), .A(n9467), .ZN(n9476) );
  AOI22_X1 U10674 ( .A1(n9471), .A2(keyinput_f43), .B1(n7990), .B2(
        keyinput_f45), .ZN(n9470) );
  OAI221_X1 U10675 ( .B1(n9471), .B2(keyinput_f43), .C1(n7990), .C2(
        keyinput_f45), .A(n9470), .ZN(n9475) );
  AOI22_X1 U10676 ( .A1(n9473), .A2(keyinput_f10), .B1(keyinput_f47), .B2(
        n7999), .ZN(n9472) );
  OAI221_X1 U10677 ( .B1(n9473), .B2(keyinput_f10), .C1(n7999), .C2(
        keyinput_f47), .A(n9472), .ZN(n9474) );
  NOR4_X1 U10678 ( .A1(n9477), .A2(n9476), .A3(n9475), .A4(n9474), .ZN(n9492)
         );
  INV_X1 U10679 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9480) );
  AOI22_X1 U10680 ( .A1(n9480), .A2(keyinput_f56), .B1(keyinput_f54), .B2(
        n9479), .ZN(n9478) );
  OAI221_X1 U10681 ( .B1(n9480), .B2(keyinput_f56), .C1(n9479), .C2(
        keyinput_f54), .A(n9478), .ZN(n9490) );
  XNOR2_X1 U10682 ( .A(n9481), .B(keyinput_f41), .ZN(n9489) );
  XNOR2_X1 U10683 ( .A(n9482), .B(keyinput_f29), .ZN(n9488) );
  XNOR2_X1 U10684 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9486) );
  XNOR2_X1 U10685 ( .A(SI_9_), .B(keyinput_f23), .ZN(n9485) );
  XNOR2_X1 U10686 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9484) );
  XNOR2_X1 U10687 ( .A(SI_18_), .B(keyinput_f14), .ZN(n9483) );
  NAND4_X1 U10688 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n9487)
         );
  NOR4_X1 U10689 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n9491)
         );
  NAND4_X1 U10690 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n9495)
         );
  OAI22_X1 U10691 ( .A1(keyinput_f26), .A2(n9592), .B1(n9496), .B2(n9495), 
        .ZN(n9497) );
  AOI21_X1 U10692 ( .B1(keyinput_f26), .B2(n9592), .A(n9497), .ZN(n9591) );
  AOI22_X1 U10693 ( .A1(n9499), .A2(keyinput_g6), .B1(keyinput_g53), .B2(n5150), .ZN(n9498) );
  OAI221_X1 U10694 ( .B1(n9499), .B2(keyinput_g6), .C1(n5150), .C2(
        keyinput_g53), .A(n9498), .ZN(n9510) );
  AOI22_X1 U10695 ( .A1(n9502), .A2(keyinput_g15), .B1(keyinput_g61), .B2(
        n9501), .ZN(n9500) );
  OAI221_X1 U10696 ( .B1(n9502), .B2(keyinput_g15), .C1(n9501), .C2(
        keyinput_g61), .A(n9500), .ZN(n9509) );
  AOI22_X1 U10697 ( .A1(n9911), .A2(keyinput_g40), .B1(n9504), .B2(
        keyinput_g51), .ZN(n9503) );
  OAI221_X1 U10698 ( .B1(n9911), .B2(keyinput_g40), .C1(n9504), .C2(
        keyinput_g51), .A(n9503), .ZN(n9508) );
  XNOR2_X1 U10699 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_g41), .ZN(n9506)
         );
  XNOR2_X1 U10700 ( .A(SI_2_), .B(keyinput_g30), .ZN(n9505) );
  NAND2_X1 U10701 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  NOR4_X1 U10702 ( .A1(n9510), .A2(n9509), .A3(n9508), .A4(n9507), .ZN(n9552)
         );
  AOI22_X1 U10703 ( .A1(SI_1_), .A2(keyinput_g31), .B1(SI_13_), .B2(
        keyinput_g19), .ZN(n9511) );
  OAI221_X1 U10704 ( .B1(SI_1_), .B2(keyinput_g31), .C1(SI_13_), .C2(
        keyinput_g19), .A(n9511), .ZN(n9520) );
  AOI22_X1 U10705 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n9512) );
  OAI221_X1 U10706 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n9512), .ZN(n9519) );
  XNOR2_X1 U10707 ( .A(n9513), .B(keyinput_g12), .ZN(n9517) );
  XNOR2_X1 U10708 ( .A(SI_31_), .B(keyinput_g1), .ZN(n9516) );
  XNOR2_X1 U10709 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9515) );
  XNOR2_X1 U10710 ( .A(SI_3_), .B(keyinput_g29), .ZN(n9514) );
  NAND4_X1 U10711 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n9514), .ZN(n9518)
         );
  NOR3_X1 U10712 ( .A1(n9520), .A2(n9519), .A3(n9518), .ZN(n9551) );
  AOI22_X1 U10713 ( .A1(n9523), .A2(keyinput_g17), .B1(keyinput_g18), .B2(
        n9522), .ZN(n9521) );
  OAI221_X1 U10714 ( .B1(n9523), .B2(keyinput_g17), .C1(n9522), .C2(
        keyinput_g18), .A(n9521), .ZN(n9535) );
  AOI22_X1 U10715 ( .A1(n9525), .A2(keyinput_g16), .B1(keyinput_g58), .B2(
        n9816), .ZN(n9524) );
  OAI221_X1 U10716 ( .B1(n9525), .B2(keyinput_g16), .C1(n9816), .C2(
        keyinput_g58), .A(n9524), .ZN(n9534) );
  INV_X1 U10717 ( .A(SI_28_), .ZN(n9528) );
  AOI22_X1 U10718 ( .A1(n9528), .A2(keyinput_g4), .B1(keyinput_g62), .B2(n9527), .ZN(n9526) );
  OAI221_X1 U10719 ( .B1(n9528), .B2(keyinput_g4), .C1(n9527), .C2(
        keyinput_g62), .A(n9526), .ZN(n9533) );
  INV_X1 U10720 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9531) );
  AOI22_X1 U10721 ( .A1(n9531), .A2(keyinput_g38), .B1(keyinput_g57), .B2(
        n9530), .ZN(n9529) );
  OAI221_X1 U10722 ( .B1(n9531), .B2(keyinput_g38), .C1(n9530), .C2(
        keyinput_g57), .A(n9529), .ZN(n9532) );
  NOR4_X1 U10723 ( .A1(n9535), .A2(n9534), .A3(n9533), .A4(n9532), .ZN(n9550)
         );
  AOI22_X1 U10724 ( .A1(n5394), .A2(keyinput_g42), .B1(n9537), .B2(keyinput_g7), .ZN(n9536) );
  OAI221_X1 U10725 ( .B1(n5394), .B2(keyinput_g42), .C1(n9537), .C2(
        keyinput_g7), .A(n9536), .ZN(n9548) );
  INV_X1 U10726 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9540) );
  INV_X1 U10727 ( .A(SI_19_), .ZN(n9539) );
  AOI22_X1 U10728 ( .A1(n9540), .A2(keyinput_g36), .B1(n9539), .B2(
        keyinput_g13), .ZN(n9538) );
  OAI221_X1 U10729 ( .B1(n9540), .B2(keyinput_g36), .C1(n9539), .C2(
        keyinput_g13), .A(n9538), .ZN(n9547) );
  AOI22_X1 U10730 ( .A1(n5421), .A2(keyinput_g2), .B1(n9542), .B2(keyinput_g39), .ZN(n9541) );
  OAI221_X1 U10731 ( .B1(n5421), .B2(keyinput_g2), .C1(n9542), .C2(
        keyinput_g39), .A(n9541), .ZN(n9546) );
  AOI22_X1 U10732 ( .A1(n9544), .A2(keyinput_g48), .B1(keyinput_g35), .B2(
        n5122), .ZN(n9543) );
  OAI221_X1 U10733 ( .B1(n9544), .B2(keyinput_g48), .C1(n5122), .C2(
        keyinput_g35), .A(n9543), .ZN(n9545) );
  NOR4_X1 U10734 ( .A1(n9548), .A2(n9547), .A3(n9546), .A4(n9545), .ZN(n9549)
         );
  NAND4_X1 U10735 ( .A1(n9552), .A2(n9551), .A3(n9550), .A4(n9549), .ZN(n9589)
         );
  AOI22_X1 U10736 ( .A1(SI_5_), .A2(keyinput_g27), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n9553) );
  OAI221_X1 U10737 ( .B1(SI_5_), .B2(keyinput_g27), .C1(SI_21_), .C2(
        keyinput_g11), .A(n9553), .ZN(n9560) );
  AOI22_X1 U10738 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g43), .ZN(n9554) );
  OAI221_X1 U10739 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P2_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n9554), .ZN(n9559) );
  AOI22_X1 U10740 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n9555) );
  OAI221_X1 U10741 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        SI_12_), .C2(keyinput_g20), .A(n9555), .ZN(n9558) );
  AOI22_X1 U10742 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        SI_18_), .B2(keyinput_g14), .ZN(n9556) );
  OAI221_X1 U10743 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        SI_18_), .C2(keyinput_g14), .A(n9556), .ZN(n9557) );
  NOR4_X1 U10744 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n9587)
         );
  XNOR2_X1 U10745 ( .A(n9847), .B(keyinput_g59), .ZN(n9567) );
  AOI22_X1 U10746 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9561) );
  OAI221_X1 U10747 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n9561), .ZN(n9566) );
  AOI22_X1 U10748 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(SI_11_), .B2(keyinput_g21), .ZN(n9562) );
  OAI221_X1 U10749 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        SI_11_), .C2(keyinput_g21), .A(n9562), .ZN(n9565) );
  AOI22_X1 U10750 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        SI_27_), .B2(keyinput_g5), .ZN(n9563) );
  OAI221_X1 U10751 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        SI_27_), .C2(keyinput_g5), .A(n9563), .ZN(n9564) );
  NOR4_X1 U10752 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n9586)
         );
  AOI22_X1 U10753 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_10_), .B2(keyinput_g22), .ZN(n9568) );
  OAI221_X1 U10754 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        SI_10_), .C2(keyinput_g22), .A(n9568), .ZN(n9575) );
  AOI22_X1 U10755 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(SI_24_), 
        .B2(keyinput_g8), .ZN(n9569) );
  OAI221_X1 U10756 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(SI_24_), 
        .C2(keyinput_g8), .A(n9569), .ZN(n9574) );
  AOI22_X1 U10757 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9570) );
  OAI221_X1 U10758 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9570), .ZN(n9573) );
  AOI22_X1 U10759 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n9571) );
  OAI221_X1 U10760 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        SI_23_), .C2(keyinput_g9), .A(n9571), .ZN(n9572) );
  NOR4_X1 U10761 ( .A1(n9575), .A2(n9574), .A3(n9573), .A4(n9572), .ZN(n9585)
         );
  AOI22_X1 U10762 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n9576) );
  OAI221_X1 U10763 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n9576), .ZN(n9583) );
  AOI22_X1 U10764 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_9_), .B2(
        keyinput_g23), .ZN(n9577) );
  OAI221_X1 U10765 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_9_), .C2(
        keyinput_g23), .A(n9577), .ZN(n9582) );
  AOI22_X1 U10766 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(SI_4_), .B2(keyinput_g28), .ZN(n9578) );
  OAI221_X1 U10767 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        SI_4_), .C2(keyinput_g28), .A(n9578), .ZN(n9581) );
  AOI22_X1 U10768 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9579) );
  OAI221_X1 U10769 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9579), .ZN(n9580) );
  NOR4_X1 U10770 ( .A1(n9583), .A2(n9582), .A3(n9581), .A4(n9580), .ZN(n9584)
         );
  NAND4_X1 U10771 ( .A1(n9587), .A2(n9586), .A3(n9585), .A4(n9584), .ZN(n9588)
         );
  OAI22_X1 U10772 ( .A1(keyinput_g26), .A2(n9592), .B1(n9589), .B2(n9588), 
        .ZN(n9590) );
  AOI211_X1 U10773 ( .C1(keyinput_g26), .C2(n9592), .A(n9591), .B(n9590), .ZN(
        n9593) );
  XNOR2_X1 U10774 ( .A(n9594), .B(n9593), .ZN(n9598) );
  NOR2_X1 U10775 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  XOR2_X1 U10776 ( .A(n9598), .B(n9597), .Z(ADD_1071_U4) );
  OAI21_X1 U10777 ( .B1(n9600), .B2(n9784), .A(n9599), .ZN(n9601) );
  INV_X1 U10778 ( .A(n9601), .ZN(n9602) );
  AND2_X1 U10779 ( .A1(n9603), .A2(n9602), .ZN(n9606) );
  INV_X1 U10780 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10781 ( .A1(n9794), .A2(n9606), .B1(n9604), .B2(n9792), .ZN(
        P1_U3484) );
  AOI22_X1 U10782 ( .A1(n9802), .A2(n9606), .B1(n9605), .B2(n9803), .ZN(
        P1_U3533) );
  NAND2_X1 U10783 ( .A1(n9608), .A2(n9607), .ZN(n9610) );
  OAI211_X1 U10784 ( .C1(n9612), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9613)
         );
  INV_X1 U10785 ( .A(n9613), .ZN(n9623) );
  NOR2_X1 U10786 ( .A1(n9614), .A2(n9784), .ZN(n9655) );
  NAND2_X1 U10787 ( .A1(n9616), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U10788 ( .B1(n9615), .B2(n9619), .A(n9618), .ZN(n9620) );
  AOI21_X1 U10789 ( .B1(n9655), .B2(n9621), .A(n9620), .ZN(n9622) );
  OAI211_X1 U10790 ( .C1(n9625), .C2(n9624), .A(n9623), .B(n9622), .ZN(
        P1_U3222) );
  OAI21_X1 U10791 ( .B1(n9626), .B2(n9784), .A(n9643), .ZN(n9627) );
  AOI21_X1 U10792 ( .B1(n9628), .B2(n9646), .A(n9627), .ZN(n9631) );
  INV_X1 U10793 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U10794 ( .A1(n9802), .A2(n9631), .B1(n9629), .B2(n9803), .ZN(
        P1_U3554) );
  INV_X1 U10795 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9630) );
  AOI22_X1 U10796 ( .A1(n9794), .A2(n9631), .B1(n9630), .B2(n9792), .ZN(
        P1_U3522) );
  OAI21_X1 U10797 ( .B1(n9844), .B2(n9633), .A(n9632), .ZN(n9634) );
  INV_X1 U10798 ( .A(n9634), .ZN(n9641) );
  OAI21_X1 U10799 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9639) );
  AOI22_X1 U10800 ( .A1(n9639), .A2(n9841), .B1(n9859), .B2(n9638), .ZN(n9640)
         );
  OAI211_X1 U10801 ( .C1(n9863), .C2(n9642), .A(n9641), .B(n9640), .ZN(
        P2_U3217) );
  OAI21_X1 U10802 ( .B1(n9644), .B2(n9784), .A(n9643), .ZN(n9645) );
  AOI21_X1 U10803 ( .B1(n9647), .B2(n9646), .A(n9645), .ZN(n9666) );
  INV_X1 U10804 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9648) );
  AOI22_X1 U10805 ( .A1(n9802), .A2(n9666), .B1(n9648), .B2(n9803), .ZN(
        P1_U3553) );
  OAI22_X1 U10806 ( .A1(n9650), .A2(n9786), .B1(n9649), .B2(n9784), .ZN(n9652)
         );
  NOR2_X1 U10807 ( .A1(n9652), .A2(n9651), .ZN(n9668) );
  AOI22_X1 U10808 ( .A1(n9802), .A2(n9668), .B1(n8995), .B2(n9803), .ZN(
        P1_U3536) );
  NOR2_X1 U10809 ( .A1(n9654), .A2(n9653), .ZN(n9658) );
  NOR4_X1 U10810 ( .A1(n9658), .A2(n9657), .A3(n9656), .A4(n9655), .ZN(n9670)
         );
  AOI22_X1 U10811 ( .A1(n9802), .A2(n9670), .B1(n9659), .B2(n9803), .ZN(
        P1_U3535) );
  OAI22_X1 U10812 ( .A1(n9661), .A2(n9786), .B1(n9660), .B2(n9784), .ZN(n9663)
         );
  NOR2_X1 U10813 ( .A1(n9663), .A2(n9662), .ZN(n9672) );
  AOI22_X1 U10814 ( .A1(n9802), .A2(n9672), .B1(n9664), .B2(n9803), .ZN(
        P1_U3534) );
  INV_X1 U10815 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10816 ( .A1(n9794), .A2(n9666), .B1(n9665), .B2(n9792), .ZN(
        P1_U3521) );
  INV_X1 U10817 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10818 ( .A1(n9794), .A2(n9668), .B1(n9667), .B2(n9792), .ZN(
        P1_U3493) );
  INV_X1 U10819 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9669) );
  AOI22_X1 U10820 ( .A1(n9794), .A2(n9670), .B1(n9669), .B2(n9792), .ZN(
        P1_U3490) );
  INV_X1 U10821 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9671) );
  AOI22_X1 U10822 ( .A1(n9794), .A2(n9672), .B1(n9671), .B2(n9792), .ZN(
        P1_U3487) );
  XNOR2_X1 U10823 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10824 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9687) );
  AOI21_X1 U10825 ( .B1(n9748), .B2(n9674), .A(n9673), .ZN(n9680) );
  AOI21_X1 U10826 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  NAND2_X1 U10827 ( .A1(n9746), .A2(n9678), .ZN(n9679) );
  AND2_X1 U10828 ( .A1(n9680), .A2(n9679), .ZN(n9686) );
  AND2_X1 U10829 ( .A1(n9682), .A2(n9681), .ZN(n9684) );
  OAI21_X1 U10830 ( .B1(n9684), .B2(n9683), .A(n9736), .ZN(n9685) );
  OAI211_X1 U10831 ( .C1(n9687), .C2(n9759), .A(n9686), .B(n9685), .ZN(
        P1_U3254) );
  INV_X1 U10832 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9702) );
  AOI21_X1 U10833 ( .B1(n9748), .B2(n9689), .A(n9688), .ZN(n9695) );
  AOI21_X1 U10834 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9693) );
  NAND2_X1 U10835 ( .A1(n9746), .A2(n9693), .ZN(n9694) );
  AND2_X1 U10836 ( .A1(n9695), .A2(n9694), .ZN(n9701) );
  AOI21_X1 U10837 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9699) );
  OR2_X1 U10838 ( .A1(n9756), .A2(n9699), .ZN(n9700) );
  OAI211_X1 U10839 ( .C1(n9702), .C2(n9759), .A(n9701), .B(n9700), .ZN(
        P1_U3255) );
  INV_X1 U10840 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9713) );
  AOI211_X1 U10841 ( .C1(n9705), .C2(n9704), .A(n9703), .B(n9715), .ZN(n9706)
         );
  AOI211_X1 U10842 ( .C1(n9748), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9712)
         );
  OAI211_X1 U10843 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9710), .A(n9736), .B(
        n9709), .ZN(n9711) );
  OAI211_X1 U10844 ( .C1(n9713), .C2(n9759), .A(n9712), .B(n9711), .ZN(
        P1_U3256) );
  INV_X1 U10845 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9726) );
  INV_X1 U10846 ( .A(n9714), .ZN(n9719) );
  AOI211_X1 U10847 ( .C1(n4384), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9718)
         );
  AOI211_X1 U10848 ( .C1(n9748), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9725)
         );
  OAI211_X1 U10849 ( .C1(n9723), .C2(n9722), .A(n9736), .B(n9721), .ZN(n9724)
         );
  OAI211_X1 U10850 ( .C1(n9726), .C2(n9759), .A(n9725), .B(n9724), .ZN(
        P1_U3257) );
  INV_X1 U10851 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9741) );
  AOI21_X1 U10852 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9730) );
  NAND2_X1 U10853 ( .A1(n9746), .A2(n9730), .ZN(n9734) );
  NAND2_X1 U10854 ( .A1(n9748), .A2(n9731), .ZN(n9733) );
  OAI211_X1 U10855 ( .C1(n9738), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9739)
         );
  OAI211_X1 U10856 ( .C1(n9741), .C2(n9759), .A(n9740), .B(n9739), .ZN(
        P1_U3258) );
  AOI21_X1 U10857 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(n9745) );
  NAND2_X1 U10858 ( .A1(n9746), .A2(n9745), .ZN(n9751) );
  NAND2_X1 U10859 ( .A1(n9748), .A2(n9747), .ZN(n9750) );
  AOI21_X1 U10860 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9755) );
  OR2_X1 U10861 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  OAI211_X1 U10862 ( .C1(n10064), .C2(n9759), .A(n9758), .B(n9757), .ZN(
        P1_U3259) );
  AND2_X1 U10863 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9760), .ZN(P1_U3292) );
  AND2_X1 U10864 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9760), .ZN(P1_U3293) );
  AND2_X1 U10865 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9760), .ZN(P1_U3294) );
  AND2_X1 U10866 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9760), .ZN(P1_U3295) );
  AND2_X1 U10867 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9760), .ZN(P1_U3296) );
  AND2_X1 U10868 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9760), .ZN(P1_U3297) );
  AND2_X1 U10869 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9760), .ZN(P1_U3298) );
  AND2_X1 U10870 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9760), .ZN(P1_U3299) );
  AND2_X1 U10871 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9760), .ZN(P1_U3300) );
  AND2_X1 U10872 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9760), .ZN(P1_U3301) );
  AND2_X1 U10873 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9760), .ZN(P1_U3302) );
  AND2_X1 U10874 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9760), .ZN(P1_U3303) );
  AND2_X1 U10875 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9760), .ZN(P1_U3304) );
  AND2_X1 U10876 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9760), .ZN(P1_U3305) );
  AND2_X1 U10877 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9760), .ZN(P1_U3306) );
  AND2_X1 U10878 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9760), .ZN(P1_U3307) );
  AND2_X1 U10879 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9760), .ZN(P1_U3308) );
  AND2_X1 U10880 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9760), .ZN(P1_U3309) );
  AND2_X1 U10881 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9760), .ZN(P1_U3310) );
  AND2_X1 U10882 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9760), .ZN(P1_U3311) );
  AND2_X1 U10883 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9760), .ZN(P1_U3312) );
  AND2_X1 U10884 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9760), .ZN(P1_U3313) );
  AND2_X1 U10885 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9760), .ZN(P1_U3314) );
  AND2_X1 U10886 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9760), .ZN(P1_U3315) );
  AND2_X1 U10887 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9760), .ZN(P1_U3316) );
  AND2_X1 U10888 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9760), .ZN(P1_U3317) );
  AND2_X1 U10889 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9760), .ZN(P1_U3318) );
  AND2_X1 U10890 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9760), .ZN(P1_U3319) );
  AND2_X1 U10891 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9760), .ZN(P1_U3320) );
  AND2_X1 U10892 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9760), .ZN(P1_U3321) );
  OAI22_X1 U10893 ( .A1(n9762), .A2(n9786), .B1(n9761), .B2(n9784), .ZN(n9764)
         );
  NOR2_X1 U10894 ( .A1(n9764), .A2(n9763), .ZN(n9795) );
  INV_X1 U10895 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9765) );
  AOI22_X1 U10896 ( .A1(n9794), .A2(n9795), .B1(n9765), .B2(n9792), .ZN(
        P1_U3463) );
  OAI211_X1 U10897 ( .C1(n9768), .C2(n9784), .A(n9767), .B(n9766), .ZN(n9769)
         );
  AOI211_X1 U10898 ( .C1(n9771), .C2(n9790), .A(n9770), .B(n9769), .ZN(n9797)
         );
  INV_X1 U10899 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10900 ( .A1(n9794), .A2(n9797), .B1(n9772), .B2(n9792), .ZN(
        P1_U3469) );
  OAI22_X1 U10901 ( .A1(n9774), .A2(n9786), .B1(n9773), .B2(n9784), .ZN(n9776)
         );
  NOR2_X1 U10902 ( .A1(n9776), .A2(n9775), .ZN(n9799) );
  INV_X1 U10903 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U10904 ( .A1(n9794), .A2(n9799), .B1(n9777), .B2(n9792), .ZN(
        P1_U3472) );
  OAI211_X1 U10905 ( .C1(n9780), .C2(n9784), .A(n9779), .B(n9778), .ZN(n9781)
         );
  AOI21_X1 U10906 ( .B1(n9782), .B2(n9790), .A(n9781), .ZN(n9801) );
  INV_X1 U10907 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9783) );
  AOI22_X1 U10908 ( .A1(n9794), .A2(n9801), .B1(n9783), .B2(n9792), .ZN(
        P1_U3475) );
  OAI22_X1 U10909 ( .A1(n9787), .A2(n9786), .B1(n9785), .B2(n9784), .ZN(n9789)
         );
  AOI211_X1 U10910 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9788), .ZN(n9805)
         );
  INV_X1 U10911 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10912 ( .A1(n9794), .A2(n9805), .B1(n9793), .B2(n9792), .ZN(
        P1_U3481) );
  AOI22_X1 U10913 ( .A1(n9802), .A2(n9795), .B1(n6522), .B2(n9803), .ZN(
        P1_U3526) );
  AOI22_X1 U10914 ( .A1(n9802), .A2(n9797), .B1(n9796), .B2(n9803), .ZN(
        P1_U3528) );
  AOI22_X1 U10915 ( .A1(n9802), .A2(n9799), .B1(n9798), .B2(n9803), .ZN(
        P1_U3529) );
  AOI22_X1 U10916 ( .A1(n9802), .A2(n9801), .B1(n9800), .B2(n9803), .ZN(
        P1_U3530) );
  AOI22_X1 U10917 ( .A1(n9802), .A2(n9805), .B1(n9804), .B2(n9803), .ZN(
        P1_U3532) );
  INV_X1 U10918 ( .A(n9806), .ZN(n9807) );
  AOI22_X1 U10919 ( .A1(n9851), .A2(n9807), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9814) );
  OAI21_X1 U10920 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9812) );
  AOI22_X1 U10921 ( .A1(n9812), .A2(n9841), .B1(n9859), .B2(n9811), .ZN(n9813)
         );
  OAI211_X1 U10922 ( .C1(n9863), .C2(n9815), .A(n9814), .B(n9813), .ZN(
        P2_U3232) );
  OAI22_X1 U10923 ( .A1(n9844), .A2(n9817), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9816), .ZN(n9818) );
  INV_X1 U10924 ( .A(n9818), .ZN(n9830) );
  INV_X1 U10925 ( .A(n9819), .ZN(n9825) );
  INV_X1 U10926 ( .A(n9820), .ZN(n9822) );
  OAI21_X1 U10927 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9824) );
  OAI21_X1 U10928 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9828) );
  AOI22_X1 U10929 ( .A1(n9828), .A2(n9841), .B1(n9859), .B2(n9827), .ZN(n9829)
         );
  OAI211_X1 U10930 ( .C1(n9863), .C2(n9831), .A(n9830), .B(n9829), .ZN(
        P2_U3238) );
  NAND2_X1 U10931 ( .A1(n9833), .A2(n9832), .ZN(n9837) );
  NAND2_X1 U10932 ( .A1(n9835), .A2(n9834), .ZN(n9836) );
  AND2_X1 U10933 ( .A1(n9837), .A2(n9836), .ZN(n9920) );
  NAND2_X1 U10934 ( .A1(n9839), .A2(n9838), .ZN(n9840) );
  NAND3_X1 U10935 ( .A1(n9841), .A2(n6937), .A3(n9840), .ZN(n9843) );
  NAND2_X1 U10936 ( .A1(n9859), .A2(n9930), .ZN(n9842) );
  OAI211_X1 U10937 ( .C1(n9920), .C2(n9844), .A(n9843), .B(n9842), .ZN(n9845)
         );
  INV_X1 U10938 ( .A(n9845), .ZN(n9846) );
  OAI21_X1 U10939 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(P2_U3239) );
  INV_X1 U10940 ( .A(n9849), .ZN(n9850) );
  AOI22_X1 U10941 ( .A1(n9851), .A2(n9850), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n9861) );
  NAND2_X1 U10942 ( .A1(n9853), .A2(n9852), .ZN(n9855) );
  AOI21_X1 U10943 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9857) );
  AOI21_X1 U10944 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9860) );
  OAI211_X1 U10945 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9860), .ZN(
        P2_U3241) );
  AOI22_X1 U10946 ( .A1(n9865), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9864), .ZN(n9874) );
  AOI22_X1 U10947 ( .A1(n9866), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9873) );
  OAI21_X1 U10948 ( .B1(n9868), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9867), .ZN(
        n9871) );
  NOR2_X1 U10949 ( .A1(n9869), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9870) );
  OAI21_X1 U10950 ( .B1(n9871), .B2(n9870), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9872) );
  OAI211_X1 U10951 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9874), .A(n9873), .B(
        n9872), .ZN(P2_U3245) );
  INV_X1 U10952 ( .A(n9875), .ZN(n9882) );
  AOI222_X1 U10953 ( .A1(n9877), .A2(n9931), .B1(n9876), .B2(n9928), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(n9942), .ZN(n9881) );
  AOI22_X1 U10954 ( .A1(n9879), .A2(n9914), .B1(n9929), .B2(n9878), .ZN(n9880)
         );
  OAI211_X1 U10955 ( .C1(n9942), .C2(n9882), .A(n9881), .B(n9880), .ZN(
        P2_U3286) );
  INV_X1 U10956 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9902) );
  XOR2_X1 U10957 ( .A(n9887), .B(n9883), .Z(n9992) );
  OAI21_X1 U10958 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9990) );
  INV_X1 U10959 ( .A(n9887), .ZN(n9888) );
  NAND3_X1 U10960 ( .A1(n4345), .A2(n9889), .A3(n9888), .ZN(n9890) );
  NAND3_X1 U10961 ( .A1(n9891), .A2(n9922), .A3(n9890), .ZN(n9989) );
  INV_X1 U10962 ( .A(n9892), .ZN(n9985) );
  NOR2_X1 U10963 ( .A1(n9894), .A2(n9893), .ZN(n9895) );
  AOI211_X1 U10964 ( .C1(n9896), .C2(n4315), .A(n9985), .B(n9895), .ZN(n9897)
         );
  OAI211_X1 U10965 ( .C1(n9898), .C2(n9990), .A(n9989), .B(n9897), .ZN(n9899)
         );
  AOI21_X1 U10966 ( .B1(n9992), .B2(n9900), .A(n9899), .ZN(n9901) );
  AOI22_X1 U10967 ( .A1(n9942), .A2(n9902), .B1(n9901), .B2(n9938), .ZN(
        P2_U3291) );
  XNOR2_X1 U10968 ( .A(n9904), .B(n9903), .ZN(n9977) );
  XNOR2_X1 U10969 ( .A(n9905), .B(n9904), .ZN(n9908) );
  OAI21_X1 U10970 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9909) );
  AOI21_X1 U10971 ( .B1(n9910), .B2(n9977), .A(n9909), .ZN(n9974) );
  AOI22_X1 U10972 ( .A1(n9942), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n9928), .B2(
        n9911), .ZN(n9918) );
  AOI21_X1 U10973 ( .B1(n9925), .B2(n4312), .A(n10004), .ZN(n9913) );
  NAND2_X1 U10974 ( .A1(n9913), .A2(n9912), .ZN(n9972) );
  INV_X1 U10975 ( .A(n9972), .ZN(n9915) );
  AOI222_X1 U10976 ( .A1(n4312), .A2(n9931), .B1(n9929), .B2(n9915), .C1(n9977), .C2(n9914), .ZN(n9917) );
  OAI211_X1 U10977 ( .C1(n9942), .C2(n9974), .A(n9918), .B(n9917), .ZN(
        P2_U3293) );
  XNOR2_X1 U10978 ( .A(n9919), .B(n9933), .ZN(n9923) );
  INV_X1 U10979 ( .A(n9920), .ZN(n9921) );
  AOI21_X1 U10980 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9967) );
  OR2_X1 U10981 ( .A1(n9924), .A2(n9968), .ZN(n9927) );
  AND3_X1 U10982 ( .A1(n9927), .A2(n9926), .A3(n9925), .ZN(n9965) );
  AOI22_X1 U10983 ( .A1(n9929), .A2(n9965), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9928), .ZN(n9941) );
  NAND2_X1 U10984 ( .A1(n9931), .A2(n9930), .ZN(n9936) );
  XNOR2_X1 U10985 ( .A(n9933), .B(n9932), .ZN(n9970) );
  NAND2_X1 U10986 ( .A1(n9934), .A2(n9970), .ZN(n9935) );
  OAI211_X1 U10987 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9939)
         );
  INV_X1 U10988 ( .A(n9939), .ZN(n9940) );
  OAI211_X1 U10989 ( .C1(n9942), .C2(n9967), .A(n9941), .B(n9940), .ZN(
        P2_U3294) );
  AND2_X1 U10990 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9947), .ZN(P2_U3297) );
  AND2_X1 U10991 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9947), .ZN(P2_U3298) );
  AND2_X1 U10992 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9947), .ZN(P2_U3299) );
  AND2_X1 U10993 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9947), .ZN(P2_U3300) );
  AND2_X1 U10994 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9947), .ZN(P2_U3301) );
  AND2_X1 U10995 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9947), .ZN(P2_U3302) );
  AND2_X1 U10996 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9947), .ZN(P2_U3303) );
  AND2_X1 U10997 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9947), .ZN(P2_U3304) );
  AND2_X1 U10998 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9947), .ZN(P2_U3305) );
  AND2_X1 U10999 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9947), .ZN(P2_U3306) );
  AND2_X1 U11000 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9947), .ZN(P2_U3307) );
  AND2_X1 U11001 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9947), .ZN(P2_U3308) );
  AND2_X1 U11002 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9947), .ZN(P2_U3309) );
  AND2_X1 U11003 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9947), .ZN(P2_U3310) );
  AND2_X1 U11004 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9947), .ZN(P2_U3311) );
  AND2_X1 U11005 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9947), .ZN(P2_U3312) );
  AND2_X1 U11006 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9947), .ZN(P2_U3313) );
  AND2_X1 U11007 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9947), .ZN(P2_U3314) );
  AND2_X1 U11008 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9947), .ZN(P2_U3315) );
  AND2_X1 U11009 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9947), .ZN(P2_U3316) );
  AND2_X1 U11010 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9947), .ZN(P2_U3317) );
  AND2_X1 U11011 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9947), .ZN(P2_U3318) );
  AND2_X1 U11012 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9947), .ZN(P2_U3319) );
  AND2_X1 U11013 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9947), .ZN(P2_U3320) );
  AND2_X1 U11014 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9947), .ZN(P2_U3321) );
  AND2_X1 U11015 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9947), .ZN(P2_U3322) );
  AND2_X1 U11016 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9947), .ZN(P2_U3323) );
  AND2_X1 U11017 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9947), .ZN(P2_U3324) );
  AND2_X1 U11018 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9947), .ZN(P2_U3325) );
  AND2_X1 U11019 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9947), .ZN(P2_U3326) );
  AOI22_X1 U11020 ( .A1(n9946), .A2(n9949), .B1(n9945), .B2(n9947), .ZN(
        P2_U3437) );
  AOI22_X1 U11021 ( .A1(n9950), .A2(n9949), .B1(n9948), .B2(n9947), .ZN(
        P2_U3438) );
  AOI22_X1 U11022 ( .A1(n9953), .A2(n10008), .B1(n9952), .B2(n9951), .ZN(n9954) );
  AND2_X1 U11023 ( .A1(n9955), .A2(n9954), .ZN(n10014) );
  INV_X1 U11024 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11025 ( .A1(n10012), .A2(n10014), .B1(n9956), .B2(n10010), .ZN(
        P2_U3451) );
  AOI21_X1 U11026 ( .B1(n9987), .B2(n9958), .A(n9957), .ZN(n9960) );
  OAI211_X1 U11027 ( .C1(n9962), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9963)
         );
  INV_X1 U11028 ( .A(n9963), .ZN(n10015) );
  INV_X1 U11029 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11030 ( .A1(n10012), .A2(n10015), .B1(n9964), .B2(n10010), .ZN(
        P2_U3454) );
  INV_X1 U11031 ( .A(n9965), .ZN(n9966) );
  OAI211_X1 U11032 ( .C1(n9968), .C2(n10002), .A(n9967), .B(n9966), .ZN(n9969)
         );
  AOI21_X1 U11033 ( .B1(n10008), .B2(n9970), .A(n9969), .ZN(n10017) );
  INV_X1 U11034 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11035 ( .A1(n10012), .A2(n10017), .B1(n9971), .B2(n10010), .ZN(
        P2_U3457) );
  OAI21_X1 U11036 ( .B1(n9973), .B2(n10002), .A(n9972), .ZN(n9976) );
  INV_X1 U11037 ( .A(n9974), .ZN(n9975) );
  AOI211_X1 U11038 ( .C1(n10000), .C2(n9977), .A(n9976), .B(n9975), .ZN(n10019) );
  INV_X1 U11039 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11040 ( .A1(n10012), .A2(n10019), .B1(n9978), .B2(n10010), .ZN(
        P2_U3460) );
  OAI22_X1 U11041 ( .A1(n9980), .A2(n10004), .B1(n9979), .B2(n10002), .ZN(
        n9982) );
  AOI211_X1 U11042 ( .C1(n10008), .C2(n9983), .A(n9982), .B(n9981), .ZN(n10021) );
  INV_X1 U11043 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11044 ( .A1(n10012), .A2(n10021), .B1(n9984), .B2(n10010), .ZN(
        P2_U3463) );
  AOI21_X1 U11045 ( .B1(n9987), .B2(n4315), .A(n9985), .ZN(n9988) );
  OAI211_X1 U11046 ( .C1(n10004), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9991)
         );
  AOI21_X1 U11047 ( .B1(n9992), .B2(n10008), .A(n9991), .ZN(n10022) );
  INV_X1 U11048 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11049 ( .A1(n10012), .A2(n10022), .B1(n9993), .B2(n10010), .ZN(
        P2_U3466) );
  INV_X1 U11050 ( .A(n9994), .ZN(n9999) );
  OAI22_X1 U11051 ( .A1(n9996), .A2(n10004), .B1(n9995), .B2(n10002), .ZN(
        n9998) );
  AOI211_X1 U11052 ( .C1(n10000), .C2(n9999), .A(n9998), .B(n9997), .ZN(n10023) );
  INV_X1 U11053 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11054 ( .A1(n10012), .A2(n10023), .B1(n10001), .B2(n10010), .ZN(
        P2_U3475) );
  OAI22_X1 U11055 ( .A1(n10005), .A2(n10004), .B1(n10003), .B2(n10002), .ZN(
        n10007) );
  AOI211_X1 U11056 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n10006), .ZN(
        n10025) );
  INV_X1 U11057 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U11058 ( .A1(n10012), .A2(n10025), .B1(n10011), .B2(n10010), .ZN(
        P2_U3487) );
  AOI22_X1 U11059 ( .A1(n10026), .A2(n10014), .B1(n10013), .B2(n10024), .ZN(
        P2_U3520) );
  AOI22_X1 U11060 ( .A1(n10026), .A2(n10015), .B1(n6705), .B2(n10024), .ZN(
        P2_U3521) );
  AOI22_X1 U11061 ( .A1(n10026), .A2(n10017), .B1(n10016), .B2(n10024), .ZN(
        P2_U3522) );
  AOI22_X1 U11062 ( .A1(n10026), .A2(n10019), .B1(n10018), .B2(n10024), .ZN(
        P2_U3523) );
  AOI22_X1 U11063 ( .A1(n10026), .A2(n10021), .B1(n10020), .B2(n10024), .ZN(
        P2_U3524) );
  AOI22_X1 U11064 ( .A1(n10026), .A2(n10022), .B1(n6822), .B2(n10024), .ZN(
        P2_U3525) );
  AOI22_X1 U11065 ( .A1(n10026), .A2(n10023), .B1(n6846), .B2(n10024), .ZN(
        P2_U3528) );
  AOI22_X1 U11066 ( .A1(n10026), .A2(n10025), .B1(n7195), .B2(n10024), .ZN(
        P2_U3532) );
  INV_X1 U11067 ( .A(n10027), .ZN(n10028) );
  NAND2_X1 U11068 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  XOR2_X1 U11069 ( .A(n10031), .B(n10030), .Z(ADD_1071_U5) );
  XOR2_X1 U11070 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11071 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(ADD_1071_U56) );
  OAI21_X1 U11072 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(ADD_1071_U57) );
  OAI21_X1 U11073 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(ADD_1071_U58) );
  OAI21_X1 U11074 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(ADD_1071_U59) );
  OAI21_X1 U11075 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(ADD_1071_U60) );
  OAI21_X1 U11076 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(ADD_1071_U61) );
  AOI21_X1 U11077 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(ADD_1071_U62) );
  AOI21_X1 U11078 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(ADD_1071_U63) );
  AOI21_X1 U11079 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(ADD_1071_U47) );
  XOR2_X1 U11080 ( .A(n10060), .B(n10059), .Z(ADD_1071_U54) );
  XOR2_X1 U11081 ( .A(n10061), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11082 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10065) );
  XNOR2_X1 U11083 ( .A(n10065), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11084 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10066), .Z(ADD_1071_U49) );
  XOR2_X1 U11085 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10067), .Z(ADD_1071_U50) );
  AOI21_X1 U11086 ( .B1(n10069), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10068), .ZN(
        n10070) );
  XOR2_X1 U11087 ( .A(n10070), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11088 ( .A(n10072), .B(n10071), .Z(ADD_1071_U53) );
  XNOR2_X1 U11089 ( .A(n10074), .B(n10073), .ZN(ADD_1071_U52) );
  AND2_X2 U4853 ( .A1(n4317), .A2(n4401), .ZN(n5204) );
  CLKBUF_X1 U4820 ( .A(n5662), .Z(n5769) );
  NAND2_X1 U4822 ( .A1(n7735), .A2(n7734), .ZN(n7733) );
endmodule

