

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837;

  CLKBUF_X3 U2373 ( .A(n4837), .Z(U4043) );
  NAND4_X1 U2374 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n3522)
         );
  BUF_X2 U2375 ( .A(n2925), .Z(n2976) );
  NOR2_X1 U2377 ( .A1(n2901), .A2(n2789), .ZN(n4837) );
  CLKBUF_X2 U2378 ( .A(n3455), .Z(n2132) );
  INV_X1 U2379 ( .A(n3455), .ZN(n3494) );
  INV_X1 U2380 ( .A(n3526), .ZN(n3518) );
  CLKBUF_X2 U2381 ( .A(n2962), .Z(n3499) );
  OR2_X1 U2382 ( .A1(n2888), .A2(n2310), .ZN(n2308) );
  AND2_X1 U2383 ( .A1(n2719), .A2(n3776), .ZN(n3930) );
  NAND2_X1 U2384 ( .A1(n4091), .A2(n3652), .ZN(n4074) );
  OR2_X1 U2385 ( .A1(n2995), .A2(n2994), .ZN(n2289) );
  NAND2_X1 U2386 ( .A1(n2690), .A2(n2733), .ZN(n3074) );
  NAND2_X1 U2387 ( .A1(n2428), .A2(n2146), .ZN(n3808) );
  MUX2_X2 U2388 ( .A(n3791), .B(n3790), .S(n2690), .Z(n3792) );
  XNOR2_X2 U2389 ( .A(n2675), .B(n2676), .ZN(n2690) );
  XNOR2_X2 U2390 ( .A(n3031), .B(n4757), .ZN(n4580) );
  NOR2_X2 U2391 ( .A1(n4568), .A2(n3029), .ZN(n3031) );
  AND2_X1 U2392 ( .A1(n3074), .A2(n2901), .ZN(n3455) );
  XNOR2_X2 U2393 ( .A(n2680), .B(n2679), .ZN(n2733) );
  NAND2_X2 U2394 ( .A1(n2387), .A2(n4493), .ZN(n2422) );
  XNOR2_X2 U2395 ( .A(n2313), .B(IR_REG_2__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U2396 ( .A1(n3884), .A2(n3883), .ZN(n3882) );
  AOI21_X1 U2397 ( .B1(n4074), .B2(n2169), .A(n2347), .ZN(n3984) );
  NAND2_X1 U2398 ( .A1(n3837), .A2(n4630), .ZN(n3838) );
  OAI22_X1 U2399 ( .A1(n3307), .A2(n2213), .B1(n2215), .B2(n2522), .ZN(n3348)
         );
  OR2_X1 U2400 ( .A1(n2422), .A2(n3870), .ZN(n2671) );
  NAND4_X1 U2401 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n3500)
         );
  NOR2_X1 U2402 ( .A1(n3248), .A2(n3247), .ZN(n3250) );
  NOR2_X1 U2403 ( .A1(n2834), .A2(n4724), .ZN(n3620) );
  XNOR2_X1 U2404 ( .A(n2846), .B(n3526), .ZN(n2915) );
  AND2_X2 U2405 ( .A1(n2387), .A2(n2389), .ZN(n2421) );
  AND2_X1 U2406 ( .A1(n4497), .A2(REG2_REG_9__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U2407 ( .A1(n2589), .A2(n2588), .ZN(n2685) );
  AND2_X1 U2408 ( .A1(n2237), .A2(n2500), .ZN(n2236) );
  AND2_X1 U2409 ( .A1(n2368), .A2(n4163), .ZN(n2237) );
  AND2_X1 U2410 ( .A1(n2377), .A2(n2554), .ZN(n2378) );
  AND2_X1 U2411 ( .A1(n2381), .A2(n2369), .ZN(n2368) );
  AND2_X1 U2412 ( .A1(n4765), .A2(n4208), .ZN(n2416) );
  INV_X1 U2413 ( .A(IR_REG_0__SCAN_IN), .ZN(n4765) );
  NOR2_X1 U2414 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2372)
         );
  INV_X1 U2415 ( .A(n2192), .ZN(n2189) );
  AOI21_X1 U2416 ( .B1(n2193), .B2(n2195), .A(n2165), .ZN(n2192) );
  AOI21_X1 U2417 ( .B1(n2207), .B2(n2205), .A(n2204), .ZN(n2203) );
  INV_X1 U2418 ( .A(n2209), .ZN(n2205) );
  NAND2_X1 U2419 ( .A1(n2288), .A2(n2160), .ZN(n2284) );
  NAND2_X1 U2420 ( .A1(n3930), .A2(n3777), .ZN(n2329) );
  NAND2_X1 U2421 ( .A1(n2350), .A2(n3721), .ZN(n2349) );
  INV_X1 U2422 ( .A(n2351), .ZN(n2350) );
  INV_X1 U2423 ( .A(n2219), .ZN(n2217) );
  INV_X1 U2424 ( .A(IR_REG_28__SCAN_IN), .ZN(n2731) );
  INV_X1 U2425 ( .A(IR_REG_27__SCAN_IN), .ZN(n2395) );
  AND4_X1 U2426 ( .A1(n2376), .A2(n2583), .A3(n2375), .A4(n2683), .ZN(n2377)
         );
  NOR2_X1 U2427 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2375)
         );
  AND3_X1 U2428 ( .A1(n4222), .A2(n4147), .A3(n4149), .ZN(n2376) );
  NOR2_X1 U2429 ( .A1(IR_REG_13__SCAN_IN), .A2(n2542), .ZN(n2554) );
  OR2_X1 U2430 ( .A1(n3539), .A2(n2259), .ZN(n2258) );
  OAI21_X1 U2431 ( .B1(n3616), .B2(n2283), .A(n2281), .ZN(n3593) );
  INV_X1 U2432 ( .A(n3074), .ZN(n2290) );
  OR2_X1 U2433 ( .A1(n2422), .A2(n3937), .ZN(n2642) );
  XNOR2_X1 U2434 ( .A(n3011), .B(n3010), .ZN(n2893) );
  AND3_X1 U2435 ( .A1(n2309), .A2(n2308), .A3(n2157), .ZN(n3027) );
  AOI21_X1 U2436 ( .B1(n4552), .B2(REG1_REG_5__SCAN_IN), .A(n4545), .ZN(n3014)
         );
  OAI21_X1 U2437 ( .B1(n3911), .B2(n2225), .A(n2222), .ZN(n3401) );
  AOI21_X1 U2438 ( .B1(n2224), .B2(n2223), .A(n2166), .ZN(n2222) );
  INV_X1 U2439 ( .A(n2230), .ZN(n2223) );
  NAND2_X1 U2440 ( .A1(n2193), .A2(n2139), .ZN(n2190) );
  NAND2_X1 U2441 ( .A1(n2189), .A2(n2139), .ZN(n2188) );
  AOI21_X1 U2442 ( .B1(n3378), .B2(n2547), .A(n2546), .ZN(n3358) );
  NAND2_X1 U2443 ( .A1(n2690), .A2(n2691), .ZN(n4783) );
  AND2_X1 U2444 ( .A1(n2822), .A2(n3794), .ZN(n2691) );
  OAI21_X2 U2445 ( .B1(n2685), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2678) );
  AND3_X1 U2446 ( .A1(n4162), .A2(n2474), .A3(n2476), .ZN(n2374) );
  INV_X1 U2447 ( .A(n3804), .ZN(n3138) );
  AOI22_X1 U2448 ( .A1(n3555), .A2(n3556), .B1(n3454), .B2(n3453), .ZN(n3608)
         );
  INV_X1 U2449 ( .A(n3419), .ZN(n2266) );
  INV_X1 U2450 ( .A(n3833), .ZN(n2301) );
  NOR2_X1 U2451 ( .A1(n2303), .A2(REG2_REG_12__SCAN_IN), .ZN(n2299) );
  NAND2_X1 U2452 ( .A1(n2270), .A2(n2135), .ZN(n2269) );
  INV_X1 U2453 ( .A(n3187), .ZN(n2270) );
  AOI21_X1 U2454 ( .B1(n3192), .B2(n2135), .A(n2155), .ZN(n2268) );
  INV_X1 U2455 ( .A(n3596), .ZN(n2280) );
  OR2_X1 U2456 ( .A1(n2285), .A2(n3486), .ZN(n2283) );
  NAND2_X1 U2457 ( .A1(n2282), .A2(n2287), .ZN(n2281) );
  INV_X1 U2458 ( .A(n2284), .ZN(n2282) );
  INV_X1 U2459 ( .A(n2387), .ZN(n2390) );
  INV_X1 U2460 ( .A(n2328), .ZN(n2327) );
  NOR2_X1 U2461 ( .A1(n3678), .A2(n2149), .ZN(n2328) );
  AND2_X1 U2462 ( .A1(n4000), .A2(n2716), .ZN(n3721) );
  NOR2_X1 U2463 ( .A1(n2712), .A2(n2352), .ZN(n2351) );
  OAI21_X1 U2464 ( .B1(n2707), .B2(n2346), .A(n3359), .ZN(n2345) );
  INV_X1 U2465 ( .A(n3724), .ZN(n2346) );
  INV_X1 U2466 ( .A(n4673), .ZN(n2216) );
  OR2_X1 U2467 ( .A1(n4678), .A2(n2367), .ZN(n3753) );
  INV_X1 U2468 ( .A(n3743), .ZN(n2358) );
  NAND2_X1 U2469 ( .A1(n2455), .A2(n2187), .ZN(n2184) );
  NOR2_X1 U2470 ( .A1(n2158), .A2(n2186), .ZN(n2185) );
  INV_X1 U2471 ( .A(n2187), .ZN(n2186) );
  AND2_X1 U2472 ( .A1(n4090), .A2(n4080), .ZN(n2365) );
  AND2_X1 U2473 ( .A1(n2141), .A2(n2367), .ZN(n2366) );
  NOR2_X1 U2474 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2583)
         );
  INV_X1 U2475 ( .A(IR_REG_9__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U2476 ( .A1(n2276), .A2(n2281), .ZN(n2275) );
  AND2_X1 U2477 ( .A1(n2283), .A2(n2280), .ZN(n2276) );
  NAND2_X1 U2478 ( .A1(n2281), .A2(n2280), .ZN(n2279) );
  NAND2_X1 U2479 ( .A1(n2291), .A2(n2292), .ZN(n3582) );
  AOI21_X1 U2480 ( .B1(n2133), .B2(n2137), .A(n2163), .ZN(n2292) );
  NAND2_X1 U2481 ( .A1(n2284), .A2(n3486), .ZN(n2278) );
  NAND2_X1 U2482 ( .A1(n2160), .A2(n2286), .ZN(n2285) );
  INV_X1 U2483 ( .A(n3617), .ZN(n2286) );
  NAND2_X1 U2484 ( .A1(n2931), .A2(n2930), .ZN(n2932) );
  AND2_X1 U2485 ( .A1(n2733), .A2(n2844), .ZN(n2827) );
  OR2_X1 U2486 ( .A1(n2422), .A2(n3880), .ZN(n2665) );
  XNOR2_X1 U2487 ( .A(n2304), .B(n4498), .ZN(n3820) );
  INV_X1 U2488 ( .A(n4498), .ZN(n2885) );
  OR2_X1 U2489 ( .A1(n4549), .A2(n4307), .ZN(n2310) );
  OR2_X1 U2490 ( .A1(n2311), .A2(n4549), .ZN(n2309) );
  NAND2_X1 U2491 ( .A1(n2252), .A2(n2251), .ZN(n3016) );
  OR2_X1 U2492 ( .A1(n4575), .A2(n4578), .ZN(n2251) );
  NAND2_X1 U2493 ( .A1(n2253), .A2(REG1_REG_7__SCAN_IN), .ZN(n2252) );
  NAND2_X1 U2494 ( .A1(n4575), .A2(n4578), .ZN(n2253) );
  NAND2_X1 U2495 ( .A1(n3241), .A2(n3240), .ZN(n3242) );
  OR2_X1 U2496 ( .A1(n3255), .A2(n3254), .ZN(n3831) );
  NAND2_X1 U2497 ( .A1(n3845), .A2(n2239), .ZN(n3847) );
  NAND2_X1 U2498 ( .A1(n4496), .A2(REG1_REG_11__SCAN_IN), .ZN(n2239) );
  AND2_X1 U2499 ( .A1(n4649), .A2(n3841), .ZN(n4667) );
  INV_X1 U2500 ( .A(n3699), .ZN(n3400) );
  INV_X1 U2501 ( .A(n2228), .ZN(n2227) );
  OAI22_X1 U2502 ( .A1(n2658), .A2(n2229), .B1(n3500), .B2(n2766), .ZN(n2228)
         );
  NAND2_X1 U2503 ( .A1(n2232), .A2(n2653), .ZN(n2229) );
  NOR2_X1 U2504 ( .A1(n2658), .A2(n2231), .ZN(n2230) );
  INV_X1 U2505 ( .A(n2232), .ZN(n2231) );
  OR2_X1 U2506 ( .A1(n3931), .A2(n3914), .ZN(n2232) );
  OAI21_X1 U2507 ( .B1(n3928), .B2(n2646), .A(n2645), .ZN(n3911) );
  OR2_X1 U2508 ( .A1(n3917), .A2(n3482), .ZN(n2645) );
  NAND2_X1 U2509 ( .A1(n2639), .A2(REG3_REG_24__SCAN_IN), .ZN(n2647) );
  INV_X1 U2510 ( .A(n3682), .ZN(n2194) );
  INV_X1 U2511 ( .A(n4016), .ZN(n2199) );
  OAI21_X1 U2512 ( .B1(n4037), .B2(n4042), .A(n2601), .ZN(n4016) );
  OR2_X1 U2513 ( .A1(n4059), .A2(n3647), .ZN(n2601) );
  NOR2_X1 U2514 ( .A1(n2569), .A2(n2211), .ZN(n2209) );
  AOI21_X1 U2515 ( .B1(n3359), .B2(n2209), .A(n2208), .ZN(n2207) );
  NOR2_X1 U2516 ( .A1(n4503), .A2(n4090), .ZN(n2208) );
  OR2_X1 U2517 ( .A1(n4094), .A2(n4093), .ZN(n4091) );
  NOR2_X1 U2518 ( .A1(n3384), .A2(n3366), .ZN(n3365) );
  OR2_X1 U2519 ( .A1(n3383), .A2(n3230), .ZN(n3384) );
  AOI21_X1 U2520 ( .B1(n3348), .B2(n2533), .A(n2532), .ZN(n3378) );
  AND2_X1 U2521 ( .A1(n2221), .A2(n2170), .ZN(n2219) );
  NAND2_X1 U2522 ( .A1(n2703), .A2(n2702), .ZN(n2704) );
  OR2_X1 U2523 ( .A1(n3138), .A2(n3310), .ZN(n2221) );
  OAI21_X1 U2524 ( .B1(n3116), .B2(n2493), .A(n2492), .ZN(n3307) );
  OR2_X1 U2525 ( .A1(n3805), .A2(n3319), .ZN(n2187) );
  OAI21_X1 U2526 ( .B1(n2697), .B2(n2337), .A(n2334), .ZN(n3318) );
  AOI21_X1 U2527 ( .B1(n2338), .B2(n2336), .A(n2335), .ZN(n2334) );
  INV_X1 U2528 ( .A(n2338), .ZN(n2337) );
  INV_X1 U2529 ( .A(n3737), .ZN(n2335) );
  INV_X1 U2530 ( .A(n2733), .ZN(n3717) );
  AND2_X1 U2531 ( .A1(n2722), .A2(n2721), .ZN(n4681) );
  AND2_X1 U2532 ( .A1(n2847), .A2(n4718), .ZN(n4707) );
  INV_X1 U2533 ( .A(IR_REG_20__SCAN_IN), .ZN(n2676) );
  INV_X1 U2534 ( .A(IR_REG_19__SCAN_IN), .ZN(n4222) );
  AND2_X1 U2535 ( .A1(n3717), .A2(n3794), .ZN(n4716) );
  NOR3_X1 U2536 ( .A1(n3922), .A2(n2363), .A3(n2361), .ZN(n4107) );
  OR2_X1 U2537 ( .A1(n3410), .A2(n2364), .ZN(n2363) );
  OR2_X1 U2538 ( .A1(n2766), .A2(n3886), .ZN(n2361) );
  OR2_X1 U2539 ( .A1(n3935), .A2(n3920), .ZN(n3922) );
  NOR2_X1 U2540 ( .A1(n2761), .A2(n3070), .ZN(n2769) );
  OR3_X1 U2541 ( .A1(n2837), .A2(n3068), .A3(n2758), .ZN(n2761) );
  NAND2_X1 U2542 ( .A1(n2687), .A2(IR_REG_31__SCAN_IN), .ZN(n2744) );
  NAND2_X1 U2543 ( .A1(n2748), .A2(n2788), .ZN(n2787) );
  XNOR2_X1 U2544 ( .A(n2385), .B(n2384), .ZN(n2389) );
  NAND2_X1 U2545 ( .A1(n2235), .A2(IR_REG_31__SCAN_IN), .ZN(n2385) );
  NAND2_X1 U2546 ( .A1(n2396), .A2(n2360), .ZN(n2235) );
  NOR2_X1 U2547 ( .A1(n2380), .A2(IR_REG_23__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U2548 ( .A1(n2555), .A2(n2378), .ZN(n2687) );
  AND2_X1 U2549 ( .A1(n2587), .A2(n4147), .ZN(n2588) );
  AND2_X1 U2550 ( .A1(n2332), .A2(n2417), .ZN(n2254) );
  INV_X1 U2551 ( .A(IR_REG_5__SCAN_IN), .ZN(n2332) );
  INV_X1 U2552 ( .A(IR_REG_3__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U2553 ( .A1(n2743), .A2(n2150), .ZN(n2901) );
  INV_X1 U2554 ( .A(n3360), .ZN(n3366) );
  OAI21_X1 U2555 ( .B1(n3493), .B2(n2258), .A(n2256), .ZN(n2262) );
  INV_X1 U2556 ( .A(n2257), .ZN(n2256) );
  OAI21_X1 U2557 ( .B1(n2258), .B2(n2260), .A(n3525), .ZN(n2257) );
  XNOR2_X1 U2558 ( .A(n2915), .B(n2916), .ZN(n2920) );
  NAND2_X1 U2559 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
  INV_X1 U2560 ( .A(n4044), .ZN(n3645) );
  INV_X1 U2561 ( .A(n2844), .ZN(n3794) );
  NAND4_X1 U2562 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n3804)
         );
  OR2_X1 U2563 ( .A1(n2724), .A2(n3018), .ZN(n2497) );
  NAND2_X1 U2564 ( .A1(n2241), .A2(n2243), .ZN(n2240) );
  INV_X1 U2565 ( .A(n4546), .ZN(n2243) );
  XNOR2_X1 U2566 ( .A(n2454), .B(IR_REG_5__SCAN_IN), .ZN(n4552) );
  INV_X1 U2567 ( .A(n2429), .ZN(n2333) );
  NOR2_X1 U2568 ( .A1(n2456), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U2569 ( .A1(n3246), .A2(n3245), .ZN(n3845) );
  XNOR2_X1 U2570 ( .A(n3847), .B(n4606), .ZN(n4603) );
  NAND2_X1 U2571 ( .A1(n2324), .A2(n2323), .ZN(n2322) );
  INV_X1 U2572 ( .A(n4668), .ZN(n2323) );
  INV_X1 U2573 ( .A(n4667), .ZN(n2324) );
  AOI21_X1 U2574 ( .B1(n2249), .B2(n2248), .A(n2247), .ZN(n2246) );
  NAND2_X1 U2575 ( .A1(n2320), .A2(n2247), .ZN(n2319) );
  INV_X1 U2576 ( .A(n4663), .ZN(n2320) );
  NOR2_X1 U2577 ( .A1(n4669), .A2(n4744), .ZN(n2317) );
  INV_X1 U2578 ( .A(n2316), .ZN(n2315) );
  AOI21_X1 U2579 ( .B1(n4671), .B2(ADDR_REG_18__SCAN_IN), .A(n4670), .ZN(n2316) );
  XNOR2_X1 U2580 ( .A(n2678), .B(n4222), .ZN(n3863) );
  AND2_X1 U2581 ( .A1(n2360), .A2(n2384), .ZN(n2359) );
  INV_X1 U2582 ( .A(n3857), .ZN(n4744) );
  NAND2_X1 U2583 ( .A1(n3426), .A2(n2294), .ZN(n2293) );
  INV_X1 U2584 ( .A(n4521), .ZN(n2294) );
  AND2_X1 U2585 ( .A1(n3222), .A2(n3223), .ZN(n3261) );
  OAI21_X1 U2586 ( .B1(n2268), .B2(n2266), .A(n2264), .ZN(n2263) );
  INV_X1 U2587 ( .A(n3418), .ZN(n2264) );
  NAND2_X1 U2588 ( .A1(n4499), .A2(REG2_REG_2__SCAN_IN), .ZN(n2883) );
  AND2_X1 U2589 ( .A1(n4758), .A2(REG2_REG_7__SCAN_IN), .ZN(n3029) );
  AND3_X1 U2590 ( .A1(n2300), .A2(n2302), .A3(n2298), .ZN(n3835) );
  NAND2_X1 U2591 ( .A1(n2301), .A2(n2299), .ZN(n2298) );
  AND2_X1 U2592 ( .A1(n3954), .A2(n2717), .ZN(n3698) );
  INV_X1 U2593 ( .A(n2207), .ZN(n2206) );
  NOR2_X1 U2594 ( .A1(n2339), .A2(n2698), .ZN(n2338) );
  INV_X1 U2595 ( .A(n3733), .ZN(n2339) );
  NAND2_X1 U2596 ( .A1(n2419), .A2(n3633), .ZN(n3727) );
  NOR2_X1 U2597 ( .A1(n3922), .A2(n2766), .ZN(n3878) );
  INV_X1 U2598 ( .A(IR_REG_26__SCAN_IN), .ZN(n2369) );
  INV_X1 U2599 ( .A(IR_REG_23__SCAN_IN), .ZN(n4223) );
  INV_X1 U2600 ( .A(IR_REG_17__SCAN_IN), .ZN(n4147) );
  INV_X1 U2601 ( .A(IR_REG_12__SCAN_IN), .ZN(n2234) );
  INV_X1 U2602 ( .A(IR_REG_10__SCAN_IN), .ZN(n2233) );
  INV_X1 U2603 ( .A(IR_REG_6__SCAN_IN), .ZN(n2474) );
  OR2_X1 U2604 ( .A1(n3548), .A2(n3549), .ZN(n2288) );
  NOR2_X1 U2605 ( .A1(n2261), .A2(n3514), .ZN(n2260) );
  INV_X1 U2606 ( .A(n3573), .ZN(n2261) );
  NOR2_X1 U2607 ( .A1(n3188), .A2(n3187), .ZN(n2267) );
  INV_X1 U2608 ( .A(n3563), .ZN(n3468) );
  AND2_X1 U2609 ( .A1(n2147), .A2(n2134), .ZN(n2297) );
  AND2_X1 U2610 ( .A1(n2297), .A2(n2296), .ZN(n4522) );
  OR2_X1 U2611 ( .A1(n2422), .A2(n3504), .ZN(n2655) );
  OR2_X1 U2612 ( .A1(n2422), .A2(n3576), .ZN(n2649) );
  NAND2_X1 U2613 ( .A1(n3814), .A2(n3813), .ZN(n3812) );
  NAND2_X1 U2614 ( .A1(n2870), .A2(n2871), .ZN(n2884) );
  NOR2_X1 U2615 ( .A1(n3820), .A2(n3821), .ZN(n3819) );
  NOR2_X1 U2616 ( .A1(n3819), .A2(n2887), .ZN(n3022) );
  NOR2_X1 U2617 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  INV_X1 U2618 ( .A(n2304), .ZN(n2886) );
  INV_X1 U2619 ( .A(n3012), .ZN(n2241) );
  NAND2_X1 U2620 ( .A1(n2893), .A2(REG1_REG_4__SCAN_IN), .ZN(n3013) );
  NOR2_X1 U2621 ( .A1(n4558), .A2(n3028), .ZN(n4570) );
  NOR2_X1 U2622 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  OAI21_X1 U2623 ( .B1(n4580), .B2(n2306), .A(n2305), .ZN(n3248) );
  NAND2_X1 U2624 ( .A1(n2307), .A2(REG2_REG_8__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2625 ( .A1(n3032), .A2(n2307), .ZN(n2305) );
  INV_X1 U2626 ( .A(n3033), .ZN(n2307) );
  NOR2_X1 U2627 ( .A1(n4580), .A2(n4581), .ZN(n4579) );
  INV_X1 U2628 ( .A(IR_REG_11__SCAN_IN), .ZN(n4161) );
  OR2_X1 U2629 ( .A1(n2543), .A2(IR_REG_10__SCAN_IN), .ZN(n2518) );
  AND2_X1 U2630 ( .A1(n3831), .A2(n3830), .ZN(n3832) );
  NOR2_X1 U2631 ( .A1(n3832), .A2(n4606), .ZN(n3833) );
  NAND2_X1 U2632 ( .A1(n4613), .A2(n2173), .ZN(n3850) );
  OAI21_X1 U2633 ( .B1(n4748), .B2(n4196), .A(n4627), .ZN(n3852) );
  OR2_X1 U2634 ( .A1(n4652), .A2(n4651), .ZN(n4649) );
  NAND2_X1 U2635 ( .A1(n2250), .A2(n3856), .ZN(n2249) );
  INV_X1 U2636 ( .A(n3854), .ZN(n2250) );
  NAND2_X1 U2637 ( .A1(n4647), .A2(n3856), .ZN(n2248) );
  OAI22_X1 U2638 ( .A1(n3930), .A2(n2153), .B1(n3701), .B2(n2325), .ZN(n3884)
         );
  AND2_X1 U2639 ( .A1(n2326), .A2(n3785), .ZN(n2325) );
  NAND2_X1 U2640 ( .A1(n2328), .A2(n3677), .ZN(n2326) );
  NAND2_X1 U2641 ( .A1(n2329), .A2(n2328), .ZN(n3895) );
  INV_X1 U2642 ( .A(n3500), .ZN(n3915) );
  AND2_X1 U2643 ( .A1(n2329), .A2(n2331), .ZN(n3913) );
  INV_X1 U2644 ( .A(n3698), .ZN(n3971) );
  NAND2_X1 U2645 ( .A1(n2349), .A2(n2348), .ZN(n2347) );
  INV_X1 U2646 ( .A(n3775), .ZN(n2348) );
  NOR2_X1 U2647 ( .A1(n2602), .A2(n4172), .ZN(n2609) );
  NAND2_X1 U2648 ( .A1(n4073), .A2(n2351), .ZN(n4001) );
  AND2_X1 U2649 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2593), .ZN(n2594) );
  NAND2_X1 U2650 ( .A1(n2594), .A2(REG3_REG_18__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U2651 ( .A1(n4073), .A2(n3766), .ZN(n4056) );
  NOR2_X2 U2652 ( .A1(n4501), .A2(n2570), .ZN(n2593) );
  NAND2_X1 U2653 ( .A1(n4074), .A2(n2204), .ZN(n4073) );
  INV_X1 U2654 ( .A(n4519), .ZN(n4090) );
  AOI21_X1 U2655 ( .B1(n2344), .B2(n2346), .A(n2342), .ZN(n2341) );
  INV_X1 U2656 ( .A(n2345), .ZN(n2344) );
  NOR2_X2 U2657 ( .A1(n2548), .A2(n4384), .ZN(n2558) );
  INV_X1 U2658 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4384) );
  NAND2_X1 U2659 ( .A1(n2343), .A2(n3724), .ZN(n3650) );
  NAND2_X1 U2660 ( .A1(n3340), .A2(n2707), .ZN(n2343) );
  NAND2_X1 U2661 ( .A1(n2218), .A2(n2220), .ZN(n2213) );
  AOI21_X1 U2662 ( .B1(n2217), .B2(n2218), .A(n2216), .ZN(n2215) );
  NAND2_X1 U2663 ( .A1(n2512), .A2(REG3_REG_11__SCAN_IN), .ZN(n2524) );
  INV_X1 U2664 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3021) );
  AOI21_X1 U2665 ( .B1(n2357), .B2(n2355), .A(n2354), .ZN(n2353) );
  INV_X1 U2666 ( .A(n2357), .ZN(n2356) );
  INV_X1 U2667 ( .A(n3751), .ZN(n2354) );
  INV_X1 U2668 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2482) );
  INV_X1 U2669 ( .A(n2181), .ZN(n2180) );
  OAI21_X1 U2670 ( .B1(n2158), .B2(n2184), .A(n2466), .ZN(n2181) );
  INV_X1 U2671 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2457) );
  OAI21_X1 U2672 ( .B1(n3318), .B2(n3317), .A(n3749), .ZN(n3057) );
  NAND2_X1 U2673 ( .A1(n2176), .A2(n2138), .ZN(n3326) );
  NAND2_X1 U2674 ( .A1(n3080), .A2(n3733), .ZN(n3144) );
  NAND2_X1 U2675 ( .A1(n2697), .A2(n3078), .ZN(n3080) );
  AND2_X1 U2676 ( .A1(n2827), .A2(n4494), .ZN(n4679) );
  NAND2_X1 U2677 ( .A1(n3727), .A2(n3729), .ZN(n3696) );
  INV_X1 U2678 ( .A(n4722), .ZN(n4696) );
  INV_X1 U2679 ( .A(n4679), .ZN(n4698) );
  INV_X1 U2680 ( .A(n2814), .ZN(n3070) );
  INV_X1 U2681 ( .A(n4695), .ZN(n4675) );
  NAND2_X1 U2682 ( .A1(n3878), .A2(n2362), .ZN(n3403) );
  NOR2_X1 U2683 ( .A1(n3886), .A2(n2364), .ZN(n2362) );
  AND2_X1 U2684 ( .A1(n3878), .A2(n3542), .ZN(n3879) );
  AND2_X1 U2685 ( .A1(n4031), .A2(n2174), .ZN(n3946) );
  NAND2_X1 U2686 ( .A1(n4031), .A2(n2144), .ZN(n3990) );
  NAND2_X1 U2687 ( .A1(n4031), .A2(n4009), .ZN(n4008) );
  AND2_X1 U2688 ( .A1(n3365), .A2(n2143), .ZN(n4039) );
  AND2_X1 U2689 ( .A1(n4039), .A2(n4029), .ZN(n4031) );
  NAND2_X1 U2690 ( .A1(n3365), .A2(n2140), .ZN(n4064) );
  NAND2_X1 U2691 ( .A1(n3365), .A2(n2365), .ZN(n4079) );
  AND2_X1 U2692 ( .A1(n3365), .A2(n4090), .ZN(n4087) );
  AND2_X1 U2693 ( .A1(n3157), .A2(n2171), .ZN(n4686) );
  NAND2_X1 U2694 ( .A1(n3157), .A2(n2141), .ZN(n3309) );
  NAND2_X1 U2695 ( .A1(n3157), .A2(n2366), .ZN(n4687) );
  INV_X1 U2696 ( .A(n3046), .ZN(n3118) );
  NAND2_X1 U2697 ( .A1(n3157), .A2(n3118), .ZN(n3308) );
  AND2_X1 U2698 ( .A1(n3159), .A2(n3165), .ZN(n3157) );
  AND2_X1 U2699 ( .A1(n4702), .A2(n4783), .ZN(n4801) );
  NAND3_X1 U2700 ( .A1(n2138), .A2(n4707), .A3(n2162), .ZN(n3327) );
  NOR2_X1 U2701 ( .A1(n3327), .A2(n3061), .ZN(n3159) );
  NAND2_X1 U2702 ( .A1(n4707), .A2(n3110), .ZN(n4777) );
  INV_X1 U2703 ( .A(n4783), .ZN(n4820) );
  AND2_X1 U2704 ( .A1(n2901), .A2(n4742), .ZN(n2833) );
  AND2_X1 U2705 ( .A1(n2395), .A2(n2731), .ZN(n2360) );
  INV_X1 U2706 ( .A(IR_REG_29__SCAN_IN), .ZN(n2384) );
  AND2_X1 U2707 ( .A1(n2396), .A2(n2395), .ZN(n2730) );
  NAND2_X1 U2708 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2858) );
  INV_X1 U2709 ( .A(n2396), .ZN(n2397) );
  INV_X1 U2710 ( .A(IR_REG_24__SCAN_IN), .ZN(n2737) );
  NOR2_X1 U2711 ( .A1(n2584), .A2(IR_REG_16__SCAN_IN), .ZN(n2587) );
  INV_X1 U2712 ( .A(IR_REG_7__SCAN_IN), .ZN(n2476) );
  NOR2_X1 U2713 ( .A1(n2416), .A2(n2729), .ZN(n2313) );
  XNOR2_X1 U2714 ( .A(n2238), .B(n4208), .ZN(n2873) );
  NAND2_X1 U2715 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2238)
         );
  NAND2_X1 U2716 ( .A1(n2289), .A2(n2152), .ZN(n3043) );
  AOI21_X1 U2717 ( .B1(n3616), .B2(n2277), .A(n2273), .ZN(n2271) );
  NAND2_X1 U2718 ( .A1(n2279), .A2(n2278), .ZN(n2277) );
  NAND2_X1 U2719 ( .A1(n2275), .A2(n2274), .ZN(n2273) );
  OAI21_X1 U2720 ( .B1(n3616), .B2(n2285), .A(n2272), .ZN(n3594) );
  INV_X1 U2721 ( .A(n2278), .ZN(n2272) );
  AND2_X1 U2722 ( .A1(n2937), .A2(n2934), .ZN(n2935) );
  NOR2_X1 U2723 ( .A1(n3616), .A2(n3617), .ZN(n3615) );
  NAND2_X1 U2724 ( .A1(n2904), .A2(STATE_REG_SCAN_IN), .ZN(n4528) );
  INV_X1 U2725 ( .A(n3626), .ZN(n4524) );
  INV_X1 U2726 ( .A(n3620), .ZN(n4518) );
  NAND4_X1 U2727 ( .A1(n2644), .A2(n2643), .A3(n2642), .A4(n2641), .ZN(n3917)
         );
  OR2_X1 U2728 ( .A1(n2724), .A2(n4300), .ZN(n2641) );
  NAND4_X1 U2729 ( .A1(n2635), .A2(n2634), .A3(n2633), .A4(n2632), .ZN(n3974)
         );
  OR2_X1 U2730 ( .A1(n2724), .A2(n2622), .ZN(n2626) );
  NAND4_X1 U2731 ( .A1(n2621), .A2(n2620), .A3(n2619), .A4(n2618), .ZN(n3973)
         );
  NAND4_X1 U2732 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n4044)
         );
  OR2_X1 U2733 ( .A1(n2724), .A2(n4422), .ZN(n2605) );
  NAND4_X1 U2734 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n4059)
         );
  NAND4_X1 U2735 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n4060)
         );
  OR2_X1 U2736 ( .A1(n2724), .A2(n4196), .ZN(n2560) );
  NAND4_X1 U2737 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n3376)
         );
  NAND4_X1 U2738 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(n4678)
         );
  OR2_X1 U2739 ( .A1(n2422), .A2(n3287), .ZN(n2508) );
  NAND4_X1 U2740 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n3120)
         );
  NAND4_X1 U2741 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n3806)
         );
  NAND2_X1 U2742 ( .A1(n3811), .A2(n3810), .ZN(n3809) );
  NAND2_X1 U2743 ( .A1(n2875), .A2(n2876), .ZN(n2890) );
  XNOR2_X1 U2744 ( .A(n2891), .B(n2885), .ZN(n3826) );
  OR2_X1 U2745 ( .A1(n2888), .A2(n4307), .ZN(n2312) );
  NAND2_X1 U2746 ( .A1(n2309), .A2(n2308), .ZN(n4548) );
  AND2_X1 U2747 ( .A1(n3013), .A2(n3012), .ZN(n4547) );
  NOR2_X1 U2748 ( .A1(n4556), .A2(n3015), .ZN(n4575) );
  XNOR2_X1 U2749 ( .A(n3016), .B(n4757), .ZN(n4586) );
  NAND2_X1 U2750 ( .A1(n4586), .A2(REG1_REG_8__SCAN_IN), .ZN(n4585) );
  XNOR2_X1 U2751 ( .A(n3250), .B(n4755), .ZN(n4590) );
  NOR2_X1 U2752 ( .A1(n4590), .A2(n4591), .ZN(n4589) );
  NAND2_X1 U2753 ( .A1(n4594), .A2(n3243), .ZN(n3246) );
  XNOR2_X1 U2754 ( .A(n3832), .B(n4606), .ZN(n4599) );
  NOR2_X1 U2755 ( .A1(n4599), .A2(n3352), .ZN(n4598) );
  NAND2_X1 U2756 ( .A1(n4602), .A2(n3848), .ZN(n4614) );
  NAND2_X1 U2757 ( .A1(n4614), .A2(n4615), .ZN(n4613) );
  XNOR2_X1 U2758 ( .A(n3850), .B(n4749), .ZN(n4619) );
  AND2_X1 U2759 ( .A1(n2796), .A2(n2869), .ZN(n4671) );
  NOR2_X1 U2760 ( .A1(n4638), .A2(n3854), .ZN(n4648) );
  AOI21_X1 U2761 ( .B1(n3401), .B2(n3400), .A(n3399), .ZN(n3402) );
  AND2_X1 U2762 ( .A1(n3887), .A2(n2364), .ZN(n3399) );
  OR2_X1 U2763 ( .A1(n2662), .A2(n2668), .ZN(n3880) );
  NAND2_X1 U2764 ( .A1(n3911), .A2(n2230), .ZN(n2226) );
  OAI21_X1 U2765 ( .B1(n3911), .B2(n2653), .A(n2232), .ZN(n3892) );
  NAND2_X1 U2766 ( .A1(n4031), .A2(n2145), .ZN(n4408) );
  NAND2_X1 U2767 ( .A1(n2191), .A2(n2193), .ZN(n3982) );
  NAND2_X1 U2768 ( .A1(n4016), .A2(n2196), .ZN(n2191) );
  NAND2_X1 U2769 ( .A1(n2197), .A2(n2200), .ZN(n3999) );
  NAND2_X1 U2770 ( .A1(n2199), .A2(n2198), .ZN(n2197) );
  NAND2_X1 U2771 ( .A1(n3358), .A2(n2209), .ZN(n2202) );
  OAI21_X1 U2772 ( .B1(n3358), .B2(n3359), .A(n2210), .ZN(n4086) );
  NAND2_X1 U2773 ( .A1(n2214), .A2(n2218), .ZN(n4672) );
  NAND2_X1 U2774 ( .A1(n3307), .A2(n2219), .ZN(n2214) );
  OAI21_X1 U2775 ( .B1(n3307), .B2(n2503), .A(n2221), .ZN(n3284) );
  NAND2_X1 U2776 ( .A1(n2183), .A2(n2187), .ZN(n3056) );
  OR2_X1 U2777 ( .A1(n3325), .A2(n2455), .ZN(n2183) );
  INV_X1 U2778 ( .A(n4689), .ZN(n4711) );
  NAND2_X1 U2779 ( .A1(n2674), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  AND2_X2 U2780 ( .A1(n2769), .A2(n2816), .ZN(n4836) );
  AOI21_X1 U2781 ( .B1(n4111), .B2(n4110), .A(n4109), .ZN(n4535) );
  AND2_X2 U2782 ( .A1(n2769), .A2(n3072), .ZN(n4824) );
  XNOR2_X1 U2783 ( .A(n2742), .B(IR_REG_25__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U2784 ( .A1(n3510), .A2(IR_REG_31__SCAN_IN), .ZN(n2383) );
  INV_X1 U2785 ( .A(n2389), .ZN(n4493) );
  INV_X1 U2786 ( .A(n2861), .ZN(n4494) );
  XNOR2_X1 U2787 ( .A(n2740), .B(IR_REG_26__SCAN_IN), .ZN(n2788) );
  INV_X1 U2788 ( .A(n2687), .ZN(n2382) );
  XNOR2_X1 U2789 ( .A(n2738), .B(n2737), .ZN(n2790) );
  NAND2_X1 U2790 ( .A1(n2746), .A2(IR_REG_31__SCAN_IN), .ZN(n2738) );
  AND2_X1 U2791 ( .A1(n2688), .A2(n2687), .ZN(n2844) );
  INV_X1 U2792 ( .A(IR_REG_21__SCAN_IN), .ZN(n2679) );
  NOR2_X1 U2793 ( .A1(n2502), .A2(n2555), .ZN(n4497) );
  INV_X1 U2794 ( .A(IR_REG_4__SCAN_IN), .ZN(n2443) );
  AND2_X1 U2795 ( .A1(n2442), .A2(n2432), .ZN(n4498) );
  INV_X1 U2796 ( .A(n2877), .ZN(n4499) );
  XNOR2_X1 U2797 ( .A(n2262), .B(n3530), .ZN(n3537) );
  NOR2_X1 U2798 ( .A1(n2317), .A2(n2315), .ZN(n2314) );
  AOI21_X1 U2799 ( .B1(n3865), .B2(n4662), .A(n3864), .ZN(n3866) );
  AND2_X1 U2800 ( .A1(n3431), .A2(n2293), .ZN(n2133) );
  OAI22_X1 U2801 ( .A1(n3358), .A2(n2168), .B1(n2203), .B2(n2142), .ZN(n4055)
         );
  MUX2_X2 U2802 ( .A(n2399), .B(n2398), .S(n2858), .Z(n2408) );
  NAND3_X1 U2803 ( .A1(n2148), .A2(n2415), .A3(n2414), .ZN(n2905) );
  NAND2_X1 U2804 ( .A1(n3965), .A2(n3971), .ZN(n3942) );
  OR2_X1 U2805 ( .A1(n3420), .A2(n3419), .ZN(n2134) );
  NOR2_X1 U2806 ( .A1(n3262), .A2(n3261), .ZN(n2135) );
  NOR2_X1 U2807 ( .A1(n2297), .A2(n2296), .ZN(n2136) );
  AND2_X1 U2808 ( .A1(n2296), .A2(n4521), .ZN(n2137) );
  NAND2_X1 U2809 ( .A1(n2333), .A2(n2372), .ZN(n2453) );
  INV_X1 U2810 ( .A(n4706), .ZN(n4089) );
  AND2_X1 U2811 ( .A1(n3076), .A2(n3110), .ZN(n2138) );
  NAND2_X1 U2812 ( .A1(n4004), .A2(n3991), .ZN(n2139) );
  AND2_X1 U2813 ( .A1(n2365), .A2(n4065), .ZN(n2140) );
  AND2_X1 U2814 ( .A1(n3118), .A2(n3310), .ZN(n2141) );
  AND2_X1 U2815 ( .A1(n4060), .A2(n4505), .ZN(n2142) );
  INV_X1 U2816 ( .A(n3694), .ZN(n2204) );
  AND2_X1 U2817 ( .A1(n2140), .A2(n4047), .ZN(n2143) );
  NOR2_X1 U2818 ( .A1(n2765), .A2(n2615), .ZN(n2144) );
  AND2_X1 U2819 ( .A1(n2144), .A2(n3977), .ZN(n2145) );
  AND3_X1 U2820 ( .A1(n2427), .A2(n2426), .A3(n2425), .ZN(n2146) );
  OR2_X1 U2821 ( .A1(n2265), .A2(n2263), .ZN(n2147) );
  XNOR2_X1 U2822 ( .A(n2383), .B(IR_REG_30__SCAN_IN), .ZN(n2387) );
  AND2_X1 U2823 ( .A1(n2411), .A2(n2410), .ZN(n2148) );
  NAND2_X1 U2824 ( .A1(n2255), .A2(n3513), .ZN(n3538) );
  AND2_X1 U2825 ( .A1(n3900), .A2(n3914), .ZN(n2149) );
  INV_X1 U2826 ( .A(IR_REG_2__SCAN_IN), .ZN(n2417) );
  AND2_X1 U2827 ( .A1(n4495), .A2(n2788), .ZN(n2150) );
  NOR2_X1 U2828 ( .A1(n4648), .A2(n4647), .ZN(n2151) );
  AND2_X1 U2829 ( .A1(n3003), .A2(n2996), .ZN(n2152) );
  OR2_X1 U2830 ( .A1(n2327), .A2(n3701), .ZN(n2153) );
  OR2_X1 U2831 ( .A1(n3615), .A2(n2288), .ZN(n2154) );
  NAND2_X1 U2832 ( .A1(n2884), .A2(n2883), .ZN(n2304) );
  NAND2_X1 U2833 ( .A1(n3268), .A2(n3267), .ZN(n2155) );
  INV_X1 U2834 ( .A(n2225), .ZN(n2224) );
  NAND2_X1 U2835 ( .A1(n2227), .A2(n2164), .ZN(n2225) );
  NAND2_X1 U2836 ( .A1(n2416), .A2(n2417), .ZN(n2429) );
  NOR2_X1 U2837 ( .A1(n4546), .A2(n2244), .ZN(n2156) );
  NAND2_X1 U2838 ( .A1(n4552), .A2(REG2_REG_5__SCAN_IN), .ZN(n2157) );
  NOR2_X1 U2839 ( .A1(n2267), .A2(n3192), .ZN(n3269) );
  NAND2_X2 U2840 ( .A1(n2390), .A2(n4493), .ZN(n2724) );
  NOR2_X1 U2841 ( .A1(n3320), .A2(n3061), .ZN(n2158) );
  NOR2_X1 U2842 ( .A1(n4598), .A2(n3833), .ZN(n2159) );
  AND2_X1 U2843 ( .A1(n2500), .A2(n4163), .ZN(n2555) );
  OR2_X1 U2844 ( .A1(n3481), .A2(n3480), .ZN(n2160) );
  AND3_X1 U2845 ( .A1(n2372), .A2(n2416), .A3(n2254), .ZN(n2464) );
  OAI21_X1 U2846 ( .B1(n3639), .B2(n3640), .A(n3641), .ZN(n3555) );
  INV_X1 U2847 ( .A(n3748), .ZN(n2355) );
  AOI21_X1 U2848 ( .B1(n4055), .B2(n2592), .A(n2371), .ZN(n4037) );
  OAI21_X1 U2849 ( .B1(n3942), .B2(n2638), .A(n2637), .ZN(n3928) );
  NAND2_X1 U2850 ( .A1(n2226), .A2(n2227), .ZN(n3877) );
  AND2_X1 U2851 ( .A1(n2464), .A2(n2374), .ZN(n2500) );
  OR2_X1 U2852 ( .A1(n3808), .A2(n3732), .ZN(n2161) );
  INV_X1 U2853 ( .A(n3359), .ZN(n2212) );
  AND2_X1 U2854 ( .A1(n3328), .A2(n3149), .ZN(n2162) );
  INV_X1 U2855 ( .A(n2608), .ZN(n2198) );
  INV_X1 U2856 ( .A(n4674), .ZN(n4688) );
  AND2_X1 U2857 ( .A1(n3433), .A2(n3432), .ZN(n2163) );
  OR2_X1 U2858 ( .A1(n3522), .A2(n3886), .ZN(n2164) );
  NAND2_X1 U2859 ( .A1(n2705), .A2(n3753), .ZN(n3340) );
  AND2_X1 U2860 ( .A1(n2555), .A2(n2554), .ZN(n2589) );
  INV_X1 U2861 ( .A(n3513), .ZN(n2259) );
  AND2_X1 U2862 ( .A1(n3973), .A2(n2765), .ZN(n2165) );
  INV_X1 U2863 ( .A(IR_REG_31__SCAN_IN), .ZN(n2729) );
  INV_X1 U2864 ( .A(n2522), .ZN(n2220) );
  INV_X1 U2865 ( .A(n2211), .ZN(n2210) );
  NOR2_X1 U2866 ( .A1(n4097), .A2(n3366), .ZN(n2211) );
  NOR2_X1 U2867 ( .A1(n3898), .A2(n3542), .ZN(n2166) );
  NOR2_X1 U2868 ( .A1(n4678), .A2(n3285), .ZN(n2167) );
  INV_X1 U2869 ( .A(n2201), .ZN(n2200) );
  NOR2_X1 U2870 ( .A1(n3645), .A2(n4029), .ZN(n2201) );
  OR2_X1 U2871 ( .A1(n2206), .A2(n2142), .ZN(n2168) );
  AOI21_X1 U2872 ( .B1(n2219), .B2(n2503), .A(n2167), .ZN(n2218) );
  INV_X1 U2873 ( .A(n3426), .ZN(n2296) );
  AOI21_X1 U2874 ( .B1(n2196), .B2(n2608), .A(n2194), .ZN(n2193) );
  OR2_X1 U2875 ( .A1(n4522), .A2(n4521), .ZN(n2295) );
  NAND2_X1 U2876 ( .A1(n2202), .A2(n2207), .ZN(n4072) );
  INV_X1 U2877 ( .A(n3701), .ZN(n2330) );
  AND2_X1 U2878 ( .A1(n3721), .A2(n2204), .ZN(n2169) );
  NAND2_X1 U2879 ( .A1(n4678), .A2(n3285), .ZN(n2170) );
  AND2_X1 U2880 ( .A1(n2366), .A2(n4674), .ZN(n2171) );
  INV_X1 U2881 ( .A(n3486), .ZN(n2287) );
  INV_X1 U2882 ( .A(n3678), .ZN(n2331) );
  NAND2_X1 U2883 ( .A1(n3073), .A2(n4050), .ZN(n4534) );
  INV_X1 U2884 ( .A(n4534), .ZN(n4706) );
  INV_X1 U2885 ( .A(n3285), .ZN(n2367) );
  INV_X1 U2886 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2244) );
  NAND2_X1 U2887 ( .A1(n3043), .A2(n3042), .ZN(n3094) );
  NAND2_X1 U2888 ( .A1(n2182), .A2(n2180), .ZN(n3156) );
  INV_X1 U2889 ( .A(n3766), .ZN(n2352) );
  INV_X1 U2890 ( .A(n3723), .ZN(n2342) );
  INV_X1 U2891 ( .A(n4065), .ZN(n3590) );
  NOR2_X1 U2892 ( .A1(n4579), .A2(n3032), .ZN(n2172) );
  AND2_X1 U2893 ( .A1(n2408), .A2(DATAI_23_), .ZN(n3947) );
  INV_X1 U2894 ( .A(n2196), .ZN(n2195) );
  NOR2_X1 U2895 ( .A1(n3681), .A2(n2201), .ZN(n2196) );
  OR2_X1 U2896 ( .A1(n4751), .A2(n2537), .ZN(n2173) );
  AND2_X1 U2897 ( .A1(n2145), .A2(n3957), .ZN(n2174) );
  INV_X1 U2898 ( .A(n4607), .ZN(n2303) );
  NAND2_X1 U2899 ( .A1(n4716), .A2(n2690), .ZN(n2823) );
  INV_X1 U2900 ( .A(n3532), .ZN(n2364) );
  AND2_X1 U2901 ( .A1(n4700), .A2(n2409), .ZN(n3104) );
  AND2_X1 U2902 ( .A1(n2138), .A2(n4707), .ZN(n2175) );
  INV_X1 U2903 ( .A(n2905), .ZN(n2419) );
  AND2_X1 U2904 ( .A1(n2914), .A2(n2921), .ZN(n3629) );
  AND2_X1 U2905 ( .A1(n4707), .A2(n3149), .ZN(n2176) );
  AND2_X1 U2906 ( .A1(n2312), .A2(n2311), .ZN(n2177) );
  INV_X1 U2907 ( .A(n4664), .ZN(n2247) );
  INV_X1 U2908 ( .A(IR_REG_1__SCAN_IN), .ZN(n4208) );
  NAND3_X1 U2909 ( .A1(n3105), .A2(n2420), .A3(n2161), .ZN(n2178) );
  NAND2_X1 U2910 ( .A1(n2178), .A2(n2433), .ZN(n3142) );
  NAND2_X1 U2911 ( .A1(n3105), .A2(n2420), .ZN(n2179) );
  XNOR2_X1 U2912 ( .A(n2179), .B(n3078), .ZN(n4784) );
  NAND2_X1 U2913 ( .A1(n3325), .A2(n2185), .ZN(n2182) );
  OAI21_X1 U2914 ( .B1(n4016), .B2(n2190), .A(n2188), .ZN(n3965) );
  NAND3_X1 U2915 ( .A1(n4161), .A2(n2234), .A3(n2233), .ZN(n2542) );
  AND2_X2 U2916 ( .A1(n2378), .A2(n2236), .ZN(n2396) );
  MUX2_X1 U2917 ( .A(n2386), .B(REG1_REG_1__SCAN_IN), .S(n2873), .Z(n3811) );
  NAND2_X1 U2918 ( .A1(n2893), .A2(n2156), .ZN(n2242) );
  NAND2_X1 U2919 ( .A1(n2242), .A2(n2240), .ZN(n4545) );
  NAND2_X1 U2920 ( .A1(n2246), .A2(n2245), .ZN(n4661) );
  NAND2_X1 U2921 ( .A1(n4638), .A2(n2248), .ZN(n2245) );
  OAI21_X1 U2922 ( .B1(n4638), .B2(n2249), .A(n2248), .ZN(n4663) );
  NAND2_X1 U2923 ( .A1(n4619), .A2(REG1_REG_14__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U2924 ( .A1(n3493), .A2(n2260), .ZN(n2255) );
  NAND2_X1 U2925 ( .A1(n3493), .A2(n3573), .ZN(n3515) );
  OAI21_X1 U2926 ( .B1(n3188), .B2(n2269), .A(n2268), .ZN(n3420) );
  NOR3_X1 U2927 ( .A1(n3188), .A2(n2266), .A3(n2269), .ZN(n2265) );
  INV_X1 U2928 ( .A(n2271), .ZN(n3574) );
  NAND3_X1 U2929 ( .A1(n2284), .A2(n2285), .A3(n3486), .ZN(n2274) );
  NAND2_X1 U2930 ( .A1(n2289), .A2(n2996), .ZN(n3001) );
  INV_X1 U2931 ( .A(n2901), .ZN(n2824) );
  NAND2_X2 U2932 ( .A1(n2290), .A2(n2901), .ZN(n3520) );
  NAND3_X1 U2933 ( .A1(n2147), .A2(n2133), .A3(n2134), .ZN(n2291) );
  INV_X1 U2934 ( .A(n2295), .ZN(n4520) );
  NAND3_X1 U2935 ( .A1(n2301), .A2(n4607), .A3(n4599), .ZN(n2300) );
  NAND2_X1 U2936 ( .A1(n4751), .A2(n3834), .ZN(n2302) );
  INV_X1 U2937 ( .A(n2312), .ZN(n3023) );
  NAND2_X1 U2938 ( .A1(n3024), .A2(n3025), .ZN(n2311) );
  NAND3_X1 U2939 ( .A1(n2321), .A2(n2318), .A3(n2314), .ZN(U3258) );
  NAND3_X1 U2940 ( .A1(n4661), .A2(n4662), .A3(n2319), .ZN(n2318) );
  NAND3_X1 U2941 ( .A1(n4665), .A2(n4666), .A3(n2322), .ZN(n2321) );
  INV_X1 U2942 ( .A(n3078), .ZN(n2336) );
  NAND2_X1 U2943 ( .A1(n3340), .A2(n2344), .ZN(n2340) );
  NAND2_X1 U2944 ( .A1(n2340), .A2(n2341), .ZN(n4094) );
  OAI21_X1 U2945 ( .B1(n3161), .B2(n2356), .A(n2353), .ZN(n3301) );
  OAI21_X1 U2946 ( .B1(n3161), .B2(n2701), .A(n3748), .ZN(n3117) );
  AOI21_X1 U2947 ( .B1(n3748), .B2(n2701), .A(n2358), .ZN(n2357) );
  NAND2_X1 U2948 ( .A1(n2396), .A2(n2359), .ZN(n3510) );
  NAND2_X1 U2949 ( .A1(n2382), .A2(n2381), .ZN(n2739) );
  XNOR2_X1 U2950 ( .A(n3022), .B(n3010), .ZN(n2888) );
  NOR2_X1 U2951 ( .A1(n4560), .A2(n4559), .ZN(n4558) );
  XNOR2_X1 U2952 ( .A(n3027), .B(n3026), .ZN(n4559) );
  NAND2_X1 U2953 ( .A1(n4686), .A2(n3349), .ZN(n3383) );
  INV_X1 U2954 ( .A(n3582), .ZN(n3586) );
  NAND2_X1 U2955 ( .A1(n3946), .A2(n3936), .ZN(n3935) );
  OR2_X1 U2956 ( .A1(n2724), .A2(n2412), .ZN(n2415) );
  OR2_X1 U2957 ( .A1(n2724), .A2(n2820), .ZN(n2404) );
  OR2_X1 U2958 ( .A1(n2724), .A2(n2386), .ZN(n2394) );
  XNOR2_X1 U2959 ( .A(n2932), .B(n3526), .ZN(n2954) );
  OR2_X1 U2960 ( .A1(n2901), .A2(n2820), .ZN(n2370) );
  AND2_X1 U2961 ( .A1(n4502), .A2(n4065), .ZN(n2371) );
  AND2_X1 U2962 ( .A1(n3466), .A2(n3604), .ZN(n2373) );
  NAND2_X1 U2963 ( .A1(n2841), .A2(n2847), .ZN(n3725) );
  INV_X1 U2964 ( .A(n4050), .ZN(n4724) );
  INV_X1 U2965 ( .A(IR_REG_25__SCAN_IN), .ZN(n2379) );
  AND2_X1 U2966 ( .A1(n2715), .A2(n4017), .ZN(n3770) );
  INV_X1 U2967 ( .A(IR_REG_16__SCAN_IN), .ZN(n4149) );
  INV_X1 U2968 ( .A(n2847), .ZN(n2401) );
  NAND2_X1 U2969 ( .A1(n3808), .A2(n2925), .ZN(n2923) );
  OR2_X1 U2970 ( .A1(n3974), .A2(n3947), .ZN(n2636) );
  INV_X1 U2971 ( .A(IR_REG_8__SCAN_IN), .ZN(n4162) );
  NOR2_X1 U2972 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2683)
         );
  NOR2_X1 U2973 ( .A1(n3584), .A2(n3583), .ZN(n3441) );
  INV_X1 U2974 ( .A(n2636), .ZN(n2638) );
  INV_X1 U2975 ( .A(n3562), .ZN(n3467) );
  OR2_X1 U2976 ( .A1(n2647), .A2(n3577), .ZN(n2661) );
  NAND2_X1 U2977 ( .A1(n2877), .A2(REG1_REG_2__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U2978 ( .A1(n3011), .A2(n3025), .ZN(n3012) );
  OR2_X1 U2979 ( .A1(n3887), .A2(n3532), .ZN(n3404) );
  OR2_X1 U2980 ( .A1(n3960), .A2(n3977), .ZN(n3954) );
  NAND2_X1 U2981 ( .A1(n2609), .A2(REG3_REG_20__SCAN_IN), .ZN(n2616) );
  OR2_X1 U2982 ( .A1(n4097), .A2(n3360), .ZN(n3723) );
  INV_X1 U2983 ( .A(n3863), .ZN(n2822) );
  AND2_X1 U2984 ( .A1(n4716), .A2(n2784), .ZN(n4695) );
  AND2_X1 U2985 ( .A1(n2817), .A2(n4708), .ZN(n4701) );
  INV_X1 U2986 ( .A(n3002), .ZN(n3003) );
  OR2_X1 U2987 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  INV_X1 U2988 ( .A(n3917), .ZN(n3958) );
  INV_X1 U2989 ( .A(n3973), .ZN(n4004) );
  INV_X1 U2990 ( .A(n3900), .ZN(n3931) );
  OR2_X1 U2991 ( .A1(n2724), .A2(n2663), .ZN(n2664) );
  OR2_X1 U2992 ( .A1(n2422), .A2(n3948), .ZN(n2632) );
  OAI21_X1 U2993 ( .B1(n2877), .B2(REG1_REG_2__SCAN_IN), .A(n2872), .ZN(n2876)
         );
  INV_X1 U2994 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4389) );
  INV_X1 U2995 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4501) );
  AND2_X1 U2996 ( .A1(n3404), .A2(n3666), .ZN(n3699) );
  INV_X1 U2997 ( .A(n3977), .ZN(n3966) );
  AND2_X1 U2998 ( .A1(n4020), .A2(n4021), .ZN(n4042) );
  AND2_X1 U2999 ( .A1(n3723), .A2(n3651), .ZN(n3359) );
  NOR2_X1 U3000 ( .A1(n2823), .A2(n2822), .ZN(n3084) );
  INV_X1 U3001 ( .A(n3684), .ZN(n4693) );
  OR2_X1 U3002 ( .A1(n2787), .A2(D_REG_0__SCAN_IN), .ZN(n2764) );
  INV_X1 U3003 ( .A(n3201), .ZN(n3349) );
  INV_X1 U3004 ( .A(n4708), .ZN(n4718) );
  INV_X1 U3005 ( .A(n2790), .ZN(n2743) );
  NAND2_X1 U3006 ( .A1(n2468), .A2(REG3_REG_7__SCAN_IN), .ZN(n2483) );
  AND2_X1 U3007 ( .A1(n2630), .A2(REG3_REG_23__SCAN_IN), .ZN(n2639) );
  OR2_X1 U3008 ( .A1(n2524), .A2(n4389), .ZN(n2535) );
  NAND2_X1 U3009 ( .A1(n2447), .A2(REG3_REG_5__SCAN_IN), .ZN(n2458) );
  OR2_X1 U3010 ( .A1(n2535), .A2(n2534), .ZN(n2548) );
  INV_X1 U3011 ( .A(n4047), .ZN(n3647) );
  INV_X1 U3012 ( .A(n4528), .ZN(n3623) );
  NAND2_X1 U3013 ( .A1(n2558), .A2(REG3_REG_15__SCAN_IN), .ZN(n2570) );
  NAND4_X1 U3014 ( .A1(n2673), .A2(n2672), .A3(n2671), .A4(n2670), .ZN(n3887)
         );
  OR2_X1 U3015 ( .A1(n2422), .A2(n3967), .ZN(n2625) );
  INV_X1 U3016 ( .A(n4659), .ZN(n4662) );
  AND2_X1 U3017 ( .A1(n4089), .A2(n3084), .ZN(n4689) );
  INV_X1 U3018 ( .A(n4681), .ZN(n4719) );
  AND2_X1 U3019 ( .A1(n2764), .A2(n2763), .ZN(n2816) );
  INV_X1 U3020 ( .A(n4801), .ZN(n4809) );
  INV_X1 U3021 ( .A(n2823), .ZN(n4812) );
  INV_X1 U3022 ( .A(n2816), .ZN(n3072) );
  AND2_X1 U3023 ( .A1(n2577), .A2(n2568), .ZN(n3844) );
  AND2_X1 U3024 ( .A1(n2490), .A2(n2478), .ZN(n4758) );
  OR2_X1 U3025 ( .A1(n2835), .A2(n2831), .ZN(n3626) );
  NAND4_X1 U3026 ( .A1(n2652), .A2(n2651), .A3(n2650), .A4(n2649), .ZN(n3900)
         );
  NAND4_X1 U3027 ( .A1(n2628), .A2(n2627), .A3(n2626), .A4(n2625), .ZN(n3960)
         );
  INV_X1 U3028 ( .A(n4758), .ZN(n4578) );
  OR2_X1 U3029 ( .A1(n4543), .A2(n4494), .ZN(n4669) );
  OR2_X1 U3030 ( .A1(n4543), .A2(n3796), .ZN(n4654) );
  AND2_X1 U3031 ( .A1(n4712), .A2(n3155), .ZN(n4101) );
  OR2_X1 U3032 ( .A1(n3869), .A2(n4435), .ZN(n2767) );
  INV_X1 U3033 ( .A(n4836), .ZN(n4834) );
  OR2_X1 U3034 ( .A1(n3869), .A2(n4489), .ZN(n2772) );
  INV_X1 U3035 ( .A(n4824), .ZN(n4822) );
  INV_X1 U3036 ( .A(n4739), .ZN(n4741) );
  AND2_X1 U3037 ( .A1(n2900), .A2(STATE_REG_SCAN_IN), .ZN(n4742) );
  INV_X1 U3038 ( .A(n3849), .ZN(n4749) );
  INV_X1 U3039 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U3040 ( .A1(n2737), .A2(n2379), .ZN(n2380) );
  INV_X1 U3041 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2386) );
  INV_X1 U3042 ( .A(n2422), .ZN(n2388) );
  NAND2_X1 U3043 ( .A1(n2388), .A2(REG3_REG_1__SCAN_IN), .ZN(n2393) );
  NAND2_X1 U3044 ( .A1(n2421), .A2(REG2_REG_1__SCAN_IN), .ZN(n2392) );
  AND2_X2 U3045 ( .A1(n2390), .A2(n2389), .ZN(n2424) );
  NAND2_X1 U3046 ( .A1(n2424), .A2(REG0_REG_1__SCAN_IN), .ZN(n2391) );
  NAND4_X2 U3047 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(n2841)
         );
  INV_X1 U3048 ( .A(n2841), .ZN(n2402) );
  INV_X1 U3049 ( .A(DATAI_1_), .ZN(n2400) );
  NAND2_X1 U3050 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2399) );
  NAND2_X1 U3051 ( .A1(n2731), .A2(n2395), .ZN(n2398) );
  MUX2_X1 U3052 ( .A(n2873), .B(n2400), .S(n2408), .Z(n2847) );
  NAND2_X1 U3053 ( .A1(n2402), .A2(n2401), .ZN(n2694) );
  NAND2_X1 U3054 ( .A1(n2694), .A2(n3725), .ZN(n2692) );
  NAND2_X1 U3055 ( .A1(n2424), .A2(REG0_REG_0__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3056 ( .A1(n2421), .A2(REG2_REG_0__SCAN_IN), .ZN(n2406) );
  INV_X1 U3057 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2403) );
  OR2_X1 U3058 ( .A1(n2422), .A2(n2403), .ZN(n2405) );
  INV_X1 U3059 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2820) );
  NAND4_X1 U3060 ( .A1(n2407), .A2(n2406), .A3(n2405), .A4(n2404), .ZN(n2817)
         );
  MUX2_X1 U3061 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2408), .Z(n4708) );
  NAND2_X1 U3062 ( .A1(n2692), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U3063 ( .A1(n2841), .A2(n2401), .ZN(n2409) );
  NAND2_X1 U3064 ( .A1(n2421), .A2(REG2_REG_2__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3065 ( .A1(n2424), .A2(REG0_REG_2__SCAN_IN), .ZN(n2410) );
  INV_X1 U3066 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2412) );
  INV_X1 U3067 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2413) );
  OR2_X1 U3068 ( .A1(n2422), .A2(n2413), .ZN(n2414) );
  INV_X1 U3069 ( .A(DATAI_2_), .ZN(n2418) );
  MUX2_X1 U3070 ( .A(n2877), .B(n2418), .S(n2408), .Z(n3110) );
  NAND2_X1 U3071 ( .A1(n2905), .A2(n3110), .ZN(n3729) );
  NAND2_X1 U3072 ( .A1(n3104), .A2(n3696), .ZN(n3105) );
  INV_X1 U3073 ( .A(n3110), .ZN(n3633) );
  OR2_X1 U3074 ( .A1(n2905), .A2(n3633), .ZN(n2420) );
  NAND2_X1 U3075 ( .A1(n2421), .A2(REG2_REG_3__SCAN_IN), .ZN(n2428) );
  OR2_X1 U3076 ( .A1(n2422), .A2(REG3_REG_3__SCAN_IN), .ZN(n2427) );
  INV_X1 U3077 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2423) );
  OR2_X1 U3078 ( .A1(n2724), .A2(n2423), .ZN(n2426) );
  NAND2_X1 U3079 ( .A1(n2424), .A2(REG0_REG_3__SCAN_IN), .ZN(n2425) );
  NAND2_X1 U3080 ( .A1(n2429), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3081 ( .A1(n2431), .A2(n2430), .ZN(n2442) );
  OR2_X1 U3082 ( .A1(n2431), .A2(n2430), .ZN(n2432) );
  MUX2_X1 U3083 ( .A(n4498), .B(DATAI_3_), .S(n2408), .Z(n3732) );
  NAND2_X1 U3084 ( .A1(n3808), .A2(n3732), .ZN(n2433) );
  NAND2_X1 U3085 ( .A1(n2424), .A2(REG0_REG_4__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3086 ( .A1(n2421), .A2(REG2_REG_4__SCAN_IN), .ZN(n2440) );
  OR2_X1 U3087 ( .A1(n2724), .A2(n2244), .ZN(n2439) );
  AND2_X2 U3088 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2447) );
  INV_X1 U3089 ( .A(n2447), .ZN(n2437) );
  INV_X1 U3090 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2435) );
  INV_X1 U3091 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3092 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3093 ( .A1(n2437), .A2(n2436), .ZN(n3150) );
  OR2_X1 U3094 ( .A1(n2422), .A2(n3150), .ZN(n2438) );
  NAND2_X1 U3095 ( .A1(n2442), .A2(IR_REG_31__SCAN_IN), .ZN(n2444) );
  XNOR2_X1 U3096 ( .A(n2444), .B(n2443), .ZN(n3010) );
  INV_X1 U3097 ( .A(DATAI_4_), .ZN(n2774) );
  MUX2_X1 U3098 ( .A(n3010), .B(n2774), .S(n2408), .Z(n3149) );
  OR2_X1 U3099 ( .A1(n3806), .A2(n3149), .ZN(n3734) );
  NAND2_X1 U3100 ( .A1(n3806), .A2(n3149), .ZN(n3737) );
  NAND2_X1 U3101 ( .A1(n3734), .A2(n3737), .ZN(n3691) );
  NAND2_X1 U3102 ( .A1(n3142), .A2(n3691), .ZN(n2446) );
  INV_X1 U3103 ( .A(n3149), .ZN(n2941) );
  NAND2_X1 U3104 ( .A1(n3806), .A2(n2941), .ZN(n2445) );
  NAND2_X1 U3105 ( .A1(n2446), .A2(n2445), .ZN(n3325) );
  NAND2_X1 U3106 ( .A1(n2421), .A2(REG2_REG_5__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3107 ( .A1(n2424), .A2(REG0_REG_5__SCAN_IN), .ZN(n2451) );
  OAI21_X1 U3108 ( .B1(n2447), .B2(REG3_REG_5__SCAN_IN), .A(n2458), .ZN(n3330)
         );
  OR2_X1 U3109 ( .A1(n2422), .A2(n3330), .ZN(n2450) );
  INV_X1 U3110 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2448) );
  OR2_X1 U3111 ( .A1(n2724), .A2(n2448), .ZN(n2449) );
  NAND4_X1 U3112 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n3805)
         );
  NAND2_X1 U3113 ( .A1(n2453), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  MUX2_X1 U3114 ( .A(n4552), .B(DATAI_5_), .S(n2408), .Z(n3319) );
  AND2_X1 U3115 ( .A1(n3805), .A2(n3319), .ZN(n2455) );
  NAND2_X1 U3116 ( .A1(n2424), .A2(REG0_REG_6__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3117 ( .A1(n2421), .A2(REG2_REG_6__SCAN_IN), .ZN(n2462) );
  INV_X1 U3118 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2456) );
  OR2_X1 U3119 ( .A1(n2724), .A2(n2456), .ZN(n2461) );
  AND2_X1 U3120 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  NOR2_X2 U3121 ( .A1(n2458), .A2(n2457), .ZN(n2468) );
  OR2_X1 U3122 ( .A1(n2459), .A2(n2468), .ZN(n3233) );
  OR2_X1 U3123 ( .A1(n2422), .A2(n3233), .ZN(n2460) );
  NAND4_X1 U3124 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n3320)
         );
  OR2_X1 U3125 ( .A1(n2464), .A2(n2729), .ZN(n2465) );
  XNOR2_X1 U3126 ( .A(n2465), .B(IR_REG_6__SCAN_IN), .ZN(n4760) );
  MUX2_X1 U3127 ( .A(n4760), .B(DATAI_6_), .S(n2408), .Z(n3061) );
  NAND2_X1 U3128 ( .A1(n3320), .A2(n3061), .ZN(n2466) );
  NAND2_X1 U3129 ( .A1(n2424), .A2(REG0_REG_7__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3130 ( .A1(n2421), .A2(REG2_REG_7__SCAN_IN), .ZN(n2472) );
  INV_X1 U3131 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2467) );
  OR2_X1 U3132 ( .A1(n2724), .A2(n2467), .ZN(n2471) );
  OR2_X1 U3133 ( .A1(n2468), .A2(REG3_REG_7__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3134 ( .A1(n2483), .A2(n2469), .ZN(n3169) );
  OR2_X1 U3135 ( .A1(n2422), .A2(n3169), .ZN(n2470) );
  NAND2_X1 U3136 ( .A1(n2464), .A2(n2474), .ZN(n2475) );
  NAND2_X1 U3137 ( .A1(n2475), .A2(IR_REG_31__SCAN_IN), .ZN(n2477) );
  NAND2_X1 U3138 ( .A1(n2477), .A2(n2476), .ZN(n2490) );
  OR2_X1 U3139 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
  INV_X1 U3140 ( .A(DATAI_7_), .ZN(n2479) );
  MUX2_X1 U3141 ( .A(n4578), .B(n2479), .S(n2408), .Z(n3165) );
  OR2_X1 U3142 ( .A1(n3120), .A2(n3165), .ZN(n3740) );
  NAND2_X1 U3143 ( .A1(n3120), .A2(n3165), .ZN(n3748) );
  NAND2_X1 U3144 ( .A1(n3740), .A2(n3748), .ZN(n3695) );
  NAND2_X1 U3145 ( .A1(n3156), .A2(n3695), .ZN(n2481) );
  INV_X1 U3146 ( .A(n3165), .ZN(n3007) );
  NAND2_X1 U3147 ( .A1(n3120), .A2(n3007), .ZN(n2480) );
  NAND2_X1 U31480 ( .A1(n2481), .A2(n2480), .ZN(n3116) );
  NAND2_X1 U31490 ( .A1(n2421), .A2(REG2_REG_8__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3150 ( .A1(n2424), .A2(REG0_REG_8__SCAN_IN), .ZN(n2488) );
  OR2_X2 U3151 ( .A1(n2483), .A2(n2482), .ZN(n2494) );
  NAND2_X1 U3152 ( .A1(n2483), .A2(n2482), .ZN(n2484) );
  NAND2_X1 U3153 ( .A1(n2494), .A2(n2484), .ZN(n3295) );
  OR2_X1 U3154 ( .A1(n2422), .A2(n3295), .ZN(n2487) );
  INV_X1 U3155 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2485) );
  OR2_X1 U3156 ( .A1(n2724), .A2(n2485), .ZN(n2486) );
  NAND4_X1 U3157 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n3162)
         );
  NAND2_X1 U3158 ( .A1(n2490), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  XNOR2_X1 U3159 ( .A(n2491), .B(IR_REG_8__SCAN_IN), .ZN(n3030) );
  MUX2_X1 U3160 ( .A(n3030), .B(DATAI_8_), .S(n2408), .Z(n3046) );
  AND2_X1 U3161 ( .A1(n3162), .A2(n3046), .ZN(n2493) );
  OR2_X1 U3162 ( .A1(n3162), .A2(n3046), .ZN(n2492) );
  NAND2_X1 U3163 ( .A1(n2424), .A2(REG0_REG_9__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U3164 ( .A1(n2421), .A2(REG2_REG_9__SCAN_IN), .ZN(n2498) );
  INV_X1 U3165 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3018) );
  AND2_X1 U3166 ( .A1(n2494), .A2(n3021), .ZN(n2495) );
  NOR2_X2 U3167 ( .A1(n2494), .A2(n3021), .ZN(n2504) );
  OR2_X1 U3168 ( .A1(n2495), .A2(n2504), .ZN(n3312) );
  OR2_X1 U3169 ( .A1(n2422), .A2(n3312), .ZN(n2496) );
  NOR2_X1 U3170 ( .A1(n2500), .A2(n2729), .ZN(n2501) );
  MUX2_X1 U3171 ( .A(n2729), .B(n2501), .S(IR_REG_9__SCAN_IN), .Z(n2502) );
  INV_X1 U3172 ( .A(n2555), .ZN(n2543) );
  MUX2_X1 U3173 ( .A(n4497), .B(DATAI_9_), .S(n2408), .Z(n3302) );
  NOR2_X1 U3174 ( .A1(n3804), .A2(n3302), .ZN(n2503) );
  INV_X1 U3175 ( .A(n3302), .ZN(n3310) );
  NAND2_X1 U3176 ( .A1(n2421), .A2(REG2_REG_10__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3177 ( .A1(n2424), .A2(REG0_REG_10__SCAN_IN), .ZN(n2509) );
  AND2_X2 U3178 ( .A1(n2504), .A2(REG3_REG_10__SCAN_IN), .ZN(n2512) );
  NOR2_X1 U3179 ( .A1(n2504), .A2(REG3_REG_10__SCAN_IN), .ZN(n2505) );
  OR2_X1 U3180 ( .A1(n2512), .A2(n2505), .ZN(n3287) );
  INV_X1 U3181 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2506) );
  OR2_X1 U3182 ( .A1(n2724), .A2(n2506), .ZN(n2507) );
  NAND2_X1 U3183 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U3184 ( .A(n2511), .B(IR_REG_10__SCAN_IN), .ZN(n3249) );
  MUX2_X1 U3185 ( .A(n3249), .B(DATAI_10_), .S(n2408), .Z(n3285) );
  NAND2_X1 U3186 ( .A1(n2424), .A2(REG0_REG_11__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U3187 ( .A1(n2421), .A2(REG2_REG_11__SCAN_IN), .ZN(n2516) );
  OR2_X1 U3188 ( .A1(n2512), .A2(REG3_REG_11__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3189 ( .A1(n2524), .A2(n2513), .ZN(n4684) );
  OR2_X1 U3190 ( .A1(n2422), .A2(n4684), .ZN(n2515) );
  INV_X1 U3191 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3244) );
  OR2_X1 U3192 ( .A1(n2724), .A2(n3244), .ZN(n2514) );
  NAND4_X1 U3193 ( .A1(n2517), .A2(n2516), .A3(n2515), .A4(n2514), .ZN(n3803)
         );
  NAND2_X1 U3194 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3195 ( .A1(n2519), .A2(n4161), .ZN(n2530) );
  OR2_X1 U3196 ( .A1(n2519), .A2(n4161), .ZN(n2520) );
  NAND2_X1 U3197 ( .A1(n2530), .A2(n2520), .ZN(n3846) );
  INV_X1 U3198 ( .A(DATAI_11_), .ZN(n2521) );
  MUX2_X1 U3199 ( .A(n3846), .B(n2521), .S(n2408), .Z(n4674) );
  OR2_X1 U3200 ( .A1(n3803), .A2(n4674), .ZN(n3341) );
  NAND2_X1 U3201 ( .A1(n3803), .A2(n4674), .ZN(n3343) );
  NAND2_X1 U3202 ( .A1(n3341), .A2(n3343), .ZN(n4673) );
  NOR2_X1 U3203 ( .A1(n3803), .A2(n4688), .ZN(n2522) );
  NAND2_X1 U3204 ( .A1(n2424), .A2(REG0_REG_12__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U3205 ( .A1(n2421), .A2(REG2_REG_12__SCAN_IN), .ZN(n2528) );
  INV_X1 U3206 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2523) );
  OR2_X1 U3207 ( .A1(n2724), .A2(n2523), .ZN(n2527) );
  NAND2_X1 U3208 ( .A1(n2524), .A2(n4389), .ZN(n2525) );
  NAND2_X1 U3209 ( .A1(n2535), .A2(n2525), .ZN(n3351) );
  OR2_X1 U32100 ( .A1(n2422), .A2(n3351), .ZN(n2526) );
  NAND4_X1 U32110 ( .A1(n2529), .A2(n2528), .A3(n2527), .A4(n2526), .ZN(n3802)
         );
  NAND2_X1 U32120 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  XNOR2_X1 U32130 ( .A(n2531), .B(IR_REG_12__SCAN_IN), .ZN(n4752) );
  MUX2_X1 U32140 ( .A(n4752), .B(DATAI_12_), .S(n2408), .Z(n3201) );
  OR2_X1 U32150 ( .A1(n3802), .A2(n3201), .ZN(n2533) );
  AND2_X1 U32160 ( .A1(n3802), .A2(n3201), .ZN(n2532) );
  NAND2_X1 U32170 ( .A1(n2421), .A2(REG2_REG_13__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32180 ( .A1(n2424), .A2(REG0_REG_13__SCAN_IN), .ZN(n2540) );
  INV_X1 U32190 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U32200 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  NAND2_X1 U32210 ( .A1(n2548), .A2(n2536), .ZN(n3387) );
  OR2_X1 U32220 ( .A1(n2422), .A2(n3387), .ZN(n2539) );
  INV_X1 U32230 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2537) );
  OR2_X1 U32240 ( .A1(n2724), .A2(n2537), .ZN(n2538) );
  NOR2_X1 U32250 ( .A1(n2543), .A2(n2542), .ZN(n2544) );
  OR2_X1 U32260 ( .A1(n2544), .A2(n2729), .ZN(n2545) );
  XNOR2_X1 U32270 ( .A(n2545), .B(IR_REG_13__SCAN_IN), .ZN(n4608) );
  MUX2_X1 U32280 ( .A(n4608), .B(DATAI_13_), .S(n2408), .Z(n3230) );
  NAND2_X1 U32290 ( .A1(n3376), .A2(n3230), .ZN(n2547) );
  NOR2_X1 U32300 ( .A1(n3376), .A2(n3230), .ZN(n2546) );
  NAND2_X1 U32310 ( .A1(n2421), .A2(REG2_REG_14__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32320 ( .A1(n2424), .A2(REG0_REG_14__SCAN_IN), .ZN(n2552) );
  AND2_X1 U32330 ( .A1(n2548), .A2(n4384), .ZN(n2549) );
  OR2_X1 U32340 ( .A1(n2549), .A2(n2558), .ZN(n3367) );
  OR2_X1 U32350 ( .A1(n2422), .A2(n3367), .ZN(n2551) );
  INV_X1 U32360 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4195) );
  OR2_X1 U32370 ( .A1(n2724), .A2(n4195), .ZN(n2550) );
  NAND4_X1 U32380 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n4097)
         );
  OR2_X1 U32390 ( .A1(n2589), .A2(n2729), .ZN(n2556) );
  XNOR2_X1 U32400 ( .A(n2556), .B(IR_REG_14__SCAN_IN), .ZN(n3849) );
  INV_X1 U32410 ( .A(DATAI_14_), .ZN(n2557) );
  MUX2_X1 U32420 ( .A(n4749), .B(n2557), .S(n2408), .Z(n3360) );
  NAND2_X1 U32430 ( .A1(n4097), .A2(n3360), .ZN(n3651) );
  NAND2_X1 U32440 ( .A1(n2421), .A2(REG2_REG_15__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32450 ( .A1(n2424), .A2(REG0_REG_15__SCAN_IN), .ZN(n2562) );
  OR2_X1 U32460 ( .A1(n2558), .A2(REG3_REG_15__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32470 ( .A1(n2570), .A2(n2559), .ZN(n4527) );
  OR2_X1 U32480 ( .A1(n2422), .A2(n4527), .ZN(n2561) );
  INV_X1 U32490 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4196) );
  NAND4_X1 U32500 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3425)
         );
  INV_X1 U32510 ( .A(IR_REG_14__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32520 ( .A1(n2589), .A2(n2564), .ZN(n2565) );
  NAND2_X1 U32530 ( .A1(n2565), .A2(IR_REG_31__SCAN_IN), .ZN(n2567) );
  INV_X1 U32540 ( .A(IR_REG_15__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32550 ( .A1(n2567), .A2(n2566), .ZN(n2577) );
  OR2_X1 U32560 ( .A1(n2567), .A2(n2566), .ZN(n2568) );
  MUX2_X1 U32570 ( .A(n3844), .B(DATAI_15_), .S(n2408), .Z(n4519) );
  NOR2_X1 U32580 ( .A1(n3425), .A2(n4519), .ZN(n2569) );
  INV_X1 U32590 ( .A(n3425), .ZN(n4503) );
  NAND2_X1 U32600 ( .A1(n2421), .A2(REG2_REG_16__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U32610 ( .A1(n2424), .A2(REG0_REG_16__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32620 ( .A1(n2570), .A2(n4501), .ZN(n2572) );
  INV_X1 U32630 ( .A(n2593), .ZN(n2571) );
  NAND2_X1 U32640 ( .A1(n2572), .A2(n2571), .ZN(n4511) );
  OR2_X1 U32650 ( .A1(n2422), .A2(n4511), .ZN(n2574) );
  INV_X1 U32660 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4433) );
  OR2_X1 U32670 ( .A1(n2724), .A2(n4433), .ZN(n2573) );
  NAND2_X1 U32680 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U32690 ( .A(n2578), .B(IR_REG_16__SCAN_IN), .ZN(n3853) );
  INV_X1 U32700 ( .A(n3853), .ZN(n4746) );
  INV_X1 U32710 ( .A(DATAI_16_), .ZN(n4745) );
  MUX2_X1 U32720 ( .A(n4746), .B(n4745), .S(n2408), .Z(n4080) );
  OR2_X1 U32730 ( .A1(n4060), .A2(n4080), .ZN(n3767) );
  NAND2_X1 U32740 ( .A1(n4060), .A2(n4080), .ZN(n3766) );
  NAND2_X1 U32750 ( .A1(n3767), .A2(n3766), .ZN(n3694) );
  INV_X1 U32760 ( .A(n4080), .ZN(n4505) );
  NAND2_X1 U32770 ( .A1(n2424), .A2(REG0_REG_17__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32780 ( .A1(n2421), .A2(REG2_REG_17__SCAN_IN), .ZN(n2581) );
  XNOR2_X1 U32790 ( .A(REG3_REG_17__SCAN_IN), .B(n2593), .ZN(n4067) );
  OR2_X1 U32800 ( .A1(n2422), .A2(n4067), .ZN(n2580) );
  INV_X1 U32810 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4429) );
  OR2_X1 U32820 ( .A1(n2724), .A2(n4429), .ZN(n2579) );
  NAND4_X1 U32830 ( .A1(n2582), .A2(n2581), .A3(n2580), .A4(n2579), .ZN(n4076)
         );
  INV_X1 U32840 ( .A(n2583), .ZN(n2584) );
  NAND2_X1 U32850 ( .A1(n2589), .A2(n2587), .ZN(n2585) );
  NAND2_X1 U32860 ( .A1(n2585), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  MUX2_X1 U32870 ( .A(IR_REG_31__SCAN_IN), .B(n2586), .S(IR_REG_17__SCAN_IN), 
        .Z(n2590) );
  NAND2_X1 U32880 ( .A1(n2590), .A2(n2685), .ZN(n4653) );
  INV_X1 U32890 ( .A(DATAI_17_), .ZN(n2591) );
  MUX2_X1 U32900 ( .A(n4653), .B(n2591), .S(n2408), .Z(n4065) );
  NAND2_X1 U32910 ( .A1(n4076), .A2(n3590), .ZN(n2592) );
  INV_X1 U32920 ( .A(n4076), .ZN(n4502) );
  NAND2_X1 U32930 ( .A1(n2421), .A2(REG2_REG_18__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U32940 ( .A1(n2424), .A2(REG0_REG_18__SCAN_IN), .ZN(n2597) );
  OAI21_X1 U32950 ( .B1(n2594), .B2(REG3_REG_18__SCAN_IN), .A(n2602), .ZN(
        n4051) );
  OR2_X1 U32960 ( .A1(n2422), .A2(n4051), .ZN(n2596) );
  INV_X1 U32970 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3858) );
  OR2_X1 U32980 ( .A1(n2724), .A2(n3858), .ZN(n2595) );
  NAND2_X1 U32990 ( .A1(n2685), .A2(IR_REG_31__SCAN_IN), .ZN(n2599) );
  XNOR2_X1 U33000 ( .A(n2599), .B(IR_REG_18__SCAN_IN), .ZN(n3857) );
  INV_X1 U33010 ( .A(DATAI_18_), .ZN(n2600) );
  MUX2_X1 U33020 ( .A(n4744), .B(n2600), .S(n2408), .Z(n4047) );
  OR2_X1 U33030 ( .A1(n4059), .A2(n4047), .ZN(n4020) );
  NAND2_X1 U33040 ( .A1(n4059), .A2(n4047), .ZN(n4021) );
  NAND2_X1 U33050 ( .A1(n2424), .A2(REG0_REG_19__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33060 ( .A1(n2421), .A2(REG2_REG_19__SCAN_IN), .ZN(n2606) );
  INV_X1 U33070 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4422) );
  INV_X1 U33080 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4172) );
  AND2_X1 U33090 ( .A1(n2602), .A2(n4172), .ZN(n2603) );
  OR2_X1 U33100 ( .A1(n2603), .A2(n2609), .ZN(n3557) );
  OR2_X1 U33110 ( .A1(n2422), .A2(n3557), .ZN(n2604) );
  INV_X1 U33120 ( .A(DATAI_19_), .ZN(n4254) );
  MUX2_X1 U33130 ( .A(n3863), .B(n4254), .S(n2408), .Z(n4029) );
  INV_X1 U33140 ( .A(n4029), .ZN(n3451) );
  NOR2_X1 U33150 ( .A1(n4044), .A2(n3451), .ZN(n2608) );
  NAND2_X1 U33160 ( .A1(n2421), .A2(REG2_REG_20__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U33170 ( .A1(n2424), .A2(REG0_REG_20__SCAN_IN), .ZN(n2613) );
  OR2_X1 U33180 ( .A1(n2609), .A2(REG3_REG_20__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33190 ( .A1(n2616), .A2(n2610), .ZN(n4010) );
  OR2_X1 U33200 ( .A1(n2422), .A2(n4010), .ZN(n2612) );
  INV_X1 U33210 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4418) );
  OR2_X1 U33220 ( .A1(n2724), .A2(n4418), .ZN(n2611) );
  NAND4_X1 U33230 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n3987)
         );
  NAND2_X1 U33240 ( .A1(n2408), .A2(DATAI_20_), .ZN(n4009) );
  INV_X1 U33250 ( .A(n4009), .ZN(n2615) );
  AND2_X1 U33260 ( .A1(n3987), .A2(n2615), .ZN(n3681) );
  OR2_X1 U33270 ( .A1(n3987), .A2(n2615), .ZN(n3682) );
  NAND2_X1 U33280 ( .A1(n2424), .A2(REG0_REG_21__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U33290 ( .A1(n2421), .A2(REG2_REG_21__SCAN_IN), .ZN(n2620) );
  INV_X1 U33300 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4414) );
  OR2_X1 U33310 ( .A1(n2724), .A2(n4414), .ZN(n2619) );
  INV_X1 U33320 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3566) );
  OR2_X2 U33330 ( .A1(n2616), .A2(n3566), .ZN(n2623) );
  NAND2_X1 U33340 ( .A1(n2616), .A2(n3566), .ZN(n2617) );
  NAND2_X1 U33350 ( .A1(n2623), .A2(n2617), .ZN(n3993) );
  OR2_X1 U33360 ( .A1(n2422), .A2(n3993), .ZN(n2618) );
  NAND2_X1 U33370 ( .A1(n2408), .A2(DATAI_21_), .ZN(n3991) );
  INV_X1 U33380 ( .A(n3991), .ZN(n2765) );
  NAND2_X1 U33390 ( .A1(n2424), .A2(REG0_REG_22__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U33400 ( .A1(n2421), .A2(REG2_REG_22__SCAN_IN), .ZN(n2627) );
  INV_X1 U33410 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2622) );
  INV_X1 U33420 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3619) );
  AND2_X1 U33430 ( .A1(n2623), .A2(n3619), .ZN(n2624) );
  NOR2_X2 U33440 ( .A1(n2623), .A2(n3619), .ZN(n2630) );
  OR2_X1 U33450 ( .A1(n2624), .A2(n2630), .ZN(n3967) );
  NAND2_X1 U33460 ( .A1(n2408), .A2(DATAI_22_), .ZN(n3977) );
  NAND2_X1 U33470 ( .A1(n3960), .A2(n3977), .ZN(n2717) );
  NAND2_X1 U33480 ( .A1(n2424), .A2(REG0_REG_23__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33490 ( .A1(n2421), .A2(REG2_REG_23__SCAN_IN), .ZN(n2634) );
  INV_X1 U33500 ( .A(REG1_REG_23__SCAN_IN), .ZN(n2629) );
  OR2_X1 U33510 ( .A1(n2724), .A2(n2629), .ZN(n2633) );
  NOR2_X1 U33520 ( .A1(n2630), .A2(REG3_REG_23__SCAN_IN), .ZN(n2631) );
  OR2_X1 U3353 ( .A1(n2639), .A2(n2631), .ZN(n3948) );
  AND2_X1 U33540 ( .A1(n3960), .A2(n3966), .ZN(n3943) );
  AOI22_X1 U3355 ( .A1(n3943), .A2(n2636), .B1(n3947), .B2(n3974), .ZN(n2637)
         );
  NAND2_X1 U3356 ( .A1(n2421), .A2(REG2_REG_24__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3357 ( .A1(n2424), .A2(REG0_REG_24__SCAN_IN), .ZN(n2643) );
  OR2_X1 U3358 ( .A1(n2639), .A2(REG3_REG_24__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3359 ( .A1(n2647), .A2(n2640), .ZN(n3937) );
  INV_X1 U3360 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U3361 ( .A1(n2408), .A2(DATAI_24_), .ZN(n3936) );
  NOR2_X1 U3362 ( .A1(n3958), .A2(n3936), .ZN(n2646) );
  INV_X1 U3363 ( .A(n3936), .ZN(n3482) );
  NAND2_X1 U3364 ( .A1(n2424), .A2(REG0_REG_25__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3365 ( .A1(n2421), .A2(REG2_REG_25__SCAN_IN), .ZN(n2651) );
  INV_X1 U3366 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4130) );
  OR2_X1 U3367 ( .A1(n2724), .A2(n4130), .ZN(n2650) );
  INV_X1 U3368 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U3369 ( .A1(n2647), .A2(n3577), .ZN(n2648) );
  NAND2_X1 U3370 ( .A1(n2661), .A2(n2648), .ZN(n3576) );
  NAND2_X1 U3371 ( .A1(n2408), .A2(DATAI_25_), .ZN(n3914) );
  INV_X1 U3372 ( .A(n3914), .ZN(n3920) );
  NOR2_X1 U3373 ( .A1(n3900), .A2(n3920), .ZN(n2653) );
  NAND2_X1 U3374 ( .A1(n2421), .A2(REG2_REG_26__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3375 ( .A1(n2424), .A2(REG0_REG_26__SCAN_IN), .ZN(n2656) );
  INV_X1 U3376 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3505) );
  XNOR2_X1 U3377 ( .A(n2661), .B(n3505), .ZN(n3504) );
  INV_X1 U3378 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4301) );
  OR2_X1 U3379 ( .A1(n2724), .A2(n4301), .ZN(n2654) );
  NAND2_X1 U3380 ( .A1(n2408), .A2(DATAI_26_), .ZN(n3904) );
  NOR2_X1 U3381 ( .A1(n3915), .A2(n3904), .ZN(n2658) );
  INV_X1 U3382 ( .A(n3904), .ZN(n2766) );
  NAND2_X1 U3383 ( .A1(n2424), .A2(REG0_REG_27__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3384 ( .A1(n2421), .A2(REG2_REG_27__SCAN_IN), .ZN(n2666) );
  INV_X1 U3385 ( .A(n2661), .ZN(n2659) );
  AOI21_X1 U3386 ( .B1(n2659), .B2(REG3_REG_26__SCAN_IN), .A(
        REG3_REG_27__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3387 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2660) );
  NOR2_X2 U3388 ( .A1(n2661), .A2(n2660), .ZN(n2668) );
  INV_X1 U3389 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3390 ( .A1(n2408), .A2(DATAI_27_), .ZN(n3542) );
  INV_X1 U3391 ( .A(n3542), .ZN(n3886) );
  INV_X1 U3392 ( .A(n3522), .ZN(n3898) );
  NAND2_X1 U3393 ( .A1(n2424), .A2(REG0_REG_28__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3394 ( .A1(n2421), .A2(REG2_REG_28__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3395 ( .A1(n2668), .A2(REG3_REG_28__SCAN_IN), .ZN(n3414) );
  OR2_X1 U3396 ( .A1(n2668), .A2(REG3_REG_28__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3397 ( .A1(n3414), .A2(n2669), .ZN(n3870) );
  OR2_X1 U3398 ( .A1(n2724), .A2(n4303), .ZN(n2670) );
  NAND2_X1 U3399 ( .A1(n2408), .A2(DATAI_28_), .ZN(n3532) );
  NAND2_X1 U3400 ( .A1(n3887), .A2(n3532), .ZN(n3666) );
  XNOR2_X1 U3401 ( .A(n3401), .B(n3699), .ZN(n3868) );
  NAND2_X1 U3402 ( .A1(n2678), .A2(n4222), .ZN(n2674) );
  NAND2_X1 U3403 ( .A1(n4222), .A2(n2676), .ZN(n2681) );
  NAND2_X1 U3404 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U3405 ( .A1(n2678), .A2(n2677), .ZN(n2680) );
  INV_X1 U3406 ( .A(n2681), .ZN(n2682) );
  NAND2_X1 U3407 ( .A1(n2683), .A2(n2682), .ZN(n2684) );
  OAI21_X1 U3408 ( .B1(n2685), .B2(n2684), .A(IR_REG_31__SCAN_IN), .ZN(n2686)
         );
  MUX2_X1 U3409 ( .A(IR_REG_31__SCAN_IN), .B(n2686), .S(IR_REG_22__SCAN_IN), 
        .Z(n2688) );
  XNOR2_X1 U3410 ( .A(n3074), .B(n2844), .ZN(n2689) );
  NAND2_X1 U3411 ( .A1(n2689), .A2(n3863), .ZN(n4702) );
  INV_X1 U3413 ( .A(n2693), .ZN(n4694) );
  OR2_X1 U3414 ( .A1(n2817), .A2(n4718), .ZN(n3684) );
  NAND2_X1 U3415 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U3416 ( .A1(n4692), .A2(n2694), .ZN(n2696) );
  INV_X1 U3417 ( .A(n3696), .ZN(n2695) );
  NAND2_X1 U3418 ( .A1(n2696), .A2(n2695), .ZN(n3077) );
  NAND2_X1 U3419 ( .A1(n3077), .A2(n3727), .ZN(n2697) );
  XNOR2_X1 U3420 ( .A(n3808), .B(n3732), .ZN(n3078) );
  INV_X1 U3421 ( .A(n3732), .ZN(n3076) );
  OR2_X1 U3422 ( .A1(n3808), .A2(n3076), .ZN(n3733) );
  INV_X1 U3423 ( .A(n3734), .ZN(n2698) );
  INV_X1 U3424 ( .A(n3319), .ZN(n3328) );
  AND2_X1 U3425 ( .A1(n3805), .A2(n3328), .ZN(n3317) );
  OR2_X1 U3426 ( .A1(n3805), .A2(n3328), .ZN(n3749) );
  INV_X1 U3427 ( .A(n3061), .ZN(n2699) );
  NAND2_X1 U3428 ( .A1(n3320), .A2(n2699), .ZN(n3750) );
  NAND2_X1 U3429 ( .A1(n3057), .A2(n3750), .ZN(n2700) );
  OR2_X1 U3430 ( .A1(n3320), .A2(n2699), .ZN(n3739) );
  NAND2_X1 U3431 ( .A1(n2700), .A2(n3739), .ZN(n3161) );
  INV_X1 U3432 ( .A(n3740), .ZN(n2701) );
  OR2_X1 U3433 ( .A1(n3162), .A2(n3118), .ZN(n3743) );
  NAND2_X1 U3434 ( .A1(n3162), .A2(n3118), .ZN(n3751) );
  INV_X1 U3435 ( .A(n3301), .ZN(n2703) );
  AND2_X1 U3436 ( .A1(n3804), .A2(n3310), .ZN(n3746) );
  INV_X1 U3437 ( .A(n3746), .ZN(n2702) );
  OR2_X1 U3438 ( .A1(n3804), .A2(n3310), .ZN(n3744) );
  NAND2_X1 U3439 ( .A1(n2704), .A2(n3744), .ZN(n3279) );
  NAND2_X1 U3440 ( .A1(n4678), .A2(n2367), .ZN(n3758) );
  NAND2_X1 U3441 ( .A1(n3279), .A2(n3758), .ZN(n2705) );
  NAND2_X1 U3442 ( .A1(n3802), .A2(n3349), .ZN(n3372) );
  INV_X1 U3443 ( .A(n3230), .ZN(n3385) );
  NAND2_X1 U3444 ( .A1(n3376), .A2(n3385), .ZN(n2706) );
  NAND2_X1 U3445 ( .A1(n3372), .A2(n2706), .ZN(n3759) );
  INV_X1 U3446 ( .A(n3343), .ZN(n3761) );
  NOR2_X1 U3447 ( .A1(n3759), .A2(n3761), .ZN(n2707) );
  INV_X1 U3448 ( .A(n3759), .ZN(n2710) );
  OR2_X1 U3449 ( .A1(n3802), .A2(n3349), .ZN(n3374) );
  NAND2_X1 U3450 ( .A1(n3341), .A2(n3374), .ZN(n2709) );
  NOR2_X1 U3451 ( .A1(n3376), .A2(n3385), .ZN(n2708) );
  AOI21_X1 U3452 ( .B1(n2710), .B2(n2709), .A(n2708), .ZN(n3724) );
  OR2_X1 U3453 ( .A1(n3425), .A2(n4090), .ZN(n3722) );
  NAND2_X1 U3454 ( .A1(n3425), .A2(n4090), .ZN(n3652) );
  NAND2_X1 U3455 ( .A1(n3722), .A2(n3652), .ZN(n4093) );
  NAND2_X1 U3456 ( .A1(n4044), .A2(n4029), .ZN(n2711) );
  AND2_X1 U3457 ( .A1(n4021), .A2(n2711), .ZN(n2715) );
  NAND2_X1 U34580 ( .A1(n4076), .A2(n4065), .ZN(n4017) );
  INV_X1 U34590 ( .A(n3770), .ZN(n2712) );
  OR2_X1 U3460 ( .A1(n4076), .A2(n4065), .ZN(n4018) );
  NAND2_X1 U3461 ( .A1(n4020), .A2(n4018), .ZN(n2714) );
  NOR2_X1 U3462 ( .A1(n4044), .A2(n4029), .ZN(n2713) );
  AOI21_X1 U3463 ( .B1(n2715), .B2(n2714), .A(n2713), .ZN(n4000) );
  OR2_X1 U3464 ( .A1(n3987), .A2(n4009), .ZN(n2716) );
  AND2_X1 U3465 ( .A1(n3987), .A2(n4009), .ZN(n3775) );
  OR2_X1 U3466 ( .A1(n3973), .A2(n3991), .ZN(n3951) );
  NAND2_X1 U34670 ( .A1(n3954), .A2(n3951), .ZN(n3720) );
  NAND2_X1 U3468 ( .A1(n3973), .A2(n3991), .ZN(n3953) );
  INV_X1 U34690 ( .A(n3953), .ZN(n2718) );
  INV_X1 U3470 ( .A(n3947), .ZN(n3957) );
  NAND2_X1 U34710 ( .A1(n3974), .A2(n3957), .ZN(n3697) );
  NAND2_X1 U3472 ( .A1(n2717), .A2(n3697), .ZN(n3772) );
  AOI21_X1 U34730 ( .B1(n2718), .B2(n3954), .A(n3772), .ZN(n3656) );
  OAI21_X1 U3474 ( .B1(n3984), .B2(n3720), .A(n3656), .ZN(n2719) );
  INV_X1 U34750 ( .A(n3974), .ZN(n3618) );
  NAND2_X1 U3476 ( .A1(n3618), .A2(n3947), .ZN(n3776) );
  OR2_X1 U34770 ( .A1(n3917), .A2(n3936), .ZN(n3777) );
  NOR2_X1 U3478 ( .A1(n3958), .A2(n3482), .ZN(n3678) );
  NOR2_X1 U34790 ( .A1(n3900), .A2(n3914), .ZN(n3893) );
  NOR2_X1 U3480 ( .A1(n3500), .A2(n3904), .ZN(n3702) );
  NOR2_X1 U34810 ( .A1(n3893), .A2(n3702), .ZN(n3785) );
  AND2_X1 U3482 ( .A1(n3500), .A2(n3904), .ZN(n3701) );
  NOR2_X1 U34830 ( .A1(n3522), .A2(n3542), .ZN(n3659) );
  AND2_X1 U3484 ( .A1(n3522), .A2(n3542), .ZN(n3783) );
  NOR2_X2 U34850 ( .A1(n3659), .A2(n3783), .ZN(n3883) );
  INV_X1 U3486 ( .A(n3659), .ZN(n2720) );
  NAND2_X1 U34870 ( .A1(n3882), .A2(n2720), .ZN(n3405) );
  XNOR2_X1 U3488 ( .A(n3405), .B(n3400), .ZN(n2736) );
  INV_X1 U34890 ( .A(n2690), .ZN(n2784) );
  NAND2_X1 U3490 ( .A1(n2784), .A2(n2733), .ZN(n2722) );
  NAND2_X1 U34910 ( .A1(n2844), .A2(n2822), .ZN(n2721) );
  NAND2_X1 U3492 ( .A1(n2421), .A2(REG2_REG_29__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U34930 ( .A1(n2424), .A2(REG0_REG_29__SCAN_IN), .ZN(n2727) );
  OR2_X1 U3494 ( .A1(n2422), .A2(n3414), .ZN(n2726) );
  INV_X1 U34950 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2723) );
  OR2_X1 U3496 ( .A1(n2724), .A2(n2723), .ZN(n2725) );
  NAND4_X1 U34970 ( .A1(n2728), .A2(n2727), .A3(n2726), .A4(n2725), .ZN(n3664)
         );
  OR2_X1 U3498 ( .A1(n2730), .A2(n2729), .ZN(n2732) );
  XNOR2_X1 U34990 ( .A(n2732), .B(n2731), .ZN(n2861) );
  NAND2_X1 U3500 ( .A1(n2861), .A2(n2827), .ZN(n4722) );
  AOI22_X1 U35010 ( .A1(n3664), .A2(n4696), .B1(n4695), .B2(n2364), .ZN(n2735)
         );
  NAND2_X1 U3502 ( .A1(n3522), .A2(n4679), .ZN(n2734) );
  OAI211_X1 U35030 ( .C1(n2736), .C2(n4681), .A(n2735), .B(n2734), .ZN(n3874)
         );
  AOI21_X1 U3504 ( .B1(n3868), .B2(n4809), .A(n3874), .ZN(n2770) );
  NAND2_X1 U35050 ( .A1(n2690), .A2(n3863), .ZN(n2828) );
  NAND2_X1 U35060 ( .A1(n2828), .A2(n2827), .ZN(n2902) );
  NAND2_X1 U35070 ( .A1(n2744), .A2(n4223), .ZN(n2746) );
  NAND2_X1 U35080 ( .A1(n2739), .A2(IR_REG_31__SCAN_IN), .ZN(n2740) );
  OAI21_X1 U35090 ( .B1(IR_REG_23__SCAN_IN), .B2(IR_REG_24__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U35100 ( .A1(n2744), .A2(n2741), .ZN(n2742) );
  INV_X1 U35110 ( .A(n2793), .ZN(n4495) );
  OR2_X1 U35120 ( .A1(n2744), .A2(n4223), .ZN(n2745) );
  NAND2_X1 U35130 ( .A1(n2746), .A2(n2745), .ZN(n2900) );
  NAND2_X1 U35140 ( .A1(n2902), .A2(n2833), .ZN(n2837) );
  NAND2_X1 U35150 ( .A1(n2790), .A2(n2793), .ZN(n2747) );
  MUX2_X1 U35160 ( .A(n2790), .B(n2747), .S(B_REG_SCAN_IN), .Z(n2748) );
  NOR4_X1 U35170 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2756) );
  NOR4_X1 U35180 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2755) );
  INV_X1 U35190 ( .A(D_REG_4__SCAN_IN), .ZN(n4738) );
  INV_X1 U35200 ( .A(D_REG_9__SCAN_IN), .ZN(n4736) );
  INV_X1 U35210 ( .A(D_REG_18__SCAN_IN), .ZN(n4732) );
  INV_X1 U35220 ( .A(D_REG_20__SCAN_IN), .ZN(n4731) );
  NAND4_X1 U35230 ( .A1(n4738), .A2(n4736), .A3(n4732), .A4(n4731), .ZN(n4169)
         );
  NOR4_X1 U35240 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2752) );
  NOR4_X1 U35250 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2751) );
  NOR4_X1 U35260 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2750) );
  NOR4_X1 U35270 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2749) );
  NAND4_X1 U35280 ( .A1(n2752), .A2(n2751), .A3(n2750), .A4(n2749), .ZN(n2753)
         );
  NOR4_X1 U35290 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n4169), 
        .A4(n2753), .ZN(n2754) );
  AND3_X1 U35300 ( .A1(n2756), .A2(n2755), .A3(n2754), .ZN(n2757) );
  NOR2_X1 U35310 ( .A1(n2787), .A2(n2757), .ZN(n3068) );
  NOR2_X1 U35320 ( .A1(n4783), .A2(n2733), .ZN(n2758) );
  OR2_X1 U35330 ( .A1(n2787), .A2(D_REG_1__SCAN_IN), .ZN(n2760) );
  INV_X1 U35340 ( .A(n2788), .ZN(n2762) );
  NAND2_X1 U35350 ( .A1(n2793), .A2(n2762), .ZN(n2759) );
  NAND2_X1 U35360 ( .A1(n2760), .A2(n2759), .ZN(n2814) );
  NAND2_X1 U35370 ( .A1(n2790), .A2(n2762), .ZN(n2763) );
  MUX2_X1 U35380 ( .A(n4303), .B(n2770), .S(n4836), .Z(n2768) );
  OAI21_X1 U35390 ( .B1(n3879), .B2(n3532), .A(n3403), .ZN(n3869) );
  NAND2_X1 U35400 ( .A1(n4836), .A2(n4812), .ZN(n4435) );
  NAND2_X1 U35410 ( .A1(n2768), .A2(n2767), .ZN(U3546) );
  INV_X1 U35420 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2771) );
  MUX2_X1 U35430 ( .A(n2771), .B(n2770), .S(n4824), .Z(n2773) );
  NAND2_X1 U35440 ( .A1(n4824), .A2(n4812), .ZN(n4489) );
  NAND2_X1 U35450 ( .A1(n2773), .A2(n2772), .ZN(U3514) );
  INV_X1 U35460 ( .A(n4742), .ZN(n2789) );
  INV_X2 U35470 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U35480 ( .A(n2774), .B(n3010), .S(STATE_REG_SCAN_IN), .Z(n2775) );
  INV_X1 U35490 ( .A(n2775), .ZN(U3348) );
  INV_X1 U35500 ( .A(n4653), .ZN(n2776) );
  NAND2_X1 U35510 ( .A1(n2776), .A2(STATE_REG_SCAN_IN), .ZN(n2777) );
  OAI21_X1 U35520 ( .B1(STATE_REG_SCAN_IN), .B2(n2591), .A(n2777), .ZN(U3335)
         );
  INV_X1 U35530 ( .A(DATAI_22_), .ZN(n2779) );
  NAND2_X1 U35540 ( .A1(n2844), .A2(STATE_REG_SCAN_IN), .ZN(n2778) );
  OAI21_X1 U35550 ( .B1(STATE_REG_SCAN_IN), .B2(n2779), .A(n2778), .ZN(U3330)
         );
  INV_X1 U35560 ( .A(DATAI_24_), .ZN(n2780) );
  MUX2_X1 U35570 ( .A(n2780), .B(n2790), .S(STATE_REG_SCAN_IN), .Z(n2781) );
  INV_X1 U35580 ( .A(n2781), .ZN(U3328) );
  INV_X1 U35590 ( .A(DATAI_26_), .ZN(n2783) );
  NAND2_X1 U35600 ( .A1(n2788), .A2(STATE_REG_SCAN_IN), .ZN(n2782) );
  OAI21_X1 U35610 ( .B1(STATE_REG_SCAN_IN), .B2(n2783), .A(n2782), .ZN(U3326)
         );
  INV_X1 U35620 ( .A(DATAI_20_), .ZN(n2786) );
  NAND2_X1 U35630 ( .A1(n2784), .A2(STATE_REG_SCAN_IN), .ZN(n2785) );
  OAI21_X1 U35640 ( .B1(STATE_REG_SCAN_IN), .B2(n2786), .A(n2785), .ZN(U3332)
         );
  NAND2_X1 U35650 ( .A1(n2833), .A2(n2787), .ZN(n4739) );
  INV_X1 U35660 ( .A(D_REG_0__SCAN_IN), .ZN(n2791) );
  NOR2_X1 U35670 ( .A1(n2789), .A2(n2788), .ZN(n2792) );
  AOI22_X1 U35680 ( .A1(n4739), .A2(n2791), .B1(n2792), .B2(n2790), .ZN(U3458)
         );
  INV_X1 U35690 ( .A(D_REG_1__SCAN_IN), .ZN(n2794) );
  AOI22_X1 U35700 ( .A1(n4739), .A2(n2794), .B1(n2793), .B2(n2792), .ZN(U3459)
         );
  NAND2_X1 U35710 ( .A1(n2827), .A2(n2900), .ZN(n2795) );
  AND2_X1 U35720 ( .A1(n2795), .A2(n2408), .ZN(n2868) );
  INV_X1 U35730 ( .A(n2868), .ZN(n2796) );
  INV_X1 U35740 ( .A(n2833), .ZN(n2832) );
  NOR2_X1 U35750 ( .A1(n2900), .A2(U3149), .ZN(n3793) );
  INV_X1 U35760 ( .A(n3793), .ZN(n3799) );
  NAND2_X1 U35770 ( .A1(n2832), .A2(n3799), .ZN(n2869) );
  NOR2_X1 U35780 ( .A1(n4671), .A2(U4043), .ZN(U3148) );
  INV_X1 U35790 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U35800 ( .A1(n3320), .A2(U4043), .ZN(n2797) );
  OAI21_X1 U35810 ( .B1(U4043), .B2(n4313), .A(n2797), .ZN(U3556) );
  INV_X1 U3582 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U3583 ( .A1(n4059), .A2(U4043), .ZN(n2798) );
  OAI21_X1 U3584 ( .B1(U4043), .B2(n4323), .A(n2798), .ZN(U3568) );
  INV_X1 U3585 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U3586 ( .A1(n3987), .A2(U4043), .ZN(n2799) );
  OAI21_X1 U3587 ( .B1(U4043), .B2(n4322), .A(n2799), .ZN(U3570) );
  INV_X1 U3588 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U3589 ( .A1(n3425), .A2(U4043), .ZN(n2800) );
  OAI21_X1 U3590 ( .B1(U4043), .B2(n4319), .A(n2800), .ZN(U3565) );
  INV_X1 U3591 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4317) );
  NAND2_X1 U3592 ( .A1(n3120), .A2(U4043), .ZN(n2801) );
  OAI21_X1 U3593 ( .B1(U4043), .B2(n4317), .A(n2801), .ZN(U3557) );
  INV_X1 U3594 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U3595 ( .A1(n3973), .A2(U4043), .ZN(n2802) );
  OAI21_X1 U3596 ( .B1(U4043), .B2(n4348), .A(n2802), .ZN(U3571) );
  INV_X1 U3597 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U3598 ( .A1(n3376), .A2(U4043), .ZN(n2803) );
  OAI21_X1 U3599 ( .B1(U4043), .B2(n4320), .A(n2803), .ZN(U3563) );
  INV_X1 U3600 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U3601 ( .A1(n2424), .A2(REG0_REG_31__SCAN_IN), .ZN(n2807) );
  NAND2_X1 U3602 ( .A1(n2421), .A2(REG2_REG_31__SCAN_IN), .ZN(n2806) );
  INV_X1 U3603 ( .A(REG1_REG_31__SCAN_IN), .ZN(n2804) );
  OR2_X1 U3604 ( .A1(n2724), .A2(n2804), .ZN(n2805) );
  AND3_X1 U3605 ( .A1(n2807), .A2(n2806), .A3(n2805), .ZN(n3704) );
  INV_X1 U3606 ( .A(n3704), .ZN(n4103) );
  NAND2_X1 U3607 ( .A1(n4103), .A2(U4043), .ZN(n2808) );
  OAI21_X1 U3608 ( .B1(U4043), .B2(n4356), .A(n2808), .ZN(U3581) );
  INV_X1 U3609 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U3610 ( .A1(n3162), .A2(U4043), .ZN(n2809) );
  OAI21_X1 U3611 ( .B1(U4043), .B2(n4316), .A(n2809), .ZN(U3558) );
  INV_X1 U3612 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4337) );
  NAND2_X1 U3613 ( .A1(n2817), .A2(U4043), .ZN(n2810) );
  OAI21_X1 U3614 ( .B1(U4043), .B2(n4337), .A(n2810), .ZN(U3550) );
  INV_X1 U3615 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U3616 ( .A1(n2905), .A2(U4043), .ZN(n2811) );
  OAI21_X1 U3617 ( .B1(U4043), .B2(n4314), .A(n2811), .ZN(U3552) );
  INV_X1 U3618 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U3619 ( .A1(n2841), .A2(U4043), .ZN(n2812) );
  OAI21_X1 U3620 ( .B1(U4043), .B2(n4336), .A(n2812), .ZN(U3551) );
  INV_X1 U3621 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4347) );
  NAND2_X1 U3622 ( .A1(n3974), .A2(U4043), .ZN(n2813) );
  OAI21_X1 U3623 ( .B1(U4043), .B2(n4347), .A(n2813), .ZN(U3573) );
  NOR2_X1 U3624 ( .A1(n3068), .A2(n2814), .ZN(n2815) );
  NAND2_X1 U3625 ( .A1(n2816), .A2(n2815), .ZN(n2835) );
  NAND4_X1 U3626 ( .A1(n2976), .A2(n2844), .A3(n4742), .A4(n3863), .ZN(n3797)
         );
  NOR2_X1 U3627 ( .A1(n2835), .A2(n3797), .ZN(n2854) );
  NAND2_X2 U3628 ( .A1(n2854), .A2(n2861), .ZN(n4514) );
  NAND2_X1 U3629 ( .A1(n2817), .A2(n2925), .ZN(n2819) );
  NAND2_X1 U3630 ( .A1(n4708), .A2(n2132), .ZN(n2818) );
  NAND2_X1 U3631 ( .A1(n2819), .A2(n2818), .ZN(n2851) );
  INV_X1 U3632 ( .A(n2851), .ZN(n2821) );
  NAND2_X1 U3633 ( .A1(n2821), .A2(n2370), .ZN(n2850) );
  NOR2_X2 U3634 ( .A1(n3084), .A2(n3494), .ZN(n2962) );
  NAND2_X1 U3635 ( .A1(n2817), .A2(n2962), .ZN(n2826) );
  AOI22_X1 U3636 ( .A1(n4708), .A2(n2925), .B1(IR_REG_0__SCAN_IN), .B2(n2824), 
        .ZN(n2825) );
  NAND2_X1 U3637 ( .A1(n2826), .A2(n2825), .ZN(n2849) );
  XOR2_X1 U3638 ( .A(n2850), .B(n2849), .Z(n2862) );
  INV_X1 U3639 ( .A(n2827), .ZN(n2830) );
  NAND2_X1 U3640 ( .A1(n2828), .A2(n4716), .ZN(n2829) );
  NAND3_X1 U3641 ( .A1(n2833), .A2(n2830), .A3(n2829), .ZN(n2831) );
  NAND2_X1 U3642 ( .A1(n2862), .A2(n4524), .ZN(n2839) );
  NOR3_X1 U3643 ( .A1(n2835), .A2(n4675), .A3(n2832), .ZN(n2834) );
  NAND3_X2 U3644 ( .A1(n4820), .A2(n3717), .A3(n2833), .ZN(n4050) );
  NAND2_X1 U3645 ( .A1(n4716), .A2(n2822), .ZN(n2836) );
  OAI21_X1 U3646 ( .B1(n4695), .B2(n2836), .A(n2835), .ZN(n2903) );
  INV_X1 U3647 ( .A(n2837), .ZN(n3069) );
  NAND2_X1 U3648 ( .A1(n2903), .A2(n3069), .ZN(n3632) );
  AOI22_X1 U3649 ( .A1(n4518), .A2(n4708), .B1(REG3_REG_0__SCAN_IN), .B2(n3632), .ZN(n2838) );
  OAI211_X1 U3650 ( .C1(n2402), .C2(n4514), .A(n2839), .B(n2838), .ZN(U3229)
         );
  INV_X1 U3651 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U3652 ( .A1(n3917), .A2(U4043), .ZN(n2840) );
  OAI21_X1 U3653 ( .B1(U4043), .B2(n4351), .A(n2840), .ZN(U3574) );
  NAND2_X1 U3654 ( .A1(n2841), .A2(n2925), .ZN(n2843) );
  NAND2_X1 U3655 ( .A1(n2401), .A2(n3455), .ZN(n2842) );
  NAND2_X1 U3656 ( .A1(n2843), .A2(n2842), .ZN(n2846) );
  NAND2_X1 U3657 ( .A1(n2844), .A2(n3863), .ZN(n2845) );
  NAND2_X2 U3658 ( .A1(n3074), .A2(n2845), .ZN(n3526) );
  NOR2_X1 U3659 ( .A1(n2847), .A2(n3520), .ZN(n2848) );
  AOI21_X1 U3660 ( .B1(n2841), .B2(n2962), .A(n2848), .ZN(n2916) );
  NAND2_X1 U3661 ( .A1(n2850), .A2(n2849), .ZN(n2853) );
  OR2_X1 U3662 ( .A1(n2851), .A2(n3526), .ZN(n2852) );
  NAND2_X1 U3663 ( .A1(n2853), .A2(n2852), .ZN(n2919) );
  XNOR2_X1 U3664 ( .A(n2920), .B(n2919), .ZN(n2857) );
  AOI22_X1 U3665 ( .A1(n4518), .A2(n2401), .B1(REG3_REG_1__SCAN_IN), .B2(n3632), .ZN(n2856) );
  NAND2_X2 U3666 ( .A1(n2854), .A2(n4494), .ZN(n4515) );
  INV_X1 U3667 ( .A(n4515), .ZN(n3635) );
  INV_X1 U3668 ( .A(n4514), .ZN(n3634) );
  AOI22_X1 U3669 ( .A1(n3635), .A2(n2817), .B1(n3634), .B2(n2905), .ZN(n2855)
         );
  OAI211_X1 U3670 ( .C1(n2857), .C2(n3626), .A(n2856), .B(n2855), .ZN(U3219)
         );
  XNOR2_X1 U3671 ( .A(n2858), .B(IR_REG_27__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U3672 ( .A1(n4494), .A2(n4540), .ZN(n3796) );
  INV_X1 U3673 ( .A(n3796), .ZN(n2865) );
  INV_X1 U3674 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U3675 ( .A1(n4765), .A2(n4727), .ZN(n3813) );
  NAND2_X1 U3676 ( .A1(n4540), .A2(n4727), .ZN(n2859) );
  NAND2_X1 U3677 ( .A1(n4494), .A2(n2859), .ZN(n4538) );
  NAND2_X1 U3678 ( .A1(n4538), .A2(n4765), .ZN(n2860) );
  NAND2_X1 U3679 ( .A1(n2860), .A2(U4043), .ZN(n2864) );
  NOR3_X1 U3680 ( .A1(n2862), .A2(n4540), .A3(n2861), .ZN(n2863) );
  AOI211_X1 U3681 ( .C1(n2865), .C2(n3813), .A(n2864), .B(n2863), .ZN(n2898)
         );
  INV_X1 U3682 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2866) );
  MUX2_X1 U3683 ( .A(n2866), .B(REG2_REG_2__SCAN_IN), .S(n2877), .Z(n2871) );
  INV_X1 U3684 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4304) );
  MUX2_X1 U3685 ( .A(n4304), .B(REG2_REG_1__SCAN_IN), .S(n2873), .Z(n3814) );
  INV_X1 U3686 ( .A(n2873), .ZN(n4500) );
  NAND2_X1 U3687 ( .A1(n4500), .A2(REG2_REG_1__SCAN_IN), .ZN(n2867) );
  NAND2_X1 U3688 ( .A1(n3812), .A2(n2867), .ZN(n2870) );
  NAND2_X1 U3689 ( .A1(n2869), .A2(n2868), .ZN(n4543) );
  INV_X1 U3690 ( .A(n4654), .ZN(n4666) );
  OAI211_X1 U3691 ( .C1(n2871), .C2(n2870), .A(n4666), .B(n2884), .ZN(n2881)
         );
  AND2_X1 U3692 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3810)
         );
  NAND2_X1 U3693 ( .A1(n4500), .A2(REG1_REG_1__SCAN_IN), .ZN(n2874) );
  NAND2_X1 U3694 ( .A1(n3809), .A2(n2874), .ZN(n2875) );
  OR2_X1 U3695 ( .A1(n4543), .A2(n4540), .ZN(n4659) );
  OAI211_X1 U3696 ( .C1(n2876), .C2(n2875), .A(n4662), .B(n2890), .ZN(n2880)
         );
  AOI22_X1 U3697 ( .A1(n4671), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2879) );
  INV_X1 U3698 ( .A(n4669), .ZN(n4563) );
  NAND2_X1 U3699 ( .A1(n4563), .A2(n4499), .ZN(n2878) );
  NAND4_X1 U3700 ( .A1(n2881), .A2(n2880), .A3(n2879), .A4(n2878), .ZN(n2882)
         );
  OR2_X1 U3701 ( .A1(n2898), .A2(n2882), .ZN(U3242) );
  INV_X1 U3702 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4307) );
  INV_X1 U3703 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3821) );
  AOI211_X1 U3704 ( .C1(n4307), .C2(n2888), .A(n3023), .B(n4654), .ZN(n2897)
         );
  NAND2_X1 U3705 ( .A1(n4499), .A2(REG1_REG_2__SCAN_IN), .ZN(n2889) );
  NAND2_X1 U3706 ( .A1(n2890), .A2(n2889), .ZN(n2891) );
  NAND2_X1 U3707 ( .A1(n3826), .A2(REG1_REG_3__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U3708 ( .A1(n2891), .A2(n4498), .ZN(n2892) );
  NAND2_X1 U3709 ( .A1(n3825), .A2(n2892), .ZN(n3011) );
  OAI211_X1 U3710 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2893), .A(n4662), .B(n3013), 
        .ZN(n2895) );
  AND2_X1 U3711 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2940) );
  AOI21_X1 U3712 ( .B1(n4671), .B2(ADDR_REG_4__SCAN_IN), .A(n2940), .ZN(n2894)
         );
  OAI211_X1 U3713 ( .C1(n4669), .C2(n3010), .A(n2895), .B(n2894), .ZN(n2896)
         );
  OR3_X1 U3714 ( .A1(n2898), .A2(n2897), .A3(n2896), .ZN(U3244) );
  INV_X1 U3715 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U3716 ( .A1(n3500), .A2(U4043), .ZN(n2899) );
  OAI21_X1 U3717 ( .B1(U4043), .B2(n4350), .A(n2899), .ZN(U3576) );
  NAND4_X1 U3718 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n2904)
         );
  NAND2_X1 U3719 ( .A1(n2905), .A2(n2925), .ZN(n2907) );
  NAND2_X1 U3720 ( .A1(n3633), .A2(n2132), .ZN(n2906) );
  NAND2_X1 U3721 ( .A1(n2907), .A2(n2906), .ZN(n2908) );
  XNOR2_X1 U3722 ( .A(n2908), .B(n3518), .ZN(n2913) );
  INV_X1 U3723 ( .A(n2913), .ZN(n2911) );
  NOR2_X1 U3724 ( .A1(n3110), .A2(n3520), .ZN(n2909) );
  AOI21_X1 U3725 ( .B1(n2905), .B2(n2962), .A(n2909), .ZN(n2912) );
  INV_X1 U3726 ( .A(n2912), .ZN(n2910) );
  NAND2_X1 U3727 ( .A1(n2911), .A2(n2910), .ZN(n2914) );
  NAND2_X1 U3728 ( .A1(n2913), .A2(n2912), .ZN(n2921) );
  INV_X1 U3729 ( .A(n2915), .ZN(n2917) );
  NOR2_X1 U3730 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  AOI21_X1 U3731 ( .B1(n2920), .B2(n2919), .A(n2918), .ZN(n3628) );
  NAND2_X1 U3732 ( .A1(n3629), .A2(n3628), .ZN(n3630) );
  NAND2_X1 U3733 ( .A1(n3630), .A2(n2921), .ZN(n2945) );
  NAND2_X1 U3734 ( .A1(n3732), .A2(n2132), .ZN(n2922) );
  NAND2_X1 U3735 ( .A1(n2923), .A2(n2922), .ZN(n2924) );
  XNOR2_X1 U3736 ( .A(n2924), .B(n3526), .ZN(n2927) );
  AND2_X1 U3737 ( .A1(n3732), .A2(n2925), .ZN(n2926) );
  AOI21_X1 U3738 ( .B1(n3808), .B2(n3499), .A(n2926), .ZN(n2928) );
  XNOR2_X1 U3739 ( .A(n2927), .B(n2928), .ZN(n2946) );
  NAND2_X1 U3740 ( .A1(n2945), .A2(n2946), .ZN(n2936) );
  INV_X1 U3741 ( .A(n2927), .ZN(n2929) );
  NAND2_X1 U3742 ( .A1(n2929), .A2(n2928), .ZN(n2934) );
  AND2_X1 U3743 ( .A1(n2936), .A2(n2934), .ZN(n2938) );
  NAND2_X1 U3744 ( .A1(n3806), .A2(n2925), .ZN(n2931) );
  NAND2_X1 U3745 ( .A1(n2941), .A2(n2132), .ZN(n2930) );
  NOR2_X1 U3746 ( .A1(n3149), .A2(n3520), .ZN(n2933) );
  AOI21_X1 U3747 ( .B1(n3806), .B2(n3499), .A(n2933), .ZN(n2955) );
  XNOR2_X1 U3748 ( .A(n2954), .B(n2955), .ZN(n2937) );
  NAND2_X1 U3749 ( .A1(n2936), .A2(n2935), .ZN(n2958) );
  OAI211_X1 U3750 ( .C1(n2938), .C2(n2937), .A(n4524), .B(n2958), .ZN(n2943)
         );
  INV_X1 U3751 ( .A(n3808), .ZN(n3731) );
  INV_X1 U3752 ( .A(n3805), .ZN(n3143) );
  OAI22_X1 U3753 ( .A1(n3731), .A2(n4515), .B1(n4514), .B2(n3143), .ZN(n2939)
         );
  AOI211_X1 U3754 ( .C1(n2941), .C2(n4518), .A(n2940), .B(n2939), .ZN(n2942)
         );
  OAI211_X1 U3755 ( .C1(n4528), .C2(n3150), .A(n2943), .B(n2942), .ZN(U3227)
         );
  INV_X1 U3756 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4357) );
  NAND2_X1 U3757 ( .A1(n3664), .A2(U4043), .ZN(n2944) );
  OAI21_X1 U3758 ( .B1(U4043), .B2(n4357), .A(n2944), .ZN(U3579) );
  OAI21_X1 U3759 ( .B1(n2946), .B2(n2945), .A(n2936), .ZN(n2947) );
  NAND2_X1 U3760 ( .A1(n2947), .A2(n4524), .ZN(n2951) );
  NAND2_X1 U3761 ( .A1(U3149), .A2(REG3_REG_3__SCAN_IN), .ZN(n3823) );
  INV_X1 U3762 ( .A(n3823), .ZN(n2949) );
  INV_X1 U3763 ( .A(n3806), .ZN(n3322) );
  OAI22_X1 U3764 ( .A1(n3322), .A2(n4514), .B1(n4515), .B2(n2419), .ZN(n2948)
         );
  AOI211_X1 U3765 ( .C1(n3732), .C2(n4518), .A(n2949), .B(n2948), .ZN(n2950)
         );
  OAI211_X1 U3766 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4528), .A(n2951), .B(n2950), 
        .ZN(U3215) );
  INV_X1 U3767 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U3768 ( .A1(n3522), .A2(U4043), .ZN(n2952) );
  OAI21_X1 U3769 ( .B1(U4043), .B2(n4354), .A(n2952), .ZN(U3577) );
  INV_X1 U3770 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U3771 ( .A1(n3887), .A2(U4043), .ZN(n2953) );
  OAI21_X1 U3772 ( .B1(U4043), .B2(n4353), .A(n2953), .ZN(U3578) );
  INV_X1 U3773 ( .A(n2955), .ZN(n2956) );
  NAND2_X1 U3774 ( .A1(n2954), .A2(n2956), .ZN(n2957) );
  NAND2_X1 U3775 ( .A1(n2958), .A2(n2957), .ZN(n2970) );
  NAND2_X1 U3776 ( .A1(n3805), .A2(n2976), .ZN(n2960) );
  NAND2_X1 U3777 ( .A1(n3319), .A2(n2132), .ZN(n2959) );
  NAND2_X1 U3778 ( .A1(n2960), .A2(n2959), .ZN(n2961) );
  XNOR2_X1 U3779 ( .A(n2961), .B(n3526), .ZN(n2973) );
  AND2_X1 U3780 ( .A1(n3319), .A2(n2976), .ZN(n2963) );
  AOI21_X1 U3781 ( .B1(n3805), .B2(n3499), .A(n2963), .ZN(n2971) );
  XNOR2_X1 U3782 ( .A(n2973), .B(n2971), .ZN(n2969) );
  XOR2_X1 U3783 ( .A(n2970), .B(n2969), .Z(n2964) );
  NAND2_X1 U3784 ( .A1(n2964), .A2(n4524), .ZN(n2968) );
  NAND2_X1 U3785 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4553) );
  INV_X1 U3786 ( .A(n4553), .ZN(n2966) );
  INV_X1 U3787 ( .A(n3320), .ZN(n3005) );
  OAI22_X1 U3788 ( .A1(n3322), .A2(n4515), .B1(n4514), .B2(n3005), .ZN(n2965)
         );
  AOI211_X1 U3789 ( .C1(n3319), .C2(n4518), .A(n2966), .B(n2965), .ZN(n2967)
         );
  OAI211_X1 U3790 ( .C1(n4528), .C2(n3330), .A(n2968), .B(n2967), .ZN(U3224)
         );
  NAND2_X1 U3791 ( .A1(n2970), .A2(n2969), .ZN(n2975) );
  INV_X1 U3792 ( .A(n2971), .ZN(n2972) );
  NAND2_X1 U3793 ( .A1(n2973), .A2(n2972), .ZN(n2974) );
  NAND2_X1 U3794 ( .A1(n2975), .A2(n2974), .ZN(n2995) );
  NAND2_X1 U3795 ( .A1(n3320), .A2(n2976), .ZN(n2978) );
  NAND2_X1 U3796 ( .A1(n3061), .A2(n2132), .ZN(n2977) );
  NAND2_X1 U3797 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
  XNOR2_X1 U3798 ( .A(n2979), .B(n3526), .ZN(n2982) );
  NAND2_X1 U3799 ( .A1(n3320), .A2(n3499), .ZN(n2981) );
  NAND2_X1 U3800 ( .A1(n3061), .A2(n2976), .ZN(n2980) );
  NAND2_X1 U3801 ( .A1(n2981), .A2(n2980), .ZN(n2983) );
  AND2_X1 U3802 ( .A1(n2982), .A2(n2983), .ZN(n2994) );
  INV_X1 U3803 ( .A(n2994), .ZN(n2986) );
  INV_X1 U3804 ( .A(n2982), .ZN(n2985) );
  INV_X1 U3805 ( .A(n2983), .ZN(n2984) );
  NAND2_X1 U3806 ( .A1(n2985), .A2(n2984), .ZN(n2996) );
  NAND2_X1 U3807 ( .A1(n2986), .A2(n2996), .ZN(n2987) );
  XNOR2_X1 U3808 ( .A(n2995), .B(n2987), .ZN(n2988) );
  NAND2_X1 U3809 ( .A1(n2988), .A2(n4524), .ZN(n2993) );
  NAND2_X1 U3810 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n4564) );
  INV_X1 U3811 ( .A(n4564), .ZN(n2991) );
  INV_X1 U3812 ( .A(n3120), .ZN(n2989) );
  OAI22_X1 U3813 ( .A1(n2989), .A2(n4514), .B1(n4515), .B2(n3143), .ZN(n2990)
         );
  AOI211_X1 U3814 ( .C1(n3061), .C2(n4518), .A(n2991), .B(n2990), .ZN(n2992)
         );
  OAI211_X1 U3815 ( .C1(n4528), .C2(n3233), .A(n2993), .B(n2992), .ZN(U3236)
         );
  NAND2_X1 U3816 ( .A1(n3120), .A2(n2976), .ZN(n2998) );
  NAND2_X1 U3817 ( .A1(n3007), .A2(n2132), .ZN(n2997) );
  NAND2_X1 U3818 ( .A1(n2998), .A2(n2997), .ZN(n2999) );
  XNOR2_X1 U3819 ( .A(n2999), .B(n3518), .ZN(n3038) );
  NOR2_X1 U3820 ( .A1(n3165), .A2(n3520), .ZN(n3000) );
  AOI21_X1 U3821 ( .B1(n3120), .B2(n3499), .A(n3000), .ZN(n3039) );
  XNOR2_X1 U3822 ( .A(n3038), .B(n3039), .ZN(n3002) );
  AOI21_X1 U3823 ( .B1(n3001), .B2(n3002), .A(n3626), .ZN(n3004) );
  NAND2_X1 U3824 ( .A1(n3004), .A2(n3043), .ZN(n3009) );
  INV_X1 U3825 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4385) );
  NOR2_X1 U3826 ( .A1(STATE_REG_SCAN_IN), .A2(n4385), .ZN(n4571) );
  INV_X1 U3827 ( .A(n3162), .ZN(n3304) );
  OAI22_X1 U3828 ( .A1(n3005), .A2(n4515), .B1(n4514), .B2(n3304), .ZN(n3006)
         );
  AOI211_X1 U3829 ( .C1(n3007), .C2(n4518), .A(n4571), .B(n3006), .ZN(n3008)
         );
  OAI211_X1 U3830 ( .C1(n4528), .C2(n3169), .A(n3009), .B(n3008), .ZN(U3210)
         );
  INV_X1 U3831 ( .A(n4497), .ZN(n3037) );
  INV_X1 U3832 ( .A(n3010), .ZN(n3025) );
  INV_X1 U3833 ( .A(n4552), .ZN(n4763) );
  AOI22_X1 U3834 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4763), .B1(n4552), .B2(n2448), .ZN(n4546) );
  INV_X1 U3835 ( .A(n4760), .ZN(n3026) );
  NOR2_X1 U3836 ( .A1(n3014), .A2(n3026), .ZN(n3015) );
  XNOR2_X1 U3837 ( .A(n3026), .B(n3014), .ZN(n4557) );
  NAND2_X1 U3838 ( .A1(n3030), .A2(n3016), .ZN(n3017) );
  INV_X1 U3839 ( .A(n3030), .ZN(n4757) );
  NAND2_X1 U3840 ( .A1(n3017), .A2(n4585), .ZN(n3020) );
  MUX2_X1 U3841 ( .A(REG1_REG_9__SCAN_IN), .B(n3018), .S(n4497), .Z(n3019) );
  NAND2_X1 U3842 ( .A1(n3019), .A2(n3020), .ZN(n3240) );
  OAI211_X1 U3843 ( .C1(n3020), .C2(n3019), .A(n4662), .B(n3240), .ZN(n3036)
         );
  NOR2_X1 U3844 ( .A1(STATE_REG_SCAN_IN), .A2(n3021), .ZN(n3099) );
  INV_X1 U3845 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4581) );
  INV_X1 U3846 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4560) );
  INV_X1 U3847 ( .A(n3022), .ZN(n3024) );
  INV_X1 U3848 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U3849 ( .A1(REG2_REG_5__SCAN_IN), .A2(n4763), .B1(n4552), .B2(n4306), .ZN(n4549) );
  NOR2_X1 U3850 ( .A1(n3027), .A2(n3026), .ZN(n3028) );
  INV_X1 U3851 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U3852 ( .A1(REG2_REG_7__SCAN_IN), .A2(n4578), .B1(n4758), .B2(n4271), .ZN(n4569) );
  NOR2_X1 U3853 ( .A1(n3031), .A2(n4757), .ZN(n3032) );
  INV_X1 U3854 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3313) );
  MUX2_X1 U3855 ( .A(n3313), .B(REG2_REG_9__SCAN_IN), .S(n4497), .Z(n3033) );
  AOI211_X1 U3856 ( .C1(n2172), .C2(n3033), .A(n3248), .B(n4654), .ZN(n3034)
         );
  AOI211_X1 U3857 ( .C1(n4671), .C2(ADDR_REG_9__SCAN_IN), .A(n3099), .B(n3034), 
        .ZN(n3035) );
  OAI211_X1 U3858 ( .C1(n4669), .C2(n3037), .A(n3036), .B(n3035), .ZN(U3249)
         );
  INV_X1 U3859 ( .A(n3038), .ZN(n3041) );
  INV_X1 U3860 ( .A(n3039), .ZN(n3040) );
  NAND2_X1 U3861 ( .A1(n3041), .A2(n3040), .ZN(n3042) );
  NAND2_X1 U3862 ( .A1(n3162), .A2(n3499), .ZN(n3045) );
  NAND2_X1 U3863 ( .A1(n3046), .A2(n2976), .ZN(n3044) );
  NAND2_X1 U3864 ( .A1(n3045), .A2(n3044), .ZN(n3093) );
  NAND2_X1 U3865 ( .A1(n3162), .A2(n2976), .ZN(n3048) );
  NAND2_X1 U3866 ( .A1(n3046), .A2(n2132), .ZN(n3047) );
  NAND2_X1 U3867 ( .A1(n3048), .A2(n3047), .ZN(n3049) );
  XNOR2_X1 U3868 ( .A(n3049), .B(n3526), .ZN(n3092) );
  XOR2_X1 U3869 ( .A(n3093), .B(n3092), .Z(n3050) );
  XNOR2_X1 U3870 ( .A(n3094), .B(n3050), .ZN(n3055) );
  INV_X1 U3871 ( .A(n3295), .ZN(n3053) );
  AOI22_X1 U3872 ( .A1(n3635), .A2(n3120), .B1(n3634), .B2(n3804), .ZN(n3051)
         );
  NAND2_X1 U3873 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4582) );
  OAI211_X1 U3874 ( .C1(n3620), .C2(n3118), .A(n3051), .B(n4582), .ZN(n3052)
         );
  AOI21_X1 U3875 ( .B1(n3053), .B2(n3623), .A(n3052), .ZN(n3054) );
  OAI21_X1 U3876 ( .B1(n3055), .B2(n3626), .A(n3054), .ZN(U3218) );
  NAND2_X1 U3877 ( .A1(n3739), .A2(n3750), .ZN(n3680) );
  XOR2_X1 U3878 ( .A(n3056), .B(n3680), .Z(n3234) );
  XOR2_X1 U3879 ( .A(n3680), .B(n3057), .Z(n3060) );
  AOI22_X1 U3880 ( .A1(n3120), .A2(n4696), .B1(n3061), .B2(n4695), .ZN(n3058)
         );
  OAI21_X1 U3881 ( .B1(n3143), .B2(n4698), .A(n3058), .ZN(n3059) );
  AOI21_X1 U3882 ( .B1(n3060), .B2(n4719), .A(n3059), .ZN(n3239) );
  OAI21_X1 U3883 ( .B1(n3234), .B2(n4801), .A(n3239), .ZN(n3065) );
  NAND2_X1 U3884 ( .A1(n3065), .A2(n4836), .ZN(n3064) );
  AND2_X1 U3885 ( .A1(n3327), .A2(n3061), .ZN(n3062) );
  NOR2_X1 U3886 ( .A1(n3159), .A2(n3062), .ZN(n3237) );
  INV_X1 U3887 ( .A(n4435), .ZN(n4112) );
  NAND2_X1 U3888 ( .A1(n3237), .A2(n4112), .ZN(n3063) );
  OAI211_X1 U3889 ( .C1(n4836), .C2(n2456), .A(n3064), .B(n3063), .ZN(U3524)
         );
  INV_X1 U3890 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4364) );
  NAND2_X1 U3891 ( .A1(n3065), .A2(n4824), .ZN(n3067) );
  INV_X1 U3892 ( .A(n4489), .ZN(n4449) );
  NAND2_X1 U3893 ( .A1(n3237), .A2(n4449), .ZN(n3066) );
  OAI211_X1 U3894 ( .C1(n4824), .C2(n4364), .A(n3067), .B(n3066), .ZN(U3479)
         );
  INV_X1 U3895 ( .A(n3068), .ZN(n3071) );
  NAND4_X1 U3896 ( .A1(n3072), .A2(n3071), .A3(n3070), .A4(n3069), .ZN(n3073)
         );
  NOR2_X1 U3897 ( .A1(n3074), .A2(n3863), .ZN(n3075) );
  NAND2_X1 U3898 ( .A1(n4089), .A2(n3075), .ZN(n4712) );
  OAI22_X1 U3899 ( .A1(n3322), .A2(n4722), .B1(n3076), .B2(n4675), .ZN(n3082)
         );
  NAND3_X1 U3900 ( .A1(n3077), .A2(n3727), .A3(n2336), .ZN(n3079) );
  AOI21_X1 U3901 ( .B1(n3080), .B2(n3079), .A(n4681), .ZN(n3081) );
  AOI211_X1 U3902 ( .C1(n4679), .C2(n2905), .A(n3082), .B(n3081), .ZN(n3083)
         );
  OAI21_X1 U3903 ( .B1(n4784), .B2(n4702), .A(n3083), .ZN(n4785) );
  NAND2_X1 U3904 ( .A1(n4785), .A2(n4534), .ZN(n3087) );
  AOI21_X1 U3905 ( .B1(n3732), .B2(n4777), .A(n2175), .ZN(n4787) );
  OAI22_X1 U3906 ( .A1(n4534), .A2(n3821), .B1(n4050), .B2(REG3_REG_3__SCAN_IN), .ZN(n3085) );
  AOI21_X1 U3907 ( .B1(n4787), .B2(n4689), .A(n3085), .ZN(n3086) );
  OAI211_X1 U3908 ( .C1(n4784), .C2(n4712), .A(n3087), .B(n3086), .ZN(U3287)
         );
  NAND2_X1 U3909 ( .A1(n3804), .A2(n2976), .ZN(n3089) );
  NAND2_X1 U3910 ( .A1(n3302), .A2(n2132), .ZN(n3088) );
  NAND2_X1 U3911 ( .A1(n3089), .A2(n3088), .ZN(n3090) );
  XNOR2_X1 U3912 ( .A(n3090), .B(n3518), .ZN(n3128) );
  AND2_X1 U3913 ( .A1(n3302), .A2(n2976), .ZN(n3091) );
  AOI21_X1 U3914 ( .B1(n3804), .B2(n3499), .A(n3091), .ZN(n3127) );
  XNOR2_X1 U3915 ( .A(n3128), .B(n3127), .ZN(n3186) );
  OAI21_X1 U3916 ( .B1(n3094), .B2(n3093), .A(n3092), .ZN(n3096) );
  NAND2_X1 U3917 ( .A1(n3094), .A2(n3093), .ZN(n3095) );
  NAND2_X1 U3918 ( .A1(n3096), .A2(n3095), .ZN(n3188) );
  OR2_X1 U3919 ( .A1(n3188), .A2(n3186), .ZN(n3134) );
  INV_X1 U3920 ( .A(n3134), .ZN(n3097) );
  AOI21_X1 U3921 ( .B1(n3186), .B2(n3188), .A(n3097), .ZN(n3103) );
  INV_X1 U3922 ( .A(n4678), .ZN(n3211) );
  OAI22_X1 U3923 ( .A1(n3304), .A2(n4515), .B1(n4514), .B2(n3211), .ZN(n3098)
         );
  AOI211_X1 U3924 ( .C1(n3302), .C2(n4518), .A(n3099), .B(n3098), .ZN(n3102)
         );
  INV_X1 U3925 ( .A(n3312), .ZN(n3100) );
  NAND2_X1 U3926 ( .A1(n3623), .A2(n3100), .ZN(n3101) );
  OAI211_X1 U3927 ( .C1(n3103), .C2(n3626), .A(n3102), .B(n3101), .ZN(U3228)
         );
  OAI21_X1 U3928 ( .B1(n3104), .B2(n3696), .A(n3105), .ZN(n4779) );
  INV_X1 U3929 ( .A(n4779), .ZN(n3115) );
  INV_X1 U3930 ( .A(n4702), .ZN(n4720) );
  AOI22_X1 U3931 ( .A1(n3808), .A2(n4696), .B1(n4695), .B2(n3633), .ZN(n3106)
         );
  OAI21_X1 U3932 ( .B1(n2402), .B2(n4698), .A(n3106), .ZN(n3109) );
  NAND3_X1 U3933 ( .A1(n4692), .A2(n3696), .A3(n2694), .ZN(n3107) );
  AOI21_X1 U3934 ( .B1(n3077), .B2(n3107), .A(n4681), .ZN(n3108) );
  AOI211_X1 U3935 ( .C1(n4720), .C2(n4779), .A(n3109), .B(n3108), .ZN(n4781)
         );
  MUX2_X1 U3936 ( .A(n2866), .B(n4781), .S(n4534), .Z(n3114) );
  INV_X1 U3937 ( .A(n4777), .ZN(n3111) );
  NOR2_X1 U3938 ( .A1(n4707), .A2(n3110), .ZN(n4776) );
  NOR3_X1 U3939 ( .A1(n4711), .A2(n3111), .A3(n4776), .ZN(n3112) );
  AOI21_X1 U3940 ( .B1(n4724), .B2(REG3_REG_2__SCAN_IN), .A(n3112), .ZN(n3113)
         );
  OAI211_X1 U3941 ( .C1(n3115), .C2(n4712), .A(n3114), .B(n3113), .ZN(U3288)
         );
  OAI21_X1 U3942 ( .B1(n3157), .B2(n3118), .A(n3308), .ZN(n3294) );
  INV_X1 U3943 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U3944 ( .A1(n3743), .A2(n3751), .ZN(n3693) );
  XOR2_X1 U3945 ( .A(n3116), .B(n3693), .Z(n3298) );
  XOR2_X1 U3946 ( .A(n3117), .B(n3693), .Z(n3122) );
  OAI22_X1 U3947 ( .A1(n3138), .A2(n4722), .B1(n4675), .B2(n3118), .ZN(n3119)
         );
  AOI21_X1 U3948 ( .B1(n4679), .B2(n3120), .A(n3119), .ZN(n3121) );
  OAI21_X1 U3949 ( .B1(n3122), .B2(n4681), .A(n3121), .ZN(n3293) );
  AOI21_X1 U3950 ( .B1(n3298), .B2(n4809), .A(n3293), .ZN(n3125) );
  MUX2_X1 U3951 ( .A(n3123), .B(n3125), .S(n4824), .Z(n3124) );
  OAI21_X1 U3952 ( .B1(n3294), .B2(n4489), .A(n3124), .ZN(U3483) );
  MUX2_X1 U3953 ( .A(n2485), .B(n3125), .S(n4836), .Z(n3126) );
  OAI21_X1 U3954 ( .B1(n3294), .B2(n4435), .A(n3126), .ZN(U3526) );
  NAND2_X1 U3955 ( .A1(n3128), .A2(n3127), .ZN(n3133) );
  AND2_X1 U3956 ( .A1(n3134), .A2(n3133), .ZN(n3136) );
  NAND2_X1 U3957 ( .A1(n4678), .A2(n2976), .ZN(n3130) );
  NAND2_X1 U3958 ( .A1(n3285), .A2(n2132), .ZN(n3129) );
  NAND2_X1 U3959 ( .A1(n3130), .A2(n3129), .ZN(n3131) );
  XNOR2_X1 U3960 ( .A(n3131), .B(n3526), .ZN(n3179) );
  AND2_X1 U3961 ( .A1(n3285), .A2(n2976), .ZN(n3132) );
  AOI21_X1 U3962 ( .B1(n4678), .B2(n3499), .A(n3132), .ZN(n3177) );
  XNOR2_X1 U3963 ( .A(n3179), .B(n3177), .ZN(n3135) );
  AND2_X1 U3964 ( .A1(n3135), .A2(n3133), .ZN(n3189) );
  NAND2_X1 U3965 ( .A1(n3134), .A2(n3189), .ZN(n3205) );
  OAI211_X1 U3966 ( .C1(n3136), .C2(n3135), .A(n4524), .B(n3205), .ZN(n3141)
         );
  INV_X1 U3967 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3137) );
  NOR2_X1 U3968 ( .A1(STATE_REG_SCAN_IN), .A2(n3137), .ZN(n4592) );
  INV_X1 U3969 ( .A(n3803), .ZN(n3280) );
  OAI22_X1 U3970 ( .A1(n3138), .A2(n4515), .B1(n4514), .B2(n3280), .ZN(n3139)
         );
  AOI211_X1 U3971 ( .C1(n3285), .C2(n4518), .A(n4592), .B(n3139), .ZN(n3140)
         );
  OAI211_X1 U3972 ( .C1(n4528), .C2(n3287), .A(n3141), .B(n3140), .ZN(U3214)
         );
  XNOR2_X1 U3973 ( .A(n3142), .B(n3691), .ZN(n3152) );
  OAI22_X1 U3974 ( .A1(n3143), .A2(n4722), .B1(n4675), .B2(n3149), .ZN(n3147)
         );
  XNOR2_X1 U3975 ( .A(n3144), .B(n3691), .ZN(n3145) );
  NOR2_X1 U3976 ( .A1(n3145), .A2(n4681), .ZN(n3146) );
  AOI211_X1 U3977 ( .C1(n4679), .C2(n3808), .A(n3147), .B(n3146), .ZN(n3148)
         );
  OAI21_X1 U3978 ( .B1(n4702), .B2(n3152), .A(n3148), .ZN(n4790) );
  OAI211_X1 U3979 ( .C1(n2175), .C2(n3149), .A(n3326), .B(n4812), .ZN(n4789)
         );
  OAI22_X1 U3980 ( .A1(n4789), .A2(n2822), .B1(n4050), .B2(n3150), .ZN(n3151)
         );
  OAI21_X1 U3981 ( .B1(n4790), .B2(n3151), .A(n4089), .ZN(n3154) );
  INV_X1 U3982 ( .A(n3152), .ZN(n4792) );
  INV_X1 U3983 ( .A(n4712), .ZN(n4725) );
  AOI22_X1 U3984 ( .A1(n4792), .A2(n4725), .B1(REG2_REG_4__SCAN_IN), .B2(n4706), .ZN(n3153) );
  NAND2_X1 U3985 ( .A1(n3154), .A2(n3153), .ZN(U3286) );
  NAND2_X1 U3986 ( .A1(n4089), .A2(n4720), .ZN(n3155) );
  XNOR2_X1 U3987 ( .A(n3156), .B(n3695), .ZN(n4802) );
  INV_X1 U3988 ( .A(n3157), .ZN(n3158) );
  OAI211_X1 U3989 ( .C1(n3159), .C2(n3165), .A(n3158), .B(n4812), .ZN(n4799)
         );
  INV_X1 U3990 ( .A(n3695), .ZN(n3160) );
  XNOR2_X1 U3991 ( .A(n3161), .B(n3160), .ZN(n3167) );
  NAND2_X1 U3992 ( .A1(n3320), .A2(n4679), .ZN(n3164) );
  NAND2_X1 U3993 ( .A1(n3162), .A2(n4696), .ZN(n3163) );
  OAI211_X1 U3994 ( .C1(n4675), .C2(n3165), .A(n3164), .B(n3163), .ZN(n3166)
         );
  AOI21_X1 U3995 ( .B1(n3167), .B2(n4719), .A(n3166), .ZN(n4800) );
  OAI21_X1 U3996 ( .B1(n2822), .B2(n4799), .A(n4800), .ZN(n3168) );
  NAND2_X1 U3997 ( .A1(n3168), .A2(n4534), .ZN(n3172) );
  INV_X1 U3998 ( .A(n3169), .ZN(n3170) );
  AOI22_X1 U3999 ( .A1(n4706), .A2(REG2_REG_7__SCAN_IN), .B1(n3170), .B2(n4724), .ZN(n3171) );
  OAI211_X1 U4000 ( .C1(n4101), .C2(n4802), .A(n3172), .B(n3171), .ZN(U3283)
         );
  NAND2_X1 U4001 ( .A1(n3803), .A2(n2976), .ZN(n3174) );
  NAND2_X1 U4002 ( .A1(n4688), .A2(n2132), .ZN(n3173) );
  NAND2_X1 U4003 ( .A1(n3174), .A2(n3173), .ZN(n3175) );
  XNOR2_X1 U4004 ( .A(n3175), .B(n3518), .ZN(n3180) );
  NOR2_X1 U4005 ( .A1(n4674), .A2(n3520), .ZN(n3176) );
  AOI21_X1 U4006 ( .B1(n3803), .B2(n3499), .A(n3176), .ZN(n3181) );
  NAND2_X1 U4007 ( .A1(n3180), .A2(n3181), .ZN(n3206) );
  INV_X1 U4008 ( .A(n3206), .ZN(n3185) );
  INV_X1 U4009 ( .A(n3177), .ZN(n3178) );
  NAND2_X1 U4010 ( .A1(n3179), .A2(n3178), .ZN(n3204) );
  INV_X1 U4011 ( .A(n3180), .ZN(n3183) );
  INV_X1 U4012 ( .A(n3181), .ZN(n3182) );
  NAND2_X1 U4013 ( .A1(n3183), .A2(n3182), .ZN(n3207) );
  AND2_X1 U4014 ( .A1(n3204), .A2(n3207), .ZN(n3184) );
  NOR2_X1 U4015 ( .A1(n3185), .A2(n3184), .ZN(n3191) );
  OR2_X1 U4016 ( .A1(n3186), .A2(n3191), .ZN(n3187) );
  AND2_X1 U4017 ( .A1(n3189), .A2(n3206), .ZN(n3190) );
  NOR2_X1 U4018 ( .A1(n3191), .A2(n3190), .ZN(n3192) );
  NAND2_X1 U4019 ( .A1(n3802), .A2(n2976), .ZN(n3194) );
  NAND2_X1 U4020 ( .A1(n3201), .A2(n2132), .ZN(n3193) );
  NAND2_X1 U4021 ( .A1(n3194), .A2(n3193), .ZN(n3195) );
  XNOR2_X1 U4022 ( .A(n3195), .B(n3526), .ZN(n3260) );
  NAND2_X1 U4023 ( .A1(n3802), .A2(n3499), .ZN(n3197) );
  NAND2_X1 U4024 ( .A1(n3201), .A2(n2976), .ZN(n3196) );
  NAND2_X1 U4025 ( .A1(n3197), .A2(n3196), .ZN(n3263) );
  XNOR2_X1 U4026 ( .A(n3260), .B(n3263), .ZN(n3198) );
  XNOR2_X1 U4027 ( .A(n3269), .B(n3198), .ZN(n3199) );
  NAND2_X1 U4028 ( .A1(n3199), .A2(n4524), .ZN(n3203) );
  NOR2_X1 U4029 ( .A1(STATE_REG_SCAN_IN), .A2(n4389), .ZN(n4600) );
  INV_X1 U4030 ( .A(n3376), .ZN(n3344) );
  OAI22_X1 U4031 ( .A1(n3280), .A2(n4515), .B1(n4514), .B2(n3344), .ZN(n3200)
         );
  AOI211_X1 U4032 ( .C1(n3201), .C2(n4518), .A(n4600), .B(n3200), .ZN(n3202)
         );
  OAI211_X1 U4033 ( .C1(n4528), .C2(n3351), .A(n3203), .B(n3202), .ZN(U3221)
         );
  NAND2_X1 U4034 ( .A1(n3205), .A2(n3204), .ZN(n3209) );
  NAND2_X1 U4035 ( .A1(n3207), .A2(n3206), .ZN(n3208) );
  XNOR2_X1 U4036 ( .A(n3209), .B(n3208), .ZN(n3210) );
  NAND2_X1 U4037 ( .A1(n3210), .A2(n4524), .ZN(n3214) );
  INV_X1 U4038 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4203) );
  NOR2_X1 U4039 ( .A1(STATE_REG_SCAN_IN), .A2(n4203), .ZN(n3257) );
  INV_X1 U4040 ( .A(n3802), .ZN(n4676) );
  OAI22_X1 U4041 ( .A1(n3211), .A2(n4515), .B1(n4514), .B2(n4676), .ZN(n3212)
         );
  AOI211_X1 U4042 ( .C1(n4688), .C2(n4518), .A(n3257), .B(n3212), .ZN(n3213)
         );
  OAI211_X1 U40430 ( .C1(n4528), .C2(n4684), .A(n3214), .B(n3213), .ZN(U3233)
         );
  INV_X1 U4044 ( .A(n3269), .ZN(n3216) );
  INV_X1 U4045 ( .A(n3260), .ZN(n3264) );
  OAI21_X1 U4046 ( .B1(n3269), .B2(n3260), .A(n3263), .ZN(n3215) );
  OAI21_X1 U4047 ( .B1(n3216), .B2(n3264), .A(n3215), .ZN(n3227) );
  NAND2_X1 U4048 ( .A1(n3376), .A2(n2976), .ZN(n3218) );
  NAND2_X1 U4049 ( .A1(n3230), .A2(n2132), .ZN(n3217) );
  NAND2_X1 U4050 ( .A1(n3218), .A2(n3217), .ZN(n3219) );
  XNOR2_X1 U4051 ( .A(n3219), .B(n3526), .ZN(n3222) );
  NAND2_X1 U4052 ( .A1(n3376), .A2(n3499), .ZN(n3221) );
  NAND2_X1 U4053 ( .A1(n3230), .A2(n2976), .ZN(n3220) );
  NAND2_X1 U4054 ( .A1(n3221), .A2(n3220), .ZN(n3223) );
  INV_X1 U4055 ( .A(n3261), .ZN(n3266) );
  INV_X1 U4056 ( .A(n3222), .ZN(n3225) );
  INV_X1 U4057 ( .A(n3223), .ZN(n3224) );
  NAND2_X1 U4058 ( .A1(n3225), .A2(n3224), .ZN(n3267) );
  NAND2_X1 U4059 ( .A1(n3266), .A2(n3267), .ZN(n3226) );
  XNOR2_X1 U4060 ( .A(n3227), .B(n3226), .ZN(n3228) );
  NAND2_X1 U4061 ( .A1(n3228), .A2(n4524), .ZN(n3232) );
  NOR2_X1 U4062 ( .A1(STATE_REG_SCAN_IN), .A2(n2534), .ZN(n4612) );
  INV_X1 U4063 ( .A(n4097), .ZN(n4516) );
  OAI22_X1 U4064 ( .A1(n4676), .A2(n4515), .B1(n4514), .B2(n4516), .ZN(n3229)
         );
  AOI211_X1 U4065 ( .C1(n3230), .C2(n4518), .A(n4612), .B(n3229), .ZN(n3231)
         );
  OAI211_X1 U4066 ( .C1(n4528), .C2(n3387), .A(n3232), .B(n3231), .ZN(U3231)
         );
  OAI22_X1 U4067 ( .A1(n4089), .A2(n4560), .B1(n3233), .B2(n4050), .ZN(n3236)
         );
  NOR2_X1 U4068 ( .A1(n3234), .A2(n4101), .ZN(n3235) );
  AOI211_X1 U4069 ( .C1(n3237), .C2(n4689), .A(n3236), .B(n3235), .ZN(n3238)
         );
  OAI21_X1 U4070 ( .B1(n4706), .B2(n3239), .A(n3238), .ZN(U3284) );
  NAND2_X1 U4071 ( .A1(n4497), .A2(REG1_REG_9__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4072 ( .A1(n3249), .A2(n3242), .ZN(n3243) );
  INV_X1 U4073 ( .A(n3249), .ZN(n4755) );
  XNOR2_X1 U4074 ( .A(n3242), .B(n4755), .ZN(n4595) );
  NAND2_X1 U4075 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4595), .ZN(n4594) );
  MUX2_X1 U4076 ( .A(n3244), .B(REG1_REG_11__SCAN_IN), .S(n3846), .Z(n3245) );
  OAI211_X1 U4077 ( .C1(n3246), .C2(n3245), .A(n3845), .B(n4662), .ZN(n3259)
         );
  NOR2_X1 U4078 ( .A1(n3250), .A2(n4755), .ZN(n3251) );
  INV_X1 U4079 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4591) );
  NOR2_X1 U4080 ( .A1(n3251), .A2(n4589), .ZN(n3255) );
  INV_X1 U4081 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3252) );
  MUX2_X1 U4082 ( .A(REG2_REG_11__SCAN_IN), .B(n3252), .S(n3846), .Z(n3254) );
  INV_X1 U4083 ( .A(n3831), .ZN(n3253) );
  AOI211_X1 U4084 ( .C1(n3255), .C2(n3254), .A(n3253), .B(n4654), .ZN(n3256)
         );
  AOI211_X1 U4085 ( .C1(n4671), .C2(ADDR_REG_11__SCAN_IN), .A(n3257), .B(n3256), .ZN(n3258) );
  OAI211_X1 U4086 ( .C1(n4669), .C2(n3846), .A(n3259), .B(n3258), .ZN(U3251)
         );
  AND2_X1 U4087 ( .A1(n3260), .A2(n3263), .ZN(n3262) );
  INV_X1 U4088 ( .A(n3263), .ZN(n3265) );
  NAND3_X1 U4089 ( .A1(n3266), .A2(n3265), .A3(n3264), .ZN(n3268) );
  NOR2_X1 U4090 ( .A1(n3360), .A2(n3520), .ZN(n3270) );
  AOI21_X1 U4091 ( .B1(n4097), .B2(n3499), .A(n3270), .ZN(n3418) );
  NAND2_X1 U4092 ( .A1(n4097), .A2(n2976), .ZN(n3272) );
  NAND2_X1 U4093 ( .A1(n3366), .A2(n2132), .ZN(n3271) );
  NAND2_X1 U4094 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  XNOR2_X1 U4095 ( .A(n3273), .B(n3518), .ZN(n3419) );
  XOR2_X1 U4096 ( .A(n3418), .B(n3419), .Z(n3274) );
  XNOR2_X1 U4097 ( .A(n3420), .B(n3274), .ZN(n3275) );
  NAND2_X1 U4098 ( .A1(n3275), .A2(n4524), .ZN(n3278) );
  NOR2_X1 U4099 ( .A1(STATE_REG_SCAN_IN), .A2(n4384), .ZN(n4625) );
  OAI22_X1 U4100 ( .A1(n3344), .A2(n4515), .B1(n4514), .B2(n4503), .ZN(n3276)
         );
  AOI211_X1 U4101 ( .C1(n3366), .C2(n4518), .A(n4625), .B(n3276), .ZN(n3277)
         );
  OAI211_X1 U4102 ( .C1(n4528), .C2(n3367), .A(n3278), .B(n3277), .ZN(U3212)
         );
  NAND2_X1 U4103 ( .A1(n3753), .A2(n3758), .ZN(n3690) );
  XNOR2_X1 U4104 ( .A(n3279), .B(n3690), .ZN(n3283) );
  OAI22_X1 U4105 ( .A1(n3280), .A2(n4722), .B1(n4675), .B2(n2367), .ZN(n3281)
         );
  AOI21_X1 U4106 ( .B1(n4679), .B2(n3804), .A(n3281), .ZN(n3282) );
  OAI21_X1 U4107 ( .B1(n3283), .B2(n4681), .A(n3282), .ZN(n3334) );
  INV_X1 U4108 ( .A(n3334), .ZN(n3292) );
  XOR2_X1 U4109 ( .A(n3284), .B(n3690), .Z(n3335) );
  INV_X1 U4110 ( .A(n4101), .ZN(n3355) );
  NAND2_X1 U4111 ( .A1(n3309), .A2(n3285), .ZN(n3286) );
  NAND2_X1 U4112 ( .A1(n4687), .A2(n3286), .ZN(n3339) );
  INV_X1 U4113 ( .A(n3287), .ZN(n3288) );
  AOI22_X1 U4114 ( .A1(n4706), .A2(REG2_REG_10__SCAN_IN), .B1(n3288), .B2(
        n4724), .ZN(n3289) );
  OAI21_X1 U4115 ( .B1(n3339), .B2(n4711), .A(n3289), .ZN(n3290) );
  AOI21_X1 U4116 ( .B1(n3335), .B2(n3355), .A(n3290), .ZN(n3291) );
  OAI21_X1 U4117 ( .B1(n4706), .B2(n3292), .A(n3291), .ZN(U3280) );
  INV_X1 U4118 ( .A(n3293), .ZN(n3300) );
  NOR2_X1 U4119 ( .A1(n3294), .A2(n4711), .ZN(n3297) );
  OAI22_X1 U4120 ( .A1(n4089), .A2(n4581), .B1(n3295), .B2(n4050), .ZN(n3296)
         );
  AOI211_X1 U4121 ( .C1(n3298), .C2(n3355), .A(n3297), .B(n3296), .ZN(n3299)
         );
  OAI21_X1 U4122 ( .B1(n3300), .B2(n4706), .A(n3299), .ZN(U3282) );
  NAND2_X1 U4123 ( .A1(n2702), .A2(n3744), .ZN(n3692) );
  XNOR2_X1 U4124 ( .A(n3301), .B(n3692), .ZN(n3306) );
  AOI22_X1 U4125 ( .A1(n4678), .A2(n4696), .B1(n4695), .B2(n3302), .ZN(n3303)
         );
  OAI21_X1 U4126 ( .B1(n3304), .B2(n4698), .A(n3303), .ZN(n3305) );
  AOI21_X1 U4127 ( .B1(n3306), .B2(n4719), .A(n3305), .ZN(n4805) );
  XNOR2_X1 U4128 ( .A(n3307), .B(n3692), .ZN(n4808) );
  INV_X1 U4129 ( .A(n3308), .ZN(n3311) );
  OAI21_X1 U4130 ( .B1(n3311), .B2(n3310), .A(n3309), .ZN(n4806) );
  NOR2_X1 U4131 ( .A1(n4806), .A2(n4711), .ZN(n3315) );
  OAI22_X1 U4132 ( .A1(n4089), .A2(n3313), .B1(n3312), .B2(n4050), .ZN(n3314)
         );
  AOI211_X1 U4133 ( .C1(n4808), .C2(n3355), .A(n3315), .B(n3314), .ZN(n3316)
         );
  OAI21_X1 U4134 ( .B1(n4706), .B2(n4805), .A(n3316), .ZN(U3281) );
  INV_X1 U4135 ( .A(n3317), .ZN(n3736) );
  NAND2_X1 U4136 ( .A1(n3736), .A2(n3749), .ZN(n3679) );
  XNOR2_X1 U4137 ( .A(n3318), .B(n3679), .ZN(n3324) );
  AOI22_X1 U4138 ( .A1(n3320), .A2(n4696), .B1(n4695), .B2(n3319), .ZN(n3321)
         );
  OAI21_X1 U4139 ( .B1(n3322), .B2(n4698), .A(n3321), .ZN(n3323) );
  AOI21_X1 U4140 ( .B1(n3324), .B2(n4719), .A(n3323), .ZN(n4794) );
  XOR2_X1 U4141 ( .A(n3679), .B(n3325), .Z(n4797) );
  INV_X1 U4142 ( .A(n3326), .ZN(n3329) );
  OAI21_X1 U4143 ( .B1(n3329), .B2(n3328), .A(n3327), .ZN(n4795) );
  NOR2_X1 U4144 ( .A1(n4795), .A2(n4711), .ZN(n3332) );
  OAI22_X1 U4145 ( .A1(n4089), .A2(n4306), .B1(n3330), .B2(n4050), .ZN(n3331)
         );
  AOI211_X1 U4146 ( .C1(n4797), .C2(n3355), .A(n3332), .B(n3331), .ZN(n3333)
         );
  OAI21_X1 U4147 ( .B1(n4706), .B2(n4794), .A(n3333), .ZN(U3285) );
  INV_X1 U4148 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4366) );
  AOI21_X1 U4149 ( .B1(n3335), .B2(n4809), .A(n3334), .ZN(n3337) );
  MUX2_X1 U4150 ( .A(n4366), .B(n3337), .S(n4824), .Z(n3336) );
  OAI21_X1 U4151 ( .B1(n3339), .B2(n4489), .A(n3336), .ZN(U3487) );
  MUX2_X1 U4152 ( .A(n2506), .B(n3337), .S(n4836), .Z(n3338) );
  OAI21_X1 U4153 ( .B1(n3339), .B2(n4435), .A(n3338), .ZN(U3528) );
  NAND2_X1 U4154 ( .A1(n3374), .A2(n3372), .ZN(n3709) );
  INV_X1 U4155 ( .A(n3341), .ZN(n3342) );
  AOI21_X1 U4156 ( .B1(n3340), .B2(n3343), .A(n3342), .ZN(n3375) );
  XOR2_X1 U4157 ( .A(n3709), .B(n3375), .Z(n3347) );
  OAI22_X1 U4158 ( .A1(n3344), .A2(n4722), .B1(n4675), .B2(n3349), .ZN(n3345)
         );
  AOI21_X1 U4159 ( .B1(n4679), .B2(n3803), .A(n3345), .ZN(n3346) );
  OAI21_X1 U4160 ( .B1(n3347), .B2(n4681), .A(n3346), .ZN(n3392) );
  INV_X1 U4161 ( .A(n3392), .ZN(n3357) );
  XOR2_X1 U4162 ( .A(n3709), .B(n3348), .Z(n3393) );
  OR2_X1 U4163 ( .A1(n4686), .A2(n3349), .ZN(n3350) );
  NAND2_X1 U4164 ( .A1(n3383), .A2(n3350), .ZN(n3398) );
  NOR2_X1 U4165 ( .A1(n3398), .A2(n4711), .ZN(n3354) );
  INV_X1 U4166 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3352) );
  OAI22_X1 U4167 ( .A1(n4089), .A2(n3352), .B1(n3351), .B2(n4050), .ZN(n3353)
         );
  AOI211_X1 U4168 ( .C1(n3393), .C2(n3355), .A(n3354), .B(n3353), .ZN(n3356)
         );
  OAI21_X1 U4169 ( .B1(n4706), .B2(n3357), .A(n3356), .ZN(U3278) );
  XNOR2_X1 U4170 ( .A(n3358), .B(n3359), .ZN(n4440) );
  XNOR2_X1 U4171 ( .A(n3650), .B(n2212), .ZN(n3363) );
  OAI22_X1 U4172 ( .A1(n4503), .A2(n4722), .B1(n4675), .B2(n3360), .ZN(n3361)
         );
  AOI21_X1 U4173 ( .B1(n4679), .B2(n3376), .A(n3361), .ZN(n3362) );
  OAI21_X1 U4174 ( .B1(n3363), .B2(n4681), .A(n3362), .ZN(n3364) );
  AOI21_X1 U4175 ( .B1(n4440), .B2(n4720), .A(n3364), .ZN(n4444) );
  INV_X1 U4176 ( .A(n3365), .ZN(n4442) );
  NAND2_X1 U4177 ( .A1(n3384), .A2(n3366), .ZN(n4441) );
  AND3_X1 U4178 ( .A1(n4442), .A2(n4689), .A3(n4441), .ZN(n3370) );
  INV_X1 U4179 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3368) );
  OAI22_X1 U4180 ( .A1(n4089), .A2(n3368), .B1(n3367), .B2(n4050), .ZN(n3369)
         );
  AOI211_X1 U4181 ( .C1(n4440), .C2(n4725), .A(n3370), .B(n3369), .ZN(n3371)
         );
  OAI21_X1 U4182 ( .B1(n4444), .B2(n4706), .A(n3371), .ZN(U3276) );
  INV_X1 U4183 ( .A(n3372), .ZN(n3373) );
  AOI21_X1 U4184 ( .B1(n3375), .B2(n3374), .A(n3373), .ZN(n3377) );
  XNOR2_X1 U4185 ( .A(n3376), .B(n3385), .ZN(n3715) );
  XNOR2_X1 U4186 ( .A(n3377), .B(n3715), .ZN(n3382) );
  XNOR2_X1 U4187 ( .A(n3378), .B(n3715), .ZN(n4821) );
  NAND2_X1 U4188 ( .A1(n4821), .A2(n4720), .ZN(n3381) );
  OAI22_X1 U4189 ( .A1(n4516), .A2(n4722), .B1(n4675), .B2(n3385), .ZN(n3379)
         );
  AOI21_X1 U4190 ( .B1(n4679), .B2(n3802), .A(n3379), .ZN(n3380) );
  OAI211_X1 U4191 ( .C1(n4681), .C2(n3382), .A(n3381), .B(n3380), .ZN(n4818)
         );
  INV_X1 U4192 ( .A(n4818), .ZN(n3391) );
  INV_X1 U4193 ( .A(n3383), .ZN(n3386) );
  OAI21_X1 U4194 ( .B1(n3386), .B2(n3385), .A(n3384), .ZN(n4817) );
  NOR2_X1 U4195 ( .A1(n4817), .A2(n4711), .ZN(n3389) );
  INV_X1 U4196 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3834) );
  OAI22_X1 U4197 ( .A1(n4089), .A2(n3834), .B1(n3387), .B2(n4050), .ZN(n3388)
         );
  AOI211_X1 U4198 ( .C1(n4821), .C2(n4725), .A(n3389), .B(n3388), .ZN(n3390)
         );
  OAI21_X1 U4199 ( .B1(n3391), .B2(n4706), .A(n3390), .ZN(U3277) );
  AOI21_X1 U4200 ( .B1(n4809), .B2(n3393), .A(n3392), .ZN(n3395) );
  MUX2_X1 U4201 ( .A(n2523), .B(n3395), .S(n4836), .Z(n3394) );
  OAI21_X1 U4202 ( .B1(n3398), .B2(n4435), .A(n3394), .ZN(U3530) );
  INV_X1 U4203 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3396) );
  MUX2_X1 U4204 ( .A(n3396), .B(n3395), .S(n4824), .Z(n3397) );
  OAI21_X1 U4205 ( .B1(n3398), .B2(n4489), .A(n3397), .ZN(U3491) );
  NAND2_X1 U4206 ( .A1(n2408), .A2(DATAI_29_), .ZN(n3663) );
  XOR2_X1 U4207 ( .A(n3663), .B(n3664), .Z(n3700) );
  XNOR2_X1 U4208 ( .A(n3402), .B(n3700), .ZN(n4120) );
  INV_X1 U4209 ( .A(n3663), .ZN(n3410) );
  AOI21_X1 U4210 ( .B1(n3410), .B2(n3403), .A(n4107), .ZN(n4118) );
  AOI22_X1 U4211 ( .A1(n4118), .A2(n4689), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4706), .ZN(n3417) );
  INV_X1 U4212 ( .A(n3404), .ZN(n3660) );
  AOI21_X1 U4213 ( .B1(n3405), .B2(n3666), .A(n3660), .ZN(n3406) );
  XNOR2_X1 U4214 ( .A(n3406), .B(n3700), .ZN(n3413) );
  INV_X1 U4215 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4216 ( .A1(n2421), .A2(REG2_REG_30__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4217 ( .A1(n2424), .A2(REG0_REG_30__SCAN_IN), .ZN(n3407) );
  OAI211_X1 U4218 ( .C1(n2724), .C2(n3409), .A(n3408), .B(n3407), .ZN(n3801)
         );
  AOI21_X1 U4219 ( .B1(n4540), .B2(B_REG_SCAN_IN), .A(n4722), .ZN(n4102) );
  AOI22_X1 U4220 ( .A1(n3801), .A2(n4102), .B1(n3410), .B2(n4695), .ZN(n3412)
         );
  NAND2_X1 U4221 ( .A1(n3887), .A2(n4679), .ZN(n3411) );
  OAI211_X1 U4222 ( .C1(n3413), .C2(n4681), .A(n3412), .B(n3411), .ZN(n4117)
         );
  NOR2_X1 U4223 ( .A1(n4050), .A2(n3414), .ZN(n3415) );
  OAI21_X1 U4224 ( .B1(n4117), .B2(n3415), .A(n4089), .ZN(n3416) );
  OAI211_X1 U4225 ( .C1(n4120), .C2(n4101), .A(n3417), .B(n3416), .ZN(U3354)
         );
  NAND2_X1 U4226 ( .A1(n3425), .A2(n2976), .ZN(n3422) );
  NAND2_X1 U4227 ( .A1(n4519), .A2(n3455), .ZN(n3421) );
  NAND2_X1 U4228 ( .A1(n3422), .A2(n3421), .ZN(n3423) );
  XNOR2_X1 U4229 ( .A(n3423), .B(n3526), .ZN(n3426) );
  AND2_X1 U4230 ( .A1(n4519), .A2(n2976), .ZN(n3424) );
  AOI21_X1 U4231 ( .B1(n3425), .B2(n3499), .A(n3424), .ZN(n4521) );
  NAND2_X1 U4232 ( .A1(n4060), .A2(n2976), .ZN(n3428) );
  NAND2_X1 U4233 ( .A1(n4505), .A2(n2132), .ZN(n3427) );
  NAND2_X1 U4234 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U4235 ( .A(n3429), .B(n3518), .ZN(n3433) );
  NOR2_X1 U4236 ( .A1(n4080), .A2(n3520), .ZN(n3430) );
  AOI21_X1 U4237 ( .B1(n4060), .B2(n3499), .A(n3430), .ZN(n3432) );
  XNOR2_X1 U4238 ( .A(n3433), .B(n3432), .ZN(n4507) );
  INV_X1 U4239 ( .A(n4507), .ZN(n3431) );
  NAND2_X1 U4240 ( .A1(n4076), .A2(n2976), .ZN(n3435) );
  NAND2_X1 U4241 ( .A1(n3590), .A2(n2132), .ZN(n3434) );
  NAND2_X1 U4242 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  XNOR2_X1 U4243 ( .A(n3436), .B(n3526), .ZN(n3584) );
  NAND2_X1 U4244 ( .A1(n4076), .A2(n3499), .ZN(n3438) );
  NAND2_X1 U4245 ( .A1(n3590), .A2(n2976), .ZN(n3437) );
  NAND2_X1 U4246 ( .A1(n3438), .A2(n3437), .ZN(n3583) );
  INV_X1 U4247 ( .A(n3584), .ZN(n3440) );
  INV_X1 U4248 ( .A(n3583), .ZN(n3439) );
  OAI22_X1 U4249 ( .A1(n3582), .A2(n3441), .B1(n3440), .B2(n3439), .ZN(n3639)
         );
  NAND2_X1 U4250 ( .A1(n4059), .A2(n2976), .ZN(n3443) );
  NAND2_X1 U4251 ( .A1(n3647), .A2(n2132), .ZN(n3442) );
  NAND2_X1 U4252 ( .A1(n3443), .A2(n3442), .ZN(n3444) );
  XNOR2_X1 U4253 ( .A(n3444), .B(n3518), .ZN(n3447) );
  NOR2_X1 U4254 ( .A1(n4047), .A2(n3520), .ZN(n3445) );
  AOI21_X1 U4255 ( .B1(n4059), .B2(n3499), .A(n3445), .ZN(n3446) );
  NOR2_X1 U4256 ( .A1(n3447), .A2(n3446), .ZN(n3640) );
  NAND2_X1 U4257 ( .A1(n3447), .A2(n3446), .ZN(n3641) );
  NAND2_X1 U4258 ( .A1(n4044), .A2(n2976), .ZN(n3449) );
  NAND2_X1 U4259 ( .A1(n3451), .A2(n2132), .ZN(n3448) );
  NAND2_X1 U4260 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  XNOR2_X1 U4261 ( .A(n3450), .B(n3526), .ZN(n3452) );
  AOI22_X1 U4262 ( .A1(n4044), .A2(n3499), .B1(n2976), .B2(n3451), .ZN(n3453)
         );
  XNOR2_X1 U4263 ( .A(n3452), .B(n3453), .ZN(n3556) );
  INV_X1 U4264 ( .A(n3452), .ZN(n3454) );
  NAND2_X1 U4265 ( .A1(n3987), .A2(n2976), .ZN(n3457) );
  OR2_X1 U4266 ( .A1(n3494), .A2(n4009), .ZN(n3456) );
  NAND2_X1 U4267 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  XNOR2_X1 U4268 ( .A(n3458), .B(n3518), .ZN(n3465) );
  NOR2_X1 U4269 ( .A1(n3520), .A2(n4009), .ZN(n3459) );
  AOI21_X1 U4270 ( .B1(n3987), .B2(n3499), .A(n3459), .ZN(n3464) );
  NOR2_X1 U4271 ( .A1(n3465), .A2(n3464), .ZN(n3606) );
  NAND2_X1 U4272 ( .A1(n3973), .A2(n2976), .ZN(n3461) );
  OR2_X1 U4273 ( .A1(n3494), .A2(n3991), .ZN(n3460) );
  NAND2_X1 U4274 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  XNOR2_X1 U4275 ( .A(n3462), .B(n3518), .ZN(n3563) );
  NOR2_X1 U4276 ( .A1(n3520), .A2(n3991), .ZN(n3463) );
  AOI21_X1 U4277 ( .B1(n3973), .B2(n3499), .A(n3463), .ZN(n3562) );
  NAND2_X1 U4278 ( .A1(n3563), .A2(n3562), .ZN(n3466) );
  NAND2_X1 U4279 ( .A1(n3465), .A2(n3464), .ZN(n3604) );
  OAI21_X1 U4280 ( .B1(n3608), .B2(n3606), .A(n2373), .ZN(n3470) );
  NAND2_X1 U4281 ( .A1(n3470), .A2(n3469), .ZN(n3616) );
  AOI22_X1 U4282 ( .A1(n3960), .A2(n2976), .B1(n3966), .B2(n3455), .ZN(n3471)
         );
  XNOR2_X1 U4283 ( .A(n3471), .B(n3526), .ZN(n3472) );
  AOI22_X1 U4284 ( .A1(n3960), .A2(n3499), .B1(n3966), .B2(n2976), .ZN(n3473)
         );
  XNOR2_X1 U4285 ( .A(n3472), .B(n3473), .ZN(n3617) );
  INV_X1 U4286 ( .A(n3472), .ZN(n3475) );
  INV_X1 U4287 ( .A(n3473), .ZN(n3474) );
  NOR2_X1 U4288 ( .A1(n3475), .A2(n3474), .ZN(n3549) );
  NAND2_X1 U4289 ( .A1(n3974), .A2(n2976), .ZN(n3477) );
  NAND2_X1 U4290 ( .A1(n3455), .A2(n3947), .ZN(n3476) );
  NAND2_X1 U4291 ( .A1(n3477), .A2(n3476), .ZN(n3478) );
  XNOR2_X1 U4292 ( .A(n3478), .B(n3518), .ZN(n3481) );
  NOR2_X1 U4293 ( .A1(n3957), .A2(n3520), .ZN(n3479) );
  AOI21_X1 U4294 ( .B1(n3974), .B2(n3499), .A(n3479), .ZN(n3480) );
  XNOR2_X1 U4295 ( .A(n3481), .B(n3480), .ZN(n3548) );
  NAND2_X1 U4296 ( .A1(n3917), .A2(n3499), .ZN(n3484) );
  NAND2_X1 U4297 ( .A1(n2976), .A2(n3482), .ZN(n3483) );
  NAND2_X1 U4298 ( .A1(n3484), .A2(n3483), .ZN(n3486) );
  OAI22_X1 U4299 ( .A1(n3958), .A2(n3520), .B1(n3936), .B2(n3494), .ZN(n3485)
         );
  XOR2_X1 U4300 ( .A(n3526), .B(n3485), .Z(n3596) );
  NAND2_X1 U4301 ( .A1(n3900), .A2(n2976), .ZN(n3488) );
  OR2_X1 U4302 ( .A1(n3494), .A2(n3914), .ZN(n3487) );
  NAND2_X1 U4303 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  XNOR2_X1 U4304 ( .A(n3489), .B(n3518), .ZN(n3492) );
  NOR2_X1 U4305 ( .A1(n3520), .A2(n3914), .ZN(n3490) );
  AOI21_X1 U4306 ( .B1(n3900), .B2(n3499), .A(n3490), .ZN(n3491) );
  NAND2_X1 U4307 ( .A1(n3492), .A2(n3491), .ZN(n3572) );
  NAND2_X1 U4308 ( .A1(n3574), .A2(n3572), .ZN(n3493) );
  OR2_X1 U4309 ( .A1(n3492), .A2(n3491), .ZN(n3573) );
  NAND2_X1 U4310 ( .A1(n3500), .A2(n2976), .ZN(n3496) );
  OR2_X1 U4311 ( .A1(n3494), .A2(n3904), .ZN(n3495) );
  NAND2_X1 U4312 ( .A1(n3496), .A2(n3495), .ZN(n3497) );
  XNOR2_X1 U4313 ( .A(n3497), .B(n3518), .ZN(n3502) );
  NOR2_X1 U4314 ( .A1(n3520), .A2(n3904), .ZN(n3498) );
  AOI21_X1 U4315 ( .B1(n3500), .B2(n3499), .A(n3498), .ZN(n3501) );
  NOR2_X1 U4316 ( .A1(n3502), .A2(n3501), .ZN(n3514) );
  NAND2_X1 U4317 ( .A1(n3502), .A2(n3501), .ZN(n3513) );
  NOR2_X1 U4318 ( .A1(n3514), .A2(n2259), .ZN(n3503) );
  XNOR2_X1 U4319 ( .A(n3515), .B(n3503), .ZN(n3509) );
  INV_X1 U4320 ( .A(n3504), .ZN(n3906) );
  OAI22_X1 U4321 ( .A1(n3931), .A2(n4515), .B1(n4514), .B2(n3898), .ZN(n3507)
         );
  OAI22_X1 U4322 ( .A1(n3620), .A2(n3904), .B1(STATE_REG_SCAN_IN), .B2(n3505), 
        .ZN(n3506) );
  AOI211_X1 U4323 ( .C1(n3906), .C2(n3623), .A(n3507), .B(n3506), .ZN(n3508)
         );
  OAI21_X1 U4324 ( .B1(n3509), .B2(n3626), .A(n3508), .ZN(U3237) );
  INV_X1 U4325 ( .A(IR_REG_30__SCAN_IN), .ZN(n4148) );
  NAND3_X1 U4326 ( .A1(n4148), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3512) );
  INV_X1 U4327 ( .A(DATAI_31_), .ZN(n3511) );
  OAI22_X1 U4328 ( .A1(n3510), .A2(n3512), .B1(STATE_REG_SCAN_IN), .B2(n3511), 
        .ZN(U3321) );
  NAND2_X1 U4329 ( .A1(n3522), .A2(n2976), .ZN(n3517) );
  OR2_X1 U4330 ( .A1(n3494), .A2(n3542), .ZN(n3516) );
  NAND2_X1 U4331 ( .A1(n3517), .A2(n3516), .ZN(n3519) );
  XNOR2_X1 U4332 ( .A(n3519), .B(n3518), .ZN(n3524) );
  NOR2_X1 U4333 ( .A1(n3520), .A2(n3542), .ZN(n3521) );
  AOI21_X1 U4334 ( .B1(n3522), .B2(n3499), .A(n3521), .ZN(n3523) );
  XNOR2_X1 U4335 ( .A(n3524), .B(n3523), .ZN(n3539) );
  AOI22_X1 U4336 ( .A1(n3887), .A2(n3499), .B1(n2364), .B2(n2976), .ZN(n3529)
         );
  AOI22_X1 U4337 ( .A1(n3887), .A2(n2976), .B1(n2364), .B2(n3455), .ZN(n3527)
         );
  XNOR2_X1 U4338 ( .A(n3527), .B(n3526), .ZN(n3528) );
  XOR2_X1 U4339 ( .A(n3529), .B(n3528), .Z(n3530) );
  INV_X1 U4340 ( .A(n3870), .ZN(n3535) );
  INV_X1 U4341 ( .A(n3664), .ZN(n3531) );
  OAI22_X1 U4342 ( .A1(n3898), .A2(n4515), .B1(n4514), .B2(n3531), .ZN(n3534)
         );
  INV_X1 U4343 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4387) );
  OAI22_X1 U4344 ( .A1(n3620), .A2(n3532), .B1(STATE_REG_SCAN_IN), .B2(n4387), 
        .ZN(n3533) );
  AOI211_X1 U4345 ( .C1(n3535), .C2(n3623), .A(n3534), .B(n3533), .ZN(n3536)
         );
  OAI21_X1 U4346 ( .B1(n3537), .B2(n3626), .A(n3536), .ZN(U3217) );
  XNOR2_X1 U4347 ( .A(n3538), .B(n3539), .ZN(n3547) );
  INV_X1 U4348 ( .A(n3880), .ZN(n3545) );
  INV_X1 U4349 ( .A(n3887), .ZN(n3540) );
  OAI22_X1 U4350 ( .A1(n3915), .A2(n4515), .B1(n4514), .B2(n3540), .ZN(n3544)
         );
  INV_X1 U4351 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3541) );
  OAI22_X1 U4352 ( .A1(n3620), .A2(n3542), .B1(STATE_REG_SCAN_IN), .B2(n3541), 
        .ZN(n3543) );
  AOI211_X1 U4353 ( .C1(n3545), .C2(n3623), .A(n3544), .B(n3543), .ZN(n3546)
         );
  OAI21_X1 U4354 ( .B1(n3547), .B2(n3626), .A(n3546), .ZN(U3211) );
  OAI21_X1 U4355 ( .B1(n3615), .B2(n3549), .A(n3548), .ZN(n3550) );
  NAND3_X1 U4356 ( .A1(n2154), .A2(n4524), .A3(n3550), .ZN(n3554) );
  INV_X1 U4357 ( .A(n3960), .ZN(n3985) );
  OAI22_X1 U4358 ( .A1(n3985), .A2(n4515), .B1(n4514), .B2(n3958), .ZN(n3552)
         );
  NOR2_X1 U4359 ( .A1(n3620), .A2(n3957), .ZN(n3551) );
  AOI211_X1 U4360 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3552), .B(n3551), .ZN(n3553) );
  OAI211_X1 U4361 ( .C1(n4528), .C2(n3948), .A(n3554), .B(n3553), .ZN(U3213)
         );
  XOR2_X1 U4362 ( .A(n3556), .B(n3555), .Z(n3561) );
  INV_X1 U4363 ( .A(n3557), .ZN(n4032) );
  AOI22_X1 U4364 ( .A1(n3635), .A2(n4059), .B1(n3634), .B2(n3987), .ZN(n3558)
         );
  NAND2_X1 U4365 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3862) );
  OAI211_X1 U4366 ( .C1(n3620), .C2(n4029), .A(n3558), .B(n3862), .ZN(n3559)
         );
  AOI21_X1 U4367 ( .B1(n4032), .B2(n3623), .A(n3559), .ZN(n3560) );
  OAI21_X1 U4368 ( .B1(n3561), .B2(n3626), .A(n3560), .ZN(U3216) );
  AOI21_X1 U4369 ( .B1(n3608), .B2(n3604), .A(n3606), .ZN(n3565) );
  XNOR2_X1 U4370 ( .A(n3563), .B(n3562), .ZN(n3564) );
  XNOR2_X1 U4371 ( .A(n3565), .B(n3564), .ZN(n3571) );
  INV_X1 U4372 ( .A(n3993), .ZN(n3569) );
  INV_X1 U4373 ( .A(n3987), .ZN(n4025) );
  OAI22_X1 U4374 ( .A1(n4025), .A2(n4515), .B1(n4514), .B2(n3985), .ZN(n3568)
         );
  OAI22_X1 U4375 ( .A1(n3620), .A2(n3991), .B1(STATE_REG_SCAN_IN), .B2(n3566), 
        .ZN(n3567) );
  AOI211_X1 U4376 ( .C1(n3569), .C2(n3623), .A(n3568), .B(n3567), .ZN(n3570)
         );
  OAI21_X1 U4377 ( .B1(n3571), .B2(n3626), .A(n3570), .ZN(U3220) );
  NAND2_X1 U4378 ( .A1(n3573), .A2(n3572), .ZN(n3575) );
  XOR2_X1 U4379 ( .A(n3575), .B(n3574), .Z(n3581) );
  INV_X1 U4380 ( .A(n3576), .ZN(n3923) );
  OAI22_X1 U4381 ( .A1(n3958), .A2(n4515), .B1(n4514), .B2(n3915), .ZN(n3579)
         );
  OAI22_X1 U4382 ( .A1(n3620), .A2(n3914), .B1(STATE_REG_SCAN_IN), .B2(n3577), 
        .ZN(n3578) );
  AOI211_X1 U4383 ( .C1(n3923), .C2(n3623), .A(n3579), .B(n3578), .ZN(n3580)
         );
  OAI21_X1 U4384 ( .B1(n3581), .B2(n3626), .A(n3580), .ZN(U3222) );
  XNOR2_X1 U4385 ( .A(n3584), .B(n3583), .ZN(n3585) );
  XNOR2_X1 U4386 ( .A(n3586), .B(n3585), .ZN(n3587) );
  NAND2_X1 U4387 ( .A1(n3587), .A2(n4524), .ZN(n3592) );
  AND2_X1 U4388 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4657) );
  INV_X1 U4389 ( .A(n4060), .ZN(n4513) );
  INV_X1 U4390 ( .A(n4059), .ZN(n3588) );
  OAI22_X1 U4391 ( .A1(n4513), .A2(n4515), .B1(n4514), .B2(n3588), .ZN(n3589)
         );
  AOI211_X1 U4392 ( .C1(n3590), .C2(n4518), .A(n4657), .B(n3589), .ZN(n3591)
         );
  OAI211_X1 U4393 ( .C1(n4528), .C2(n4067), .A(n3592), .B(n3591), .ZN(U3225)
         );
  INV_X1 U4394 ( .A(n3593), .ZN(n3595) );
  NAND2_X1 U4395 ( .A1(n3595), .A2(n3594), .ZN(n3597) );
  XNOR2_X1 U4396 ( .A(n3597), .B(n3596), .ZN(n3603) );
  INV_X1 U4397 ( .A(n3937), .ZN(n3601) );
  OAI22_X1 U4398 ( .A1(n3618), .A2(n4515), .B1(n4514), .B2(n3931), .ZN(n3600)
         );
  INV_X1 U4399 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3598) );
  OAI22_X1 U4400 ( .A1(n3620), .A2(n3936), .B1(STATE_REG_SCAN_IN), .B2(n3598), 
        .ZN(n3599) );
  AOI211_X1 U4401 ( .C1(n3601), .C2(n3623), .A(n3600), .B(n3599), .ZN(n3602)
         );
  OAI21_X1 U4402 ( .B1(n3603), .B2(n3626), .A(n3602), .ZN(U3226) );
  INV_X1 U4403 ( .A(n3604), .ZN(n3605) );
  NOR2_X1 U4404 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U4405 ( .A(n3608), .B(n3607), .ZN(n3614) );
  INV_X1 U4406 ( .A(n4010), .ZN(n3612) );
  OAI22_X1 U4407 ( .A1(n4004), .A2(n4514), .B1(n4515), .B2(n3645), .ZN(n3611)
         );
  INV_X1 U4408 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3609) );
  OAI22_X1 U4409 ( .A1(n3620), .A2(n4009), .B1(STATE_REG_SCAN_IN), .B2(n3609), 
        .ZN(n3610) );
  AOI211_X1 U4410 ( .C1(n3612), .C2(n3623), .A(n3611), .B(n3610), .ZN(n3613)
         );
  OAI21_X1 U4411 ( .B1(n3614), .B2(n3626), .A(n3613), .ZN(U3230) );
  AOI21_X1 U4412 ( .B1(n3617), .B2(n3616), .A(n3615), .ZN(n3627) );
  INV_X1 U4413 ( .A(n3967), .ZN(n3624) );
  OAI22_X1 U4414 ( .A1(n4004), .A2(n4515), .B1(n4514), .B2(n3618), .ZN(n3622)
         );
  OAI22_X1 U4415 ( .A1(n3620), .A2(n3977), .B1(STATE_REG_SCAN_IN), .B2(n3619), 
        .ZN(n3621) );
  AOI211_X1 U4416 ( .C1(n3624), .C2(n3623), .A(n3622), .B(n3621), .ZN(n3625)
         );
  OAI21_X1 U4417 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(U3232) );
  OAI21_X1 U4418 ( .B1(n3628), .B2(n3629), .A(n3630), .ZN(n3631) );
  NAND2_X1 U4419 ( .A1(n3631), .A2(n4524), .ZN(n3638) );
  AOI22_X1 U4420 ( .A1(n4518), .A2(n3633), .B1(REG3_REG_2__SCAN_IN), .B2(n3632), .ZN(n3637) );
  AOI22_X1 U4421 ( .A1(n3635), .A2(n2841), .B1(n3634), .B2(n3808), .ZN(n3636)
         );
  NAND3_X1 U4422 ( .A1(n3638), .A2(n3637), .A3(n3636), .ZN(U3234) );
  INV_X1 U4423 ( .A(n3640), .ZN(n3642) );
  NAND2_X1 U4424 ( .A1(n3642), .A2(n3641), .ZN(n3643) );
  XNOR2_X1 U4425 ( .A(n3639), .B(n3643), .ZN(n3644) );
  NAND2_X1 U4426 ( .A1(n3644), .A2(n4524), .ZN(n3649) );
  INV_X1 U4427 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4207) );
  NOR2_X1 U4428 ( .A1(STATE_REG_SCAN_IN), .A2(n4207), .ZN(n4670) );
  OAI22_X1 U4429 ( .A1(n4502), .A2(n4515), .B1(n4514), .B2(n3645), .ZN(n3646)
         );
  AOI211_X1 U4430 ( .C1(n3647), .C2(n4518), .A(n4670), .B(n3646), .ZN(n3648)
         );
  OAI211_X1 U4431 ( .C1(n4528), .C2(n4051), .A(n3649), .B(n3648), .ZN(U3235)
         );
  NOR2_X1 U4432 ( .A1(n3678), .A2(n2149), .ZN(n3778) );
  NOR2_X1 U4433 ( .A1(n3650), .A2(n2342), .ZN(n3653) );
  NAND2_X1 U4434 ( .A1(n3652), .A2(n3651), .ZN(n3747) );
  OAI211_X1 U4435 ( .C1(n3653), .C2(n3747), .A(n3767), .B(n3722), .ZN(n3654)
         );
  NAND3_X1 U4436 ( .A1(n3654), .A2(n3770), .A3(n3766), .ZN(n3655) );
  AOI21_X1 U4437 ( .B1(n3721), .B2(n3655), .A(n3775), .ZN(n3657) );
  OAI21_X1 U4438 ( .B1(n3657), .B2(n3720), .A(n3656), .ZN(n3658) );
  NAND3_X1 U4439 ( .A1(n3777), .A2(n3776), .A3(n3658), .ZN(n3662) );
  OR2_X1 U4440 ( .A1(n3660), .A2(n3659), .ZN(n3669) );
  AND2_X1 U4441 ( .A1(n2408), .A2(DATAI_31_), .ZN(n3705) );
  INV_X1 U4442 ( .A(n3705), .ZN(n4104) );
  AND2_X1 U4443 ( .A1(n4103), .A2(n4104), .ZN(n3787) );
  AND2_X1 U4444 ( .A1(n2408), .A2(DATAI_30_), .ZN(n4111) );
  INV_X1 U4445 ( .A(n4111), .ZN(n4114) );
  NOR2_X1 U4446 ( .A1(n3801), .A2(n4114), .ZN(n3661) );
  NOR2_X1 U4447 ( .A1(n3787), .A2(n3661), .ZN(n3706) );
  OAI21_X1 U4448 ( .B1(n3664), .B2(n3663), .A(n3706), .ZN(n3667) );
  AOI211_X1 U4449 ( .C1(n3778), .C2(n3662), .A(n3669), .B(n3667), .ZN(n3672)
         );
  NAND2_X1 U4450 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  AND2_X1 U4451 ( .A1(n3666), .A2(n3665), .ZN(n3668) );
  AND2_X1 U4452 ( .A1(n3668), .A2(n2330), .ZN(n3781) );
  AOI21_X1 U4453 ( .B1(n3669), .B2(n3668), .A(n3667), .ZN(n3670) );
  INV_X1 U4454 ( .A(n3670), .ZN(n3788) );
  AOI21_X1 U4455 ( .B1(n3883), .B2(n3781), .A(n3788), .ZN(n3671) );
  AOI21_X1 U4456 ( .B1(n3672), .B2(n3785), .A(n3671), .ZN(n3676) );
  NOR2_X1 U4457 ( .A1(n4103), .A2(n4114), .ZN(n3675) );
  INV_X1 U4458 ( .A(n3801), .ZN(n3673) );
  NOR2_X1 U4459 ( .A1(n3673), .A2(n4111), .ZN(n3703) );
  OAI21_X1 U4460 ( .B1(n3703), .B2(n3704), .A(n3705), .ZN(n3674) );
  OAI21_X1 U4461 ( .B1(n3676), .B2(n3675), .A(n3674), .ZN(n3719) );
  OR2_X1 U4462 ( .A1(n3893), .A2(n2149), .ZN(n3912) );
  INV_X1 U4463 ( .A(n3912), .ZN(n3689) );
  INV_X1 U4464 ( .A(n3777), .ZN(n3677) );
  NOR2_X1 U4465 ( .A1(n3678), .A2(n3677), .ZN(n3929) );
  NOR2_X1 U4466 ( .A1(n3680), .A2(n3679), .ZN(n3688) );
  XNOR2_X1 U4467 ( .A(n4044), .B(n4029), .ZN(n4015) );
  INV_X1 U4468 ( .A(n4015), .ZN(n4023) );
  INV_X1 U4469 ( .A(n3681), .ZN(n3683) );
  NAND2_X1 U4470 ( .A1(n3683), .A2(n3682), .ZN(n4003) );
  NAND2_X1 U4471 ( .A1(n4018), .A2(n4017), .ZN(n4057) );
  INV_X1 U4472 ( .A(n4057), .ZN(n3686) );
  NAND2_X1 U4473 ( .A1(n2817), .A2(n4718), .ZN(n3726) );
  NAND2_X1 U4474 ( .A1(n3684), .A2(n3726), .ZN(n4768) );
  INV_X1 U4475 ( .A(n4768), .ZN(n3685) );
  AND4_X1 U4476 ( .A1(n4023), .A2(n4003), .A3(n3686), .A4(n3685), .ZN(n3687)
         );
  NAND4_X1 U4477 ( .A1(n3689), .A2(n3929), .A3(n3688), .A4(n3687), .ZN(n3716)
         );
  INV_X1 U4478 ( .A(n4042), .ZN(n4038) );
  NOR4_X1 U4479 ( .A1(n4038), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3713)
         );
  NOR4_X1 U4480 ( .A1(n2212), .A2(n3694), .A3(n4673), .A4(n3693), .ZN(n3712)
         );
  NOR4_X1 U4481 ( .A1(n3696), .A2(n3695), .A3(n4093), .A4(n2693), .ZN(n3711)
         );
  NAND2_X1 U4482 ( .A1(n3953), .A2(n3951), .ZN(n3983) );
  AND2_X1 U4483 ( .A1(n3776), .A2(n3697), .ZN(n3956) );
  NAND4_X1 U4484 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3956), .ZN(n3708)
         );
  NOR2_X1 U4485 ( .A1(n3702), .A2(n3701), .ZN(n3897) );
  AOI21_X1 U4486 ( .B1(n3705), .B2(n3704), .A(n3703), .ZN(n3786) );
  NAND4_X1 U4487 ( .A1(n3883), .A2(n3897), .A3(n3786), .A4(n3706), .ZN(n3707)
         );
  NOR4_X1 U4488 ( .A1(n3983), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3710)
         );
  NAND4_X1 U4489 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3714)
         );
  OR4_X1 U4490 ( .A1(n3716), .A2(n2336), .A3(n3715), .A4(n3714), .ZN(n3718) );
  MUX2_X1 U4491 ( .A(n3719), .B(n3718), .S(n3717), .Z(n3791) );
  INV_X1 U4492 ( .A(n3720), .ZN(n3774) );
  INV_X1 U4493 ( .A(n3721), .ZN(n3771) );
  NAND2_X1 U4494 ( .A1(n3747), .A2(n3722), .ZN(n3765) );
  NAND3_X1 U4495 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3764) );
  OAI211_X1 U4496 ( .C1(n4693), .C2(n2733), .A(n3725), .B(n3726), .ZN(n3728)
         );
  NAND3_X1 U4497 ( .A1(n3728), .A2(n3727), .A3(n2694), .ZN(n3730) );
  OAI211_X1 U4498 ( .C1(n3732), .C2(n3731), .A(n3730), .B(n3729), .ZN(n3735)
         );
  NAND3_X1 U4499 ( .A1(n3735), .A2(n3734), .A3(n3733), .ZN(n3738) );
  NAND4_X1 U4500 ( .A1(n3738), .A2(n3737), .A3(n3750), .A4(n3736), .ZN(n3741)
         );
  NAND3_X1 U4501 ( .A1(n3741), .A2(n3740), .A3(n3739), .ZN(n3742) );
  NAND3_X1 U4502 ( .A1(n3742), .A2(n3748), .A3(n3751), .ZN(n3745) );
  NAND3_X1 U4503 ( .A1(n3745), .A2(n3744), .A3(n3743), .ZN(n3757) );
  NOR2_X1 U4504 ( .A1(n3747), .A2(n3746), .ZN(n3756) );
  NOR2_X1 U4505 ( .A1(n2355), .A2(n3749), .ZN(n3752) );
  NAND4_X1 U4506 ( .A1(n3752), .A2(n2702), .A3(n3751), .A4(n3750), .ZN(n3754)
         );
  NAND2_X1 U4507 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  AOI22_X1 U4508 ( .A1(n3757), .A2(n3756), .B1(n3765), .B2(n3755), .ZN(n3762)
         );
  INV_X1 U4509 ( .A(n3758), .ZN(n3760) );
  NOR4_X1 U4510 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3763)
         );
  AOI21_X1 U4511 ( .B1(n3765), .B2(n3764), .A(n3763), .ZN(n3768) );
  OAI21_X1 U4512 ( .B1(n3768), .B2(n2352), .A(n3767), .ZN(n3769) );
  OAI221_X1 U4513 ( .B1(n3771), .B2(n3770), .C1(n3771), .C2(n3769), .A(n3953), 
        .ZN(n3773) );
  AOI221_X1 U4514 ( .B1(n3775), .B2(n3774), .C1(n3773), .C2(n3774), .A(n3772), 
        .ZN(n3780) );
  NAND2_X1 U4515 ( .A1(n3777), .A2(n3776), .ZN(n3779) );
  OAI21_X1 U4516 ( .B1(n3780), .B2(n3779), .A(n3778), .ZN(n3784) );
  INV_X1 U4517 ( .A(n3781), .ZN(n3782) );
  AOI211_X1 U4518 ( .C1(n3785), .C2(n3784), .A(n3783), .B(n3782), .ZN(n3789)
         );
  OAI22_X1 U4519 ( .A1(n3789), .A2(n3788), .B1(n3787), .B2(n3786), .ZN(n3790)
         );
  XNOR2_X1 U4520 ( .A(n3792), .B(n3863), .ZN(n3800) );
  NAND2_X1 U4521 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  OAI211_X1 U4522 ( .C1(n3797), .C2(n3796), .A(B_REG_SCAN_IN), .B(n3795), .ZN(
        n3798) );
  OAI21_X1 U4523 ( .B1(n3800), .B2(n3799), .A(n3798), .ZN(U3239) );
  MUX2_X1 U4524 ( .A(DATAO_REG_30__SCAN_IN), .B(n3801), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4525 ( .A(DATAO_REG_25__SCAN_IN), .B(n3900), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4526 ( .A(DATAO_REG_22__SCAN_IN), .B(n3960), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4527 ( .A(DATAO_REG_19__SCAN_IN), .B(n4044), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4528 ( .A(DATAO_REG_17__SCAN_IN), .B(n4076), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4529 ( .A(DATAO_REG_16__SCAN_IN), .B(n4060), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4530 ( .A(DATAO_REG_14__SCAN_IN), .B(n4097), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4531 ( .A(DATAO_REG_12__SCAN_IN), .B(n3802), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4532 ( .A(DATAO_REG_11__SCAN_IN), .B(n3803), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4533 ( .A(DATAO_REG_10__SCAN_IN), .B(n4678), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4534 ( .A(DATAO_REG_9__SCAN_IN), .B(n3804), .S(U4043), .Z(U3559) );
  MUX2_X1 U4535 ( .A(DATAO_REG_5__SCAN_IN), .B(n3805), .S(U4043), .Z(U3555) );
  MUX2_X1 U4536 ( .A(DATAO_REG_4__SCAN_IN), .B(n3806), .S(U4043), .Z(U3554) );
  MUX2_X1 U4537 ( .A(DATAO_REG_3__SCAN_IN), .B(n3808), .S(U4043), .Z(U3553) );
  OAI211_X1 U4538 ( .C1(n3811), .C2(n3810), .A(n4662), .B(n3809), .ZN(n3818)
         );
  OAI211_X1 U4539 ( .C1(n3814), .C2(n3813), .A(n4666), .B(n3812), .ZN(n3817)
         );
  AOI22_X1 U4540 ( .A1(n4671), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3816) );
  NAND2_X1 U4541 ( .A1(n4563), .A2(n4500), .ZN(n3815) );
  NAND4_X1 U4542 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(U3241)
         );
  AOI211_X1 U4543 ( .C1(n3821), .C2(n3820), .A(n3819), .B(n4654), .ZN(n3822)
         );
  INV_X1 U4544 ( .A(n3822), .ZN(n3829) );
  INV_X1 U4545 ( .A(n4671), .ZN(n4567) );
  INV_X1 U4546 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4333) );
  OAI21_X1 U4547 ( .B1(n4567), .B2(n4333), .A(n3823), .ZN(n3824) );
  AOI21_X1 U4548 ( .B1(n4498), .B2(n4563), .A(n3824), .ZN(n3828) );
  OAI211_X1 U4549 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3826), .A(n4662), .B(n3825), 
        .ZN(n3827) );
  NAND3_X1 U4550 ( .A1(n3829), .A2(n3828), .A3(n3827), .ZN(U3243) );
  INV_X1 U4551 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U4552 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3844), .ZN(n3837) );
  INV_X1 U4553 ( .A(n3844), .ZN(n4748) );
  INV_X1 U4554 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4555 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3844), .B1(n4748), .B2(
        n4088), .ZN(n4632) );
  INV_X1 U4556 ( .A(n3846), .ZN(n4496) );
  NAND2_X1 U4557 ( .A1(n4496), .A2(REG2_REG_11__SCAN_IN), .ZN(n3830) );
  INV_X1 U4558 ( .A(n4752), .ZN(n4606) );
  NAND2_X1 U4559 ( .A1(n4608), .A2(REG2_REG_13__SCAN_IN), .ZN(n4607) );
  INV_X1 U4560 ( .A(n4608), .ZN(n4751) );
  NAND2_X1 U4561 ( .A1(n3849), .A2(n3835), .ZN(n3836) );
  XNOR2_X1 U4562 ( .A(n4749), .B(n3835), .ZN(n4621) );
  NAND2_X1 U4563 ( .A1(REG2_REG_14__SCAN_IN), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U4564 ( .A1(n3836), .A2(n4620), .ZN(n4631) );
  NAND2_X1 U4565 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  XNOR2_X1 U4566 ( .A(n3853), .B(n3838), .ZN(n4641) );
  NOR2_X1 U4567 ( .A1(REG2_REG_16__SCAN_IN), .A2(n4641), .ZN(n4640) );
  NOR2_X1 U4568 ( .A1(n3853), .A2(n3838), .ZN(n3839) );
  NOR2_X1 U4569 ( .A1(n4640), .A2(n3839), .ZN(n4652) );
  INV_X1 U4570 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U4571 ( .A1(n4653), .A2(n4275), .ZN(n3841) );
  OR2_X1 U4572 ( .A1(n4653), .A2(n4275), .ZN(n3840) );
  NAND2_X1 U4573 ( .A1(n3841), .A2(n3840), .ZN(n4651) );
  AOI22_X1 U4574 ( .A1(n3857), .A2(REG2_REG_18__SCAN_IN), .B1(n4285), .B2(
        n4744), .ZN(n4668) );
  NAND2_X1 U4575 ( .A1(n4667), .A2(n4668), .ZN(n4665) );
  OAI21_X1 U4576 ( .B1(n4285), .B2(n4744), .A(n4665), .ZN(n3843) );
  INV_X1 U4577 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4286) );
  MUX2_X1 U4578 ( .A(n4286), .B(REG2_REG_19__SCAN_IN), .S(n3863), .Z(n3842) );
  XNOR2_X1 U4579 ( .A(n3843), .B(n3842), .ZN(n3867) );
  AOI22_X1 U4580 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3844), .B1(n4748), .B2(
        n4196), .ZN(n4629) );
  AOI22_X1 U4581 ( .A1(n4608), .A2(REG1_REG_13__SCAN_IN), .B1(n2537), .B2(
        n4751), .ZN(n4615) );
  NAND2_X1 U4582 ( .A1(n4752), .A2(n3847), .ZN(n3848) );
  NAND2_X1 U4583 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U4584 ( .A1(n3849), .A2(n3850), .ZN(n3851) );
  NAND2_X1 U4585 ( .A1(n3851), .A2(n4618), .ZN(n4628) );
  NAND2_X1 U4586 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  XNOR2_X1 U4587 ( .A(n3853), .B(n3852), .ZN(n4639) );
  NOR2_X1 U4588 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4639), .ZN(n4638) );
  NOR2_X1 U4589 ( .A1(n3853), .A2(n3852), .ZN(n3854) );
  NAND2_X1 U4590 ( .A1(n4653), .A2(n4429), .ZN(n3856) );
  OR2_X1 U4591 ( .A1(n4653), .A2(n4429), .ZN(n3855) );
  NAND2_X1 U4592 ( .A1(n3856), .A2(n3855), .ZN(n4647) );
  AOI22_X1 U4593 ( .A1(n3857), .A2(REG1_REG_18__SCAN_IN), .B1(n3858), .B2(
        n4744), .ZN(n4664) );
  OAI21_X1 U4594 ( .B1(n3858), .B2(n4744), .A(n4661), .ZN(n3860) );
  XNOR2_X1 U4595 ( .A(n3863), .B(n4422), .ZN(n3859) );
  XNOR2_X1 U4596 ( .A(n3860), .B(n3859), .ZN(n3865) );
  NAND2_X1 U4597 ( .A1(n4671), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3861) );
  OAI211_X1 U4598 ( .C1(n4669), .C2(n3863), .A(n3862), .B(n3861), .ZN(n3864)
         );
  OAI21_X1 U4599 ( .B1(n3867), .B2(n4654), .A(n3866), .ZN(U3259) );
  INV_X1 U4600 ( .A(n3868), .ZN(n3876) );
  NOR2_X1 U4601 ( .A1(n3869), .A2(n4711), .ZN(n3873) );
  INV_X1 U4602 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3871) );
  OAI22_X1 U4603 ( .A1(n4089), .A2(n3871), .B1(n3870), .B2(n4050), .ZN(n3872)
         );
  AOI211_X1 U4604 ( .C1(n3874), .C2(n4089), .A(n3873), .B(n3872), .ZN(n3875)
         );
  OAI21_X1 U4605 ( .B1(n3876), .B2(n4101), .A(n3875), .ZN(U3262) );
  XNOR2_X1 U4606 ( .A(n3877), .B(n3883), .ZN(n4124) );
  INV_X1 U4607 ( .A(n3878), .ZN(n3903) );
  AOI21_X1 U4608 ( .B1(n3886), .B2(n3903), .A(n3879), .ZN(n4122) );
  INV_X1 U4609 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4291) );
  OAI22_X1 U4610 ( .A1(n4534), .A2(n4291), .B1(n3880), .B2(n4050), .ZN(n3881)
         );
  AOI21_X1 U4611 ( .B1(n4122), .B2(n4689), .A(n3881), .ZN(n3891) );
  OAI21_X1 U4612 ( .B1(n3884), .B2(n3883), .A(n3882), .ZN(n3885) );
  NAND2_X1 U4613 ( .A1(n3885), .A2(n4719), .ZN(n3889) );
  AOI22_X1 U4614 ( .A1(n3887), .A2(n4696), .B1(n4695), .B2(n3886), .ZN(n3888)
         );
  OAI211_X1 U4615 ( .C1(n3915), .C2(n4698), .A(n3889), .B(n3888), .ZN(n4121)
         );
  NAND2_X1 U4616 ( .A1(n4121), .A2(n4534), .ZN(n3890) );
  OAI211_X1 U4617 ( .C1(n4124), .C2(n4101), .A(n3891), .B(n3890), .ZN(U3263)
         );
  XNOR2_X1 U4618 ( .A(n3892), .B(n3897), .ZN(n4126) );
  INV_X1 U4619 ( .A(n4126), .ZN(n3910) );
  INV_X1 U4620 ( .A(n3893), .ZN(n3894) );
  NAND2_X1 U4621 ( .A1(n3895), .A2(n3894), .ZN(n3896) );
  XOR2_X1 U4622 ( .A(n3897), .B(n3896), .Z(n3902) );
  OAI22_X1 U4623 ( .A1(n3898), .A2(n4722), .B1(n4675), .B2(n3904), .ZN(n3899)
         );
  AOI21_X1 U4624 ( .B1(n4679), .B2(n3900), .A(n3899), .ZN(n3901) );
  OAI21_X1 U4625 ( .B1(n3902), .B2(n4681), .A(n3901), .ZN(n4125) );
  INV_X1 U4626 ( .A(n3922), .ZN(n3905) );
  OAI21_X1 U4627 ( .B1(n3905), .B2(n3904), .A(n3903), .ZN(n4458) );
  AOI22_X1 U4628 ( .A1(n4706), .A2(REG2_REG_26__SCAN_IN), .B1(n3906), .B2(
        n4724), .ZN(n3907) );
  OAI21_X1 U4629 ( .B1(n4458), .B2(n4711), .A(n3907), .ZN(n3908) );
  AOI21_X1 U4630 ( .B1(n4125), .B2(n4534), .A(n3908), .ZN(n3909) );
  OAI21_X1 U4631 ( .B1(n3910), .B2(n4101), .A(n3909), .ZN(U3264) );
  XNOR2_X1 U4632 ( .A(n3911), .B(n3912), .ZN(n4129) );
  INV_X1 U4633 ( .A(n4129), .ZN(n3927) );
  XNOR2_X1 U4634 ( .A(n3913), .B(n3912), .ZN(n3919) );
  OAI22_X1 U4635 ( .A1(n3915), .A2(n4722), .B1(n4675), .B2(n3914), .ZN(n3916)
         );
  AOI21_X1 U4636 ( .B1(n4679), .B2(n3917), .A(n3916), .ZN(n3918) );
  OAI21_X1 U4637 ( .B1(n3919), .B2(n4681), .A(n3918), .ZN(n4128) );
  NAND2_X1 U4638 ( .A1(n3935), .A2(n3920), .ZN(n3921) );
  NAND2_X1 U4639 ( .A1(n3922), .A2(n3921), .ZN(n4462) );
  AOI22_X1 U4640 ( .A1(n4706), .A2(REG2_REG_25__SCAN_IN), .B1(n3923), .B2(
        n4724), .ZN(n3924) );
  OAI21_X1 U4641 ( .B1(n4462), .B2(n4711), .A(n3924), .ZN(n3925) );
  AOI21_X1 U4642 ( .B1(n4128), .B2(n4534), .A(n3925), .ZN(n3926) );
  OAI21_X1 U4643 ( .B1(n3927), .B2(n4101), .A(n3926), .ZN(U3265) );
  XNOR2_X1 U4644 ( .A(n3928), .B(n3929), .ZN(n4133) );
  INV_X1 U4645 ( .A(n4133), .ZN(n3941) );
  XNOR2_X1 U4646 ( .A(n3930), .B(n3929), .ZN(n3934) );
  OAI22_X1 U4647 ( .A1(n3931), .A2(n4722), .B1(n4675), .B2(n3936), .ZN(n3932)
         );
  AOI21_X1 U4648 ( .B1(n4679), .B2(n3974), .A(n3932), .ZN(n3933) );
  OAI21_X1 U4649 ( .B1(n3934), .B2(n4681), .A(n3933), .ZN(n4132) );
  OAI21_X1 U4650 ( .B1(n3946), .B2(n3936), .A(n3935), .ZN(n4466) );
  NOR2_X1 U4651 ( .A1(n4466), .A2(n4711), .ZN(n3939) );
  INV_X1 U4652 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4289) );
  OAI22_X1 U4653 ( .A1(n4089), .A2(n4289), .B1(n3937), .B2(n4050), .ZN(n3938)
         );
  AOI211_X1 U4654 ( .C1(n4132), .C2(n4089), .A(n3939), .B(n3938), .ZN(n3940)
         );
  OAI21_X1 U4655 ( .B1(n3941), .B2(n4101), .A(n3940), .ZN(U3266) );
  INV_X1 U4656 ( .A(n3942), .ZN(n3944) );
  NOR2_X1 U4657 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  XNOR2_X1 U4658 ( .A(n3945), .B(n3956), .ZN(n4138) );
  AOI21_X1 U4659 ( .B1(n3947), .B2(n4408), .A(n3946), .ZN(n4136) );
  INV_X1 U4660 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3949) );
  OAI22_X1 U4661 ( .A1(n4534), .A2(n3949), .B1(n3948), .B2(n4050), .ZN(n3950)
         );
  AOI21_X1 U4662 ( .B1(n4136), .B2(n4689), .A(n3950), .ZN(n3964) );
  INV_X1 U4663 ( .A(n3951), .ZN(n3952) );
  AOI21_X1 U4664 ( .B1(n3984), .B2(n3953), .A(n3952), .ZN(n3972) );
  OAI21_X1 U4665 ( .B1(n3972), .B2(n3971), .A(n3954), .ZN(n3955) );
  XOR2_X1 U4666 ( .A(n3956), .B(n3955), .Z(n3962) );
  OAI22_X1 U4667 ( .A1(n3958), .A2(n4722), .B1(n4675), .B2(n3957), .ZN(n3959)
         );
  AOI21_X1 U4668 ( .B1(n4679), .B2(n3960), .A(n3959), .ZN(n3961) );
  OAI21_X1 U4669 ( .B1(n3962), .B2(n4681), .A(n3961), .ZN(n4135) );
  NAND2_X1 U4670 ( .A1(n4135), .A2(n4534), .ZN(n3963) );
  OAI211_X1 U4671 ( .C1(n4138), .C2(n4101), .A(n3964), .B(n3963), .ZN(U3267)
         );
  OAI21_X1 U4672 ( .B1(n3965), .B2(n3971), .A(n3942), .ZN(n4411) );
  NAND2_X1 U4673 ( .A1(n3990), .A2(n3966), .ZN(n4407) );
  AND2_X1 U4674 ( .A1(n4407), .A2(n4689), .ZN(n3970) );
  INV_X1 U4675 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3968) );
  OAI22_X1 U4676 ( .A1(n4534), .A2(n3968), .B1(n3967), .B2(n4050), .ZN(n3969)
         );
  AOI21_X1 U4677 ( .B1(n3970), .B2(n4408), .A(n3969), .ZN(n3981) );
  XNOR2_X1 U4678 ( .A(n3972), .B(n3971), .ZN(n3979) );
  NAND2_X1 U4679 ( .A1(n3973), .A2(n4679), .ZN(n3976) );
  NAND2_X1 U4680 ( .A1(n3974), .A2(n4696), .ZN(n3975) );
  OAI211_X1 U4681 ( .C1(n4675), .C2(n3977), .A(n3976), .B(n3975), .ZN(n3978)
         );
  AOI21_X1 U4682 ( .B1(n3979), .B2(n4719), .A(n3978), .ZN(n4410) );
  OR2_X1 U4683 ( .A1(n4410), .A2(n4706), .ZN(n3980) );
  OAI211_X1 U4684 ( .C1(n4411), .C2(n4101), .A(n3981), .B(n3980), .ZN(U3268)
         );
  XNOR2_X1 U4685 ( .A(n3982), .B(n3983), .ZN(n4413) );
  INV_X1 U4686 ( .A(n4413), .ZN(n3998) );
  XNOR2_X1 U4687 ( .A(n3984), .B(n3983), .ZN(n3989) );
  OAI22_X1 U4688 ( .A1(n3985), .A2(n4722), .B1(n4675), .B2(n3991), .ZN(n3986)
         );
  AOI21_X1 U4689 ( .B1(n4679), .B2(n3987), .A(n3986), .ZN(n3988) );
  OAI21_X1 U4690 ( .B1(n3989), .B2(n4681), .A(n3988), .ZN(n4412) );
  INV_X1 U4691 ( .A(n4008), .ZN(n3992) );
  OAI21_X1 U4692 ( .B1(n3992), .B2(n3991), .A(n3990), .ZN(n4472) );
  NOR2_X1 U4693 ( .A1(n4472), .A2(n4711), .ZN(n3996) );
  INV_X1 U4694 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3994) );
  OAI22_X1 U4695 ( .A1(n4089), .A2(n3994), .B1(n3993), .B2(n4050), .ZN(n3995)
         );
  AOI211_X1 U4696 ( .C1(n4412), .C2(n4089), .A(n3996), .B(n3995), .ZN(n3997)
         );
  OAI21_X1 U4697 ( .B1(n3998), .B2(n4101), .A(n3997), .ZN(U3269) );
  XNOR2_X1 U4698 ( .A(n3999), .B(n4003), .ZN(n4417) );
  INV_X1 U4699 ( .A(n4417), .ZN(n4014) );
  NAND2_X1 U4700 ( .A1(n4001), .A2(n4000), .ZN(n4002) );
  XOR2_X1 U4701 ( .A(n4003), .B(n4002), .Z(n4007) );
  OAI22_X1 U4702 ( .A1(n4004), .A2(n4722), .B1(n4009), .B2(n4675), .ZN(n4005)
         );
  AOI21_X1 U4703 ( .B1(n4679), .B2(n4044), .A(n4005), .ZN(n4006) );
  OAI21_X1 U4704 ( .B1(n4007), .B2(n4681), .A(n4006), .ZN(n4416) );
  OAI21_X1 U4705 ( .B1(n4031), .B2(n4009), .A(n4008), .ZN(n4476) );
  NOR2_X1 U4706 ( .A1(n4476), .A2(n4711), .ZN(n4012) );
  INV_X1 U4707 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4288) );
  OAI22_X1 U4708 ( .A1(n4089), .A2(n4288), .B1(n4010), .B2(n4050), .ZN(n4011)
         );
  AOI211_X1 U4709 ( .C1(n4416), .C2(n4089), .A(n4012), .B(n4011), .ZN(n4013)
         );
  OAI21_X1 U4710 ( .B1(n4014), .B2(n4101), .A(n4013), .ZN(U3270) );
  XNOR2_X1 U4711 ( .A(n4016), .B(n4015), .ZN(n4421) );
  INV_X1 U4712 ( .A(n4421), .ZN(n4036) );
  INV_X1 U4713 ( .A(n4017), .ZN(n4019) );
  OAI21_X1 U4714 ( .B1(n4056), .B2(n4019), .A(n4018), .ZN(n4043) );
  INV_X1 U4715 ( .A(n4020), .ZN(n4022) );
  OAI21_X1 U4716 ( .B1(n4043), .B2(n4022), .A(n4021), .ZN(n4024) );
  XNOR2_X1 U4717 ( .A(n4024), .B(n4023), .ZN(n4028) );
  OAI22_X1 U4718 ( .A1(n4025), .A2(n4722), .B1(n4675), .B2(n4029), .ZN(n4026)
         );
  AOI21_X1 U4719 ( .B1(n4679), .B2(n4059), .A(n4026), .ZN(n4027) );
  OAI21_X1 U4720 ( .B1(n4028), .B2(n4681), .A(n4027), .ZN(n4420) );
  NOR2_X1 U4721 ( .A1(n4039), .A2(n4029), .ZN(n4030) );
  OR2_X1 U4722 ( .A1(n4031), .A2(n4030), .ZN(n4480) );
  AOI22_X1 U4723 ( .A1(n4706), .A2(REG2_REG_19__SCAN_IN), .B1(n4032), .B2(
        n4724), .ZN(n4033) );
  OAI21_X1 U4724 ( .B1(n4480), .B2(n4711), .A(n4033), .ZN(n4034) );
  AOI21_X1 U4725 ( .B1(n4420), .B2(n4534), .A(n4034), .ZN(n4035) );
  OAI21_X1 U4726 ( .B1(n4036), .B2(n4101), .A(n4035), .ZN(U3271) );
  XNOR2_X1 U4727 ( .A(n4037), .B(n4038), .ZN(n4426) );
  INV_X1 U4728 ( .A(n4064), .ZN(n4041) );
  INV_X1 U4729 ( .A(n4039), .ZN(n4040) );
  OAI211_X1 U4730 ( .C1(n4041), .C2(n4047), .A(n4040), .B(n4812), .ZN(n4424)
         );
  XNOR2_X1 U4731 ( .A(n4043), .B(n4042), .ZN(n4049) );
  NAND2_X1 U4732 ( .A1(n4076), .A2(n4679), .ZN(n4046) );
  NAND2_X1 U4733 ( .A1(n4044), .A2(n4696), .ZN(n4045) );
  OAI211_X1 U4734 ( .C1(n4675), .C2(n4047), .A(n4046), .B(n4045), .ZN(n4048)
         );
  AOI21_X1 U4735 ( .B1(n4049), .B2(n4719), .A(n4048), .ZN(n4425) );
  OAI21_X1 U4736 ( .B1(n2822), .B2(n4424), .A(n4425), .ZN(n4053) );
  OAI22_X1 U4737 ( .A1(n4534), .A2(n4285), .B1(n4051), .B2(n4050), .ZN(n4052)
         );
  AOI21_X1 U4738 ( .B1(n4053), .B2(n4534), .A(n4052), .ZN(n4054) );
  OAI21_X1 U4739 ( .B1(n4426), .B2(n4101), .A(n4054), .ZN(U3272) );
  XNOR2_X1 U4740 ( .A(n4055), .B(n4057), .ZN(n4428) );
  INV_X1 U4741 ( .A(n4428), .ZN(n4071) );
  XOR2_X1 U4742 ( .A(n4057), .B(n4056), .Z(n4063) );
  NOR2_X1 U4743 ( .A1(n4065), .A2(n4675), .ZN(n4058) );
  AOI21_X1 U4744 ( .B1(n4059), .B2(n4696), .A(n4058), .ZN(n4062) );
  NAND2_X1 U4745 ( .A1(n4060), .A2(n4679), .ZN(n4061) );
  OAI211_X1 U4746 ( .C1(n4063), .C2(n4681), .A(n4062), .B(n4061), .ZN(n4427)
         );
  INV_X1 U4747 ( .A(n4079), .ZN(n4066) );
  OAI21_X1 U4748 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4485) );
  NOR2_X1 U4749 ( .A1(n4485), .A2(n4711), .ZN(n4069) );
  OAI22_X1 U4750 ( .A1(n4534), .A2(n4275), .B1(n4067), .B2(n4050), .ZN(n4068)
         );
  AOI211_X1 U4751 ( .C1(n4427), .C2(n4534), .A(n4069), .B(n4068), .ZN(n4070)
         );
  OAI21_X1 U4752 ( .B1(n4071), .B2(n4101), .A(n4070), .ZN(U3273) );
  XNOR2_X1 U4753 ( .A(n4072), .B(n2204), .ZN(n4432) );
  INV_X1 U4754 ( .A(n4432), .ZN(n4085) );
  OAI211_X1 U4755 ( .C1(n4074), .C2(n2204), .A(n4073), .B(n4719), .ZN(n4078)
         );
  NOR2_X1 U4756 ( .A1(n4080), .A2(n4675), .ZN(n4075) );
  AOI21_X1 U4757 ( .B1(n4076), .B2(n4696), .A(n4075), .ZN(n4077) );
  OAI211_X1 U4758 ( .C1(n4503), .C2(n4698), .A(n4078), .B(n4077), .ZN(n4431)
         );
  OAI21_X1 U4759 ( .B1(n4087), .B2(n4080), .A(n4079), .ZN(n4490) );
  NOR2_X1 U4760 ( .A1(n4490), .A2(n4711), .ZN(n4083) );
  INV_X1 U4761 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4081) );
  OAI22_X1 U4762 ( .A1(n4089), .A2(n4081), .B1(n4511), .B2(n4050), .ZN(n4082)
         );
  AOI211_X1 U4763 ( .C1(n4431), .C2(n4089), .A(n4083), .B(n4082), .ZN(n4084)
         );
  OAI21_X1 U4764 ( .B1(n4085), .B2(n4101), .A(n4084), .ZN(U3274) );
  XOR2_X1 U4765 ( .A(n4086), .B(n4093), .Z(n4439) );
  AOI21_X1 U4766 ( .B1(n4519), .B2(n4442), .A(n4087), .ZN(n4436) );
  OAI22_X1 U4767 ( .A1(n4089), .A2(n4088), .B1(n4527), .B2(n4050), .ZN(n4099)
         );
  OAI22_X1 U4768 ( .A1(n4513), .A2(n4722), .B1(n4675), .B2(n4090), .ZN(n4096)
         );
  INV_X1 U4769 ( .A(n4091), .ZN(n4092) );
  AOI211_X1 U4770 ( .C1(n4094), .C2(n4093), .A(n4681), .B(n4092), .ZN(n4095)
         );
  AOI211_X1 U4771 ( .C1(n4679), .C2(n4097), .A(n4096), .B(n4095), .ZN(n4438)
         );
  NOR2_X1 U4772 ( .A1(n4438), .A2(n4706), .ZN(n4098) );
  AOI211_X1 U4773 ( .C1(n4436), .C2(n4689), .A(n4099), .B(n4098), .ZN(n4100)
         );
  OAI21_X1 U4774 ( .B1(n4101), .B2(n4439), .A(n4100), .ZN(U3275) );
  NAND2_X1 U4775 ( .A1(n4107), .A2(n4114), .ZN(n4108) );
  XNOR2_X1 U4776 ( .A(n4108), .B(n4104), .ZN(n4530) );
  NAND2_X1 U4777 ( .A1(n4530), .A2(n4112), .ZN(n4106) );
  NAND2_X1 U4778 ( .A1(n4103), .A2(n4102), .ZN(n4113) );
  OAI21_X1 U4779 ( .B1(n4104), .B2(n4675), .A(n4113), .ZN(n4529) );
  NAND2_X1 U4780 ( .A1(n4529), .A2(n4836), .ZN(n4105) );
  OAI211_X1 U4781 ( .C1(n4836), .C2(n2804), .A(n4106), .B(n4105), .ZN(U3549)
         );
  INV_X1 U4782 ( .A(n4107), .ZN(n4110) );
  INV_X1 U4783 ( .A(n4108), .ZN(n4109) );
  NAND2_X1 U4784 ( .A1(n4535), .A2(n4112), .ZN(n4116) );
  OAI21_X1 U4785 ( .B1(n4114), .B2(n4675), .A(n4113), .ZN(n4533) );
  NAND2_X1 U4786 ( .A1(n4533), .A2(n4836), .ZN(n4115) );
  OAI211_X1 U4787 ( .C1(n4836), .C2(n3409), .A(n4116), .B(n4115), .ZN(U3548)
         );
  AOI21_X1 U4788 ( .B1(n4812), .B2(n4118), .A(n4117), .ZN(n4119) );
  OAI21_X1 U4789 ( .B1(n4120), .B2(n4801), .A(n4119), .ZN(n4453) );
  MUX2_X1 U4790 ( .A(REG1_REG_29__SCAN_IN), .B(n4453), .S(n4836), .Z(U3547) );
  AOI21_X1 U4791 ( .B1(n4812), .B2(n4122), .A(n4121), .ZN(n4123) );
  OAI21_X1 U4792 ( .B1(n4124), .B2(n4801), .A(n4123), .ZN(n4454) );
  MUX2_X1 U4793 ( .A(REG1_REG_27__SCAN_IN), .B(n4454), .S(n4836), .Z(U3545) );
  AOI21_X1 U4794 ( .B1(n4126), .B2(n4809), .A(n4125), .ZN(n4455) );
  MUX2_X1 U4795 ( .A(n4301), .B(n4455), .S(n4836), .Z(n4127) );
  OAI21_X1 U4796 ( .B1(n4435), .B2(n4458), .A(n4127), .ZN(U3544) );
  AOI21_X1 U4797 ( .B1(n4129), .B2(n4809), .A(n4128), .ZN(n4459) );
  MUX2_X1 U4798 ( .A(n4130), .B(n4459), .S(n4836), .Z(n4131) );
  OAI21_X1 U4799 ( .B1(n4435), .B2(n4462), .A(n4131), .ZN(U3543) );
  AOI21_X1 U4800 ( .B1(n4133), .B2(n4809), .A(n4132), .ZN(n4463) );
  MUX2_X1 U4801 ( .A(n4300), .B(n4463), .S(n4836), .Z(n4134) );
  OAI21_X1 U4802 ( .B1(n4435), .B2(n4466), .A(n4134), .ZN(U3542) );
  AOI21_X1 U4803 ( .B1(n4812), .B2(n4136), .A(n4135), .ZN(n4137) );
  OAI21_X1 U4804 ( .B1(n4138), .B2(n4801), .A(n4137), .ZN(n4467) );
  MUX2_X1 U4805 ( .A(REG1_REG_23__SCAN_IN), .B(n4467), .S(n4836), .Z(n4406) );
  NAND4_X1 U4806 ( .A1(REG2_REG_1__SCAN_IN), .A2(REG0_REG_1__SCAN_IN), .A3(
        n2413), .A4(n2400), .ZN(n4139) );
  NOR3_X1 U4807 ( .A1(REG2_REG_5__SCAN_IN), .A2(REG0_REG_4__SCAN_IN), .A3(
        n4139), .ZN(n4145) );
  NAND4_X1 U4808 ( .A1(REG1_REG_8__SCAN_IN), .A2(DATAI_8_), .A3(
        REG2_REG_7__SCAN_IN), .A4(n4581), .ZN(n4143) );
  NAND4_X1 U4809 ( .A1(REG0_REG_10__SCAN_IN), .A2(REG0_REG_9__SCAN_IN), .A3(
        REG2_REG_9__SCAN_IN), .A4(n4591), .ZN(n4142) );
  INV_X1 U4810 ( .A(DATAI_9_), .ZN(n4220) );
  INV_X1 U4811 ( .A(DATAI_10_), .ZN(n4754) );
  NAND4_X1 U4812 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4364), .A3(n4220), .A4(n4754), .ZN(n4141) );
  INV_X1 U4813 ( .A(DATAI_0_), .ZN(n4764) );
  NAND4_X1 U4814 ( .A1(REG0_REG_0__SCAN_IN), .A2(REG1_REG_3__SCAN_IN), .A3(
        REG1_REG_6__SCAN_IN), .A4(n4764), .ZN(n4140) );
  NOR4_X1 U4815 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4144)
         );
  NAND4_X1 U4816 ( .A1(REG2_REG_4__SCAN_IN), .A2(DATAI_2_), .A3(n4145), .A4(
        n4144), .ZN(n4171) );
  NOR4_X1 U4817 ( .A1(REG1_REG_12__SCAN_IN), .A2(REG2_REG_12__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(DATAO_REG_1__SCAN_IN), .ZN(n4146) );
  INV_X1 U4818 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4464) );
  NAND3_X1 U4819 ( .A1(REG1_REG_24__SCAN_IN), .A2(n4146), .A3(n4464), .ZN(
        n4170) );
  NAND4_X1 U4820 ( .A1(n4222), .A2(n4147), .A3(n4208), .A4(IR_REG_18__SCAN_IN), 
        .ZN(n4151) );
  INV_X1 U4821 ( .A(DATAI_23_), .ZN(n4743) );
  NAND4_X1 U4822 ( .A1(n4149), .A2(n4148), .A3(n4743), .A4(IR_REG_27__SCAN_IN), 
        .ZN(n4150) );
  NOR2_X1 U4823 ( .A1(n4151), .A2(n4150), .ZN(n4167) );
  AND4_X1 U4824 ( .A1(n4289), .A2(REG0_REG_22__SCAN_IN), .A3(IR_REG_3__SCAN_IN), .A4(IR_REG_0__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U4825 ( .A1(REG0_REG_14__SCAN_IN), .A2(DATAI_13_), .A3(
        REG0_REG_13__SCAN_IN), .A4(n4195), .ZN(n4153) );
  NAND4_X1 U4826 ( .A1(REG1_REG_11__SCAN_IN), .A2(DATAI_11_), .A3(
        REG1_REG_10__SCAN_IN), .A4(n3252), .ZN(n4152) );
  NOR2_X1 U4827 ( .A1(n4153), .A2(n4152), .ZN(n4159) );
  INV_X1 U4828 ( .A(DATAI_21_), .ZN(n4255) );
  NAND4_X1 U4829 ( .A1(REG0_REG_21__SCAN_IN), .A2(REG1_REG_20__SCAN_IN), .A3(
        n4255), .A4(n4288), .ZN(n4155) );
  NAND4_X1 U4830 ( .A1(DATAI_19_), .A2(DATAI_18_), .A3(REG2_REG_18__SCAN_IN), 
        .A4(n4286), .ZN(n4154) );
  NOR2_X1 U4831 ( .A1(n4155), .A2(n4154), .ZN(n4158) );
  NOR4_X1 U4832 ( .A1(IR_REG_29__SCAN_IN), .A2(REG3_REG_5__SCAN_IN), .A3(
        REG3_REG_3__SCAN_IN), .A4(n4385), .ZN(n4157) );
  NOR4_X1 U4833 ( .A1(REG2_REG_17__SCAN_IN), .A2(REG1_REG_16__SCAN_IN), .A3(
        REG0_REG_16__SCAN_IN), .A4(n4745), .ZN(n4156) );
  NAND4_X1 U4834 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4160)
         );
  NOR3_X1 U4835 ( .A1(IR_REG_23__SCAN_IN), .A2(ADDR_REG_5__SCAN_IN), .A3(n4160), .ZN(n4165) );
  AND4_X1 U4836 ( .A1(n4163), .A2(n4162), .A3(n4161), .A4(IR_REG_4__SCAN_IN), 
        .ZN(n4164) );
  NAND4_X1 U4837 ( .A1(n4167), .A2(n4166), .A3(n4165), .A4(n4164), .ZN(n4168)
         );
  NOR4_X1 U4838 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4190)
         );
  NAND4_X1 U4839 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_0__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U4840 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n4175) );
  NAND4_X1 U4841 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_12__SCAN_IN), .A3(
        n2534), .A4(n4203), .ZN(n4174) );
  INV_X1 U4842 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4512) );
  NAND4_X1 U4843 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG3_REG_16__SCAN_IN), .A3(
        n4172), .A4(n4512), .ZN(n4173) );
  NOR4_X1 U4844 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4189)
         );
  NOR4_X1 U4845 ( .A1(REG1_REG_15__SCAN_IN), .A2(REG0_REG_15__SCAN_IN), .A3(
        DATAI_15_), .A4(n2557), .ZN(n4188) );
  NOR4_X1 U4846 ( .A1(REG3_REG_28__SCAN_IN), .A2(DATAO_REG_26__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n4186) );
  NOR4_X1 U4847 ( .A1(DATAO_REG_6__SCAN_IN), .A2(DATAO_REG_8__SCAN_IN), .A3(
        DATAO_REG_20__SCAN_IN), .A4(DATAO_REG_24__SCAN_IN), .ZN(n4185) );
  NOR4_X1 U4848 ( .A1(REG2_REG_30__SCAN_IN), .A2(ADDR_REG_1__SCAN_IN), .A3(
        DATAI_30_), .A4(REG2_REG_31__SCAN_IN), .ZN(n4177) );
  NAND3_X1 U4849 ( .A1(DATAO_REG_2__SCAN_IN), .A2(DATAO_REG_15__SCAN_IN), .A3(
        n4177), .ZN(n4178) );
  NOR3_X1 U4850 ( .A1(REG1_REG_26__SCAN_IN), .A2(REG0_REG_25__SCAN_IN), .A3(
        n4178), .ZN(n4184) );
  NAND4_X1 U4851 ( .A1(ADDR_REG_18__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(
        DATAO_REG_28__SCAN_IN), .A4(DATAO_REG_21__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U4852 ( .A1(DATAO_REG_0__SCAN_IN), .A2(DATAO_REG_18__SCAN_IN), .A3(
        DATAO_REG_13__SCAN_IN), .A4(ADDR_REG_6__SCAN_IN), .ZN(n4181) );
  NAND4_X1 U4853 ( .A1(REG1_REG_28__SCAN_IN), .A2(REG2_REG_27__SCAN_IN), .A3(
        REG2_REG_25__SCAN_IN), .A4(ADDR_REG_13__SCAN_IN), .ZN(n4180) );
  NAND4_X1 U4854 ( .A1(REG0_REG_26__SCAN_IN), .A2(DATAO_REG_23__SCAN_IN), .A3(
        REG0_REG_31__SCAN_IN), .A4(DATAO_REG_7__SCAN_IN), .ZN(n4179) );
  NOR4_X1 U4855 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4183)
         );
  AND4_X1 U4856 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4187)
         );
  NAND4_X1 U4857 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4404)
         );
  AOI22_X1 U4858 ( .A1(n2423), .A2(keyinput14), .B1(keyinput76), .B2(n2456), 
        .ZN(n4191) );
  OAI221_X1 U4859 ( .B1(n2423), .B2(keyinput14), .C1(n2456), .C2(keyinput76), 
        .A(n4191), .ZN(n4200) );
  AOI22_X1 U4860 ( .A1(n2485), .A2(keyinput90), .B1(n2506), .B2(keyinput28), 
        .ZN(n4192) );
  OAI221_X1 U4861 ( .B1(n2485), .B2(keyinput90), .C1(n2506), .C2(keyinput28), 
        .A(n4192), .ZN(n4199) );
  AOI22_X1 U4862 ( .A1(n3244), .A2(keyinput39), .B1(keyinput5), .B2(n2523), 
        .ZN(n4193) );
  OAI221_X1 U4863 ( .B1(n3244), .B2(keyinput39), .C1(n2523), .C2(keyinput5), 
        .A(n4193), .ZN(n4198) );
  AOI22_X1 U4864 ( .A1(n4196), .A2(keyinput27), .B1(keyinput37), .B2(n4195), 
        .ZN(n4194) );
  OAI221_X1 U4865 ( .B1(n4196), .B2(keyinput27), .C1(n4195), .C2(keyinput37), 
        .A(n4194), .ZN(n4197) );
  NOR4_X1 U4866 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4250)
         );
  AOI22_X1 U4867 ( .A1(n2400), .A2(keyinput122), .B1(keyinput10), .B2(n4764), 
        .ZN(n4201) );
  OAI221_X1 U4868 ( .B1(n2400), .B2(keyinput122), .C1(n4764), .C2(keyinput10), 
        .A(n4201), .ZN(n4205) );
  AOI22_X1 U4869 ( .A1(n4203), .A2(keyinput58), .B1(keyinput21), .B2(n2413), 
        .ZN(n4202) );
  OAI221_X1 U4870 ( .B1(n4203), .B2(keyinput58), .C1(n2413), .C2(keyinput21), 
        .A(n4202), .ZN(n4204) );
  NOR2_X1 U4871 ( .A1(n4205), .A2(n4204), .ZN(n4249) );
  AOI22_X1 U4872 ( .A1(n4207), .A2(keyinput103), .B1(keyinput70), .B2(n4512), 
        .ZN(n4206) );
  OAI221_X1 U4873 ( .B1(n4207), .B2(keyinput103), .C1(n4512), .C2(keyinput70), 
        .A(n4206), .ZN(n4218) );
  XNOR2_X1 U4874 ( .A(IR_REG_3__SCAN_IN), .B(keyinput54), .ZN(n4212) );
  XNOR2_X1 U4875 ( .A(IR_REG_1__SCAN_IN), .B(keyinput56), .ZN(n4211) );
  XNOR2_X1 U4876 ( .A(IR_REG_8__SCAN_IN), .B(keyinput30), .ZN(n4210) );
  XNOR2_X1 U4877 ( .A(IR_REG_4__SCAN_IN), .B(keyinput4), .ZN(n4209) );
  AND4_X1 U4878 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4216)
         );
  XNOR2_X1 U4879 ( .A(keyinput117), .B(DATAI_8_), .ZN(n4215) );
  XNOR2_X1 U4880 ( .A(DATAI_2_), .B(keyinput84), .ZN(n4214) );
  XNOR2_X1 U4881 ( .A(IR_REG_0__SCAN_IN), .B(keyinput7), .ZN(n4213) );
  NAND4_X1 U4882 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  NOR2_X1 U4883 ( .A1(n4218), .A2(n4217), .ZN(n4248) );
  AOI22_X1 U4884 ( .A1(n4754), .A2(keyinput45), .B1(n4220), .B2(keyinput29), 
        .ZN(n4219) );
  OAI221_X1 U4885 ( .B1(n4754), .B2(keyinput45), .C1(n4220), .C2(keyinput29), 
        .A(n4219), .ZN(n4228) );
  AOI22_X1 U4886 ( .A1(n4223), .A2(keyinput57), .B1(n4222), .B2(keyinput71), 
        .ZN(n4221) );
  OAI221_X1 U4887 ( .B1(n4223), .B2(keyinput57), .C1(n4222), .C2(keyinput71), 
        .A(n4221), .ZN(n4227) );
  XNOR2_X1 U4888 ( .A(IR_REG_30__SCAN_IN), .B(keyinput19), .ZN(n4225) );
  XNOR2_X1 U4889 ( .A(keyinput20), .B(D_REG_0__SCAN_IN), .ZN(n4224) );
  NAND2_X1 U4890 ( .A1(n4225), .A2(n4224), .ZN(n4226) );
  NOR3_X1 U4891 ( .A1(n4228), .A2(n4227), .A3(n4226), .ZN(n4246) );
  XNOR2_X1 U4892 ( .A(n4736), .B(keyinput99), .ZN(n4239) );
  XNOR2_X1 U4893 ( .A(IR_REG_11__SCAN_IN), .B(keyinput127), .ZN(n4232) );
  XNOR2_X1 U4894 ( .A(IR_REG_9__SCAN_IN), .B(keyinput86), .ZN(n4231) );
  XNOR2_X1 U4895 ( .A(IR_REG_16__SCAN_IN), .B(keyinput98), .ZN(n4230) );
  XNOR2_X1 U4896 ( .A(IR_REG_18__SCAN_IN), .B(keyinput18), .ZN(n4229) );
  NAND4_X1 U4897 ( .A1(n4232), .A2(n4231), .A3(n4230), .A4(n4229), .ZN(n4238)
         );
  XNOR2_X1 U4898 ( .A(IR_REG_17__SCAN_IN), .B(keyinput64), .ZN(n4236) );
  XNOR2_X1 U4899 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput63), .ZN(n4235) );
  XNOR2_X1 U4900 ( .A(IR_REG_27__SCAN_IN), .B(keyinput51), .ZN(n4234) );
  XNOR2_X1 U4901 ( .A(IR_REG_29__SCAN_IN), .B(keyinput123), .ZN(n4233) );
  NAND4_X1 U4902 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4237)
         );
  NOR3_X1 U4903 ( .A1(n4239), .A2(n4238), .A3(n4237), .ZN(n4245) );
  INV_X1 U4904 ( .A(DATAI_13_), .ZN(n4750) );
  AOI22_X1 U4905 ( .A1(n4750), .A2(keyinput91), .B1(keyinput94), .B2(n2521), 
        .ZN(n4240) );
  OAI221_X1 U4906 ( .B1(n4750), .B2(keyinput91), .C1(n2521), .C2(keyinput94), 
        .A(n4240), .ZN(n4243) );
  INV_X1 U4907 ( .A(D_REG_2__SCAN_IN), .ZN(n4740) );
  AOI22_X1 U4908 ( .A1(n4738), .A2(keyinput95), .B1(keyinput32), .B2(n4740), 
        .ZN(n4241) );
  OAI221_X1 U4909 ( .B1(n4738), .B2(keyinput95), .C1(n4740), .C2(keyinput32), 
        .A(n4241), .ZN(n4242) );
  NOR2_X1 U4910 ( .A1(n4243), .A2(n4242), .ZN(n4244) );
  AND3_X1 U4911 ( .A1(n4246), .A2(n4245), .A3(n4244), .ZN(n4247) );
  AND4_X1 U4912 ( .A1(n4250), .A2(n4249), .A3(n4248), .A4(n4247), .ZN(n4283)
         );
  INV_X1 U4913 ( .A(DATAI_30_), .ZN(n4252) );
  AOI22_X1 U4914 ( .A1(n4252), .A2(keyinput66), .B1(n4743), .B2(keyinput111), 
        .ZN(n4251) );
  OAI221_X1 U4915 ( .B1(n4252), .B2(keyinput66), .C1(n4743), .C2(keyinput111), 
        .A(n4251), .ZN(n4261) );
  AOI22_X1 U4916 ( .A1(n4255), .A2(keyinput53), .B1(keyinput33), .B2(n4254), 
        .ZN(n4253) );
  OAI221_X1 U4917 ( .B1(n4255), .B2(keyinput53), .C1(n4254), .C2(keyinput33), 
        .A(n4253), .ZN(n4260) );
  AOI22_X1 U4918 ( .A1(n2600), .A2(keyinput46), .B1(keyinput52), .B2(n4745), 
        .ZN(n4256) );
  OAI221_X1 U4919 ( .B1(n2600), .B2(keyinput46), .C1(n4745), .C2(keyinput52), 
        .A(n4256), .ZN(n4259) );
  INV_X1 U4920 ( .A(DATAI_15_), .ZN(n4747) );
  AOI22_X1 U4921 ( .A1(n4747), .A2(keyinput97), .B1(keyinput34), .B2(n2557), 
        .ZN(n4257) );
  OAI221_X1 U4922 ( .B1(n4747), .B2(keyinput97), .C1(n2557), .C2(keyinput34), 
        .A(n4257), .ZN(n4258) );
  NOR4_X1 U4923 ( .A1(n4261), .A2(n4260), .A3(n4259), .A4(n4258), .ZN(n4282)
         );
  INV_X1 U4924 ( .A(D_REG_11__SCAN_IN), .ZN(n4735) );
  INV_X1 U4925 ( .A(D_REG_6__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U4926 ( .A1(n4735), .A2(keyinput82), .B1(n4737), .B2(keyinput116), 
        .ZN(n4262) );
  OAI221_X1 U4927 ( .B1(n4735), .B2(keyinput82), .C1(n4737), .C2(keyinput116), 
        .A(n4262), .ZN(n4269) );
  INV_X1 U4928 ( .A(D_REG_15__SCAN_IN), .ZN(n4733) );
  INV_X1 U4929 ( .A(D_REG_14__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U4930 ( .A1(n4733), .A2(keyinput26), .B1(n4734), .B2(keyinput0), 
        .ZN(n4263) );
  OAI221_X1 U4931 ( .B1(n4733), .B2(keyinput26), .C1(n4734), .C2(keyinput0), 
        .A(n4263), .ZN(n4268) );
  AOI22_X1 U4932 ( .A1(n4732), .A2(keyinput2), .B1(keyinput40), .B2(n4731), 
        .ZN(n4264) );
  OAI221_X1 U4933 ( .B1(n4732), .B2(keyinput2), .C1(n4731), .C2(keyinput40), 
        .A(n4264), .ZN(n4267) );
  INV_X1 U4934 ( .A(D_REG_29__SCAN_IN), .ZN(n4729) );
  INV_X1 U4935 ( .A(D_REG_26__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U4936 ( .A1(n4729), .A2(keyinput17), .B1(keyinput83), .B2(n4730), 
        .ZN(n4265) );
  OAI221_X1 U4937 ( .B1(n4729), .B2(keyinput17), .C1(n4730), .C2(keyinput83), 
        .A(n4265), .ZN(n4266) );
  NOR4_X1 U4938 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n4281)
         );
  AOI22_X1 U4939 ( .A1(n4560), .A2(keyinput23), .B1(n4271), .B2(keyinput114), 
        .ZN(n4270) );
  OAI221_X1 U4940 ( .B1(n4560), .B2(keyinput23), .C1(n4271), .C2(keyinput114), 
        .A(n4270), .ZN(n4279) );
  AOI22_X1 U4941 ( .A1(n4581), .A2(keyinput106), .B1(n3313), .B2(keyinput55), 
        .ZN(n4272) );
  OAI221_X1 U4942 ( .B1(n4581), .B2(keyinput106), .C1(n3313), .C2(keyinput55), 
        .A(n4272), .ZN(n4278) );
  AOI22_X1 U4943 ( .A1(n4591), .A2(keyinput75), .B1(n3252), .B2(keyinput92), 
        .ZN(n4273) );
  OAI221_X1 U4944 ( .B1(n4591), .B2(keyinput75), .C1(n3252), .C2(keyinput92), 
        .A(n4273), .ZN(n4277) );
  AOI22_X1 U4945 ( .A1(n4275), .A2(keyinput3), .B1(keyinput24), .B2(n3352), 
        .ZN(n4274) );
  OAI221_X1 U4946 ( .B1(n4275), .B2(keyinput3), .C1(n3352), .C2(keyinput24), 
        .A(n4274), .ZN(n4276) );
  NOR4_X1 U4947 ( .A1(n4279), .A2(n4278), .A3(n4277), .A4(n4276), .ZN(n4280)
         );
  NAND4_X1 U4948 ( .A1(n4283), .A2(n4282), .A3(n4281), .A4(n4280), .ZN(n4402)
         );
  AOI22_X1 U4949 ( .A1(n4286), .A2(keyinput93), .B1(keyinput11), .B2(n4285), 
        .ZN(n4284) );
  OAI221_X1 U4950 ( .B1(n4286), .B2(keyinput93), .C1(n4285), .C2(keyinput11), 
        .A(n4284), .ZN(n4297) );
  AOI22_X1 U4951 ( .A1(n4289), .A2(keyinput35), .B1(keyinput38), .B2(n4288), 
        .ZN(n4287) );
  OAI221_X1 U4952 ( .B1(n4289), .B2(keyinput35), .C1(n4288), .C2(keyinput38), 
        .A(n4287), .ZN(n4296) );
  INV_X1 U4953 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4954 ( .A1(n4292), .A2(keyinput126), .B1(n4291), .B2(keyinput77), 
        .ZN(n4290) );
  OAI221_X1 U4955 ( .B1(n4292), .B2(keyinput126), .C1(n4291), .C2(keyinput77), 
        .A(n4290), .ZN(n4295) );
  INV_X1 U4956 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4532) );
  INV_X1 U4957 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U4958 ( .A1(n4532), .A2(keyinput96), .B1(n4537), .B2(keyinput109), 
        .ZN(n4293) );
  OAI221_X1 U4959 ( .B1(n4532), .B2(keyinput96), .C1(n4537), .C2(keyinput109), 
        .A(n4293), .ZN(n4294) );
  NOR4_X1 U4960 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(n4345)
         );
  AOI22_X1 U4961 ( .A1(n4433), .A2(keyinput8), .B1(n4418), .B2(keyinput105), 
        .ZN(n4298) );
  OAI221_X1 U4962 ( .B1(n4433), .B2(keyinput8), .C1(n4418), .C2(keyinput105), 
        .A(n4298), .ZN(n4311) );
  AOI22_X1 U4963 ( .A1(n4301), .A2(keyinput112), .B1(keyinput16), .B2(n4300), 
        .ZN(n4299) );
  OAI221_X1 U4964 ( .B1(n4301), .B2(keyinput112), .C1(n4300), .C2(keyinput16), 
        .A(n4299), .ZN(n4310) );
  AOI22_X1 U4965 ( .A1(n4304), .A2(keyinput67), .B1(n4303), .B2(keyinput79), 
        .ZN(n4302) );
  OAI221_X1 U4966 ( .B1(n4304), .B2(keyinput67), .C1(n4303), .C2(keyinput79), 
        .A(n4302), .ZN(n4309) );
  AOI22_X1 U4967 ( .A1(n4307), .A2(keyinput107), .B1(n4306), .B2(keyinput80), 
        .ZN(n4305) );
  OAI221_X1 U4968 ( .B1(n4307), .B2(keyinput107), .C1(n4306), .C2(keyinput80), 
        .A(n4305), .ZN(n4308) );
  NOR4_X1 U4969 ( .A1(n4311), .A2(n4310), .A3(n4309), .A4(n4308), .ZN(n4344)
         );
  AOI22_X1 U4970 ( .A1(n4314), .A2(keyinput125), .B1(n4313), .B2(keyinput49), 
        .ZN(n4312) );
  OAI221_X1 U4971 ( .B1(n4314), .B2(keyinput125), .C1(n4313), .C2(keyinput49), 
        .A(n4312), .ZN(n4327) );
  AOI22_X1 U4972 ( .A1(n4317), .A2(keyinput42), .B1(n4316), .B2(keyinput101), 
        .ZN(n4315) );
  OAI221_X1 U4973 ( .B1(n4317), .B2(keyinput42), .C1(n4316), .C2(keyinput101), 
        .A(n4315), .ZN(n4326) );
  AOI22_X1 U4974 ( .A1(n4320), .A2(keyinput113), .B1(n4319), .B2(keyinput102), 
        .ZN(n4318) );
  OAI221_X1 U4975 ( .B1(n4320), .B2(keyinput113), .C1(n4319), .C2(keyinput102), 
        .A(n4318), .ZN(n4325) );
  AOI22_X1 U4976 ( .A1(n4323), .A2(keyinput89), .B1(n4322), .B2(keyinput110), 
        .ZN(n4321) );
  OAI221_X1 U4977 ( .B1(n4323), .B2(keyinput89), .C1(n4322), .C2(keyinput110), 
        .A(n4321), .ZN(n4324) );
  NOR4_X1 U4978 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(n4343)
         );
  INV_X1 U4979 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4330) );
  INV_X1 U4980 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4981 ( .A1(n4330), .A2(keyinput15), .B1(n4329), .B2(keyinput85), 
        .ZN(n4328) );
  OAI221_X1 U4982 ( .B1(n4330), .B2(keyinput15), .C1(n4329), .C2(keyinput85), 
        .A(n4328), .ZN(n4341) );
  INV_X1 U4983 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4566) );
  INV_X1 U4984 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U4985 ( .A1(n4566), .A2(keyinput62), .B1(n4555), .B2(keyinput88), 
        .ZN(n4331) );
  OAI221_X1 U4986 ( .B1(n4566), .B2(keyinput62), .C1(n4555), .C2(keyinput88), 
        .A(n4331), .ZN(n4340) );
  INV_X1 U4987 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4988 ( .A1(n4334), .A2(keyinput47), .B1(n4333), .B2(keyinput6), 
        .ZN(n4332) );
  OAI221_X1 U4989 ( .B1(n4334), .B2(keyinput47), .C1(n4333), .C2(keyinput6), 
        .A(n4332), .ZN(n4339) );
  AOI22_X1 U4990 ( .A1(n4337), .A2(keyinput41), .B1(n4336), .B2(keyinput60), 
        .ZN(n4335) );
  OAI221_X1 U4991 ( .B1(n4337), .B2(keyinput41), .C1(n4336), .C2(keyinput60), 
        .A(n4335), .ZN(n4338) );
  NOR4_X1 U4992 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n4342)
         );
  NAND4_X1 U4993 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4401)
         );
  AOI22_X1 U4994 ( .A1(n4348), .A2(keyinput68), .B1(keyinput104), .B2(n4347), 
        .ZN(n4346) );
  OAI221_X1 U4995 ( .B1(n4348), .B2(keyinput68), .C1(n4347), .C2(keyinput104), 
        .A(n4346), .ZN(n4361) );
  AOI22_X1 U4996 ( .A1(n4351), .A2(keyinput100), .B1(keyinput115), .B2(n4350), 
        .ZN(n4349) );
  OAI221_X1 U4997 ( .B1(n4351), .B2(keyinput100), .C1(n4350), .C2(keyinput115), 
        .A(n4349), .ZN(n4360) );
  AOI22_X1 U4998 ( .A1(n4354), .A2(keyinput78), .B1(keyinput81), .B2(n4353), 
        .ZN(n4352) );
  OAI221_X1 U4999 ( .B1(n4354), .B2(keyinput78), .C1(n4353), .C2(keyinput81), 
        .A(n4352), .ZN(n4359) );
  AOI22_X1 U5000 ( .A1(n4357), .A2(keyinput13), .B1(keyinput118), .B2(n4356), 
        .ZN(n4355) );
  OAI221_X1 U5001 ( .B1(n4357), .B2(keyinput13), .C1(n4356), .C2(keyinput118), 
        .A(n4355), .ZN(n4358) );
  NOR4_X1 U5002 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4399)
         );
  INV_X1 U5003 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4775) );
  INV_X1 U5004 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U5005 ( .A1(n4775), .A2(keyinput61), .B1(keyinput22), .B2(n4769), 
        .ZN(n4362) );
  OAI221_X1 U5006 ( .B1(n4775), .B2(keyinput61), .C1(n4769), .C2(keyinput22), 
        .A(n4362), .ZN(n4372) );
  INV_X1 U5007 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4793) );
  AOI22_X1 U5008 ( .A1(n4793), .A2(keyinput87), .B1(keyinput59), .B2(n4364), 
        .ZN(n4363) );
  OAI221_X1 U5009 ( .B1(n4793), .B2(keyinput87), .C1(n4364), .C2(keyinput59), 
        .A(n4363), .ZN(n4371) );
  INV_X1 U5010 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5011 ( .A1(n4810), .A2(keyinput108), .B1(n4366), .B2(keyinput25), 
        .ZN(n4365) );
  OAI221_X1 U5012 ( .B1(n4810), .B2(keyinput108), .C1(n4366), .C2(keyinput25), 
        .A(n4365), .ZN(n4370) );
  INV_X1 U5013 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4368) );
  INV_X1 U5014 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4823) );
  AOI22_X1 U5015 ( .A1(n4368), .A2(keyinput72), .B1(keyinput74), .B2(n4823), 
        .ZN(n4367) );
  OAI221_X1 U5016 ( .B1(n4368), .B2(keyinput72), .C1(n4823), .C2(keyinput74), 
        .A(n4367), .ZN(n4369) );
  NOR4_X1 U5017 ( .A1(n4372), .A2(n4371), .A3(n4370), .A4(n4369), .ZN(n4398)
         );
  INV_X1 U5018 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4487) );
  INV_X1 U5019 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U5020 ( .A1(n4487), .A2(keyinput9), .B1(keyinput36), .B2(n4374), 
        .ZN(n4373) );
  OAI221_X1 U5021 ( .B1(n4487), .B2(keyinput9), .C1(n4374), .C2(keyinput36), 
        .A(n4373), .ZN(n4382) );
  INV_X1 U5022 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4470) );
  INV_X1 U5023 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5024 ( .A1(n4470), .A2(keyinput124), .B1(keyinput44), .B2(n4376), 
        .ZN(n4375) );
  OAI221_X1 U5025 ( .B1(n4470), .B2(keyinput124), .C1(n4376), .C2(keyinput44), 
        .A(n4375), .ZN(n4381) );
  INV_X1 U5026 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U5027 ( .A1(n4460), .A2(keyinput119), .B1(keyinput50), .B2(n4464), 
        .ZN(n4377) );
  OAI221_X1 U5028 ( .B1(n4460), .B2(keyinput119), .C1(n4464), .C2(keyinput50), 
        .A(n4377), .ZN(n4380) );
  INV_X1 U5029 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4456) );
  INV_X1 U5030 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U5031 ( .A1(n4456), .A2(keyinput73), .B1(keyinput69), .B2(n4448), 
        .ZN(n4378) );
  OAI221_X1 U5032 ( .B1(n4456), .B2(keyinput73), .C1(n4448), .C2(keyinput69), 
        .A(n4378), .ZN(n4379) );
  NOR4_X1 U5033 ( .A1(n4382), .A2(n4381), .A3(n4380), .A4(n4379), .ZN(n4397)
         );
  AOI22_X1 U5034 ( .A1(n4385), .A2(keyinput120), .B1(n4384), .B2(keyinput43), 
        .ZN(n4383) );
  OAI221_X1 U5035 ( .B1(n4385), .B2(keyinput120), .C1(n4384), .C2(keyinput43), 
        .A(n4383), .ZN(n4395) );
  AOI22_X1 U5036 ( .A1(n2435), .A2(keyinput65), .B1(n4387), .B2(keyinput1), 
        .ZN(n4386) );
  OAI221_X1 U5037 ( .B1(n2435), .B2(keyinput65), .C1(n4387), .C2(keyinput1), 
        .A(n4386), .ZN(n4394) );
  AOI22_X1 U5038 ( .A1(n4389), .A2(keyinput121), .B1(n4501), .B2(keyinput48), 
        .ZN(n4388) );
  OAI221_X1 U5039 ( .B1(n4389), .B2(keyinput121), .C1(n4501), .C2(keyinput48), 
        .A(n4388), .ZN(n4393) );
  INV_X1 U5040 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5041 ( .A1(n4391), .A2(keyinput31), .B1(n2534), .B2(keyinput12), 
        .ZN(n4390) );
  OAI221_X1 U5042 ( .B1(n4391), .B2(keyinput31), .C1(n2534), .C2(keyinput12), 
        .A(n4390), .ZN(n4392) );
  NOR4_X1 U5043 ( .A1(n4395), .A2(n4394), .A3(n4393), .A4(n4392), .ZN(n4396)
         );
  NAND4_X1 U5044 ( .A1(n4399), .A2(n4398), .A3(n4397), .A4(n4396), .ZN(n4400)
         );
  NOR3_X1 U5045 ( .A1(n4402), .A2(n4401), .A3(n4400), .ZN(n4403) );
  XOR2_X1 U5046 ( .A(n4404), .B(n4403), .Z(n4405) );
  XNOR2_X1 U5047 ( .A(n4406), .B(n4405), .ZN(U3541) );
  NAND3_X1 U5048 ( .A1(n4408), .A2(n4812), .A3(n4407), .ZN(n4409) );
  OAI211_X1 U5049 ( .C1(n4411), .C2(n4801), .A(n4410), .B(n4409), .ZN(n4468)
         );
  MUX2_X1 U5050 ( .A(REG1_REG_22__SCAN_IN), .B(n4468), .S(n4836), .Z(U3540) );
  AOI21_X1 U5051 ( .B1(n4413), .B2(n4809), .A(n4412), .ZN(n4469) );
  MUX2_X1 U5052 ( .A(n4414), .B(n4469), .S(n4836), .Z(n4415) );
  OAI21_X1 U5053 ( .B1(n4435), .B2(n4472), .A(n4415), .ZN(U3539) );
  AOI21_X1 U5054 ( .B1(n4417), .B2(n4809), .A(n4416), .ZN(n4473) );
  MUX2_X1 U5055 ( .A(n4418), .B(n4473), .S(n4836), .Z(n4419) );
  OAI21_X1 U5056 ( .B1(n4435), .B2(n4476), .A(n4419), .ZN(U3538) );
  AOI21_X1 U5057 ( .B1(n4421), .B2(n4809), .A(n4420), .ZN(n4477) );
  MUX2_X1 U5058 ( .A(n4422), .B(n4477), .S(n4836), .Z(n4423) );
  OAI21_X1 U5059 ( .B1(n4435), .B2(n4480), .A(n4423), .ZN(U3537) );
  OAI211_X1 U5060 ( .C1(n4426), .C2(n4801), .A(n4425), .B(n4424), .ZN(n4481)
         );
  MUX2_X1 U5061 ( .A(REG1_REG_18__SCAN_IN), .B(n4481), .S(n4836), .Z(U3536) );
  AOI21_X1 U5062 ( .B1(n4428), .B2(n4809), .A(n4427), .ZN(n4482) );
  MUX2_X1 U5063 ( .A(n4429), .B(n4482), .S(n4836), .Z(n4430) );
  OAI21_X1 U5064 ( .B1(n4435), .B2(n4485), .A(n4430), .ZN(U3535) );
  AOI21_X1 U5065 ( .B1(n4432), .B2(n4809), .A(n4431), .ZN(n4486) );
  MUX2_X1 U5066 ( .A(n4433), .B(n4486), .S(n4836), .Z(n4434) );
  OAI21_X1 U5067 ( .B1(n4435), .B2(n4490), .A(n4434), .ZN(U3534) );
  NAND2_X1 U5068 ( .A1(n4436), .A2(n4812), .ZN(n4437) );
  OAI211_X1 U5069 ( .C1(n4439), .C2(n4801), .A(n4438), .B(n4437), .ZN(n4491)
         );
  MUX2_X1 U5070 ( .A(REG1_REG_15__SCAN_IN), .B(n4491), .S(n4836), .Z(U3533) );
  INV_X1 U5071 ( .A(n4440), .ZN(n4445) );
  NAND3_X1 U5072 ( .A1(n4442), .A2(n4812), .A3(n4441), .ZN(n4443) );
  OAI211_X1 U5073 ( .C1(n4445), .C2(n4783), .A(n4444), .B(n4443), .ZN(n4492)
         );
  MUX2_X1 U5074 ( .A(REG1_REG_14__SCAN_IN), .B(n4492), .S(n4836), .Z(U3532) );
  NAND2_X1 U5075 ( .A1(n4530), .A2(n4449), .ZN(n4447) );
  NAND2_X1 U5076 ( .A1(n4529), .A2(n4824), .ZN(n4446) );
  OAI211_X1 U5077 ( .C1(n4824), .C2(n4448), .A(n4447), .B(n4446), .ZN(U3517)
         );
  INV_X1 U5078 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5079 ( .A1(n4535), .A2(n4449), .ZN(n4451) );
  NAND2_X1 U5080 ( .A1(n4533), .A2(n4824), .ZN(n4450) );
  OAI211_X1 U5081 ( .C1(n4824), .C2(n4452), .A(n4451), .B(n4450), .ZN(U3516)
         );
  MUX2_X1 U5082 ( .A(REG0_REG_29__SCAN_IN), .B(n4453), .S(n4824), .Z(U3515) );
  MUX2_X1 U5083 ( .A(REG0_REG_27__SCAN_IN), .B(n4454), .S(n4824), .Z(U3513) );
  MUX2_X1 U5084 ( .A(n4456), .B(n4455), .S(n4824), .Z(n4457) );
  OAI21_X1 U5085 ( .B1(n4458), .B2(n4489), .A(n4457), .ZN(U3512) );
  MUX2_X1 U5086 ( .A(n4460), .B(n4459), .S(n4824), .Z(n4461) );
  OAI21_X1 U5087 ( .B1(n4462), .B2(n4489), .A(n4461), .ZN(U3511) );
  MUX2_X1 U5088 ( .A(n4464), .B(n4463), .S(n4824), .Z(n4465) );
  OAI21_X1 U5089 ( .B1(n4466), .B2(n4489), .A(n4465), .ZN(U3510) );
  MUX2_X1 U5090 ( .A(REG0_REG_23__SCAN_IN), .B(n4467), .S(n4824), .Z(U3509) );
  MUX2_X1 U5091 ( .A(REG0_REG_22__SCAN_IN), .B(n4468), .S(n4824), .Z(U3508) );
  MUX2_X1 U5092 ( .A(n4470), .B(n4469), .S(n4824), .Z(n4471) );
  OAI21_X1 U5093 ( .B1(n4472), .B2(n4489), .A(n4471), .ZN(U3507) );
  INV_X1 U5094 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U5095 ( .A(n4474), .B(n4473), .S(n4824), .Z(n4475) );
  OAI21_X1 U5096 ( .B1(n4476), .B2(n4489), .A(n4475), .ZN(U3506) );
  INV_X1 U5097 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4478) );
  MUX2_X1 U5098 ( .A(n4478), .B(n4477), .S(n4824), .Z(n4479) );
  OAI21_X1 U5099 ( .B1(n4480), .B2(n4489), .A(n4479), .ZN(U3505) );
  MUX2_X1 U5100 ( .A(REG0_REG_18__SCAN_IN), .B(n4481), .S(n4824), .Z(U3503) );
  INV_X1 U5101 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4483) );
  MUX2_X1 U5102 ( .A(n4483), .B(n4482), .S(n4824), .Z(n4484) );
  OAI21_X1 U5103 ( .B1(n4485), .B2(n4489), .A(n4484), .ZN(U3501) );
  MUX2_X1 U5104 ( .A(n4487), .B(n4486), .S(n4824), .Z(n4488) );
  OAI21_X1 U5105 ( .B1(n4490), .B2(n4489), .A(n4488), .ZN(U3499) );
  MUX2_X1 U5106 ( .A(REG0_REG_15__SCAN_IN), .B(n4491), .S(n4824), .Z(U3497) );
  MUX2_X1 U5107 ( .A(REG0_REG_14__SCAN_IN), .B(n4492), .S(n4824), .Z(U3495) );
  MUX2_X1 U5108 ( .A(n2387), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5109 ( .A(DATAI_29_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5110 ( .A(n4494), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5111 ( .A(n4540), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5112 ( .A(DATAI_25_), .B(n4495), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5113 ( .A(n2733), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5114 ( .A(n2822), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5115 ( .A(n4496), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5116 ( .A(DATAI_9_), .B(n4497), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5117 ( .A(n4498), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5118 ( .A(n4499), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5119 ( .A(n4500), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  NOR2_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .ZN(n4644) );
  OAI22_X1 U5121 ( .A1(n4503), .A2(n4515), .B1(n4514), .B2(n4502), .ZN(n4504)
         );
  AOI211_X1 U5122 ( .C1(n4505), .C2(n4518), .A(n4644), .B(n4504), .ZN(n4510)
         );
  NOR2_X1 U5123 ( .A1(n4520), .A2(n2136), .ZN(n4506) );
  XOR2_X1 U5124 ( .A(n4507), .B(n4506), .Z(n4508) );
  NAND2_X1 U5125 ( .A1(n4508), .A2(n4524), .ZN(n4509) );
  OAI211_X1 U5126 ( .C1(n4528), .C2(n4511), .A(n4510), .B(n4509), .ZN(U3223)
         );
  NOR2_X1 U5127 ( .A1(STATE_REG_SCAN_IN), .A2(n4512), .ZN(n4636) );
  OAI22_X1 U5128 ( .A1(n4516), .A2(n4515), .B1(n4514), .B2(n4513), .ZN(n4517)
         );
  AOI211_X1 U5129 ( .C1(n4519), .C2(n4518), .A(n4636), .B(n4517), .ZN(n4526)
         );
  OAI21_X1 U5130 ( .B1(n4522), .B2(n2136), .A(n4521), .ZN(n4523) );
  OAI211_X1 U5131 ( .C1(n2295), .C2(n2136), .A(n4524), .B(n4523), .ZN(n4525)
         );
  OAI211_X1 U5132 ( .C1(n4528), .C2(n4527), .A(n4526), .B(n4525), .ZN(U3238)
         );
  AOI22_X1 U5133 ( .A1(n4530), .A2(n4689), .B1(n4534), .B2(n4529), .ZN(n4531)
         );
  OAI21_X1 U5134 ( .B1(n4534), .B2(n4532), .A(n4531), .ZN(U3260) );
  AOI22_X1 U5135 ( .A1(n4535), .A2(n4689), .B1(n4534), .B2(n4533), .ZN(n4536)
         );
  OAI21_X1 U5136 ( .B1(n4537), .B2(n4534), .A(n4536), .ZN(U3261) );
  INV_X1 U5137 ( .A(n4538), .ZN(n4539) );
  OAI21_X1 U5138 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4540), .A(n4539), .ZN(n4541)
         );
  XNOR2_X1 U5139 ( .A(n4541), .B(n4765), .ZN(n4544) );
  AOI22_X1 U5140 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4671), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4542) );
  OAI21_X1 U5141 ( .B1(n4544), .B2(n4543), .A(n4542), .ZN(U3240) );
  AOI211_X1 U5142 ( .C1(n4547), .C2(n4546), .A(n4545), .B(n4659), .ZN(n4551)
         );
  AOI211_X1 U5143 ( .C1(n2177), .C2(n4549), .A(n4548), .B(n4654), .ZN(n4550)
         );
  AOI211_X1 U5144 ( .C1(n4563), .C2(n4552), .A(n4551), .B(n4550), .ZN(n4554)
         );
  OAI211_X1 U5145 ( .C1(n4567), .C2(n4555), .A(n4554), .B(n4553), .ZN(U3245)
         );
  AOI211_X1 U5146 ( .C1(n2456), .C2(n4557), .A(n4556), .B(n4659), .ZN(n4562)
         );
  AOI211_X1 U5147 ( .C1(n4560), .C2(n4559), .A(n4558), .B(n4654), .ZN(n4561)
         );
  AOI211_X1 U5148 ( .C1(n4563), .C2(n4760), .A(n4562), .B(n4561), .ZN(n4565)
         );
  OAI211_X1 U5149 ( .C1(n4567), .C2(n4566), .A(n4565), .B(n4564), .ZN(U3246)
         );
  AOI211_X1 U5150 ( .C1(n4570), .C2(n4569), .A(n4568), .B(n4654), .ZN(n4572)
         );
  AOI211_X1 U5151 ( .C1(n4671), .C2(ADDR_REG_7__SCAN_IN), .A(n4572), .B(n4571), 
        .ZN(n4577) );
  AOI22_X1 U5152 ( .A1(REG1_REG_7__SCAN_IN), .A2(n4578), .B1(n4758), .B2(n2467), .ZN(n4574) );
  AOI21_X1 U5153 ( .B1(n4575), .B2(n4574), .A(n4659), .ZN(n4573) );
  OAI21_X1 U5154 ( .B1(n4575), .B2(n4574), .A(n4573), .ZN(n4576) );
  OAI211_X1 U5155 ( .C1(n4669), .C2(n4578), .A(n4577), .B(n4576), .ZN(U3247)
         );
  AOI211_X1 U5156 ( .C1(n4581), .C2(n4580), .A(n4579), .B(n4654), .ZN(n4584)
         );
  INV_X1 U5157 ( .A(n4582), .ZN(n4583) );
  AOI211_X1 U5158 ( .C1(n4671), .C2(ADDR_REG_8__SCAN_IN), .A(n4584), .B(n4583), 
        .ZN(n4588) );
  OAI211_X1 U5159 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4586), .A(n4662), .B(n4585), 
        .ZN(n4587) );
  OAI211_X1 U5160 ( .C1(n4669), .C2(n4757), .A(n4588), .B(n4587), .ZN(U3248)
         );
  AOI211_X1 U5161 ( .C1(n4591), .C2(n4590), .A(n4589), .B(n4654), .ZN(n4593)
         );
  AOI211_X1 U5162 ( .C1(n4671), .C2(ADDR_REG_10__SCAN_IN), .A(n4593), .B(n4592), .ZN(n4597) );
  OAI211_X1 U5163 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4595), .A(n4662), .B(n4594), .ZN(n4596) );
  OAI211_X1 U5164 ( .C1(n4669), .C2(n4755), .A(n4597), .B(n4596), .ZN(U3250)
         );
  AOI211_X1 U5165 ( .C1(n3352), .C2(n4599), .A(n4598), .B(n4654), .ZN(n4601)
         );
  AOI211_X1 U5166 ( .C1(n4671), .C2(ADDR_REG_12__SCAN_IN), .A(n4601), .B(n4600), .ZN(n4605) );
  OAI211_X1 U5167 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4603), .A(n4662), .B(n4602), .ZN(n4604) );
  OAI211_X1 U5168 ( .C1(n4669), .C2(n4606), .A(n4605), .B(n4604), .ZN(U3252)
         );
  OAI21_X1 U5169 ( .B1(n4608), .B2(REG2_REG_13__SCAN_IN), .A(n4607), .ZN(n4610) );
  OAI21_X1 U5170 ( .B1(n2159), .B2(n4610), .A(n4666), .ZN(n4609) );
  AOI21_X1 U5171 ( .B1(n2159), .B2(n4610), .A(n4609), .ZN(n4611) );
  AOI211_X1 U5172 ( .C1(n4671), .C2(ADDR_REG_13__SCAN_IN), .A(n4612), .B(n4611), .ZN(n4617) );
  OAI211_X1 U5173 ( .C1(n4615), .C2(n4614), .A(n4662), .B(n4613), .ZN(n4616)
         );
  OAI211_X1 U5174 ( .C1(n4669), .C2(n4751), .A(n4617), .B(n4616), .ZN(U3253)
         );
  OAI211_X1 U5175 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4619), .A(n4662), .B(n4618), .ZN(n4623) );
  OAI211_X1 U5176 ( .C1(REG2_REG_14__SCAN_IN), .C2(n4621), .A(n4666), .B(n4620), .ZN(n4622) );
  OAI211_X1 U5177 ( .C1(n4669), .C2(n4749), .A(n4623), .B(n4622), .ZN(n4624)
         );
  AOI211_X1 U5178 ( .C1(n4671), .C2(ADDR_REG_14__SCAN_IN), .A(n4625), .B(n4624), .ZN(n4626) );
  INV_X1 U5179 ( .A(n4626), .ZN(U3254) );
  OAI211_X1 U5180 ( .C1(n4629), .C2(n4628), .A(n4662), .B(n4627), .ZN(n4634)
         );
  OAI211_X1 U5181 ( .C1(n4632), .C2(n4631), .A(n4666), .B(n4630), .ZN(n4633)
         );
  OAI211_X1 U5182 ( .C1(n4669), .C2(n4748), .A(n4634), .B(n4633), .ZN(n4635)
         );
  AOI211_X1 U5183 ( .C1(n4671), .C2(ADDR_REG_15__SCAN_IN), .A(n4636), .B(n4635), .ZN(n4637) );
  INV_X1 U5184 ( .A(n4637), .ZN(U3255) );
  AOI21_X1 U5185 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4639), .A(n4638), .ZN(n4646) );
  AOI21_X1 U5186 ( .B1(REG2_REG_16__SCAN_IN), .B2(n4641), .A(n4640), .ZN(n4642) );
  OAI22_X1 U5187 ( .A1(n4642), .A2(n4654), .B1(n4746), .B2(n4669), .ZN(n4643)
         );
  AOI211_X1 U5188 ( .C1(n4671), .C2(ADDR_REG_16__SCAN_IN), .A(n4644), .B(n4643), .ZN(n4645) );
  OAI21_X1 U5189 ( .B1(n4646), .B2(n4659), .A(n4645), .ZN(U3256) );
  AOI21_X1 U5190 ( .B1(n4648), .B2(n4647), .A(n2151), .ZN(n4660) );
  INV_X1 U5191 ( .A(n4649), .ZN(n4650) );
  AOI21_X1 U5192 ( .B1(n4652), .B2(n4651), .A(n4650), .ZN(n4655) );
  OAI22_X1 U5193 ( .A1(n4655), .A2(n4654), .B1(n4653), .B2(n4669), .ZN(n4656)
         );
  AOI211_X1 U5194 ( .C1(n4671), .C2(ADDR_REG_17__SCAN_IN), .A(n4657), .B(n4656), .ZN(n4658) );
  OAI21_X1 U5195 ( .B1(n4660), .B2(n4659), .A(n4658), .ZN(U3257) );
  XNOR2_X1 U5196 ( .A(n4672), .B(n4673), .ZN(n4813) );
  XNOR2_X1 U5197 ( .A(n3340), .B(n4673), .ZN(n4682) );
  OAI22_X1 U5198 ( .A1(n4676), .A2(n4722), .B1(n4675), .B2(n4674), .ZN(n4677)
         );
  AOI21_X1 U5199 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n4680) );
  OAI21_X1 U5200 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4683) );
  AOI21_X1 U5201 ( .B1(n4720), .B2(n4813), .A(n4683), .ZN(n4815) );
  OAI22_X1 U5202 ( .A1(n4684), .A2(n4050), .B1(n3252), .B2(n4089), .ZN(n4685)
         );
  INV_X1 U5203 ( .A(n4685), .ZN(n4691) );
  AOI21_X1 U5204 ( .B1(n4688), .B2(n4687), .A(n4686), .ZN(n4811) );
  AOI22_X1 U5205 ( .A1(n4813), .A2(n4725), .B1(n4689), .B2(n4811), .ZN(n4690)
         );
  OAI211_X1 U5206 ( .C1(n4706), .C2(n4815), .A(n4691), .B(n4690), .ZN(U3279)
         );
  OAI21_X1 U5207 ( .B1(n4694), .B2(n4693), .A(n4692), .ZN(n4705) );
  INV_X1 U5208 ( .A(n2817), .ZN(n4699) );
  AOI22_X1 U5209 ( .A1(n2905), .A2(n4696), .B1(n4695), .B2(n2401), .ZN(n4697)
         );
  OAI21_X1 U5210 ( .B1(n4699), .B2(n4698), .A(n4697), .ZN(n4704) );
  OAI21_X1 U5211 ( .B1(n2693), .B2(n4701), .A(n4700), .ZN(n4772) );
  NOR2_X1 U5212 ( .A1(n4772), .A2(n4702), .ZN(n4703) );
  AOI211_X1 U5213 ( .C1(n4719), .C2(n4705), .A(n4704), .B(n4703), .ZN(n4770)
         );
  AOI22_X1 U5214 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4724), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4706), .ZN(n4715) );
  INV_X1 U5215 ( .A(n4707), .ZN(n4710) );
  NAND2_X1 U5216 ( .A1(n2401), .A2(n4708), .ZN(n4709) );
  NAND2_X1 U5217 ( .A1(n4710), .A2(n4709), .ZN(n4771) );
  OAI22_X1 U5218 ( .A1(n4772), .A2(n4712), .B1(n4711), .B2(n4771), .ZN(n4713)
         );
  INV_X1 U5219 ( .A(n4713), .ZN(n4714) );
  OAI211_X1 U5220 ( .C1(n4706), .C2(n4770), .A(n4715), .B(n4714), .ZN(U3289)
         );
  INV_X1 U5221 ( .A(n4716), .ZN(n4717) );
  NOR2_X1 U5222 ( .A1(n4718), .A2(n4717), .ZN(n4767) );
  NAND2_X1 U5223 ( .A1(n2690), .A2(n2822), .ZN(n4723) );
  OAI21_X1 U5224 ( .B1(n4720), .B2(n4719), .A(n4768), .ZN(n4721) );
  OAI21_X1 U5225 ( .B1(n2402), .B2(n4722), .A(n4721), .ZN(n4766) );
  AOI21_X1 U5226 ( .B1(n4767), .B2(n4723), .A(n4766), .ZN(n4728) );
  AOI22_X1 U5227 ( .A1(n4725), .A2(n4768), .B1(REG3_REG_0__SCAN_IN), .B2(n4724), .ZN(n4726) );
  OAI221_X1 U5228 ( .B1(n4706), .B2(n4728), .C1(n4534), .C2(n4727), .A(n4726), 
        .ZN(U3290) );
  AND2_X1 U5229 ( .A1(D_REG_31__SCAN_IN), .A2(n4739), .ZN(U3291) );
  AND2_X1 U5230 ( .A1(D_REG_30__SCAN_IN), .A2(n4739), .ZN(U3292) );
  NOR2_X1 U5231 ( .A1(n4741), .A2(n4729), .ZN(U3293) );
  AND2_X1 U5232 ( .A1(D_REG_28__SCAN_IN), .A2(n4739), .ZN(U3294) );
  AND2_X1 U5233 ( .A1(D_REG_27__SCAN_IN), .A2(n4739), .ZN(U3295) );
  NOR2_X1 U5234 ( .A1(n4741), .A2(n4730), .ZN(U3296) );
  AND2_X1 U5235 ( .A1(D_REG_25__SCAN_IN), .A2(n4739), .ZN(U3297) );
  AND2_X1 U5236 ( .A1(D_REG_24__SCAN_IN), .A2(n4739), .ZN(U3298) );
  AND2_X1 U5237 ( .A1(D_REG_23__SCAN_IN), .A2(n4739), .ZN(U3299) );
  AND2_X1 U5238 ( .A1(D_REG_22__SCAN_IN), .A2(n4739), .ZN(U3300) );
  AND2_X1 U5239 ( .A1(D_REG_21__SCAN_IN), .A2(n4739), .ZN(U3301) );
  NOR2_X1 U5240 ( .A1(n4741), .A2(n4731), .ZN(U3302) );
  AND2_X1 U5241 ( .A1(D_REG_19__SCAN_IN), .A2(n4739), .ZN(U3303) );
  NOR2_X1 U5242 ( .A1(n4741), .A2(n4732), .ZN(U3304) );
  AND2_X1 U5243 ( .A1(D_REG_17__SCAN_IN), .A2(n4739), .ZN(U3305) );
  AND2_X1 U5244 ( .A1(D_REG_16__SCAN_IN), .A2(n4739), .ZN(U3306) );
  NOR2_X1 U5245 ( .A1(n4741), .A2(n4733), .ZN(U3307) );
  NOR2_X1 U5246 ( .A1(n4741), .A2(n4734), .ZN(U3308) );
  AND2_X1 U5247 ( .A1(D_REG_13__SCAN_IN), .A2(n4739), .ZN(U3309) );
  AND2_X1 U5248 ( .A1(D_REG_12__SCAN_IN), .A2(n4739), .ZN(U3310) );
  NOR2_X1 U5249 ( .A1(n4741), .A2(n4735), .ZN(U3311) );
  AND2_X1 U5250 ( .A1(D_REG_10__SCAN_IN), .A2(n4739), .ZN(U3312) );
  NOR2_X1 U5251 ( .A1(n4741), .A2(n4736), .ZN(U3313) );
  AND2_X1 U5252 ( .A1(D_REG_8__SCAN_IN), .A2(n4739), .ZN(U3314) );
  AND2_X1 U5253 ( .A1(D_REG_7__SCAN_IN), .A2(n4739), .ZN(U3315) );
  NOR2_X1 U5254 ( .A1(n4741), .A2(n4737), .ZN(U3316) );
  AND2_X1 U5255 ( .A1(D_REG_5__SCAN_IN), .A2(n4739), .ZN(U3317) );
  NOR2_X1 U5256 ( .A1(n4741), .A2(n4738), .ZN(U3318) );
  AND2_X1 U5257 ( .A1(D_REG_3__SCAN_IN), .A2(n4739), .ZN(U3319) );
  NOR2_X1 U5258 ( .A1(n4741), .A2(n4740), .ZN(U3320) );
  AOI21_X1 U5259 ( .B1(U3149), .B2(n4743), .A(n4742), .ZN(U3329) );
  AOI22_X1 U5260 ( .A1(STATE_REG_SCAN_IN), .A2(n4744), .B1(n2600), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5261 ( .A1(STATE_REG_SCAN_IN), .A2(n4746), .B1(n4745), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5262 ( .A1(STATE_REG_SCAN_IN), .A2(n4748), .B1(n4747), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5263 ( .A1(STATE_REG_SCAN_IN), .A2(n4749), .B1(n2557), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5264 ( .A1(STATE_REG_SCAN_IN), .A2(n4751), .B1(n4750), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5265 ( .A1(U3149), .A2(n4752), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4753) );
  INV_X1 U5266 ( .A(n4753), .ZN(U3340) );
  AOI22_X1 U5267 ( .A1(STATE_REG_SCAN_IN), .A2(n4755), .B1(n4754), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5268 ( .A(DATAI_8_), .ZN(n4756) );
  AOI22_X1 U5269 ( .A1(STATE_REG_SCAN_IN), .A2(n4757), .B1(n4756), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U5270 ( .A1(U3149), .A2(n4758), .B1(DATAI_7_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4759) );
  INV_X1 U5271 ( .A(n4759), .ZN(U3345) );
  OAI22_X1 U5272 ( .A1(U3149), .A2(n4760), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4761) );
  INV_X1 U5273 ( .A(n4761), .ZN(U3346) );
  INV_X1 U5274 ( .A(DATAI_5_), .ZN(n4762) );
  AOI22_X1 U5275 ( .A1(STATE_REG_SCAN_IN), .A2(n4763), .B1(n4762), .B2(U3149), 
        .ZN(U3347) );
  AOI22_X1 U5276 ( .A1(STATE_REG_SCAN_IN), .A2(n4765), .B1(n4764), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5277 ( .C1(n4820), .C2(n4768), .A(n4767), .B(n4766), .ZN(n4825)
         );
  AOI22_X1 U5278 ( .A1(n4824), .A2(n4825), .B1(n4769), .B2(n4822), .ZN(U3467)
         );
  INV_X1 U5279 ( .A(n4770), .ZN(n4774) );
  OAI22_X1 U5280 ( .A1(n4772), .A2(n4783), .B1(n2823), .B2(n4771), .ZN(n4773)
         );
  NOR2_X1 U5281 ( .A1(n4774), .A2(n4773), .ZN(n4826) );
  AOI22_X1 U5282 ( .A1(n4824), .A2(n4826), .B1(n4775), .B2(n4822), .ZN(U3469)
         );
  NOR2_X1 U5283 ( .A1(n4776), .A2(n2823), .ZN(n4778) );
  AOI22_X1 U5284 ( .A1(n4779), .A2(n4820), .B1(n4778), .B2(n4777), .ZN(n4780)
         );
  AND2_X1 U5285 ( .A1(n4781), .A2(n4780), .ZN(n4827) );
  INV_X1 U5286 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5287 ( .A1(n4824), .A2(n4827), .B1(n4782), .B2(n4822), .ZN(U3471)
         );
  NOR2_X1 U5288 ( .A1(n4784), .A2(n4783), .ZN(n4786) );
  AOI211_X1 U5289 ( .C1(n4812), .C2(n4787), .A(n4786), .B(n4785), .ZN(n4828)
         );
  INV_X1 U5290 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5291 ( .A1(n4824), .A2(n4828), .B1(n4788), .B2(n4822), .ZN(U3473)
         );
  INV_X1 U5292 ( .A(n4789), .ZN(n4791) );
  AOI211_X1 U5293 ( .C1(n4792), .C2(n4820), .A(n4791), .B(n4790), .ZN(n4829)
         );
  AOI22_X1 U5294 ( .A1(n4824), .A2(n4829), .B1(n4793), .B2(n4822), .ZN(U3475)
         );
  OAI21_X1 U5295 ( .B1(n2823), .B2(n4795), .A(n4794), .ZN(n4796) );
  AOI21_X1 U5296 ( .B1(n4797), .B2(n4809), .A(n4796), .ZN(n4830) );
  INV_X1 U5297 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5298 ( .A1(n4824), .A2(n4830), .B1(n4798), .B2(n4822), .ZN(U3477)
         );
  OAI211_X1 U5299 ( .C1(n4802), .C2(n4801), .A(n4800), .B(n4799), .ZN(n4803)
         );
  INV_X1 U5300 ( .A(n4803), .ZN(n4831) );
  INV_X1 U5301 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4804) );
  AOI22_X1 U5302 ( .A1(n4824), .A2(n4831), .B1(n4804), .B2(n4822), .ZN(U3481)
         );
  OAI21_X1 U5303 ( .B1(n2823), .B2(n4806), .A(n4805), .ZN(n4807) );
  AOI21_X1 U5304 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4832) );
  AOI22_X1 U5305 ( .A1(n4824), .A2(n4832), .B1(n4810), .B2(n4822), .ZN(U3485)
         );
  AOI22_X1 U5306 ( .A1(n4813), .A2(n4820), .B1(n4812), .B2(n4811), .ZN(n4814)
         );
  AND2_X1 U5307 ( .A1(n4815), .A2(n4814), .ZN(n4833) );
  INV_X1 U5308 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4816) );
  AOI22_X1 U5309 ( .A1(n4824), .A2(n4833), .B1(n4816), .B2(n4822), .ZN(U3489)
         );
  NOR2_X1 U5310 ( .A1(n4817), .A2(n2823), .ZN(n4819) );
  AOI211_X1 U5311 ( .C1(n4821), .C2(n4820), .A(n4819), .B(n4818), .ZN(n4835)
         );
  AOI22_X1 U5312 ( .A1(n4824), .A2(n4835), .B1(n4823), .B2(n4822), .ZN(U3493)
         );
  AOI22_X1 U5313 ( .A1(n4836), .A2(n4825), .B1(n2820), .B2(n4834), .ZN(U3518)
         );
  AOI22_X1 U5314 ( .A1(n4836), .A2(n4826), .B1(n2386), .B2(n4834), .ZN(U3519)
         );
  AOI22_X1 U5315 ( .A1(n4836), .A2(n4827), .B1(n2412), .B2(n4834), .ZN(U3520)
         );
  AOI22_X1 U5316 ( .A1(n4836), .A2(n4828), .B1(n2423), .B2(n4834), .ZN(U3521)
         );
  AOI22_X1 U5317 ( .A1(n4836), .A2(n4829), .B1(n2244), .B2(n4834), .ZN(U3522)
         );
  AOI22_X1 U5318 ( .A1(n4836), .A2(n4830), .B1(n2448), .B2(n4834), .ZN(U3523)
         );
  AOI22_X1 U5319 ( .A1(n4836), .A2(n4831), .B1(n2467), .B2(n4834), .ZN(U3525)
         );
  AOI22_X1 U5320 ( .A1(n4836), .A2(n4832), .B1(n3018), .B2(n4834), .ZN(U3527)
         );
  AOI22_X1 U5321 ( .A1(n4836), .A2(n4833), .B1(n3244), .B2(n4834), .ZN(U3529)
         );
  AOI22_X1 U5322 ( .A1(n4836), .A2(n4835), .B1(n2537), .B2(n4834), .ZN(U3531)
         );
  INV_X2 U2376 ( .A(n3520), .ZN(n2925) );
  CLKBUF_X1 U3412 ( .A(n2692), .Z(n2693) );
endmodule

