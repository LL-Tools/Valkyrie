

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481;

  CLKBUF_X1 U3393 ( .A(n4221), .Z(n2945) );
  CLKBUF_X1 U3394 ( .A(n3838), .Z(n2978) );
  CLKBUF_X2 U3395 ( .A(n3145), .Z(n3774) );
  CLKBUF_X2 U3396 ( .A(n3150), .Z(n3806) );
  CLKBUF_X1 U3397 ( .A(n3203), .Z(n4030) );
  CLKBUF_X2 U3398 ( .A(n3158), .Z(n3804) );
  CLKBUF_X2 U3399 ( .A(n3137), .Z(n3796) );
  CLKBUF_X2 U3400 ( .A(n3152), .Z(n4339) );
  INV_X1 U3402 ( .A(n3296), .ZN(n3320) );
  AND2_X1 U3403 ( .A1(n4348), .A2(n3045), .ZN(n3221) );
  AND2_X1 U3404 ( .A1(n4344), .A2(n3002), .ZN(n3207) );
  CLKBUF_X2 U3405 ( .A(n3139), .Z(n3775) );
  CLKBUF_X2 U3406 ( .A(n2973), .Z(n3807) );
  AOI22_X1 U3407 ( .A1(n6392), .A2(keyinput36), .B1(keyinput20), .B2(n4794), 
        .ZN(n6391) );
  AOI22_X1 U3408 ( .A1(n6339), .A2(keyinput31), .B1(keyinput38), .B2(n6338), 
        .ZN(n6337) );
  NAND2_X1 U3409 ( .A1(n3201), .A2(n2980), .ZN(n4221) );
  NAND2_X1 U3410 ( .A1(n3267), .A2(n3266), .ZN(n3349) );
  OAI221_X1 U3411 ( .B1(n6392), .B2(keyinput36), .C1(n4794), .C2(keyinput20), 
        .A(n6391), .ZN(n6405) );
  OAI221_X1 U3412 ( .B1(n6339), .B2(keyinput31), .C1(n6338), .C2(keyinput38), 
        .A(n6337), .ZN(n6340) );
  NOR2_X1 U3413 ( .A1(n3302), .A2(n5766), .ZN(n3303) );
  INV_X1 U3414 ( .A(n3821), .ZN(n3763) );
  AND2_X2 U3415 ( .A1(n3037), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3044)
         );
  XNOR2_X1 U3416 ( .A(n3349), .B(n3295), .ZN(n4451) );
  INV_X1 U3417 ( .A(n4605), .ZN(n5295) );
  XOR2_X1 U3418 ( .A(n4144), .B(n4226), .Z(n2983) );
  AND2_X2 U3419 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4340) );
  INV_X1 U3420 ( .A(n3201), .ZN(n5619) );
  AND2_X1 U3421 ( .A1(n4605), .A2(n4604), .ZN(n5374) );
  AND2_X1 U3422 ( .A1(n2968), .A2(n2969), .ZN(n4542) );
  OR2_X1 U3423 ( .A1(n4385), .A2(n4297), .ZN(n6319) );
  AOI22_X1 U3424 ( .A1(n4990), .A2(n5369), .B1(REIP_REG_30__SCAN_IN), .B2(
        n4989), .ZN(n4991) );
  INV_X1 U3425 ( .A(n5374), .ZN(n5359) );
  INV_X2 U3427 ( .A(n3185), .ZN(n3216) );
  AND4_X2 U3428 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n3060)
         );
  AND2_X4 U3429 ( .A1(n3044), .A2(n4357), .ZN(n3160) );
  AND2_X4 U3430 ( .A1(n4338), .A2(n3042), .ZN(n3159) );
  AND2_X4 U3431 ( .A1(n3042), .A2(n4434), .ZN(n3150) );
  NAND2_X2 U3432 ( .A1(n4864), .A2(n4254), .ZN(n4878) );
  OAI22_X2 U3433 ( .A1(n3939), .A2(n3970), .B1(n3938), .B2(n6309), .ZN(n3940)
         );
  NAND2_X2 U3434 ( .A1(n3882), .A2(n3881), .ZN(n6157) );
  NOR2_X1 U3435 ( .A1(n4381), .A2(n4456), .ZN(n4405) );
  NAND2_X1 U3436 ( .A1(n3009), .A2(n3008), .ZN(n4381) );
  AND2_X1 U3437 ( .A1(n4382), .A2(n3007), .ZN(n3008) );
  AND2_X1 U3438 ( .A1(n2954), .A2(n3084), .ZN(n3886) );
  CLKBUF_X2 U3439 ( .A(n3887), .Z(n2977) );
  BUF_X2 U3441 ( .A(n4140), .Z(n2946) );
  CLKBUF_X2 U3442 ( .A(n3144), .Z(n3795) );
  CLKBUF_X2 U3443 ( .A(n3138), .Z(n3358) );
  INV_X1 U3444 ( .A(n3011), .ZN(n3222) );
  CLKBUF_X2 U34450 ( .A(n3161), .Z(n3805) );
  NAND2_X1 U34460 ( .A1(n4259), .A2(n4258), .ZN(n4261) );
  AOI21_X1 U34470 ( .B1(n4018), .B2(n4858), .A(n4017), .ZN(n4019) );
  AOI21_X1 U34480 ( .B1(n4878), .B2(n4877), .A(n4256), .ZN(n5127) );
  INV_X1 U3449 ( .A(n4000), .ZN(n3999) );
  NAND2_X1 U3450 ( .A1(n3016), .A2(n3020), .ZN(n4000) );
  AOI211_X1 U34510 ( .C1(EBX_REG_27__SCAN_IN), .C2(n5353), .A(n5016), .B(n5015), .ZN(n5017) );
  AOI211_X1 U34520 ( .C1(n5082), .C2(n5328), .A(n4997), .B(n4996), .ZN(n4999)
         );
  NAND2_X1 U34530 ( .A1(n4020), .A2(n4803), .ZN(n5086) );
  NAND2_X1 U3454 ( .A1(n4021), .A2(n4287), .ZN(n4289) );
  OR2_X1 U34550 ( .A1(n4021), .A2(n4287), .ZN(n4288) );
  CLKBUF_X1 U34560 ( .A(n4745), .Z(n4804) );
  NOR2_X2 U3457 ( .A1(n4727), .A2(n4832), .ZN(n4737) );
  AND2_X1 U3458 ( .A1(n4652), .A2(n3004), .ZN(n4726) );
  NAND2_X1 U34590 ( .A1(n4225), .A2(n2984), .ZN(n4144) );
  NAND2_X1 U34600 ( .A1(n3001), .A2(n3000), .ZN(n4773) );
  NOR2_X1 U34610 ( .A1(n4543), .A2(n4596), .ZN(n2965) );
  NOR2_X1 U34620 ( .A1(n4406), .A2(n4516), .ZN(n4515) );
  NOR2_X1 U34630 ( .A1(n4406), .A2(n4516), .ZN(n2968) );
  AOI21_X1 U34640 ( .B1(n5120), .B2(n3021), .A(n2991), .ZN(n3020) );
  AOI21_X1 U34650 ( .B1(n3398), .B2(n3531), .A(n3397), .ZN(n4456) );
  OAI21_X1 U3466 ( .B1(n3417), .B2(n3421), .A(n3416), .ZN(n4407) );
  OAI21_X1 U3467 ( .B1(n3965), .B2(n3970), .A(n3964), .ZN(n3966) );
  OAI21_X1 U34680 ( .B1(n3948), .B2(n3970), .A(n3947), .ZN(n3950) );
  CLKBUF_X1 U34690 ( .A(n3907), .Z(n5407) );
  OAI21_X1 U34700 ( .B1(n4379), .B2(n3329), .A(n4380), .ZN(n4372) );
  XNOR2_X1 U34710 ( .A(n3934), .B(n6463), .ZN(n4398) );
  NAND2_X1 U34720 ( .A1(n3006), .A2(n2990), .ZN(n3969) );
  NOR2_X2 U34730 ( .A1(n5766), .A2(n5295), .ZN(n4608) );
  NOR2_X1 U34740 ( .A1(n4713), .A2(n4714), .ZN(n4691) );
  NAND2_X1 U3475 ( .A1(n3370), .A2(n3369), .ZN(n3393) );
  NAND2_X2 U3476 ( .A1(n4215), .A2(n4214), .ZN(n4605) );
  CLKBUF_X1 U3477 ( .A(n4447), .Z(n5926) );
  CLKBUF_X1 U3478 ( .A(n4341), .Z(n6029) );
  NOR2_X1 U3479 ( .A1(n4506), .A2(n4469), .ZN(n4565) );
  OR2_X1 U3480 ( .A1(n2961), .A2(n2962), .ZN(n4506) );
  INV_X1 U3481 ( .A(n5921), .ZN(n6288) );
  INV_X1 U3482 ( .A(n2998), .ZN(n4682) );
  NAND2_X1 U3483 ( .A1(n3335), .A2(n3334), .ZN(n5966) );
  NOR2_X1 U3484 ( .A1(n4754), .A2(n4741), .ZN(n4115) );
  AND2_X1 U3485 ( .A1(n3116), .A2(n3003), .ZN(n3827) );
  OR2_X1 U3486 ( .A1(n4057), .A2(EBX_REG_1__SCAN_IN), .ZN(n2999) );
  NOR2_X1 U3487 ( .A1(n3917), .A2(n3971), .ZN(n3259) );
  AOI21_X1 U3488 ( .B1(n4244), .B2(n4030), .A(n6273), .ZN(n3206) );
  OR2_X1 U3489 ( .A1(n3890), .A2(n3258), .ZN(n3971) );
  AND2_X1 U3490 ( .A1(n3913), .A2(n3083), .ZN(n2954) );
  INV_X2 U3491 ( .A(n4221), .ZN(n4052) );
  CLKBUF_X2 U3492 ( .A(n3202), .Z(n4244) );
  OR2_X1 U3493 ( .A1(n3228), .A2(n3227), .ZN(n3912) );
  OR2_X1 U3494 ( .A1(n3257), .A2(n3256), .ZN(n3917) );
  NAND4_X1 U3495 ( .A1(n3320), .A2(n3889), .A3(n3302), .A4(n4046), .ZN(n4029)
         );
  BUF_X2 U3496 ( .A(n3114), .Z(n3839) );
  INV_X1 U3497 ( .A(n3889), .ZN(n4492) );
  NAND2_X1 U3498 ( .A1(n3190), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3336) );
  INV_X4 U3499 ( .A(n3190), .ZN(n3843) );
  AND2_X1 U3500 ( .A1(n3157), .A2(n3156), .ZN(n3167) );
  AND4_X2 U3501 ( .A1(n3135), .A2(n3136), .A3(n3133), .A4(n3134), .ZN(n3190)
         );
  OR2_X2 U3502 ( .A1(n3081), .A2(n3080), .ZN(n3302) );
  NAND2_X1 U3503 ( .A1(n3051), .A2(n3050), .ZN(n3185) );
  AND4_X2 U3504 ( .A1(n3113), .A2(n2982), .A3(n3112), .A4(n3111), .ZN(n3889)
         );
  AND4_X1 U3505 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3168)
         );
  AND3_X1 U3506 ( .A1(n3155), .A2(n3154), .A3(n3153), .ZN(n3157) );
  AND4_X1 U3507 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3166)
         );
  AND4_X1 U3508 ( .A1(n3041), .A2(n3040), .A3(n3039), .A4(n3038), .ZN(n3051)
         );
  AND4_X1 U3509 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3112)
         );
  AND4_X1 U3510 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3113)
         );
  AND4_X1 U3511 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3111)
         );
  AND4_X1 U3512 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n3061)
         );
  AND4_X1 U3513 ( .A1(n3069), .A2(n3068), .A3(n3067), .A4(n3066), .ZN(n3070)
         );
  AND4_X1 U3514 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(n3135)
         );
  AND4_X1 U3515 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n3136)
         );
  AND4_X1 U3516 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3071)
         );
  AND4_X1 U3517 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3133)
         );
  AND4_X1 U3518 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3134)
         );
  AND4_X1 U3519 ( .A1(n3049), .A2(n3048), .A3(n3047), .A4(n3046), .ZN(n3050)
         );
  AND4_X1 U3520 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n3169)
         );
  BUF_X2 U3521 ( .A(n3160), .Z(n3797) );
  BUF_X2 U3522 ( .A(n3159), .Z(n3798) );
  BUF_X2 U3523 ( .A(n3231), .Z(n3247) );
  AND2_X2 U3525 ( .A1(n4361), .A2(n4434), .ZN(n3279) );
  AND2_X2 U3526 ( .A1(n4357), .A2(n4338), .ZN(n3138) );
  AND2_X2 U3527 ( .A1(n4357), .A2(n3043), .ZN(n3161) );
  AND2_X2 U3528 ( .A1(n3036), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4338)
         );
  AND2_X2 U3529 ( .A1(n4357), .A2(n4434), .ZN(n3139) );
  AND2_X2 U3530 ( .A1(n4340), .A2(n3043), .ZN(n3145) );
  INV_X2 U3531 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5766) );
  AND2_X2 U3532 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4434) );
  NOR2_X2 U3533 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3043) );
  AND2_X1 U3534 ( .A1(n4729), .A2(n3004), .ZN(n2947) );
  AND2_X1 U3535 ( .A1(n4289), .A2(n4288), .ZN(n5082) );
  NAND2_X1 U3536 ( .A1(n4542), .A2(n4545), .ZN(n4543) );
  NAND2_X1 U3537 ( .A1(n4636), .A2(n2951), .ZN(n2948) );
  AND2_X2 U3538 ( .A1(n2948), .A2(n2949), .ZN(n4707) );
  OR2_X1 U3539 ( .A1(n2950), .A2(n3024), .ZN(n2949) );
  INV_X1 U3540 ( .A(n3986), .ZN(n2950) );
  AND2_X1 U3541 ( .A1(n3026), .A2(n3986), .ZN(n2951) );
  NAND2_X1 U3542 ( .A1(n3983), .A2(n5478), .ZN(n2952) );
  NAND2_X1 U3543 ( .A1(n3983), .A2(n5478), .ZN(n5469) );
  NOR2_X1 U3544 ( .A1(n4543), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U3545 ( .A1(n3979), .A2(n3978), .ZN(n2953) );
  NAND2_X1 U3546 ( .A1(n3979), .A2(n3978), .ZN(n4560) );
  AND2_X1 U3547 ( .A1(n3084), .A2(n3083), .ZN(n4154) );
  CLKBUF_X1 U3548 ( .A(n4574), .Z(n2955) );
  NAND2_X1 U3549 ( .A1(n3936), .A2(n3935), .ZN(n4458) );
  NAND2_X1 U3550 ( .A1(n3968), .A2(n3967), .ZN(n4574) );
  AND2_X2 U3551 ( .A1(n4361), .A2(n3044), .ZN(n3144) );
  AND2_X2 U3552 ( .A1(n3044), .A2(n4340), .ZN(n3152) );
  NAND2_X1 U3553 ( .A1(n4753), .A2(n4831), .ZN(n2956) );
  OR2_X1 U3555 ( .A1(n4115), .A2(n4114), .ZN(n2957) );
  NAND2_X1 U3556 ( .A1(n4649), .A2(n4650), .ZN(n2958) );
  OR2_X2 U3557 ( .A1(n2958), .A2(n2959), .ZN(n5191) );
  OR2_X1 U3558 ( .A1(n2960), .A2(n4714), .ZN(n2959) );
  INV_X1 U3559 ( .A(n4692), .ZN(n2960) );
  NAND2_X1 U3560 ( .A1(n4758), .A2(n4759), .ZN(n2961) );
  OR2_X1 U3561 ( .A1(n2963), .A2(n4554), .ZN(n2962) );
  INV_X1 U3562 ( .A(n4505), .ZN(n2963) );
  NAND2_X1 U3563 ( .A1(n5469), .A2(n5470), .ZN(n3984) );
  OR2_X1 U3564 ( .A1(n5135), .A2(n2992), .ZN(n3016) );
  OAI21_X1 U3565 ( .B1(n3920), .B2(n3970), .A(n3919), .ZN(n5526) );
  OR2_X1 U3566 ( .A1(n5511), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3927)
         );
  NAND2_X2 U3567 ( .A1(n3319), .A2(n3318), .ZN(n3920) );
  NAND2_X4 U3568 ( .A1(n3969), .A2(n3972), .ZN(n3980) );
  NAND2_X2 U3569 ( .A1(n5127), .A2(n5126), .ZN(n5125) );
  XNOR2_X1 U3570 ( .A(n3977), .B(n4078), .ZN(n4575) );
  NAND2_X2 U3571 ( .A1(n3984), .A2(n5471), .ZN(n4636) );
  NAND2_X2 U3572 ( .A1(n3372), .A2(n3352), .ZN(n3933) );
  NOR2_X2 U3573 ( .A1(n4823), .A2(n4822), .ZN(n4816) );
  NOR2_X2 U3574 ( .A1(n4666), .A2(n4667), .ZN(n4649) );
  NOR2_X1 U3575 ( .A1(n4381), .A2(n4456), .ZN(n2964) );
  AND2_X2 U3576 ( .A1(n2965), .A2(n2966), .ZN(n4622) );
  AND2_X1 U3577 ( .A1(n2967), .A2(n4600), .ZN(n2966) );
  INV_X1 U3578 ( .A(n4623), .ZN(n2967) );
  AND2_X1 U3579 ( .A1(n2970), .A2(n4518), .ZN(n2969) );
  INV_X1 U3580 ( .A(n4547), .ZN(n2970) );
  NOR2_X1 U3581 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3045) );
  AND2_X1 U3582 ( .A1(n3044), .A2(n4357), .ZN(n2971) );
  AND2_X1 U3583 ( .A1(n4434), .A2(n4340), .ZN(n2972) );
  AND2_X1 U3584 ( .A1(n4434), .A2(n4340), .ZN(n2973) );
  AND2_X1 U3585 ( .A1(n3044), .A2(n4340), .ZN(n2974) );
  AND2_X1 U3586 ( .A1(n3044), .A2(n4340), .ZN(n2975) );
  AND2_X1 U3587 ( .A1(n4340), .A2(n3043), .ZN(n2976) );
  AND2_X1 U3588 ( .A1(n2979), .A2(n3179), .ZN(n3838) );
  NAND2_X1 U3589 ( .A1(n3297), .A2(n3689), .ZN(n4379) );
  NOR2_X1 U3590 ( .A1(n4553), .A2(n4554), .ZN(n4555) );
  AND2_X2 U3591 ( .A1(n4745), .A2(n4748), .ZN(n4746) );
  NOR2_X2 U3592 ( .A1(n4263), .A2(n4805), .ZN(n4745) );
  NAND2_X1 U3593 ( .A1(n5619), .A2(n3843), .ZN(n4140) );
  OAI211_X2 U3594 ( .C1(n3939), .C2(n3421), .A(n3380), .B(n3379), .ZN(n4382)
         );
  NAND4_X1 U3595 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n2979)
         );
  NAND4_X1 U3596 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n2980)
         );
  AND2_X2 U3597 ( .A1(n4819), .A2(n3010), .ZN(n4262) );
  NOR2_X2 U3598 ( .A1(n4826), .A2(n4825), .ZN(n4819) );
  NOR2_X4 U3599 ( .A1(n4625), .A2(n4653), .ZN(n4652) );
  OR2_X1 U3600 ( .A1(n4029), .A2(n6180), .ZN(n3823) );
  INV_X1 U3601 ( .A(n3823), .ZN(n2981) );
  NAND2_X1 U3602 ( .A1(n3843), .A2(n3035), .ZN(n3242) );
  AND2_X1 U3603 ( .A1(n4046), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3035) );
  XNOR2_X1 U3604 ( .A(n3301), .B(n3300), .ZN(n4447) );
  NAND2_X2 U3605 ( .A1(n3216), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3890) );
  OR2_X1 U3606 ( .A1(n4326), .A2(n4165), .ZN(n4347) );
  AND2_X1 U3607 ( .A1(n6157), .A2(n6181), .ZN(n4298) );
  NAND2_X1 U3608 ( .A1(n3031), .A2(n4658), .ZN(n3030) );
  NAND2_X1 U3609 ( .A1(n4637), .A2(n4638), .ZN(n3031) );
  AND2_X1 U3610 ( .A1(n5530), .A2(n4009), .ZN(n5483) );
  AND2_X1 U3611 ( .A1(n3888), .A2(n3302), .ZN(n3084) );
  OR2_X1 U3612 ( .A1(n3346), .A2(n3345), .ZN(n3931) );
  NAND3_X1 U3613 ( .A1(n4003), .A2(n4151), .A3(n4492), .ZN(n3187) );
  NAND2_X1 U3614 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  XNOR2_X1 U3615 ( .A(n3969), .B(n3420), .ZN(n3965) );
  AND2_X1 U3616 ( .A1(n3115), .A2(n3843), .ZN(n3003) );
  INV_X1 U3617 ( .A(n4153), .ZN(n3913) );
  NAND2_X1 U3618 ( .A1(n3843), .A2(n3180), .ZN(n4058) );
  XNOR2_X1 U3619 ( .A(n4056), .B(n4550), .ZN(n4629) );
  AOI21_X1 U3620 ( .B1(n3197), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3194), 
        .ZN(n3195) );
  OR2_X1 U3621 ( .A1(n3890), .A2(n3245), .ZN(n3229) );
  NAND2_X2 U3622 ( .A1(n3890), .A2(n3336), .ZN(n3861) );
  NAND2_X1 U3623 ( .A1(n2997), .A2(n3889), .ZN(n4163) );
  NAND2_X1 U3624 ( .A1(n3246), .A2(n6180), .ZN(n3261) );
  INV_X1 U3625 ( .A(n5275), .ZN(n5346) );
  INV_X1 U3626 ( .A(n4771), .ZN(n3000) );
  OR2_X1 U3627 ( .A1(n4347), .A2(n6157), .ZN(n4335) );
  NOR2_X1 U3628 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6026), .ZN(n4207) );
  NAND2_X1 U3629 ( .A1(n5125), .A2(n3032), .ZN(n4873) );
  AOI21_X1 U3630 ( .B1(n3029), .B2(n3027), .A(n2988), .ZN(n3026) );
  INV_X1 U3631 ( .A(n4638), .ZN(n3027) );
  OR2_X1 U3632 ( .A1(n4636), .A2(n4637), .ZN(n3028) );
  INV_X1 U3633 ( .A(n3030), .ZN(n3029) );
  CLKBUF_X1 U3634 ( .A(n3827), .Z(n3828) );
  NAND2_X1 U3635 ( .A1(n4045), .A2(n4044), .ZN(n4173) );
  CLKBUF_X1 U3636 ( .A(n4418), .Z(n4419) );
  OR2_X1 U3637 ( .A1(n3933), .A2(n4452), .ZN(n5928) );
  AND2_X1 U3638 ( .A1(n4839), .A2(n4370), .ZN(n5397) );
  OR2_X1 U3639 ( .A1(n5533), .A2(n4006), .ZN(n5530) );
  AND2_X1 U3640 ( .A1(n6151), .A2(n4298), .ZN(n5533) );
  INV_X1 U3641 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6026) );
  CLKBUF_X1 U3642 ( .A(n4356), .Z(n5764) );
  NAND2_X1 U3643 ( .A1(n3839), .A2(n3843), .ZN(n3844) );
  NAND2_X1 U3644 ( .A1(n3006), .A2(n3391), .ZN(n3418) );
  INV_X1 U3645 ( .A(n3997), .ZN(n3021) );
  INV_X1 U3646 ( .A(n3392), .ZN(n3391) );
  INV_X1 U3647 ( .A(n3393), .ZN(n3006) );
  OR2_X1 U3648 ( .A1(n3408), .A2(n3407), .ZN(n3961) );
  OR2_X1 U3649 ( .A1(n3390), .A2(n3389), .ZN(n3945) );
  INV_X1 U3650 ( .A(n3880), .ZN(n3876) );
  AOI22_X1 U3651 ( .A1(n3159), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2974), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3652 ( .A1(n3144), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3653 ( .A1(n3158), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3654 ( .A1(n3144), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3089) );
  AOI22_X1 U3655 ( .A1(n3222), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3150), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3067) );
  NAND2_X1 U3656 ( .A1(n3239), .A2(n3034), .ZN(n3240) );
  AND2_X1 U3657 ( .A1(n3913), .A2(n3839), .ZN(n3115) );
  AND2_X1 U3658 ( .A1(n3612), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3628)
         );
  INV_X1 U3659 ( .A(n4207), .ZN(n3689) );
  INV_X1 U3660 ( .A(n4140), .ZN(n4125) );
  NAND2_X1 U3661 ( .A1(n3906), .A2(n3190), .ZN(n3885) );
  OR2_X1 U3662 ( .A1(n3290), .A2(n3289), .ZN(n3291) );
  NAND2_X1 U3663 ( .A1(n4150), .A2(n2993), .ZN(n4152) );
  AND2_X1 U3664 ( .A1(n3872), .A2(n2978), .ZN(n3880) );
  AND2_X1 U3665 ( .A1(n3836), .A2(n3835), .ZN(n3894) );
  OR2_X1 U3666 ( .A1(n3837), .A2(n3834), .ZN(n3836) );
  NAND2_X1 U3667 ( .A1(n3348), .A2(n3347), .ZN(n5706) );
  AOI21_X1 U3668 ( .B1(n3210), .B2(n3292), .A(n3191), .ZN(n3192) );
  AND2_X1 U3669 ( .A1(n3331), .A2(n6071), .ZN(n5828) );
  OAI21_X1 U3670 ( .B1(n6310), .B2(n6285), .A(n4785), .ZN(n4476) );
  INV_X1 U3671 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6145) );
  AND2_X1 U3672 ( .A1(n5619), .A2(n3190), .ZN(n3172) );
  NOR2_X1 U3673 ( .A1(n6230), .A2(n5241), .ZN(n5231) );
  INV_X1 U3674 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5258) );
  INV_X1 U3675 ( .A(n5368), .ZN(n5330) );
  AND2_X1 U3676 ( .A1(n3180), .A2(n3190), .ZN(n2997) );
  OAI21_X1 U3677 ( .B1(n4629), .B2(n4231), .A(n4056), .ZN(n2998) );
  INV_X1 U3678 ( .A(n6319), .ZN(n4215) );
  AND2_X1 U3679 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4608), .ZN(n4245) );
  NAND2_X1 U3680 ( .A1(n4649), .A2(n4650), .ZN(n4713) );
  AND2_X1 U3681 ( .A1(n4764), .A2(n4820), .ZN(n3010) );
  NOR2_X1 U3682 ( .A1(n2980), .A2(n3843), .ZN(n3887) );
  AND4_X1 U3683 ( .A1(n3893), .A2(n3892), .A3(n3303), .A4(n3891), .ZN(n4201)
         );
  AND2_X1 U3684 ( .A1(n3826), .A2(n5115), .ZN(n3723) );
  AND2_X1 U3685 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3692)
         );
  NAND2_X1 U3686 ( .A1(n3628), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3646)
         );
  NAND2_X1 U3687 ( .A1(n3581), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3611)
         );
  CLKBUF_X1 U3688 ( .A(n4727), .Z(n4728) );
  AND2_X1 U3689 ( .A1(n3551), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3552)
         );
  NAND2_X1 U3690 ( .A1(n3552), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3566)
         );
  NOR2_X1 U3691 ( .A1(n5147), .A2(n3005), .ZN(n3004) );
  INV_X1 U3692 ( .A(n4695), .ZN(n3005) );
  NOR2_X1 U3693 ( .A1(n3538), .A2(n4722), .ZN(n3551) );
  CLKBUF_X1 U3694 ( .A(n4625), .Z(n4626) );
  OR2_X1 U3695 ( .A1(n3483), .A2(n3479), .ZN(n3484) );
  NOR2_X1 U3696 ( .A1(n6392), .A2(n3484), .ZN(n3510) );
  INV_X1 U3697 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U3698 ( .A1(n3980), .A2(n4643), .ZN(n5470) );
  NAND2_X1 U3699 ( .A1(n3480), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3483)
         );
  NOR2_X1 U3700 ( .A1(n3455), .A2(n3454), .ZN(n3480) );
  CLKBUF_X1 U3701 ( .A(n4543), .Z(n4544) );
  NAND2_X1 U3702 ( .A1(n3451), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3455)
         );
  NAND2_X1 U3703 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  NOR2_X1 U3704 ( .A1(n3395), .A2(n5509), .ZN(n3412) );
  NAND2_X1 U3705 ( .A1(n3412), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3422)
         );
  NAND2_X1 U3706 ( .A1(n3378), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3395)
         );
  INV_X1 U3707 ( .A(n4374), .ZN(n3007) );
  INV_X1 U3708 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6453) );
  INV_X1 U3709 ( .A(n4773), .ZN(n4223) );
  NOR2_X1 U3710 ( .A1(n4269), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4270)
         );
  INV_X1 U3711 ( .A(n3001), .ZN(n4801) );
  AOI21_X1 U3712 ( .B1(n3998), .B2(n3997), .A(n3018), .ZN(n3017) );
  NAND2_X1 U3713 ( .A1(n5135), .A2(n3997), .ZN(n3019) );
  OR2_X1 U3714 ( .A1(n5135), .A2(n3998), .ZN(n3022) );
  NAND2_X1 U3715 ( .A1(n4811), .A2(n4812), .ZN(n4807) );
  NOR2_X2 U3716 ( .A1(n4807), .A2(n4806), .ZN(n4749) );
  NOR2_X1 U3717 ( .A1(n4255), .A2(n3980), .ZN(n4256) );
  NAND2_X1 U3718 ( .A1(n4753), .A2(n4831), .ZN(n4739) );
  OR2_X1 U3719 ( .A1(n3980), .A2(n4253), .ZN(n4254) );
  AOI21_X1 U3720 ( .B1(n3026), .B2(n3030), .A(n2986), .ZN(n3024) );
  AND2_X1 U3721 ( .A1(n3980), .A2(n4960), .ZN(n4708) );
  NAND2_X1 U3722 ( .A1(n4590), .A2(n4588), .ZN(n5284) );
  INV_X1 U3723 ( .A(n5580), .ZN(n4949) );
  NAND2_X1 U3724 ( .A1(n4447), .A2(n2978), .ZN(n3916) );
  INV_X1 U3725 ( .A(n5706), .ZN(n5797) );
  CLKBUF_X1 U3726 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4784) );
  AND2_X1 U3727 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U3728 ( .A1(n4336), .A2(n4335), .ZN(n6138) );
  AND2_X1 U3729 ( .A1(n5607), .A2(n4481), .ZN(n5643) );
  CLKBUF_X1 U3730 ( .A(n3179), .Z(n4477) );
  INV_X1 U3731 ( .A(n5629), .ZN(n4777) );
  OR2_X1 U3732 ( .A1(n5928), .A2(n5888), .ZN(n5889) );
  INV_X1 U3733 ( .A(n5736), .ZN(n6082) );
  NAND2_X1 U3734 ( .A1(n6180), .A2(n4476), .ZN(n5630) );
  AND2_X1 U3735 ( .A1(n6395), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3883) );
  INV_X1 U3736 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6209) );
  INV_X1 U3737 ( .A(n4266), .ZN(n5036) );
  NOR2_X1 U3738 ( .A1(n5075), .A2(n5224), .ZN(n5068) );
  NAND2_X1 U3739 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5231), .ZN(n5224) );
  NAND2_X1 U3740 ( .A1(n4235), .A2(n4234), .ZN(n5275) );
  AND2_X1 U3741 ( .A1(n4608), .A2(n2997), .ZN(n5351) );
  AND2_X1 U3742 ( .A1(n4609), .A2(n4608), .ZN(n5353) );
  NAND2_X1 U3743 ( .A1(n3843), .A2(n2994), .ZN(n4606) );
  INV_X1 U3744 ( .A(n5369), .ZN(n5367) );
  INV_X1 U3745 ( .A(n5343), .ZN(n5375) );
  NOR2_X2 U3746 ( .A1(n4231), .A2(n4230), .ZN(n5369) );
  NAND2_X1 U3747 ( .A1(n6168), .A2(n4245), .ZN(n4230) );
  INV_X1 U3748 ( .A(n4838), .ZN(n5392) );
  NAND2_X1 U3749 ( .A1(n4833), .A2(n4840), .ZN(n4838) );
  AND2_X1 U3750 ( .A1(n4839), .A2(n4371), .ZN(n4654) );
  INV_X1 U3751 ( .A(n5397), .ZN(n5403) );
  INV_X1 U3752 ( .A(n4654), .ZN(n4457) );
  AND3_X1 U3753 ( .A1(n4299), .A2(n4329), .A3(n4298), .ZN(n5426) );
  CLKBUF_X1 U3754 ( .A(n6307), .Z(n6170) );
  INV_X2 U3755 ( .A(n5436), .ZN(n5437) );
  INV_X1 U3756 ( .A(n5426), .ZN(n5439) );
  INV_X1 U3757 ( .A(n6440), .ZN(n5459) );
  INV_X1 U3758 ( .A(n4522), .ZN(n6438) );
  INV_X1 U3759 ( .A(n4403), .ZN(n6437) );
  XNOR2_X1 U3760 ( .A(n4218), .B(n4217), .ZN(n4854) );
  OR2_X1 U3761 ( .A1(n4216), .A2(n4011), .ZN(n4218) );
  INV_X1 U3762 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5509) );
  INV_X1 U3763 ( .A(n5533), .ZN(n5503) );
  OR2_X1 U3764 ( .A1(n5182), .A2(n4190), .ZN(n5161) );
  AND2_X1 U3765 ( .A1(n4935), .A2(n4189), .ZN(n5168) );
  XNOR2_X1 U3766 ( .A(n4261), .B(n4260), .ZN(n4926) );
  OR2_X1 U3767 ( .A1(n4636), .A2(n3030), .ZN(n3023) );
  NAND2_X1 U3768 ( .A1(n3025), .A2(n3029), .ZN(n4657) );
  NAND2_X1 U3769 ( .A1(n3028), .A2(n4638), .ZN(n4659) );
  NAND2_X1 U3770 ( .A1(n4636), .A2(n4638), .ZN(n3025) );
  CLKBUF_X1 U3771 ( .A(n4464), .Z(n4465) );
  CLKBUF_X1 U3772 ( .A(n4968), .Z(n4969) );
  INV_X1 U3773 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6293) );
  CLKBUF_X1 U3774 ( .A(n4451), .Z(n4452) );
  INV_X1 U3775 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6284) );
  INV_X1 U3776 ( .A(n6029), .ZN(n6279) );
  INV_X1 U3777 ( .A(n6289), .ZN(n6275) );
  INV_X1 U3778 ( .A(n6291), .ZN(n6294) );
  INV_X1 U3779 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6445) );
  AND2_X2 U3780 ( .A1(n4363), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4361)
         );
  NAND2_X1 U3781 ( .A1(n6157), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4785) );
  INV_X1 U3782 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5200) );
  INV_X1 U3783 ( .A(n4792), .ZN(n6269) );
  OAI21_X1 U3784 ( .B1(n5691), .B2(n5675), .A(n5895), .ZN(n5692) );
  INV_X1 U3785 ( .A(n5734), .ZN(n5726) );
  OAI21_X1 U3786 ( .B1(n5730), .B2(n6034), .A(n5713), .ZN(n5731) );
  INV_X1 U3787 ( .A(n5763), .ZN(n5748) );
  INV_X1 U3788 ( .A(n5889), .ZN(n5954) );
  OR4_X1 U3789 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n5988) );
  OR2_X1 U3790 ( .A1(n5999), .A2(n6290), .ZN(n6020) );
  INV_X1 U3791 ( .A(n5601), .ZN(n6075) );
  INV_X1 U3792 ( .A(n5613), .ZN(n6088) );
  INV_X1 U3793 ( .A(n5616), .ZN(n6094) );
  INV_X1 U3794 ( .A(n5626), .ZN(n6112) );
  INV_X1 U3795 ( .A(n5634), .ZN(n6126) );
  AND2_X1 U3796 ( .A1(n3883), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6181) );
  AOI21_X1 U3797 ( .B1(DATAI_30_), .B2(n5396), .A(n3909), .ZN(n3910) );
  INV_X1 U3798 ( .A(n4012), .ZN(n3014) );
  NAND2_X1 U3799 ( .A1(n4200), .A2(n5631), .ZN(n3015) );
  AOI21_X1 U3800 ( .B1(n4023), .B2(n5631), .A(n4026), .ZN(n4027) );
  AOI21_X1 U3801 ( .B1(n4990), .B2(n5590), .A(n4197), .ZN(n4198) );
  INV_X1 U3802 ( .A(n4196), .ZN(n4197) );
  NAND2_X1 U3803 ( .A1(n3019), .A2(n3017), .ZN(n4847) );
  NAND2_X1 U3804 ( .A1(n4262), .A2(n4264), .ZN(n4263) );
  NAND2_X1 U3805 ( .A1(n4652), .A2(n4695), .ZN(n4694) );
  AND4_X1 U3806 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n2982)
         );
  INV_X1 U3807 ( .A(n4023), .ZN(n5003) );
  INV_X1 U3808 ( .A(n3980), .ZN(n3981) );
  AND2_X2 U3809 ( .A1(n4434), .A2(n4340), .ZN(n3151) );
  NAND2_X1 U3810 ( .A1(n3022), .A2(n3997), .ZN(n4015) );
  AND2_X1 U3811 ( .A1(n4819), .A2(n4820), .ZN(n4763) );
  NAND2_X1 U3812 ( .A1(n3023), .A2(n3026), .ZN(n4697) );
  NAND2_X1 U3813 ( .A1(n3199), .A2(n3198), .ZN(n3308) );
  OR2_X1 U3814 ( .A1(n4773), .A2(n4222), .ZN(n2984) );
  INV_X1 U3815 ( .A(n3179), .ZN(n3114) );
  OR2_X1 U3816 ( .A1(n3194), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2985)
         );
  INV_X1 U3817 ( .A(n2996), .ZN(n4160) );
  NAND2_X1 U3818 ( .A1(n3201), .A2(n3190), .ZN(n2996) );
  NOR2_X1 U3819 ( .A1(n3980), .A2(n4705), .ZN(n2986) );
  NOR2_X1 U3820 ( .A1(n3980), .A2(n5565), .ZN(n2987) );
  AND2_X1 U3821 ( .A1(n3980), .A2(n4166), .ZN(n2988) );
  NAND2_X1 U3822 ( .A1(n2999), .A2(n4055), .ZN(n4056) );
  AND2_X1 U3823 ( .A1(n4816), .A2(n4817), .ZN(n4766) );
  AND2_X1 U3824 ( .A1(n3212), .A2(n3190), .ZN(n2989) );
  INV_X1 U3825 ( .A(n3303), .ZN(n3821) );
  INV_X1 U3826 ( .A(n5120), .ZN(n3018) );
  OAI21_X1 U3827 ( .B1(n4560), .B2(n2987), .A(n3982), .ZN(n5477) );
  AND2_X1 U3828 ( .A1(n3391), .A2(n3419), .ZN(n2990) );
  AND2_X1 U3829 ( .A1(n3980), .A2(n5167), .ZN(n2991) );
  OR2_X1 U3830 ( .A1(n3018), .A2(n3998), .ZN(n2992) );
  INV_X1 U3831 ( .A(n5541), .ZN(n5591) );
  INV_X1 U3832 ( .A(n5590), .ZN(n5540) );
  AND2_X1 U3833 ( .A1(n4173), .A2(n4148), .ZN(n5590) );
  NOR2_X1 U3834 ( .A1(n5284), .A2(n5285), .ZN(n4619) );
  AND2_X1 U3835 ( .A1(n4151), .A2(n3190), .ZN(n2993) );
  INV_X1 U3836 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3012) );
  INV_X1 U3837 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3013) );
  AND2_X1 U3838 ( .A1(n4794), .A2(n6168), .ZN(n2994) );
  AND2_X1 U3839 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n2995) );
  INV_X1 U3840 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4363) );
  NOR2_X2 U3841 ( .A1(n3296), .A2(n5766), .ZN(n3531) );
  NOR2_X1 U3842 ( .A1(n4233), .A2(n3190), .ZN(n4235) );
  NOR2_X2 U3843 ( .A1(n4799), .A2(n4798), .ZN(n3001) );
  AND2_X2 U3844 ( .A1(n4766), .A2(n4767), .ZN(n4811) );
  NOR2_X2 U3845 ( .A1(n5191), .A2(n5192), .ZN(n4753) );
  NOR2_X2 U3846 ( .A1(n4567), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U3847 ( .A1(n4565), .A2(n4566), .ZN(n4567) );
  NAND2_X1 U3848 ( .A1(n4031), .A2(n3202), .ZN(n3002) );
  NOR2_X1 U3849 ( .A1(n3190), .A2(n3180), .ZN(n3202) );
  NAND2_X1 U3850 ( .A1(n3211), .A2(n3201), .ZN(n4344) );
  NAND2_X1 U3852 ( .A1(n3116), .A2(n3115), .ZN(n4041) );
  NAND2_X1 U3853 ( .A1(n2947), .A2(n4652), .ZN(n4727) );
  INV_X1 U3854 ( .A(n4372), .ZN(n3009) );
  NOR2_X1 U3855 ( .A1(n4372), .A2(n4374), .ZN(n4373) );
  NAND4_X1 U3856 ( .A1(n4363), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n3013), .A4(n3012), .ZN(n3011) );
  NAND2_X1 U3857 ( .A1(n3222), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3156) );
  NAND3_X1 U3858 ( .A1(n4013), .A2(n3015), .A3(n3014), .ZN(U2956) );
  XNOR2_X1 U3859 ( .A(n4289), .B(n4205), .ZN(n4200) );
  OAI211_X1 U3860 ( .C1(n4273), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4272), .B(n4271), .ZN(n4286) );
  NOR2_X1 U3861 ( .A1(n4369), .A2(n3328), .ZN(n3329) );
  INV_X1 U3862 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U3863 ( .A1(n4853), .A2(n5328), .ZN(n4252) );
  NAND2_X1 U3864 ( .A1(n3926), .A2(n3925), .ZN(n5510) );
  NOR2_X1 U3865 ( .A1(n4343), .A2(n3186), .ZN(n4146) );
  INV_X1 U3866 ( .A(n3187), .ZN(n3171) );
  OR2_X1 U3867 ( .A1(n3277), .A2(n3276), .ZN(n3278) );
  INV_X1 U3868 ( .A(n3180), .ZN(n4149) );
  NAND2_X1 U3869 ( .A1(n3999), .A2(n4014), .ZN(n4018) );
  NAND2_X1 U3870 ( .A1(n3319), .A2(n3971), .ZN(n3299) );
  XNOR2_X1 U3871 ( .A(n4438), .B(n5966), .ZN(n4341) );
  NAND2_X1 U3872 ( .A1(n4286), .A2(n5533), .ZN(n4294) );
  OAI21_X2 U3873 ( .B1(n4707), .B2(n4708), .A(n4709), .ZN(n4953) );
  NAND2_X2 U3874 ( .A1(n3993), .A2(n3992), .ZN(n5135) );
  OR2_X1 U3875 ( .A1(n3981), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3032)
         );
  AND3_X1 U3876 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3033) );
  AND2_X1 U3877 ( .A1(n4833), .A2(n3302), .ZN(n5393) );
  NAND2_X1 U3878 ( .A1(n2977), .A2(n5619), .ZN(n4343) );
  INV_X1 U3879 ( .A(n4057), .ZN(n4065) );
  NAND2_X1 U3880 ( .A1(n3201), .A2(n3889), .ZN(n4153) );
  INV_X1 U3881 ( .A(n3531), .ZN(n3421) );
  INV_X1 U3882 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4260) );
  AND3_X1 U3883 ( .A1(n3238), .A2(n3237), .A3(n3236), .ZN(n3034) );
  AND2_X1 U3884 ( .A1(n6293), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3842)
         );
  INV_X1 U3885 ( .A(n4154), .ZN(n4155) );
  INV_X1 U3886 ( .A(n3912), .ZN(n3245) );
  INV_X1 U3887 ( .A(n3291), .ZN(n3923) );
  OR2_X1 U3888 ( .A1(n3368), .A2(n3367), .ZN(n3937) );
  INV_X1 U3889 ( .A(n4848), .ZN(n4001) );
  NAND2_X1 U3890 ( .A1(n4052), .A2(n5207), .ZN(n4057) );
  AND2_X1 U3891 ( .A1(n6445), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3834)
         );
  NAND2_X1 U3892 ( .A1(n3159), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3164)
         );
  INV_X1 U3893 ( .A(n3883), .ZN(n3332) );
  AOI22_X1 U3894 ( .A1(n3158), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2973), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3038) );
  AND2_X1 U3895 ( .A1(n4756), .A2(n4741), .ZN(n4114) );
  INV_X1 U3896 ( .A(n3371), .ZN(n3369) );
  NOR2_X1 U3897 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  NAND2_X1 U3898 ( .A1(n4207), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3424)
         );
  INV_X1 U3899 ( .A(n3242), .ZN(n3872) );
  OR3_X1 U3900 ( .A1(n3837), .A2(n6445), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n3900) );
  NOR2_X1 U3901 ( .A1(n3786), .A2(n4025), .ZN(n3787) );
  NAND2_X1 U3902 ( .A1(n3277), .A2(n3276), .ZN(n4438) );
  NOR2_X1 U3903 ( .A1(n4231), .A2(n4052), .ZN(n4136) );
  INV_X1 U3904 ( .A(n4030), .ZN(n3906) );
  AND2_X1 U3905 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3743), .ZN(n3744)
         );
  INV_X1 U3906 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3454) );
  AND4_X1 U3907 ( .A1(n4334), .A2(n4333), .A3(n4332), .A4(n4331), .ZN(n4336)
         );
  INV_X1 U3908 ( .A(n5630), .ZN(n5831) );
  AND2_X1 U3909 ( .A1(n5765), .A2(n5764), .ZN(n6072) );
  AND2_X1 U3910 ( .A1(n3901), .A2(n3900), .ZN(n6153) );
  NAND2_X1 U3911 ( .A1(n3744), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3786)
         );
  NAND2_X1 U3912 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5068), .ZN(n5055) );
  OR2_X1 U3913 ( .A1(n3535), .A2(n5258), .ZN(n3538) );
  NOR2_X1 U3914 ( .A1(n3422), .A2(n5493), .ZN(n3451) );
  NAND2_X1 U3915 ( .A1(n4758), .A2(n4759), .ZN(n4553) );
  AND2_X1 U3916 ( .A1(n4854), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U3917 ( .A1(n2946), .A2(n2945), .ZN(n4227) );
  NOR2_X1 U3918 ( .A1(n3646), .A2(n3645), .ZN(n3675) );
  NOR2_X1 U3919 ( .A1(n6339), .A2(n3566), .ZN(n3581) );
  NAND2_X1 U3920 ( .A1(n3510), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3535)
         );
  NOR2_X1 U3921 ( .A1(n6453), .A2(n3353), .ZN(n3378) );
  AOI211_X1 U3922 ( .C1(n4889), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4195), .B(n4194), .ZN(n4196) );
  NAND2_X1 U3923 ( .A1(n4873), .A2(n4257), .ZN(n4258) );
  OR2_X1 U3924 ( .A1(n3980), .A2(n4960), .ZN(n4709) );
  AND2_X1 U3925 ( .A1(n5595), .A2(n4661), .ZN(n4468) );
  OR2_X1 U3926 ( .A1(n5891), .A2(n6029), .ZN(n5673) );
  INV_X1 U3927 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6140) );
  OR2_X1 U3928 ( .A1(n5928), .A2(n5927), .ZN(n5964) );
  NAND2_X1 U3929 ( .A1(n6265), .A2(n4476), .ZN(n5629) );
  NOR2_X1 U3930 ( .A1(n5275), .A2(n4236), .ZN(n5251) );
  INV_X1 U3931 ( .A(n5336), .ZN(n5328) );
  NAND2_X1 U3932 ( .A1(n4619), .A2(n4620), .ZN(n4666) );
  INV_X1 U3933 ( .A(n4833), .ZN(n4774) );
  INV_X1 U3934 ( .A(n3908), .ZN(n3909) );
  AND2_X1 U3935 ( .A1(n4839), .A2(n4151), .ZN(n5396) );
  INV_X1 U3936 ( .A(n5435), .ZN(n6307) );
  AND2_X1 U3937 ( .A1(n3828), .A2(n4298), .ZN(n4385) );
  AOI21_X1 U3938 ( .B1(n4385), .B2(n4384), .A(n5459), .ZN(n5458) );
  NAND2_X1 U3939 ( .A1(n3692), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3742)
         );
  NAND2_X1 U3940 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3353) );
  INV_X1 U3941 ( .A(n5530), .ZN(n5517) );
  INV_X1 U3942 ( .A(n2983), .ZN(n4990) );
  AND2_X1 U3943 ( .A1(n4937), .A2(n5175), .ZN(n4935) );
  OR3_X1 U3944 ( .A1(n5581), .A2(n4183), .A3(n4182), .ZN(n5190) );
  OR2_X1 U3945 ( .A1(n4468), .A2(n4186), .ZN(n5568) );
  INV_X1 U3946 ( .A(n4662), .ZN(n5582) );
  INV_X1 U3947 ( .A(n5669), .ZN(n5657) );
  INV_X1 U3948 ( .A(n5695), .ZN(n5672) );
  OR2_X1 U3949 ( .A1(n4488), .A2(n4452), .ZN(n4489) );
  INV_X1 U3950 ( .A(n5775), .ZN(n5822) );
  INV_X1 U3951 ( .A(n5858), .ZN(n5850) );
  INV_X1 U3952 ( .A(n5875), .ZN(n5882) );
  NOR2_X1 U3953 ( .A1(n5928), .A2(n5926), .ZN(n5859) );
  INV_X1 U3954 ( .A(n5964), .ZN(n5987) );
  INV_X1 U3955 ( .A(n3920), .ZN(n6290) );
  INV_X1 U3956 ( .A(n6027), .ZN(n6065) );
  INV_X1 U3957 ( .A(n5640), .ZN(n6127) );
  AND2_X1 U3958 ( .A1(n5202), .A2(n6181), .ZN(n4297) );
  INV_X1 U3959 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6180) );
  AOI21_X1 U3960 ( .B1(n4888), .B2(n5369), .A(n4250), .ZN(n4251) );
  INV_X1 U3961 ( .A(n5353), .ZN(n5370) );
  NAND2_X1 U3962 ( .A1(n4605), .A2(n4219), .ZN(n5336) );
  INV_X1 U3963 ( .A(n5393), .ZN(n4835) );
  NAND2_X1 U3964 ( .A1(n4403), .A2(n3905), .ZN(n4839) );
  NAND2_X1 U3965 ( .A1(n5426), .A2(n3843), .ZN(n5410) );
  OR2_X1 U3966 ( .A1(n6170), .A2(n5426), .ZN(n5436) );
  NAND2_X1 U3967 ( .A1(n4385), .A2(n3884), .ZN(n4403) );
  INV_X1 U3968 ( .A(n5458), .ZN(n4522) );
  OR2_X1 U3969 ( .A1(n6169), .A2(n4383), .ZN(n6440) );
  INV_X1 U3970 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5493) );
  INV_X1 U3971 ( .A(n5483), .ZN(n5525) );
  AND2_X1 U3972 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  OR2_X1 U3973 ( .A1(n4471), .A2(n4470), .ZN(n5552) );
  NAND2_X1 U3974 ( .A1(n4173), .A2(n4050), .ZN(n5541) );
  OR2_X1 U3975 ( .A1(n6316), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5599) );
  OR2_X1 U3976 ( .A1(n6021), .A2(n3920), .ZN(n5640) );
  NAND2_X1 U3977 ( .A1(n5643), .A2(n6290), .ZN(n5695) );
  OR2_X1 U3978 ( .A1(n4489), .A2(n3920), .ZN(n5734) );
  OR2_X1 U3979 ( .A1(n5735), .A2(n6290), .ZN(n5763) );
  OR2_X1 U3980 ( .A1(n5735), .A2(n3920), .ZN(n5795) );
  OR2_X1 U3981 ( .A1(n5806), .A2(n3920), .ZN(n5858) );
  NAND2_X1 U3982 ( .A1(n5859), .A2(n6290), .ZN(n5918) );
  OR2_X1 U3983 ( .A1(n5999), .A2(n3920), .ZN(n6027) );
  NAND2_X1 U3984 ( .A1(n6077), .A2(n3920), .ZN(n6132) );
  INV_X1 U3985 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6395) );
  INV_X1 U3986 ( .A(n6263), .ZN(n6261) );
  INV_X1 U3987 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6199) );
  INV_X1 U3988 ( .A(n6255), .ZN(n6253) );
  NAND2_X1 U3989 ( .A1(n4252), .A2(n4251), .ZN(U2796) );
  OAI21_X1 U3990 ( .B1(n4993), .B2(n4835), .A(n4204), .ZN(U2829) );
  AND2_X2 U3991 ( .A1(n3312), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3042)
         );
  AND2_X2 U3992 ( .A1(n3042), .A2(n3043), .ZN(n3137) );
  INV_X1 U3993 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3036) );
  AND2_X2 U3994 ( .A1(n4338), .A2(n4340), .ZN(n3231) );
  AOI22_X1 U3995 ( .A1(n3137), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3041) );
  INV_X1 U3996 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3037) );
  AOI22_X1 U3997 ( .A1(n3279), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2975), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3040) );
  NOR2_X4 U3998 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U3999 ( .A1(n3159), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3039) );
  AND2_X2 U4000 ( .A1(n4361), .A2(n4338), .ZN(n3158) );
  AOI22_X1 U4001 ( .A1(n3150), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3049) );
  AOI22_X1 U4002 ( .A1(n3138), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3048) );
  AOI22_X1 U4003 ( .A1(n3161), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U4004 ( .A1(n3144), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3046) );
  AOI22_X1 U4005 ( .A1(n3139), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U4006 ( .A1(n3279), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U4007 ( .A1(n3137), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U4008 ( .A1(n3231), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U4009 ( .A1(n3150), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3057) );
  NAND2_X2 U4010 ( .A1(n3061), .A2(n3060), .ZN(n3179) );
  AOI22_X1 U4011 ( .A1(n3137), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U4012 ( .A1(n3158), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U4013 ( .A1(n3159), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U4014 ( .A1(n3279), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U4015 ( .A1(n3161), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U4016 ( .A1(n3144), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U4017 ( .A1(n3138), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3066) );
  NAND2_X2 U4018 ( .A1(n3071), .A2(n3070), .ZN(n3296) );
  NOR2_X2 U4019 ( .A1(n3114), .A2(n3296), .ZN(n3082) );
  NAND2_X1 U4020 ( .A1(n3296), .A2(n3114), .ZN(n3888) );
  AOI22_X1 U4021 ( .A1(n3137), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3075) );
  AOI22_X1 U4022 ( .A1(n3159), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3074) );
  AOI22_X1 U4023 ( .A1(n3139), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3073) );
  AOI22_X1 U4024 ( .A1(n3222), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3072) );
  NAND4_X1 U4025 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(n3081)
         );
  AOI22_X1 U4026 ( .A1(n3144), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U4027 ( .A1(n3158), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U4028 ( .A1(n3150), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3221), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U4029 ( .A1(n3279), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3076) );
  NAND4_X1 U4030 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3080)
         );
  NAND2_X1 U4031 ( .A1(n3082), .A2(n3216), .ZN(n3083) );
  OAI21_X1 U4032 ( .B1(n3216), .B2(n3203), .A(n4154), .ZN(n3200) );
  INV_X1 U4033 ( .A(n3200), .ZN(n3116) );
  AOI22_X1 U4034 ( .A1(n3137), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3088) );
  AOI22_X1 U4035 ( .A1(n3279), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3152), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3087) );
  AOI22_X1 U4036 ( .A1(n3159), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3086) );
  AOI22_X1 U4037 ( .A1(n3158), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2972), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3085) );
  NAND4_X1 U4038 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3094)
         );
  AOI22_X1 U4039 ( .A1(n3161), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3139), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U4040 ( .A1(n3138), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3091) );
  AOI22_X1 U4041 ( .A1(n3150), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3090) );
  NAND4_X1 U4042 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), .ZN(n3093)
         );
  NAND2_X1 U4044 ( .A1(n3137), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U4045 ( .A1(n3158), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U4046 ( .A1(n3231), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3096)
         );
  NAND2_X1 U4047 ( .A1(n3151), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3095)
         );
  NAND2_X1 U4048 ( .A1(n3222), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4049 ( .A1(n3150), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3101)
         );
  NAND2_X1 U4050 ( .A1(n3161), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U4051 ( .A1(n3139), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3099)
         );
  NAND2_X1 U4052 ( .A1(n3144), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U4053 ( .A1(n3138), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U4054 ( .A1(n3221), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U4055 ( .A1(n3145), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U4056 ( .A1(n2975), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U4057 ( .A1(n3159), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3109)
         );
  NAND2_X1 U4058 ( .A1(n3279), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3108)
         );
  NAND2_X1 U4059 ( .A1(n2971), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4060 ( .A1(n3150), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3120)
         );
  NAND2_X1 U4061 ( .A1(n3222), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U4062 ( .A1(n3161), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U4063 ( .A1(n3139), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3117)
         );
  NAND2_X1 U4064 ( .A1(n3137), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U4065 ( .A1(n3158), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4066 ( .A1(n3231), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3122)
         );
  NAND2_X1 U4067 ( .A1(n3151), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3121)
         );
  NAND2_X1 U4068 ( .A1(n3279), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3128)
         );
  NAND2_X1 U4069 ( .A1(n3159), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3127)
         );
  NAND2_X1 U4070 ( .A1(n2975), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3126) );
  NAND2_X1 U4071 ( .A1(n3160), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U4072 ( .A1(n3144), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U4073 ( .A1(n3138), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4074 ( .A1(n3221), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4075 ( .A1(n3145), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U4076 ( .A1(n3137), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4077 ( .A1(n3138), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4078 ( .A1(n3221), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U4079 ( .A1(n3139), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U4080 ( .A1(n3279), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3149)
         );
  NAND2_X1 U4081 ( .A1(n3144), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4082 ( .A1(n3231), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U4083 ( .A1(n3145), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4084 ( .A1(n3150), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3155)
         );
  NAND2_X1 U4085 ( .A1(n3151), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3154)
         );
  NAND2_X1 U4086 ( .A1(n3152), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4087 ( .A1(n3158), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4088 ( .A1(n3160), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4089 ( .A1(n3161), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3162) );
  NAND4_X4 U4090 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3180)
         );
  NOR2_X1 U4091 ( .A1(n6199), .A2(n6209), .ZN(n6202) );
  INV_X1 U4092 ( .A(n6202), .ZN(n3170) );
  OAI21_X1 U4093 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n3170), .ZN(n4035) );
  NAND2_X1 U4094 ( .A1(n4149), .A2(n4035), .ZN(n3181) );
  NAND2_X1 U4095 ( .A1(n3827), .A2(n3181), .ZN(n3174) );
  AND2_X2 U4096 ( .A1(n3296), .A2(n3302), .ZN(n4151) );
  NAND3_X1 U4097 ( .A1(n4151), .A2(n3839), .A3(n3889), .ZN(n3186) );
  AND2_X2 U4098 ( .A1(n3216), .A2(n3179), .ZN(n4003) );
  NAND2_X1 U4099 ( .A1(n3172), .A2(n3171), .ZN(n4033) );
  NOR2_X2 U4100 ( .A1(n4033), .A2(n3180), .ZN(n4440) );
  NOR2_X1 U4101 ( .A1(n4146), .A2(n4440), .ZN(n3173) );
  NAND2_X1 U4102 ( .A1(n3174), .A2(n3173), .ZN(n3175) );
  NAND2_X1 U4103 ( .A1(n3175), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3196) );
  INV_X1 U4104 ( .A(n3196), .ZN(n3178) );
  NOR2_X1 U4105 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6182) );
  NAND2_X1 U4106 ( .A1(n6182), .A2(n6180), .ZN(n4005) );
  INV_X1 U4107 ( .A(n4005), .ZN(n3333) );
  XNOR2_X1 U4108 ( .A(n6140), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6022)
         );
  NAND2_X1 U4109 ( .A1(n3333), .A2(n6022), .ZN(n3177) );
  NAND2_X1 U4110 ( .A1(n3332), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4111 ( .A1(n3177), .A2(n3176), .ZN(n3194) );
  NAND2_X1 U4112 ( .A1(n3178), .A2(n2985), .ZN(n3269) );
  NAND3_X1 U4113 ( .A1(n3888), .A2(n3302), .A3(n3216), .ZN(n4031) );
  NAND2_X1 U4114 ( .A1(n3181), .A2(n3839), .ZN(n3182) );
  NAND3_X1 U4115 ( .A1(n3886), .A2(n3207), .A3(n3182), .ZN(n3183) );
  NAND2_X1 U4116 ( .A1(n3183), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3193) );
  OAI21_X1 U4117 ( .B1(n3203), .B2(n5619), .A(n4149), .ZN(n3184) );
  INV_X1 U4118 ( .A(n3184), .ZN(n3189) );
  NAND3_X1 U4119 ( .A1(n3187), .A2(n4029), .A3(n3186), .ZN(n3188) );
  NAND2_X1 U4120 ( .A1(n3189), .A2(n3188), .ZN(n3210) );
  INV_X1 U4121 ( .A(n3336), .ZN(n3292) );
  NOR2_X1 U4122 ( .A1(n3242), .A2(n3203), .ZN(n3191) );
  NAND2_X1 U4123 ( .A1(n3193), .A2(n3192), .ZN(n3197) );
  NAND2_X1 U4124 ( .A1(n3196), .A2(n3195), .ZN(n3268) );
  NAND2_X1 U4125 ( .A1(n3269), .A2(n3268), .ZN(n3215) );
  NAND2_X1 U4126 ( .A1(n3197), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3199) );
  MUX2_X1 U4127 ( .A(n3883), .B(n4005), .S(n6293), .Z(n3198) );
  OAI21_X1 U4128 ( .B1(n3200), .B2(n5619), .A(n3180), .ZN(n3214) );
  INV_X1 U4129 ( .A(n6182), .ZN(n6273) );
  NAND2_X1 U4130 ( .A1(n3913), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4131 ( .A1(n3204), .A2(n3336), .ZN(n3205) );
  OAI211_X1 U4132 ( .C1(n3201), .C2(n4029), .A(n3206), .B(n3205), .ZN(n3209)
         );
  INV_X1 U4133 ( .A(n3207), .ZN(n3208) );
  NOR2_X1 U4134 ( .A1(n3209), .A2(n3208), .ZN(n3213) );
  INV_X1 U4135 ( .A(n3211), .ZN(n3212) );
  NAND2_X1 U4136 ( .A1(n3210), .A2(n2989), .ZN(n4159) );
  NAND3_X1 U4137 ( .A1(n3214), .A2(n3213), .A3(n4159), .ZN(n3309) );
  AND2_X2 U4138 ( .A1(n3308), .A2(n3309), .ZN(n3311) );
  XNOR2_X1 U4139 ( .A(n3215), .B(n3311), .ZN(n4356) );
  NAND2_X1 U4140 ( .A1(n4356), .A2(n6180), .ZN(n3230) );
  AOI22_X1 U4141 ( .A1(n3808), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4142 ( .A1(n3796), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4143 ( .A1(n4339), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4144 ( .A1(n3161), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3217) );
  NAND4_X1 U4145 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3228)
         );
  AOI22_X1 U4146 ( .A1(n3806), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3804), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4147 ( .A1(n3798), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3225) );
  INV_X1 U4148 ( .A(n3221), .ZN(n3600) );
  AOI22_X1 U4149 ( .A1(n3775), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4150 ( .A1(n3794), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3223) );
  NAND4_X1 U4151 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3227)
         );
  NAND2_X1 U4152 ( .A1(n3230), .A2(n3229), .ZN(n3301) );
  AOI22_X1 U4153 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n3159), .B1(n3144), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4154 ( .A1(n3247), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4155 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n3796), .B1(n3145), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4156 ( .A1(n3804), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3232) );
  NAND4_X1 U4157 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3241)
         );
  AOI22_X1 U4158 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n3794), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3239) );
  INV_X2 U4159 ( .A(n3600), .ZN(n3799) );
  AOI22_X1 U4160 ( .A1(n3150), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4161 ( .A1(n4339), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4162 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n3808), .B1(n3160), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3236) );
  OR2_X2 U4163 ( .A1(n3241), .A2(n3240), .ZN(n3973) );
  NOR2_X1 U4164 ( .A1(n3890), .A2(n3973), .ZN(n3260) );
  INV_X1 U4165 ( .A(n3260), .ZN(n3244) );
  NAND2_X1 U4166 ( .A1(n3872), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3243) );
  OAI211_X1 U4167 ( .C1(n3245), .C2(n3336), .A(n3244), .B(n3243), .ZN(n3298)
         );
  INV_X1 U4168 ( .A(n3308), .ZN(n3246) );
  AOI22_X1 U4169 ( .A1(n3137), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4170 ( .A1(n3247), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3138), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4171 ( .A1(n4339), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4172 ( .A1(n3794), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3248) );
  NAND4_X1 U4173 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3257)
         );
  AOI22_X1 U4174 ( .A1(n3806), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3145), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4175 ( .A1(n3798), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4176 ( .A1(n3804), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4177 ( .A1(n3144), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3252) );
  NAND4_X1 U4178 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3256)
         );
  INV_X1 U4179 ( .A(n3973), .ZN(n3258) );
  AOI21_X1 U4180 ( .B1(n3260), .B2(n3917), .A(n3259), .ZN(n3317) );
  NAND2_X1 U4181 ( .A1(n3261), .A2(n3317), .ZN(n3265) );
  INV_X1 U4182 ( .A(n3917), .ZN(n3264) );
  NAND2_X1 U4183 ( .A1(n3872), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3263) );
  AOI21_X1 U4184 ( .B1(n3216), .B2(n3973), .A(n6180), .ZN(n3262) );
  OAI211_X1 U4185 ( .C1(n3843), .C2(n3264), .A(n3263), .B(n3262), .ZN(n3315)
         );
  NAND2_X1 U4186 ( .A1(n3265), .A2(n3315), .ZN(n3319) );
  OAI21_X1 U4187 ( .B1(n3301), .B2(n3298), .A(n3299), .ZN(n3267) );
  NAND2_X1 U4188 ( .A1(n3301), .A2(n3298), .ZN(n3266) );
  NAND2_X1 U4189 ( .A1(n3268), .A2(n3311), .ZN(n3270) );
  NAND2_X1 U4190 ( .A1(n3270), .A2(n3269), .ZN(n3277) );
  NAND2_X1 U4191 ( .A1(n3197), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3275) );
  AND2_X1 U4192 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4193 ( .A1(n3271), .A2(n6145), .ZN(n4475) );
  INV_X1 U4194 ( .A(n3271), .ZN(n3272) );
  NAND2_X1 U4195 ( .A1(n3272), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4196 ( .A1(n4475), .A2(n3273), .ZN(n5767) );
  AOI22_X1 U4197 ( .A1(n3333), .A2(n5767), .B1(n3332), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4198 ( .A1(n3278), .A2(n4438), .ZN(n4418) );
  AOI22_X1 U4199 ( .A1(n3796), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3284) );
  INV_X1 U4200 ( .A(n3279), .ZN(n3280) );
  INV_X2 U4201 ( .A(n3280), .ZN(n3808) );
  AOI22_X1 U4202 ( .A1(n3808), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4203 ( .A1(n3798), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4204 ( .A1(n3804), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4205 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3290)
         );
  AOI22_X1 U4206 ( .A1(n3806), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4207 ( .A1(n3138), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2976), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3287) );
  INV_X1 U4208 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6442) );
  AOI22_X1 U4209 ( .A1(n3161), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4210 ( .A1(n3795), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4211 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3289)
         );
  OAI22_X2 U4212 ( .A1(n4418), .A2(STATE2_REG_0__SCAN_IN), .B1(n3923), .B2(
        n3890), .ZN(n3294) );
  AOI22_X1 U4213 ( .A1(n3292), .A2(n3291), .B1(n3872), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3293) );
  XNOR2_X2 U4214 ( .A(n3294), .B(n3293), .ZN(n3350) );
  INV_X1 U4215 ( .A(n3350), .ZN(n3295) );
  NAND2_X1 U4216 ( .A1(n4451), .A2(n3531), .ZN(n3297) );
  XNOR2_X1 U4217 ( .A(n3299), .B(n3298), .ZN(n3300) );
  NAND2_X1 U4218 ( .A1(n4447), .A2(n3531), .ZN(n3307) );
  AOI22_X1 U4219 ( .A1(n3763), .A2(EAX_REG_1__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3305) );
  AND2_X1 U4220 ( .A1(n4151), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4221 ( .A1(n3327), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3304) );
  AND2_X1 U4222 ( .A1(n3305), .A2(n3304), .ZN(n3306) );
  NAND2_X1 U4223 ( .A1(n3307), .A2(n3306), .ZN(n4367) );
  NOR2_X1 U4224 ( .A1(n3308), .A2(n3309), .ZN(n3310) );
  OR2_X1 U4225 ( .A1(n3311), .A2(n3310), .ZN(n5921) );
  INV_X1 U4226 ( .A(n3327), .ZN(n3375) );
  AOI22_X1 U4227 ( .A1(n3763), .A2(EAX_REG_0__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3313) );
  OAI21_X1 U4228 ( .B1(n3375), .B2(n3312), .A(n3313), .ZN(n3314) );
  AOI21_X1 U4229 ( .B1(n6288), .B2(n3531), .A(n3314), .ZN(n4377) );
  NOR2_X2 U4230 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3826) );
  INV_X1 U4231 ( .A(n3315), .ZN(n3316) );
  NAND2_X1 U4232 ( .A1(n3317), .A2(n3316), .ZN(n3318) );
  NAND3_X1 U4233 ( .A1(n3920), .A2(n3320), .A3(n3302), .ZN(n3321) );
  NAND2_X1 U4234 ( .A1(n3321), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4376) );
  NOR2_X1 U4235 ( .A1(n4377), .A2(n4376), .ZN(n4375) );
  AOI21_X1 U4236 ( .B1(n4377), .B2(n3826), .A(n4375), .ZN(n3322) );
  INV_X1 U4237 ( .A(n3322), .ZN(n4366) );
  NAND2_X1 U4238 ( .A1(n4367), .A2(n4366), .ZN(n4369) );
  INV_X1 U4239 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4240 ( .A1(n3763), .A2(EAX_REG_2__SCAN_IN), .ZN(n3324) );
  OAI21_X1 U4241 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3353), .ZN(n5516) );
  NAND2_X1 U4242 ( .A1(n3826), .A2(n5516), .ZN(n3323) );
  OAI211_X1 U4243 ( .C1(n3689), .C2(n3325), .A(n3324), .B(n3323), .ZN(n3326)
         );
  AOI21_X1 U4244 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n3327), .A(n3326), 
        .ZN(n3328) );
  NAND2_X1 U4245 ( .A1(n4369), .A2(n3328), .ZN(n4380) );
  NAND2_X1 U4246 ( .A1(n3197), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3335) );
  NOR3_X1 U4247 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6145), .A3(n6140), 
        .ZN(n5805) );
  NAND2_X1 U4248 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5805), .ZN(n5800) );
  NAND2_X1 U4249 ( .A1(n6284), .A2(n5800), .ZN(n3331) );
  NAND3_X1 U4250 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6078) );
  INV_X1 U4251 ( .A(n6078), .ZN(n3330) );
  NAND2_X1 U4252 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3330), .ZN(n6071) );
  AOI22_X1 U4253 ( .A1(n3333), .A2(n5828), .B1(n3332), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4254 ( .A1(n4341), .A2(n6180), .ZN(n3348) );
  AOI22_X1 U4255 ( .A1(n3796), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4256 ( .A1(n3808), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4257 ( .A1(n3798), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4258 ( .A1(n3804), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4259 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3346)
         );
  AOI22_X1 U4260 ( .A1(n3806), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4261 ( .A1(n3138), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4262 ( .A1(n3805), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4263 ( .A1(n3795), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3341) );
  NAND4_X1 U4264 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3345)
         );
  AOI22_X1 U4265 ( .A1(n3861), .A2(n3931), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3872), .ZN(n3347) );
  NAND3_X1 U4266 ( .A1(n3349), .A2(n3350), .A3(n5706), .ZN(n3372) );
  NAND2_X1 U4267 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  NAND2_X1 U4268 ( .A1(n3351), .A2(n5797), .ZN(n3352) );
  INV_X1 U4269 ( .A(n3933), .ZN(n3357) );
  AOI21_X1 U4270 ( .B1(n6453), .B2(n3353), .A(n3378), .ZN(n4616) );
  INV_X2 U4271 ( .A(n3826), .ZN(n4211) );
  OAI22_X1 U4272 ( .A1(n4616), .A2(n4211), .B1(n6453), .B2(n3689), .ZN(n3354)
         );
  AOI21_X1 U4273 ( .B1(n3763), .B2(EAX_REG_3__SCAN_IN), .A(n3354), .ZN(n3355)
         );
  OAI21_X1 U4274 ( .B1(n3012), .B2(n3375), .A(n3355), .ZN(n3356) );
  AOI21_X1 U4275 ( .B1(n3357), .B2(n3531), .A(n3356), .ZN(n4374) );
  INV_X1 U4276 ( .A(n3372), .ZN(n3370) );
  AOI22_X1 U4277 ( .A1(n3806), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4278 ( .A1(n3798), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3160), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4279 ( .A1(n3796), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4280 ( .A1(n3358), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4281 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3368)
         );
  AOI22_X1 U4282 ( .A1(n3804), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4283 ( .A1(n3794), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4284 ( .A1(n3795), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4285 ( .A1(n4339), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4286 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3367)
         );
  AOI22_X1 U4287 ( .A1(n3861), .A2(n3937), .B1(n3872), .B2(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4288 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  NAND2_X1 U4289 ( .A1(n3393), .A2(n3373), .ZN(n3939) );
  INV_X1 U4290 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6441) );
  INV_X1 U4291 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3374) );
  OAI22_X1 U4292 ( .A1(n3821), .A2(n6441), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3374), .ZN(n3377) );
  NOR2_X1 U4293 ( .A1(n3375), .A2(n5200), .ZN(n3376) );
  OAI21_X1 U4294 ( .B1(n3377), .B2(n3376), .A(n4211), .ZN(n3380) );
  OAI21_X1 U4295 ( .B1(n3378), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3395), 
        .ZN(n5360) );
  NAND2_X1 U4296 ( .A1(n5360), .A2(n3826), .ZN(n3379) );
  AOI22_X1 U4297 ( .A1(n3796), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3384) );
  INV_X1 U4298 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6333) );
  AOI22_X1 U4299 ( .A1(n3808), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4300 ( .A1(n3798), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4301 ( .A1(n3804), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4302 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4303 ( .A1(n3806), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4304 ( .A1(n3358), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4305 ( .A1(n3805), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4306 ( .A1(n3795), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4307 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  AOI22_X1 U4308 ( .A1(n3861), .A2(n3945), .B1(n3872), .B2(
        INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U4309 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  NAND2_X1 U4310 ( .A1(n3418), .A2(n3394), .ZN(n3948) );
  INV_X1 U4311 ( .A(n3948), .ZN(n3398) );
  AOI21_X1 U4312 ( .B1(n3395), .B2(n5509), .A(n3412), .ZN(n5341) );
  AOI22_X1 U4313 ( .A1(n3763), .A2(EAX_REG_5__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3396) );
  OAI21_X1 U4314 ( .B1(n4211), .B2(n5341), .A(n3396), .ZN(n3397) );
  AOI22_X1 U4315 ( .A1(n3798), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4316 ( .A1(n3804), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4317 ( .A1(n3808), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4318 ( .A1(n3796), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3399) );
  NAND4_X1 U4319 ( .A1(n3402), .A2(n3401), .A3(n3400), .A4(n3399), .ZN(n3408)
         );
  AOI22_X1 U4320 ( .A1(n3247), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4321 ( .A1(n3794), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4322 ( .A1(n3806), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4323 ( .A1(n3805), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3403) );
  NAND4_X1 U4324 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3407)
         );
  NAND2_X1 U4325 ( .A1(n3861), .A2(n3961), .ZN(n3410) );
  NAND2_X1 U4326 ( .A1(n3872), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4327 ( .A1(n3410), .A2(n3409), .ZN(n3419) );
  INV_X1 U4328 ( .A(n3419), .ZN(n3411) );
  NAND2_X1 U4329 ( .A1(n3418), .A2(n3411), .ZN(n3953) );
  INV_X1 U4330 ( .A(n3953), .ZN(n3417) );
  INV_X1 U4331 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3414) );
  OAI21_X1 U4332 ( .B1(n3412), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3422), 
        .ZN(n5495) );
  NAND2_X1 U4333 ( .A1(n3826), .A2(n5495), .ZN(n3413) );
  OAI21_X1 U4334 ( .B1(n3414), .B2(n3689), .A(n3413), .ZN(n3415) );
  AOI21_X1 U4335 ( .B1(n3763), .B2(EAX_REG_6__SCAN_IN), .A(n3415), .ZN(n3416)
         );
  NAND2_X1 U4336 ( .A1(n4405), .A2(n4407), .ZN(n4406) );
  AOI22_X1 U4337 ( .A1(n3861), .A2(n3973), .B1(INSTQUEUE_REG_0__7__SCAN_IN), 
        .B2(n3872), .ZN(n3420) );
  INV_X1 U4338 ( .A(n3965), .ZN(n3427) );
  AOI21_X1 U4339 ( .B1(n3422), .B2(n5493), .A(n3451), .ZN(n3423) );
  INV_X1 U4340 ( .A(n3423), .ZN(n5487) );
  AOI22_X1 U4341 ( .A1(n5487), .A2(n3826), .B1(n3763), .B2(EAX_REG_7__SCAN_IN), 
        .ZN(n3425) );
  AOI21_X1 U4342 ( .B1(n3427), .B2(n3531), .A(n3426), .ZN(n4516) );
  XOR2_X1 U4343 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3451), .Z(n5318) );
  AOI22_X1 U4344 ( .A1(n3763), .A2(EAX_REG_8__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4345 ( .A1(n3804), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4346 ( .A1(n3794), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4347 ( .A1(n3358), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4348 ( .A1(n3796), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4349 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3437)
         );
  AOI22_X1 U4350 ( .A1(n3806), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4351 ( .A1(n3798), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4352 ( .A1(n3795), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4353 ( .A1(n3805), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3432) );
  NAND4_X1 U4354 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3436)
         );
  OAI21_X1 U4355 ( .B1(n3437), .B2(n3436), .A(n3531), .ZN(n3438) );
  OAI211_X1 U4356 ( .C1(n5318), .C2(n4211), .A(n3439), .B(n3438), .ZN(n4518)
         );
  NAND2_X1 U4357 ( .A1(n4515), .A2(n4518), .ZN(n4548) );
  AOI22_X1 U4358 ( .A1(n3808), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4359 ( .A1(n3794), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4360 ( .A1(n3775), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4361 ( .A1(n3798), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4362 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3449)
         );
  AOI22_X1 U4363 ( .A1(n3806), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4364 ( .A1(n3796), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4365 ( .A1(n3804), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4366 ( .A1(n3247), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4367 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3448)
         );
  OAI21_X1 U4368 ( .B1(n3449), .B2(n3448), .A(n3531), .ZN(n3450) );
  OAI21_X1 U4369 ( .B1(n3454), .B2(n3689), .A(n3450), .ZN(n3453) );
  XNOR2_X1 U4370 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3455), .ZN(n5308) );
  NOR2_X1 U4371 ( .A1(n5308), .A2(n4211), .ZN(n3452) );
  AOI211_X1 U4372 ( .C1(n3763), .C2(EAX_REG_9__SCAN_IN), .A(n3453), .B(n3452), 
        .ZN(n4547) );
  XOR2_X1 U4373 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3480), .Z(n5482) );
  AOI22_X1 U4374 ( .A1(n3763), .A2(EAX_REG_10__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4375 ( .A1(n3358), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4376 ( .A1(n3796), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4377 ( .A1(n3805), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4378 ( .A1(n4339), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4379 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3465)
         );
  AOI22_X1 U4380 ( .A1(n3804), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4381 ( .A1(n3798), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4382 ( .A1(n3795), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4383 ( .A1(n3806), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3460) );
  NAND4_X1 U4384 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(n3464)
         );
  OAI21_X1 U4385 ( .B1(n3465), .B2(n3464), .A(n3531), .ZN(n3466) );
  OAI211_X1 U4386 ( .C1(n5482), .C2(n4211), .A(n3467), .B(n3466), .ZN(n4545)
         );
  INV_X1 U4387 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4388 ( .A1(n3804), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4389 ( .A1(n3796), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4390 ( .A1(n3775), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4391 ( .A1(n3806), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4392 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3477)
         );
  AOI22_X1 U4393 ( .A1(n3798), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4394 ( .A1(n3795), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4395 ( .A1(n3808), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4396 ( .A1(n3247), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4397 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3476)
         );
  OAI21_X1 U4398 ( .B1(n3477), .B2(n3476), .A(n3531), .ZN(n3478) );
  OAI21_X1 U4399 ( .B1(n3479), .B2(n3689), .A(n3478), .ZN(n3482) );
  XNOR2_X1 U4400 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3483), .ZN(n5474)
         );
  NOR2_X1 U4401 ( .A1(n5474), .A2(n4211), .ZN(n3481) );
  AOI211_X1 U4402 ( .C1(n3303), .C2(EAX_REG_11__SCAN_IN), .A(n3482), .B(n3481), 
        .ZN(n4596) );
  AOI21_X1 U4403 ( .B1(n6392), .B2(n3484), .A(n3510), .ZN(n5464) );
  AOI22_X1 U4404 ( .A1(n3303), .A2(EAX_REG_12__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4405 ( .A1(n3796), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4406 ( .A1(n3798), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4407 ( .A1(n3247), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4408 ( .A1(n3806), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3485) );
  NAND4_X1 U4409 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3494)
         );
  AOI22_X1 U4410 ( .A1(n4339), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4411 ( .A1(n3808), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4412 ( .A1(n3358), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4413 ( .A1(n3804), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3489) );
  NAND4_X1 U4414 ( .A1(n3492), .A2(n3491), .A3(n3490), .A4(n3489), .ZN(n3493)
         );
  OAI21_X1 U4415 ( .B1(n3494), .B2(n3493), .A(n3531), .ZN(n3495) );
  OAI211_X1 U4416 ( .C1(n5464), .C2(n4211), .A(n3496), .B(n3495), .ZN(n4600)
         );
  NAND2_X1 U4417 ( .A1(n4595), .A2(n4600), .ZN(n4599) );
  INV_X1 U4418 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U4419 ( .A1(n3806), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4420 ( .A1(n3796), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4421 ( .A1(n3795), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4422 ( .A1(n3358), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4423 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3506)
         );
  AOI22_X1 U4424 ( .A1(n3804), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4425 ( .A1(n3798), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4426 ( .A1(n3247), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4427 ( .A1(n3808), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4428 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3505)
         );
  OAI21_X1 U4429 ( .B1(n3506), .B2(n3505), .A(n3531), .ZN(n3507) );
  OAI21_X1 U4430 ( .B1(n4675), .B2(n3689), .A(n3507), .ZN(n3509) );
  XOR2_X1 U4431 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3510), .Z(n5271) );
  NOR2_X1 U4432 ( .A1(n5271), .A2(n4211), .ZN(n3508) );
  AOI211_X1 U4433 ( .C1(n3303), .C2(EAX_REG_13__SCAN_IN), .A(n3509), .B(n3508), 
        .ZN(n4623) );
  XNOR2_X1 U4434 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3535), .ZN(n5262)
         );
  AOI22_X1 U4435 ( .A1(n3303), .A2(EAX_REG_14__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4436 ( .A1(n3798), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4437 ( .A1(n3804), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4438 ( .A1(n3794), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4439 ( .A1(n3775), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4440 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3520)
         );
  AOI22_X1 U4441 ( .A1(n3796), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4442 ( .A1(n3806), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4443 ( .A1(n4339), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4444 ( .A1(n3358), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4445 ( .A1(n3518), .A2(n3517), .A3(n3516), .A4(n3515), .ZN(n3519)
         );
  OAI21_X1 U4446 ( .B1(n3520), .B2(n3519), .A(n3531), .ZN(n3521) );
  OAI211_X1 U4447 ( .C1(n5262), .C2(n4211), .A(n3522), .B(n3521), .ZN(n4627)
         );
  NAND2_X1 U4448 ( .A1(n4622), .A2(n4627), .ZN(n4625) );
  INV_X1 U4449 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U4450 ( .A1(n3806), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4451 ( .A1(n3796), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4452 ( .A1(n3358), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4453 ( .A1(n3797), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3523) );
  NAND4_X1 U4454 ( .A1(n3526), .A2(n3525), .A3(n3524), .A4(n3523), .ZN(n3533)
         );
  AOI22_X1 U4455 ( .A1(n3795), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4456 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n3804), .B1(n4339), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4457 ( .A1(n3247), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4458 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3798), .B1(n3775), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3527) );
  NAND4_X1 U4459 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3532)
         );
  OAI21_X1 U4460 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3534) );
  OAI21_X1 U4461 ( .B1(n4722), .B2(n3689), .A(n3534), .ZN(n3537) );
  XNOR2_X1 U4462 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3538), .ZN(n5250)
         );
  NOR2_X1 U4463 ( .A1(n5250), .A2(n4211), .ZN(n3536) );
  AOI211_X1 U4464 ( .C1(n3763), .C2(EAX_REG_15__SCAN_IN), .A(n3537), .B(n3536), 
        .ZN(n4653) );
  XOR2_X1 U4465 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3551), .Z(n5244) );
  AOI22_X1 U4466 ( .A1(n3303), .A2(EAX_REG_16__SCAN_IN), .B1(n4207), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4467 ( .A1(n3804), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4468 ( .A1(n3247), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4469 ( .A1(n3794), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4470 ( .A1(n3358), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4471 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3548)
         );
  AOI22_X1 U4472 ( .A1(n3806), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4473 ( .A1(n3798), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4474 ( .A1(n3795), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4475 ( .A1(n4339), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4476 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3547)
         );
  OAI21_X1 U4477 ( .B1(n3548), .B2(n3547), .A(n2981), .ZN(n3549) );
  OAI211_X1 U4478 ( .C1(n5244), .C2(n4211), .A(n3550), .B(n3549), .ZN(n4695)
         );
  OAI21_X1 U4479 ( .B1(n3552), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n3566), 
        .ZN(n5238) );
  AOI22_X1 U4480 ( .A1(n3303), .A2(EAX_REG_17__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4481 ( .A1(n3358), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4482 ( .A1(n4339), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4483 ( .A1(n3796), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4484 ( .A1(n3795), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4485 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3562)
         );
  AOI22_X1 U4486 ( .A1(n3798), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4487 ( .A1(n3247), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4488 ( .A1(n3806), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4489 ( .A1(n3804), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3557) );
  NAND4_X1 U4490 ( .A1(n3560), .A2(n3559), .A3(n3558), .A4(n3557), .ZN(n3561)
         );
  OAI21_X1 U4491 ( .B1(n3562), .B2(n3561), .A(n2981), .ZN(n3563) );
  NAND3_X1 U4492 ( .A1(n4211), .A2(n3564), .A3(n3563), .ZN(n3565) );
  OAI21_X1 U4493 ( .B1(n4211), .B2(n5238), .A(n3565), .ZN(n5147) );
  INV_X1 U4494 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6339) );
  AOI21_X1 U4495 ( .B1(n6339), .B2(n3566), .A(n3581), .ZN(n5227) );
  AOI22_X1 U4496 ( .A1(n3303), .A2(EAX_REG_18__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4497 ( .A1(n3796), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4498 ( .A1(n3798), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4499 ( .A1(n3795), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4500 ( .A1(n4339), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4501 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3578)
         );
  INV_X1 U4502 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3571) );
  NOR2_X1 U4503 ( .A1(n3280), .A2(n3571), .ZN(n3572) );
  AOI211_X1 U4504 ( .C1(INSTQUEUE_REG_9__2__SCAN_IN), .C2(n3799), .A(n3826), 
        .B(n3572), .ZN(n3576) );
  AOI22_X1 U4505 ( .A1(n3806), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4506 ( .A1(n3794), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4507 ( .A1(n3804), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4508 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  OR2_X1 U4509 ( .A1(n2981), .A2(n3826), .ZN(n3640) );
  OAI21_X1 U4510 ( .B1(n3578), .B2(n3577), .A(n3640), .ZN(n3579) );
  AOI22_X1 U4511 ( .A1(n3826), .A2(n5227), .B1(n3580), .B2(n3579), .ZN(n4729)
         );
  OAI21_X1 U4512 ( .B1(n3581), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3611), 
        .ZN(n5136) );
  AOI22_X1 U4513 ( .A1(n3303), .A2(EAX_REG_19__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4514 ( .A1(n3804), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4515 ( .A1(n3797), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4516 ( .A1(n3806), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4517 ( .A1(n3775), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4518 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3591)
         );
  AOI22_X1 U4519 ( .A1(n3795), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4520 ( .A1(n3798), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4521 ( .A1(n3796), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4522 ( .A1(n3794), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4523 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3590)
         );
  OAI21_X1 U4524 ( .B1(n3591), .B2(n3590), .A(n2981), .ZN(n3592) );
  NAND3_X1 U4525 ( .A1(n4211), .A2(n3593), .A3(n3592), .ZN(n3594) );
  OAI21_X1 U4526 ( .B1(n4211), .B2(n5136), .A(n3594), .ZN(n4832) );
  XNOR2_X1 U4527 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3611), .ZN(n5069)
         );
  AOI22_X1 U4528 ( .A1(n3303), .A2(EAX_REG_20__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4529 ( .A1(n3795), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4530 ( .A1(n3798), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3804), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4531 ( .A1(n3247), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4532 ( .A1(n3796), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4533 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3607)
         );
  INV_X1 U4534 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3599) );
  OAI21_X1 U4535 ( .B1(n3600), .B2(n3599), .A(n4211), .ZN(n3601) );
  AOI21_X1 U4536 ( .B1(n3797), .B2(INSTQUEUE_REG_7__4__SCAN_IN), .A(n3601), 
        .ZN(n3605) );
  AOI22_X1 U4537 ( .A1(n3775), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4538 ( .A1(n3806), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4539 ( .A1(n4339), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4540 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3606)
         );
  OAI21_X1 U4541 ( .B1(n3607), .B2(n3606), .A(n3640), .ZN(n3608) );
  AOI22_X1 U4542 ( .A1(n3826), .A2(n5069), .B1(n3609), .B2(n3608), .ZN(n4738)
         );
  NAND2_X1 U4543 ( .A1(n4737), .A2(n4738), .ZN(n4826) );
  INV_X1 U4544 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3610) );
  INV_X1 U4545 ( .A(n3628), .ZN(n3627) );
  OR2_X1 U4546 ( .A1(n3612), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3613)
         );
  NAND2_X1 U4547 ( .A1(n3627), .A2(n3613), .ZN(n5129) );
  INV_X1 U4548 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U4549 ( .A1(n3795), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4550 ( .A1(n3808), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4551 ( .A1(n3805), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4552 ( .A1(n3797), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3614) );
  NAND4_X1 U4553 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(n3623)
         );
  AOI22_X1 U4554 ( .A1(n3798), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3804), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4555 ( .A1(n3796), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4556 ( .A1(n4339), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4557 ( .A1(n3806), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4558 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3622)
         );
  OAI21_X1 U4559 ( .B1(n3623), .B2(n3622), .A(n2981), .ZN(n3625) );
  OAI21_X1 U4560 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6026), .A(n5766), 
        .ZN(n3624) );
  OAI211_X1 U4561 ( .C1(n4304), .C2(n3821), .A(n3625), .B(n3624), .ZN(n3626)
         );
  OAI21_X1 U4562 ( .B1(n5129), .B2(n4211), .A(n3626), .ZN(n4825) );
  INV_X1 U4563 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U4564 ( .A1(n3627), .A2(n6412), .ZN(n3629) );
  AND2_X1 U4565 ( .A1(n3629), .A2(n3646), .ZN(n5052) );
  AOI22_X1 U4566 ( .A1(n3763), .A2(EAX_REG_22__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4567 ( .A1(n3796), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4568 ( .A1(n3804), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4569 ( .A1(n3798), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3795), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4570 ( .A1(n3808), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3630) );
  NAND4_X1 U4571 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3642)
         );
  AOI22_X1 U4572 ( .A1(n3806), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4573 ( .A1(n3358), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4574 ( .A1(n3805), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4575 ( .A1(n3807), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3635) );
  NAND2_X1 U4576 ( .A1(n3799), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3634) );
  AND3_X1 U4577 ( .A1(n3635), .A2(n3634), .A3(n4211), .ZN(n3636) );
  NAND4_X1 U4578 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3641)
         );
  OAI21_X1 U4579 ( .B1(n3642), .B2(n3641), .A(n3640), .ZN(n3643) );
  AOI22_X1 U4580 ( .A1(n5052), .A2(n3826), .B1(n3644), .B2(n3643), .ZN(n4820)
         );
  INV_X1 U4581 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3645) );
  AND2_X1 U4582 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  OR2_X1 U4583 ( .A1(n3647), .A2(n3675), .ZN(n5042) );
  AOI22_X1 U4584 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n3796), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4585 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3808), .B1(n4339), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4586 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3798), .B1(n3797), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4587 ( .A1(n3804), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4588 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3657)
         );
  AOI22_X1 U4589 ( .A1(n3806), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4590 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n3358), .B1(n3774), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4591 ( .A1(n3805), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3653) );
  INV_X1 U4592 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6446) );
  AOI22_X1 U4593 ( .A1(n3795), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3652) );
  NAND4_X1 U4594 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3656)
         );
  OR2_X1 U4595 ( .A1(n3657), .A2(n3656), .ZN(n3669) );
  AOI22_X1 U4596 ( .A1(n3796), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4597 ( .A1(n3808), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4598 ( .A1(n3798), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4599 ( .A1(n3804), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3658) );
  NAND4_X1 U4600 ( .A1(n3661), .A2(n3660), .A3(n3659), .A4(n3658), .ZN(n3667)
         );
  AOI22_X1 U4601 ( .A1(n3806), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4602 ( .A1(n3358), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4603 ( .A1(n3805), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4604 ( .A1(n3795), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4605 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3666)
         );
  OR2_X1 U4606 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  NAND2_X1 U4607 ( .A1(n3669), .A2(n3668), .ZN(n3703) );
  OAI211_X1 U4608 ( .C1(n3669), .C2(n3668), .A(n2981), .B(n3703), .ZN(n3672)
         );
  AOI21_X1 U4609 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5766), .A(n3826), 
        .ZN(n3671) );
  NAND2_X1 U4610 ( .A1(n3763), .A2(EAX_REG_23__SCAN_IN), .ZN(n3670) );
  NAND3_X1 U4611 ( .A1(n3672), .A2(n3671), .A3(n3670), .ZN(n3673) );
  OAI21_X1 U4612 ( .B1(n5042), .B2(n4211), .A(n3673), .ZN(n3674) );
  INV_X1 U4613 ( .A(n3674), .ZN(n4764) );
  NOR2_X1 U4614 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3676)
         );
  OR2_X1 U4615 ( .A1(n3692), .A2(n3676), .ZN(n4266) );
  INV_X1 U4616 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6426) );
  AOI22_X1 U4617 ( .A1(n3796), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3798), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4618 ( .A1(n3806), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4619 ( .A1(n3358), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4620 ( .A1(n3805), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3677) );
  NAND4_X1 U4621 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3686)
         );
  AOI22_X1 U4622 ( .A1(n3804), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4623 ( .A1(n4339), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4624 ( .A1(n3794), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4625 ( .A1(n3795), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4626 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3685)
         );
  NOR2_X1 U4627 ( .A1(n3686), .A2(n3685), .ZN(n3704) );
  AOI21_X1 U4628 ( .B1(n3704), .B2(n3703), .A(n3823), .ZN(n3687) );
  OAI21_X1 U4629 ( .B1(n3704), .B2(n3703), .A(n3687), .ZN(n3688) );
  OAI21_X1 U4630 ( .B1(n6426), .B2(n3689), .A(n3688), .ZN(n3690) );
  AOI21_X1 U4631 ( .B1(n3763), .B2(EAX_REG_24__SCAN_IN), .A(n3690), .ZN(n3691)
         );
  OAI21_X1 U4632 ( .B1(n5036), .B2(n4211), .A(n3691), .ZN(n4264) );
  OAI21_X1 U4633 ( .B1(n3692), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n3742), 
        .ZN(n5124) );
  AOI22_X1 U4634 ( .A1(n3796), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4635 ( .A1(n3808), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4636 ( .A1(n3798), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4637 ( .A1(n3804), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4638 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3702)
         );
  AOI22_X1 U4639 ( .A1(n3806), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4640 ( .A1(n3358), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4641 ( .A1(n3805), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4642 ( .A1(n3795), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4643 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3701)
         );
  OR2_X1 U4644 ( .A1(n3702), .A2(n3701), .ZN(n3708) );
  NOR2_X1 U4645 ( .A1(n3704), .A2(n3703), .ZN(n3709) );
  XNOR2_X1 U4646 ( .A(n3708), .B(n3709), .ZN(n3706) );
  AOI22_X1 U4647 ( .A1(n3763), .A2(EAX_REG_25__SCAN_IN), .B1(n5766), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3705) );
  OAI21_X1 U4648 ( .B1(n3823), .B2(n3706), .A(n3705), .ZN(n3707) );
  AOI22_X1 U4649 ( .A1(n3826), .A2(n5124), .B1(n3707), .B2(n4211), .ZN(n4805)
         );
  NAND2_X1 U4650 ( .A1(n3709), .A2(n3708), .ZN(n3726) );
  AOI22_X1 U4651 ( .A1(n3798), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4652 ( .A1(n3804), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4653 ( .A1(n3794), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4654 ( .A1(n3775), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3710) );
  NAND4_X1 U4655 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3719)
         );
  AOI22_X1 U4656 ( .A1(n3795), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3358), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4657 ( .A1(n3806), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3796), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4658 ( .A1(n4339), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4659 ( .A1(n3231), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4660 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3718)
         );
  NOR2_X1 U4661 ( .A1(n3719), .A2(n3718), .ZN(n3727) );
  XOR2_X1 U4662 ( .A(n3726), .B(n3727), .Z(n3720) );
  NAND2_X1 U4663 ( .A1(n3720), .A2(n2981), .ZN(n3725) );
  OAI21_X1 U4664 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6026), .A(n5766), 
        .ZN(n3721) );
  INV_X1 U4665 ( .A(n3721), .ZN(n3722) );
  AOI21_X1 U4666 ( .B1(n3763), .B2(EAX_REG_26__SCAN_IN), .A(n3722), .ZN(n3724)
         );
  XNOR2_X1 U4667 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3742), .ZN(n5115)
         );
  AOI21_X1 U4668 ( .B1(n3725), .B2(n3724), .A(n3723), .ZN(n4748) );
  NOR2_X1 U4669 ( .A1(n3727), .A2(n3726), .ZN(n3749) );
  AOI22_X1 U4670 ( .A1(n3796), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4671 ( .A1(n3808), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4672 ( .A1(n3798), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4673 ( .A1(n3804), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3728) );
  NAND4_X1 U4674 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3737)
         );
  AOI22_X1 U4675 ( .A1(n3806), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4676 ( .A1(n3358), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4677 ( .A1(n3805), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4678 ( .A1(n3795), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4679 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3736)
         );
  OR2_X1 U4680 ( .A1(n3737), .A2(n3736), .ZN(n3748) );
  INV_X1 U4681 ( .A(n3748), .ZN(n3738) );
  XNOR2_X1 U4682 ( .A(n3749), .B(n3738), .ZN(n3739) );
  NAND2_X1 U4683 ( .A1(n3739), .A2(n2981), .ZN(n3747) );
  NAND2_X1 U4684 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5766), .ZN(n3740)
         );
  NAND2_X1 U4685 ( .A1(n3740), .A2(n4211), .ZN(n3741) );
  AOI21_X1 U4686 ( .B1(n3763), .B2(EAX_REG_27__SCAN_IN), .A(n3741), .ZN(n3746)
         );
  INV_X1 U4687 ( .A(n3742), .ZN(n3743) );
  OAI21_X1 U4688 ( .B1(n3744), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n3786), 
        .ZN(n5013) );
  NOR2_X1 U4689 ( .A1(n5013), .A2(n4211), .ZN(n3745) );
  AOI21_X1 U4690 ( .B1(n3747), .B2(n3746), .A(n3745), .ZN(n4802) );
  NAND2_X1 U4691 ( .A1(n4746), .A2(n4802), .ZN(n4020) );
  NAND2_X1 U4692 ( .A1(n3749), .A2(n3748), .ZN(n3768) );
  AOI22_X1 U4693 ( .A1(n3806), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3808), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4694 ( .A1(n4339), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4695 ( .A1(n3231), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4696 ( .A1(n3795), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4697 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4698 ( .A1(n3804), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4699 ( .A1(n3796), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4700 ( .A1(n3358), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4701 ( .A1(n3798), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4702 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4703 ( .A1(n3759), .A2(n3758), .ZN(n3769) );
  XOR2_X1 U4704 ( .A(n3768), .B(n3769), .Z(n3760) );
  NAND2_X1 U4705 ( .A1(n3760), .A2(n2981), .ZN(n3765) );
  NAND2_X1 U4706 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5766), .ZN(n3761)
         );
  NAND2_X1 U4707 ( .A1(n3761), .A2(n4211), .ZN(n3762) );
  AOI21_X1 U4708 ( .B1(n3763), .B2(EAX_REG_28__SCAN_IN), .A(n3762), .ZN(n3764)
         );
  NAND2_X1 U4709 ( .A1(n3765), .A2(n3764), .ZN(n3767) );
  XNOR2_X1 U4710 ( .A(n3786), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5001)
         );
  NAND2_X1 U4711 ( .A1(n5001), .A2(n3826), .ZN(n3766) );
  NAND2_X1 U4712 ( .A1(n3767), .A2(n3766), .ZN(n4022) );
  NOR2_X2 U4713 ( .A1(n4020), .A2(n4022), .ZN(n4021) );
  NOR2_X1 U4714 ( .A1(n3769), .A2(n3768), .ZN(n3816) );
  AOI22_X1 U4715 ( .A1(n3796), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4716 ( .A1(n3808), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4339), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4717 ( .A1(n3798), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4718 ( .A1(n3804), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4719 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3781)
         );
  AOI22_X1 U4720 ( .A1(n3806), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4721 ( .A1(n3358), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4722 ( .A1(n3805), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3775), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4723 ( .A1(n3795), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4724 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  OR2_X1 U4725 ( .A1(n3781), .A2(n3780), .ZN(n3815) );
  INV_X1 U4726 ( .A(n3815), .ZN(n3782) );
  XNOR2_X1 U4727 ( .A(n3816), .B(n3782), .ZN(n3783) );
  NAND2_X1 U4728 ( .A1(n3783), .A2(n2981), .ZN(n3793) );
  NAND2_X1 U4729 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n5766), .ZN(n3784)
         );
  NAND2_X1 U4730 ( .A1(n3784), .A2(n4211), .ZN(n3785) );
  AOI21_X1 U4731 ( .B1(n3763), .B2(EAX_REG_29__SCAN_IN), .A(n3785), .ZN(n3792)
         );
  INV_X1 U4732 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U4733 ( .A1(n3787), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4216)
         );
  INV_X1 U4734 ( .A(n3787), .ZN(n3789) );
  INV_X1 U4735 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4736 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  NAND2_X1 U4737 ( .A1(n4216), .A2(n3790), .ZN(n4995) );
  NOR2_X1 U4738 ( .A1(n4995), .A2(n4211), .ZN(n3791) );
  AOI21_X1 U4739 ( .B1(n3793), .B2(n3792), .A(n3791), .ZN(n4287) );
  XNOR2_X1 U4740 ( .A(n4216), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4988)
         );
  AOI22_X1 U4741 ( .A1(n3795), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n3796), .B1(n4339), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4743 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n3798), .B1(n3797), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4744 ( .A1(n3775), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4745 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3814)
         );
  AOI22_X1 U4746 ( .A1(n3804), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4747 ( .A1(n3806), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3805), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4748 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n3358), .B1(n3774), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4749 ( .A1(n3808), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3807), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4750 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  NOR2_X1 U4751 ( .A1(n3814), .A2(n3813), .ZN(n3818) );
  NAND2_X1 U4752 ( .A1(n3816), .A2(n3815), .ZN(n3817) );
  XOR2_X1 U4753 ( .A(n3818), .B(n3817), .Z(n3824) );
  INV_X1 U4754 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3820) );
  OAI21_X1 U4755 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6026), .A(n5766), 
        .ZN(n3819) );
  OAI21_X1 U4756 ( .B1(n3821), .B2(n3820), .A(n3819), .ZN(n3822) );
  AOI21_X1 U4757 ( .B1(n3824), .B2(n2981), .A(n3822), .ZN(n3825) );
  AOI21_X1 U4758 ( .B1(n3826), .B2(n4988), .A(n3825), .ZN(n4205) );
  XNOR2_X1 U4759 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4760 ( .A1(n3841), .A2(n3842), .ZN(n3840) );
  NAND2_X1 U4761 ( .A1(n6140), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4762 ( .A1(n3840), .A2(n3829), .ZN(n3859) );
  XNOR2_X1 U4763 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4764 ( .A1(n3859), .A2(n3857), .ZN(n3831) );
  NAND2_X1 U4765 ( .A1(n6145), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4766 ( .A1(n3831), .A2(n3830), .ZN(n3864) );
  XNOR2_X1 U4767 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4768 ( .A1(n3864), .A2(n3862), .ZN(n3833) );
  NAND2_X1 U4769 ( .A1(n6284), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4770 ( .A1(n3833), .A2(n3832), .ZN(n3837) );
  NAND2_X1 U4771 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5200), .ZN(n3835) );
  NAND2_X1 U4772 ( .A1(n3861), .A2(n3894), .ZN(n3879) );
  AOI21_X1 U4773 ( .B1(n3861), .B2(n3180), .A(n3839), .ZN(n3848) );
  OAI21_X1 U4774 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3847) );
  NOR3_X1 U4775 ( .A1(n3848), .A2(n6180), .A3(n3847), .ZN(n3855) );
  XNOR2_X1 U4776 ( .A(n3312), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3846)
         );
  OAI21_X1 U4777 ( .B1(n4003), .B2(n3846), .A(n3843), .ZN(n3845) );
  NAND2_X1 U4778 ( .A1(n3844), .A2(n4149), .ZN(n3856) );
  NAND2_X1 U4779 ( .A1(n3845), .A2(n3856), .ZN(n3850) );
  INV_X1 U4780 ( .A(n3850), .ZN(n3853) );
  INV_X1 U4781 ( .A(n3847), .ZN(n3895) );
  INV_X1 U4782 ( .A(n3846), .ZN(n3851) );
  NAND2_X1 U4783 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  NAND4_X1 U4784 ( .A1(n3861), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3852)
         );
  AOI22_X1 U4785 ( .A1(n3853), .A2(n3895), .B1(n3876), .B2(n3852), .ZN(n3854)
         );
  NOR2_X1 U4786 ( .A1(n3855), .A2(n3854), .ZN(n3868) );
  INV_X1 U4787 ( .A(n3856), .ZN(n3860) );
  INV_X1 U4788 ( .A(n3857), .ZN(n3858) );
  XNOR2_X1 U4789 ( .A(n3859), .B(n3858), .ZN(n3896) );
  NAND3_X1 U4790 ( .A1(n3860), .A2(n3896), .A3(n3861), .ZN(n3867) );
  AOI21_X1 U4791 ( .B1(n3896), .B2(n3861), .A(n3860), .ZN(n3866) );
  INV_X1 U4792 ( .A(n3862), .ZN(n3863) );
  XNOR2_X1 U4793 ( .A(n3864), .B(n3863), .ZN(n3897) );
  INV_X1 U4794 ( .A(n3897), .ZN(n3865) );
  AOI211_X1 U4795 ( .C1(n3868), .C2(n3867), .A(n3866), .B(n3865), .ZN(n3874)
         );
  INV_X1 U4796 ( .A(n3868), .ZN(n3870) );
  INV_X1 U4797 ( .A(n3896), .ZN(n3869) );
  NAND3_X1 U4798 ( .A1(n3872), .A2(n3870), .A3(n3869), .ZN(n3871) );
  OAI21_X1 U4799 ( .B1(n3897), .B2(n3876), .A(n3871), .ZN(n3873) );
  OAI22_X1 U4800 ( .A1(n3874), .A2(n3873), .B1(n3872), .B2(n3900), .ZN(n3875)
         );
  OAI21_X1 U4801 ( .B1(n3900), .B2(n3876), .A(n3875), .ZN(n3877) );
  AOI21_X1 U4802 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6180), .A(n3877), 
        .ZN(n3878) );
  NAND2_X1 U4803 ( .A1(n3879), .A2(n3878), .ZN(n3882) );
  NAND2_X1 U4804 ( .A1(n3880), .A2(n3894), .ZN(n3881) );
  INV_X1 U4805 ( .A(READY_N), .ZN(n4384) );
  AND2_X1 U4806 ( .A1(n3180), .A2(n4384), .ZN(n3884) );
  AND2_X1 U4807 ( .A1(n3886), .A2(n3885), .ZN(n4032) );
  NAND2_X1 U4808 ( .A1(n4032), .A2(n2977), .ZN(n6150) );
  INV_X1 U4809 ( .A(n4298), .ZN(n4383) );
  INV_X1 U4810 ( .A(n3888), .ZN(n3893) );
  AND3_X1 U4811 ( .A1(n5619), .A2(n3889), .A3(n6395), .ZN(n3892) );
  INV_X1 U4812 ( .A(n3890), .ZN(n3891) );
  NAND2_X1 U4813 ( .A1(n4201), .A2(n2977), .ZN(n3903) );
  INV_X1 U4814 ( .A(n3894), .ZN(n3899) );
  NAND3_X1 U4815 ( .A1(n3897), .A2(n3896), .A3(n3895), .ZN(n3898) );
  NAND2_X1 U4816 ( .A1(n3899), .A2(n3898), .ZN(n3901) );
  NOR2_X1 U4817 ( .A1(READY_N), .A2(n6153), .ZN(n4037) );
  NAND2_X1 U4818 ( .A1(n4440), .A2(n4037), .ZN(n4333) );
  INV_X1 U4819 ( .A(n6181), .ZN(n6178) );
  OR2_X1 U4820 ( .A1(n4333), .A2(n6178), .ZN(n3902) );
  OAI211_X1 U4821 ( .C1(n6150), .C2(n4383), .A(n3903), .B(n3902), .ZN(n3904)
         );
  INV_X1 U4822 ( .A(n3904), .ZN(n3905) );
  NAND2_X1 U4823 ( .A1(n3906), .A2(n3302), .ZN(n4370) );
  NAND2_X1 U4824 ( .A1(n4200), .A2(n5397), .ZN(n3911) );
  INV_X2 U4825 ( .A(n4839), .ZN(n5406) );
  INV_X1 U4826 ( .A(n3302), .ZN(n4840) );
  NOR3_X1 U4827 ( .A1(n5406), .A2(n4840), .A3(n4477), .ZN(n3907) );
  AOI22_X1 U4828 ( .A1(n5407), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5406), .ZN(n3908) );
  NAND2_X1 U4829 ( .A1(n3911), .A2(n3910), .ZN(U2861) );
  NAND2_X1 U4830 ( .A1(n3917), .A2(n3912), .ZN(n3922) );
  OAI211_X1 U4831 ( .C1(n3917), .C2(n3912), .A(n4244), .B(n3922), .ZN(n3914)
         );
  AND3_X1 U4832 ( .A1(n3914), .A2(n3913), .A3(n4477), .ZN(n3915) );
  NAND2_X1 U4833 ( .A1(n3916), .A2(n3915), .ZN(n5520) );
  INV_X1 U4834 ( .A(n2978), .ZN(n3970) );
  INV_X1 U4835 ( .A(n4244), .ZN(n6309) );
  OAI21_X1 U4836 ( .B1(n6309), .B2(n3917), .A(n2996), .ZN(n3918) );
  INV_X1 U4837 ( .A(n3918), .ZN(n3919) );
  NAND2_X1 U4838 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5527)
         );
  XNOR2_X1 U4839 ( .A(n5527), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5519)
         );
  NAND2_X1 U4840 ( .A1(n5520), .A2(n5519), .ZN(n5518) );
  INV_X1 U4841 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5587) );
  OR2_X1 U4842 ( .A1(n5527), .A2(n5587), .ZN(n3921) );
  NAND2_X1 U4843 ( .A1(n5518), .A2(n3921), .ZN(n5511) );
  NAND2_X1 U4844 ( .A1(n4451), .A2(n2978), .ZN(n3926) );
  NAND2_X1 U4845 ( .A1(n3922), .A2(n3923), .ZN(n3930) );
  OAI21_X1 U4846 ( .B1(n3923), .B2(n3922), .A(n3930), .ZN(n3924) );
  AOI21_X1 U4847 ( .B1(n3924), .B2(n4244), .A(n4160), .ZN(n3925) );
  NAND2_X1 U4848 ( .A1(n3927), .A2(n5510), .ZN(n3929) );
  NAND2_X1 U4849 ( .A1(n5511), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3928)
         );
  NAND2_X1 U4850 ( .A1(n3929), .A2(n3928), .ZN(n4399) );
  NAND2_X1 U4851 ( .A1(n3930), .A2(n3931), .ZN(n3944) );
  OAI211_X1 U4852 ( .C1(n3931), .C2(n3930), .A(n3944), .B(n4244), .ZN(n3932)
         );
  OAI21_X2 U4853 ( .B1(n3933), .B2(n3970), .A(n3932), .ZN(n3934) );
  INV_X1 U4854 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U4855 ( .A1(n4399), .A2(n4398), .ZN(n3936) );
  NAND2_X1 U4856 ( .A1(n3934), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3935)
         );
  INV_X1 U4857 ( .A(n3937), .ZN(n3943) );
  XNOR2_X1 U4858 ( .A(n3944), .B(n3943), .ZN(n3938) );
  INV_X1 U4859 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4067) );
  XNOR2_X1 U4860 ( .A(n3940), .B(n4067), .ZN(n4459) );
  NAND2_X1 U4861 ( .A1(n4458), .A2(n4459), .ZN(n3942) );
  NAND2_X1 U4862 ( .A1(n3940), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3941)
         );
  NAND2_X1 U4863 ( .A1(n3942), .A2(n3941), .ZN(n4968) );
  NOR2_X1 U4864 ( .A1(n3944), .A2(n3943), .ZN(n3946) );
  NAND2_X1 U4865 ( .A1(n3946), .A2(n3945), .ZN(n3960) );
  OAI211_X1 U4866 ( .C1(n3946), .C2(n3945), .A(n3960), .B(n4244), .ZN(n3947)
         );
  INV_X1 U4867 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3949) );
  XNOR2_X1 U4868 ( .A(n3950), .B(n3949), .ZN(n4967) );
  NAND2_X1 U4869 ( .A1(n4968), .A2(n4967), .ZN(n3952) );
  NAND2_X1 U4870 ( .A1(n3950), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3951)
         );
  NAND2_X1 U4871 ( .A1(n3952), .A2(n3951), .ZN(n4503) );
  NAND3_X1 U4872 ( .A1(n3969), .A2(n2978), .A3(n3953), .ZN(n3956) );
  XNOR2_X1 U4873 ( .A(n3960), .B(n3961), .ZN(n3954) );
  NAND2_X1 U4874 ( .A1(n3954), .A2(n4244), .ZN(n3955) );
  NAND2_X1 U4875 ( .A1(n3956), .A2(n3955), .ZN(n3957) );
  INV_X1 U4876 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4513) );
  XNOR2_X1 U4877 ( .A(n3957), .B(n4513), .ZN(n4504) );
  NAND2_X1 U4878 ( .A1(n4503), .A2(n4504), .ZN(n3959) );
  NAND2_X1 U4879 ( .A1(n3957), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3958)
         );
  NAND2_X1 U4880 ( .A1(n3959), .A2(n3958), .ZN(n4464) );
  INV_X1 U4881 ( .A(n3960), .ZN(n3962) );
  NAND2_X1 U4882 ( .A1(n3962), .A2(n3961), .ZN(n3975) );
  XNOR2_X1 U4883 ( .A(n3975), .B(n3973), .ZN(n3963) );
  NAND2_X1 U4884 ( .A1(n3963), .A2(n4244), .ZN(n3964) );
  INV_X1 U4885 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6462) );
  XNOR2_X1 U4886 ( .A(n3966), .B(n6462), .ZN(n4463) );
  NAND2_X1 U4887 ( .A1(n4464), .A2(n4463), .ZN(n3968) );
  NAND2_X1 U4888 ( .A1(n3966), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3967)
         );
  NOR2_X1 U4889 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  NAND2_X1 U4890 ( .A1(n4244), .A2(n3973), .ZN(n3974) );
  OR2_X1 U4891 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  NAND2_X1 U4892 ( .A1(n3980), .A2(n3976), .ZN(n3977) );
  INV_X1 U4893 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4078) );
  NAND2_X1 U4894 ( .A1(n4574), .A2(n4575), .ZN(n3979) );
  NAND2_X1 U4895 ( .A1(n3977), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3978)
         );
  INV_X1 U4896 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U4897 ( .A1(n3980), .A2(n5565), .ZN(n3982) );
  INV_X1 U4898 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6398) );
  AND2_X1 U4899 ( .A1(n3980), .A2(n6398), .ZN(n5479) );
  OR2_X2 U4900 ( .A1(n5477), .A2(n5479), .ZN(n3983) );
  OR2_X1 U4901 ( .A1(n3980), .A2(n6398), .ZN(n5478) );
  INV_X1 U4902 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4643) );
  OR2_X1 U4903 ( .A1(n3980), .A2(n4643), .ZN(n5471) );
  INV_X1 U4904 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3985) );
  NOR2_X1 U4905 ( .A1(n3980), .A2(n3985), .ZN(n4637) );
  NAND2_X1 U4906 ( .A1(n3980), .A2(n3985), .ZN(n4638) );
  XNOR2_X1 U4907 ( .A(n3980), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4658)
         );
  INV_X1 U4908 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4166) );
  INV_X1 U4909 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U4910 ( .A1(n3980), .A2(n4705), .ZN(n3986) );
  INV_X1 U4911 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4960) );
  INV_X1 U4912 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U4913 ( .A1(n3980), .A2(n3987), .ZN(n3988) );
  NAND2_X1 U4914 ( .A1(n4953), .A2(n3988), .ZN(n5141) );
  NOR3_X1 U4915 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n3989) );
  NAND2_X1 U4916 ( .A1(n5141), .A2(n3989), .ZN(n3990) );
  NAND2_X1 U4917 ( .A1(n3990), .A2(n3981), .ZN(n3993) );
  INV_X1 U4918 ( .A(n5141), .ZN(n3991) );
  NAND2_X1 U4919 ( .A1(n3991), .A2(n2995), .ZN(n3992) );
  NOR2_X1 U4920 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4944) );
  NOR2_X1 U4921 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3994) );
  INV_X1 U4922 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6354) );
  INV_X1 U4923 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6455) );
  AND4_X1 U4924 ( .A1(n4944), .A2(n3994), .A3(n6354), .A4(n6455), .ZN(n3995)
         );
  NOR2_X1 U4925 ( .A1(n3980), .A2(n3995), .ZN(n3998) );
  AND2_X1 U4926 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4945) );
  AND2_X1 U4927 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3996) );
  AND2_X1 U4928 ( .A1(n4945), .A2(n3996), .ZN(n4927) );
  AND2_X1 U4929 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U4930 ( .A1(n4927), .A2(n4187), .ZN(n4190) );
  NAND2_X1 U4931 ( .A1(n3980), .A2(n4190), .ZN(n3997) );
  XNOR2_X1 U4932 ( .A(n3980), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5120)
         );
  INV_X1 U4933 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5167) );
  INV_X1 U4934 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4919) );
  NOR2_X1 U4935 ( .A1(n3981), .A2(n4919), .ZN(n4912) );
  NAND2_X1 U4936 ( .A1(n3999), .A2(n4912), .ZN(n4859) );
  NAND2_X1 U4937 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4192) );
  NOR2_X2 U4938 ( .A1(n4859), .A2(n4192), .ZN(n4850) );
  NOR2_X1 U4939 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4911)
         );
  NOR2_X1 U4940 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U4941 ( .A1(n4911), .A2(n4896), .ZN(n4848) );
  NAND2_X1 U4942 ( .A1(n4000), .A2(n4001), .ZN(n4269) );
  AOI21_X1 U4943 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4850), .A(n4270), 
        .ZN(n4002) );
  XNOR2_X1 U4944 ( .A(n4002), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4051)
         );
  AND2_X1 U4945 ( .A1(n4003), .A2(n4032), .ZN(n6151) );
  NAND2_X1 U4946 ( .A1(n4051), .A2(n5533), .ZN(n4013) );
  NAND3_X1 U4947 ( .A1(n6180), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6192) );
  INV_X1 U4948 ( .A(n6192), .ZN(n4004) );
  NOR2_X2 U4949 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6289) );
  AND2_X2 U4950 ( .A1(n4004), .A2(n6289), .ZN(n5631) );
  INV_X1 U4951 ( .A(n5631), .ZN(n6076) );
  NAND2_X1 U4952 ( .A1(n6275), .A2(n4005), .ZN(n6306) );
  AND2_X1 U4953 ( .A1(n6306), .A2(n6180), .ZN(n4006) );
  INV_X1 U4954 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U4955 ( .A1(n6180), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U4956 ( .A1(n6026), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4007) );
  AND2_X1 U4957 ( .A1(n4008), .A2(n4007), .ZN(n5531) );
  INV_X1 U4958 ( .A(n5531), .ZN(n4009) );
  NAND2_X1 U4959 ( .A1(n5483), .A2(n4988), .ZN(n4010) );
  NAND2_X1 U4960 ( .A1(n6289), .A2(n6395), .ZN(n6316) );
  INV_X2 U4961 ( .A(n5599), .ZN(n5585) );
  NAND2_X1 U4962 ( .A1(n5585), .A2(REIP_REG_30__SCAN_IN), .ZN(n4193) );
  OAI211_X1 U4963 ( .C1(n5530), .C2(n4011), .A(n4010), .B(n4193), .ZN(n4012)
         );
  AND2_X1 U4964 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4014)
         );
  AND2_X1 U4965 ( .A1(n4911), .A2(n5167), .ZN(n4016) );
  NAND2_X1 U4966 ( .A1(n4015), .A2(n4016), .ZN(n4858) );
  AND2_X1 U4967 ( .A1(n4919), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4017)
         );
  INV_X1 U4968 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4139) );
  XNOR2_X1 U4969 ( .A(n4019), .B(n4139), .ZN(n4893) );
  NAND2_X1 U4970 ( .A1(n4893), .A2(n5533), .ZN(n4028) );
  AOI21_X1 U4971 ( .B1(n4022), .B2(n4020), .A(n4021), .ZN(n4023) );
  NAND2_X1 U4972 ( .A1(n5483), .A2(n5001), .ZN(n4024) );
  NAND2_X1 U4973 ( .A1(n5585), .A2(REIP_REG_28__SCAN_IN), .ZN(n4894) );
  OAI211_X1 U4974 ( .C1(n5530), .C2(n4025), .A(n4024), .B(n4894), .ZN(n4026)
         );
  NAND2_X1 U4975 ( .A1(n4028), .A2(n4027), .ZN(U2958) );
  INV_X1 U4976 ( .A(n4029), .ZN(n6134) );
  NAND2_X1 U4977 ( .A1(n6134), .A2(n3180), .ZN(n4039) );
  NAND2_X1 U4978 ( .A1(n2978), .A2(n3320), .ZN(n4165) );
  OAI211_X1 U4979 ( .C1(n4031), .C2(n4030), .A(n3843), .B(n4165), .ZN(n4158)
         );
  NAND2_X1 U4980 ( .A1(n4032), .A2(n4158), .ZN(n4034) );
  NAND2_X1 U4981 ( .A1(n4034), .A2(n4033), .ZN(n4164) );
  INV_X1 U4982 ( .A(n4035), .ZN(n4036) );
  INV_X1 U4983 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U4984 ( .A1(n4036), .A2(n6200), .ZN(n6198) );
  INV_X1 U4985 ( .A(n6198), .ZN(n4329) );
  OAI211_X1 U4986 ( .C1(n4149), .C2(n4329), .A(n4492), .B(n4037), .ZN(n4038)
         );
  OAI211_X1 U4987 ( .C1(n6157), .C2(n4039), .A(n4164), .B(n4038), .ZN(n4040)
         );
  NAND2_X1 U4988 ( .A1(n4040), .A2(n6181), .ZN(n4045) );
  NAND2_X1 U4989 ( .A1(n4149), .A2(n6198), .ZN(n4234) );
  NAND2_X1 U4990 ( .A1(n4234), .A2(n4384), .ZN(n4327) );
  INV_X1 U4991 ( .A(n4151), .ZN(n4042) );
  OAI211_X1 U4992 ( .C1(n4041), .C2(n4327), .A(n3843), .B(n4042), .ZN(n4043)
         );
  NAND3_X1 U4993 ( .A1(n4043), .A2(n4298), .A3(n3889), .ZN(n4044) );
  INV_X1 U4994 ( .A(n6151), .ZN(n6162) );
  AND2_X1 U4995 ( .A1(n4146), .A2(n4046), .ZN(n4047) );
  NOR2_X1 U4996 ( .A1(n4440), .A2(n4047), .ZN(n4049) );
  NAND2_X1 U4997 ( .A1(n3828), .A2(n3180), .ZN(n4048) );
  NAND4_X1 U4998 ( .A1(n6162), .A2(n4049), .A3(n4048), .A4(n6150), .ZN(n4050)
         );
  NAND2_X1 U4999 ( .A1(n4051), .A2(n5591), .ZN(n4199) );
  INV_X2 U5000 ( .A(n4058), .ZN(n5207) );
  INV_X1 U5001 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U5002 ( .A1(n5207), .A2(n4053), .ZN(n4054) );
  OAI211_X1 U5003 ( .C1(n4125), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4054), 
        .B(n2945), .ZN(n4055) );
  INV_X1 U5004 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5371) );
  AOI22_X1 U5005 ( .A1(n2945), .A2(n5371), .B1(n2946), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4550) );
  INV_X1 U5006 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U5007 ( .A1(n4065), .A2(n5395), .ZN(n4062) );
  INV_X1 U5008 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U5009 ( .A1(n2946), .A2(n4059), .ZN(n4060) );
  OAI211_X1 U5010 ( .C1(n4231), .C2(EBX_REG_2__SCAN_IN), .A(n4060), .B(n2945), 
        .ZN(n4061) );
  NAND2_X1 U5011 ( .A1(n4062), .A2(n4061), .ZN(n4683) );
  NAND2_X1 U5012 ( .A1(n4682), .A2(n4683), .ZN(n4412) );
  INV_X1 U5013 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U5014 ( .A1(n4136), .A2(n4573), .ZN(n4064) );
  NAND2_X1 U5015 ( .A1(n4052), .A2(EBX_REG_3__SCAN_IN), .ZN(n4063) );
  OAI211_X1 U5016 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n4227), .A(n4064), 
        .B(n4063), .ZN(n4413) );
  NOR2_X2 U5017 ( .A1(n4412), .A2(n4413), .ZN(n4758) );
  INV_X1 U5018 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4066) );
  NAND2_X1 U5019 ( .A1(n4065), .A2(n4066), .ZN(n4070) );
  NAND2_X1 U5020 ( .A1(n2946), .A2(n4067), .ZN(n4068) );
  OAI211_X1 U5021 ( .C1(n4231), .C2(EBX_REG_4__SCAN_IN), .A(n4068), .B(n2945), 
        .ZN(n4069) );
  NAND2_X1 U5022 ( .A1(n4070), .A2(n4069), .ZN(n4759) );
  INV_X1 U5023 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5024 ( .A1(n4136), .A2(n4559), .ZN(n4072) );
  NAND2_X1 U5025 ( .A1(n4052), .A2(EBX_REG_5__SCAN_IN), .ZN(n4071) );
  OAI211_X1 U5026 ( .C1(INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n4227), .A(n4072), 
        .B(n4071), .ZN(n4554) );
  INV_X1 U5027 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U5028 ( .A1(n4065), .A2(n6454), .ZN(n4075) );
  NAND2_X1 U5029 ( .A1(n2946), .A2(n4513), .ZN(n4073) );
  OAI211_X1 U5030 ( .C1(n4231), .C2(EBX_REG_6__SCAN_IN), .A(n4073), .B(n2945), 
        .ZN(n4074) );
  NAND2_X1 U5031 ( .A1(n4075), .A2(n4074), .ZN(n4505) );
  INV_X1 U5032 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5033 ( .A1(n4136), .A2(n4520), .ZN(n4077) );
  NAND2_X1 U5034 ( .A1(n4052), .A2(EBX_REG_7__SCAN_IN), .ZN(n4076) );
  OAI211_X1 U5035 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n4227), .A(n4077), 
        .B(n4076), .ZN(n4469) );
  INV_X1 U5036 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U5037 ( .A1(n4065), .A2(n5315), .ZN(n4081) );
  NAND2_X1 U5038 ( .A1(n2946), .A2(n4078), .ZN(n4079) );
  OAI211_X1 U5039 ( .C1(n4231), .C2(EBX_REG_8__SCAN_IN), .A(n4079), .B(n2945), 
        .ZN(n4080) );
  NAND2_X1 U5040 ( .A1(n4081), .A2(n4080), .ZN(n4566) );
  INV_X1 U5041 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4593) );
  INV_X1 U5042 ( .A(n4227), .ZN(n4551) );
  AOI22_X1 U5043 ( .A1(n4136), .A2(n4593), .B1(n4551), .B2(n5565), .ZN(n4082)
         );
  OAI21_X1 U5044 ( .B1(n2945), .B2(n4593), .A(n4082), .ZN(n4591) );
  INV_X1 U5045 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4083) );
  NAND2_X1 U5046 ( .A1(n4065), .A2(n4083), .ZN(n4086) );
  NAND2_X1 U5047 ( .A1(n4125), .A2(n4231), .ZN(n4128) );
  NAND2_X1 U5048 ( .A1(n4125), .A2(EBX_REG_10__SCAN_IN), .ZN(n4085) );
  NAND2_X1 U5049 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4231), .ZN(n4084) );
  NAND4_X1 U5050 ( .A1(n4086), .A2(n4128), .A3(n4085), .A4(n4084), .ZN(n4588)
         );
  INV_X1 U5051 ( .A(n4136), .ZN(n4107) );
  INV_X1 U5052 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U5053 ( .A1(n5207), .A2(n5390), .ZN(n4087) );
  OAI211_X1 U5054 ( .C1(n4052), .C2(n4643), .A(n4087), .B(n2946), .ZN(n4088)
         );
  OAI21_X1 U5055 ( .B1(n4107), .B2(EBX_REG_11__SCAN_IN), .A(n4088), .ZN(n5285)
         );
  INV_X1 U5056 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U5057 ( .A1(n4065), .A2(n4089), .ZN(n4092) );
  NAND2_X1 U5058 ( .A1(n4125), .A2(EBX_REG_12__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5059 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4231), .ZN(n4090) );
  NAND4_X1 U5060 ( .A1(n4092), .A2(n4128), .A3(n4091), .A4(n4090), .ZN(n4620)
         );
  INV_X1 U5061 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U5062 ( .A1(n5207), .A2(n5388), .ZN(n4093) );
  OAI211_X1 U5063 ( .C1(n4052), .C2(n4166), .A(n4093), .B(n2946), .ZN(n4094)
         );
  OAI21_X1 U5064 ( .B1(n4107), .B2(EBX_REG_13__SCAN_IN), .A(n4094), .ZN(n4667)
         );
  INV_X1 U5065 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4095) );
  NAND2_X1 U5066 ( .A1(n4065), .A2(n4095), .ZN(n4098) );
  NAND2_X1 U5067 ( .A1(n4125), .A2(EBX_REG_14__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U5068 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4231), .ZN(n4096) );
  NAND4_X1 U5069 ( .A1(n4098), .A2(n4128), .A3(n4097), .A4(n4096), .ZN(n4650)
         );
  INV_X1 U5070 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U5071 ( .A1(n5207), .A2(n6378), .ZN(n4099) );
  OAI211_X1 U5072 ( .C1(n4052), .C2(n4960), .A(n4099), .B(n2946), .ZN(n4100)
         );
  OAI21_X1 U5073 ( .B1(n4107), .B2(EBX_REG_15__SCAN_IN), .A(n4100), .ZN(n4714)
         );
  INV_X1 U5074 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U5075 ( .A1(n4065), .A2(n4101), .ZN(n4104) );
  NAND2_X1 U5076 ( .A1(n4125), .A2(EBX_REG_16__SCAN_IN), .ZN(n4103) );
  NAND2_X1 U5077 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4231), .ZN(n4102) );
  NAND4_X1 U5078 ( .A1(n4104), .A2(n4128), .A3(n4103), .A4(n4102), .ZN(n4692)
         );
  INV_X1 U5079 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5183) );
  INV_X1 U5080 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U5081 ( .A1(n5207), .A2(n5381), .ZN(n4105) );
  OAI211_X1 U5082 ( .C1(n4052), .C2(n5183), .A(n4105), .B(n2946), .ZN(n4106)
         );
  OAI21_X1 U5083 ( .B1(n4107), .B2(EBX_REG_17__SCAN_IN), .A(n4106), .ZN(n5192)
         );
  INV_X1 U5084 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U5085 ( .A1(n4065), .A2(n5081), .ZN(n4110) );
  INV_X1 U5086 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5087 ( .A1(n2946), .A2(n4253), .ZN(n4108) );
  OAI211_X1 U5088 ( .C1(n4231), .C2(EBX_REG_19__SCAN_IN), .A(n4108), .B(n2945), 
        .ZN(n4109) );
  NAND2_X1 U5089 ( .A1(n4110), .A2(n4109), .ZN(n4831) );
  NAND2_X1 U5090 ( .A1(n4227), .A2(EBX_REG_18__SCAN_IN), .ZN(n4112) );
  NAND2_X1 U5091 ( .A1(n4231), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U5092 ( .A1(n4112), .A2(n4111), .ZN(n4740) );
  INV_X1 U5093 ( .A(n4740), .ZN(n4113) );
  NAND2_X1 U5094 ( .A1(n4113), .A2(n4052), .ZN(n4756) );
  OAI22_X1 U5095 ( .A1(n4227), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4231), .ZN(n4741) );
  AND2_X1 U5096 ( .A1(n4740), .A2(n2945), .ZN(n4754) );
  INV_X1 U5097 ( .A(EBX_REG_21__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U5098 ( .A1(n4136), .A2(n4828), .ZN(n4117) );
  NAND2_X1 U5099 ( .A1(n4052), .A2(EBX_REG_21__SCAN_IN), .ZN(n4116) );
  OAI211_X1 U5100 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n4227), .A(n4117), .B(n4116), .ZN(n4822) );
  INV_X1 U5101 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U5102 ( .A1(n4065), .A2(n4118), .ZN(n4121) );
  NAND2_X1 U5103 ( .A1(n4125), .A2(EBX_REG_22__SCAN_IN), .ZN(n4120) );
  NAND2_X1 U5104 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n4231), .ZN(n4119) );
  NAND4_X1 U5105 ( .A1(n4121), .A2(n4120), .A3(n4128), .A4(n4119), .ZN(n4817)
         );
  INV_X1 U5106 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U5107 ( .A1(n4136), .A2(n5043), .ZN(n4124) );
  NAND2_X1 U5108 ( .A1(n2945), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4122) );
  OAI211_X1 U5109 ( .C1(n4231), .C2(EBX_REG_23__SCAN_IN), .A(n4122), .B(n2946), 
        .ZN(n4123) );
  AND2_X1 U5110 ( .A1(n4124), .A2(n4123), .ZN(n4767) );
  INV_X1 U5111 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5112 ( .A1(n4065), .A2(n4813), .ZN(n4129) );
  NAND2_X1 U5113 ( .A1(n4125), .A2(EBX_REG_24__SCAN_IN), .ZN(n4127) );
  NAND2_X1 U5114 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4231), .ZN(n4126) );
  NAND4_X1 U5115 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4812)
         );
  INV_X1 U5116 ( .A(EBX_REG_25__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5117 ( .A1(n4136), .A2(n4809), .ZN(n4131) );
  NAND2_X1 U5118 ( .A1(n4052), .A2(EBX_REG_25__SCAN_IN), .ZN(n4130) );
  OAI211_X1 U5119 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n4227), .A(n4131), .B(n4130), .ZN(n4806) );
  INV_X1 U5120 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U5121 ( .A1(n4065), .A2(n5026), .ZN(n4134) );
  NAND2_X1 U5122 ( .A1(n2946), .A2(n4919), .ZN(n4132) );
  OAI211_X1 U5123 ( .C1(n4231), .C2(EBX_REG_26__SCAN_IN), .A(n4132), .B(n2945), 
        .ZN(n4133) );
  NAND2_X1 U5124 ( .A1(n4134), .A2(n4133), .ZN(n4750) );
  NAND2_X1 U5125 ( .A1(n4749), .A2(n4750), .ZN(n4799) );
  INV_X1 U5126 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4135) );
  NAND2_X1 U5127 ( .A1(n4136), .A2(n4135), .ZN(n4138) );
  NAND2_X1 U5128 ( .A1(n4052), .A2(EBX_REG_27__SCAN_IN), .ZN(n4137) );
  OAI211_X1 U5129 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n4227), .A(n4138), .B(n4137), .ZN(n4798) );
  INV_X1 U5130 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5004) );
  NAND2_X1 U5131 ( .A1(n4065), .A2(n5004), .ZN(n4143) );
  NAND2_X1 U5132 ( .A1(n2946), .A2(n4139), .ZN(n4141) );
  OAI211_X1 U5133 ( .C1(n4231), .C2(EBX_REG_28__SCAN_IN), .A(n4141), .B(n2945), 
        .ZN(n4142) );
  AND2_X1 U5134 ( .A1(n4143), .A2(n4142), .ZN(n4771) );
  NAND2_X1 U5135 ( .A1(n4773), .A2(n4052), .ZN(n4225) );
  OAI22_X1 U5136 ( .A1(n4227), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4231), .ZN(n4222) );
  AOI22_X1 U5137 ( .A1(n4227), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n4231), .ZN(n4226) );
  INV_X1 U5138 ( .A(n4041), .ZN(n4145) );
  NAND2_X1 U5139 ( .A1(n4145), .A2(n4244), .ZN(n6169) );
  NAND2_X1 U5140 ( .A1(n4146), .A2(n3216), .ZN(n4147) );
  NAND2_X1 U5141 ( .A1(n6169), .A2(n4147), .ZN(n4148) );
  AND2_X1 U5142 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4883) );
  NOR2_X1 U5143 ( .A1(n4033), .A2(n4149), .ZN(n6136) );
  NAND2_X1 U5144 ( .A1(n4173), .A2(n6136), .ZN(n5595) );
  NAND2_X1 U5145 ( .A1(n3889), .A2(n3180), .ZN(n4150) );
  NAND2_X1 U5146 ( .A1(n4153), .A2(n4152), .ZN(n4157) );
  NAND2_X1 U5147 ( .A1(n4155), .A2(n4052), .ZN(n4156) );
  NAND4_X1 U5148 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4342)
         );
  AND2_X1 U5149 ( .A1(n4160), .A2(n2978), .ZN(n4161) );
  OR2_X1 U5150 ( .A1(n4342), .A2(n4161), .ZN(n4162) );
  NAND2_X1 U5151 ( .A1(n4173), .A2(n4162), .ZN(n4661) );
  NAND2_X1 U5152 ( .A1(n4164), .A2(n4163), .ZN(n4326) );
  INV_X1 U5153 ( .A(n4347), .ZN(n6158) );
  NAND2_X1 U5154 ( .A1(n6158), .A2(n4173), .ZN(n4662) );
  NAND2_X1 U5155 ( .A1(n4468), .A2(n4662), .ZN(n5580) );
  AND2_X1 U5156 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U5157 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5158 ( .A1(n4166), .A2(n4669), .ZN(n4701) );
  NAND2_X1 U5159 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4701), .ZN(n4958) );
  NAND2_X1 U5160 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4961) );
  NOR2_X1 U5161 ( .A1(n4958), .A2(n4961), .ZN(n4179) );
  NAND2_X1 U5162 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U5163 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5554) );
  NOR2_X1 U5164 ( .A1(n5553), .A2(n5554), .ZN(n4168) );
  NAND2_X1 U5165 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4167) );
  NOR2_X1 U5166 ( .A1(n4059), .A2(n5587), .ZN(n5574) );
  NAND3_X1 U5167 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n5574), .ZN(n4966) );
  NOR2_X1 U5168 ( .A1(n4167), .A2(n4966), .ZN(n4467) );
  NAND2_X1 U5169 ( .A1(n4168), .A2(n4467), .ZN(n4177) );
  NOR2_X1 U5170 ( .A1(n4661), .A2(n4177), .ZN(n4169) );
  AOI21_X1 U5171 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4411) );
  NAND2_X1 U5172 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U5173 ( .A1(n4411), .A2(n4976), .ZN(n4972) );
  NAND3_X1 U5174 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4972), .ZN(n4471) );
  INV_X1 U5175 ( .A(n4168), .ZN(n4641) );
  NOR2_X1 U5176 ( .A1(n4471), .A2(n4641), .ZN(n4180) );
  AOI22_X1 U5177 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4169), .B1(n5582), 
        .B2(n4180), .ZN(n4660) );
  OR2_X1 U5178 ( .A1(n5595), .A2(n4177), .ZN(n4668) );
  NAND2_X1 U5179 ( .A1(n4660), .A2(n4668), .ZN(n4642) );
  NAND2_X1 U5180 ( .A1(n4179), .A2(n4642), .ZN(n5196) );
  INV_X1 U5181 ( .A(n5196), .ZN(n4170) );
  NAND2_X1 U5182 ( .A1(n4170), .A2(n2995), .ZN(n5182) );
  INV_X1 U5183 ( .A(n4945), .ZN(n4171) );
  NOR2_X1 U5184 ( .A1(n5182), .A2(n4171), .ZN(n5172) );
  NAND2_X1 U5185 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4172) );
  NAND2_X1 U5186 ( .A1(n5172), .A2(n4172), .ZN(n4937) );
  OR2_X1 U5187 ( .A1(n4661), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4175)
         );
  OR2_X1 U5188 ( .A1(n4173), .A2(n5585), .ZN(n4174) );
  NAND2_X1 U5189 ( .A1(n4175), .A2(n4174), .ZN(n5581) );
  INV_X1 U5190 ( .A(n4179), .ZN(n4176) );
  NOR2_X1 U5191 ( .A1(n4177), .A2(n4176), .ZN(n4178) );
  NOR2_X1 U5192 ( .A1(n4468), .A2(n4178), .ZN(n4183) );
  AND2_X1 U5193 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  NOR2_X1 U5194 ( .A1(n4662), .A2(n4181), .ZN(n4182) );
  NAND2_X1 U5195 ( .A1(n2995), .A2(n4945), .ZN(n4184) );
  AND2_X1 U5196 ( .A1(n5580), .A2(n4184), .ZN(n4185) );
  NOR2_X1 U5197 ( .A1(n5190), .A2(n4185), .ZN(n5175) );
  INV_X1 U5198 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U5199 ( .A1(n6461), .A2(n5595), .ZN(n5579) );
  INV_X1 U5200 ( .A(n5579), .ZN(n4186) );
  NAND2_X1 U5201 ( .A1(n5568), .A2(n4662), .ZN(n4948) );
  INV_X1 U5202 ( .A(n4187), .ZN(n4188) );
  NAND2_X1 U5203 ( .A1(n4948), .A2(n4188), .ZN(n4189) );
  OAI21_X1 U5204 ( .B1(n4949), .B2(n4914), .A(n5168), .ZN(n4908) );
  AOI21_X1 U5205 ( .B1(n4192), .B2(n5580), .A(n4908), .ZN(n4281) );
  OAI21_X1 U5206 ( .B1(n4883), .B2(n4949), .A(n4281), .ZN(n4889) );
  INV_X1 U5207 ( .A(n4914), .ZN(n4191) );
  NOR2_X1 U5208 ( .A1(n5161), .A2(n4191), .ZN(n4904) );
  INV_X1 U5209 ( .A(n4192), .ZN(n4895) );
  NAND2_X1 U5210 ( .A1(n4904), .A2(n4895), .ZN(n4885) );
  INV_X1 U5211 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4280) );
  NOR3_X1 U5212 ( .A1(n4885), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4280), 
        .ZN(n4195) );
  INV_X1 U5213 ( .A(n4193), .ZN(n4194) );
  NAND2_X1 U5214 ( .A1(n4199), .A2(n4198), .ZN(U2988) );
  INV_X1 U5215 ( .A(n4200), .ZN(n4993) );
  NAND2_X1 U5216 ( .A1(n4201), .A2(n5207), .ZN(n4202) );
  OAI21_X4 U5217 ( .B1(n4335), .B2(n6178), .A(n4202), .ZN(n4833) );
  INV_X1 U5218 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4985) );
  OAI22_X1 U5219 ( .A1(n2983), .A2(n4838), .B1(n4833), .B2(n4985), .ZN(n4203)
         );
  INV_X1 U5220 ( .A(n4203), .ZN(n4204) );
  INV_X1 U5221 ( .A(n4289), .ZN(n4206) );
  NAND2_X1 U5222 ( .A1(n4206), .A2(n4205), .ZN(n4210) );
  AOI22_X1 U5223 ( .A1(n3763), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4207), .ZN(n4208) );
  INV_X1 U5224 ( .A(n4208), .ZN(n4209) );
  XNOR2_X2 U5225 ( .A(n4210), .B(n4209), .ZN(n4853) );
  NOR2_X1 U5226 ( .A1(n4033), .A2(n6153), .ZN(n5202) );
  INV_X1 U5227 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U5228 ( .A1(n6395), .A2(n5766), .ZN(n6188) );
  NOR3_X1 U5229 ( .A1(n6180), .A2(n6034), .A3(n6188), .ZN(n6176) );
  NOR3_X1 U5230 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6395), .A3(n4211), .ZN(
        n6185) );
  INV_X1 U5231 ( .A(n6185), .ZN(n4212) );
  NAND2_X1 U5232 ( .A1(n5599), .A2(n4212), .ZN(n4213) );
  NOR2_X1 U5233 ( .A1(n6176), .A2(n4213), .ZN(n4214) );
  INV_X1 U5234 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4217) );
  NOR2_X1 U5235 ( .A1(n4854), .A2(n6395), .ZN(n4219) );
  NAND2_X1 U5236 ( .A1(n4052), .A2(EBX_REG_29__SCAN_IN), .ZN(n4220) );
  INV_X1 U5237 ( .A(n4220), .ZN(n4224) );
  AOI21_X1 U5238 ( .B1(n4222), .B2(n2945), .A(n4224), .ZN(n4274) );
  NAND2_X1 U5239 ( .A1(n4223), .A2(n4274), .ZN(n4277) );
  OAI211_X1 U5240 ( .C1(n4277), .C2(n4226), .A(n4220), .B(n4225), .ZN(n4229)
         );
  OAI22_X1 U5241 ( .A1(n4227), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4231), .ZN(n4228) );
  XNOR2_X1 U5242 ( .A(n4229), .B(n4228), .ZN(n4888) );
  NOR2_X1 U5243 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4232) );
  INV_X1 U5244 ( .A(n4232), .ZN(n6168) );
  NAND2_X1 U5245 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4239) );
  NAND3_X1 U5246 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4237) );
  NAND2_X1 U5247 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5075) );
  INV_X1 U5248 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U5249 ( .A1(n4608), .A2(n4232), .ZN(n4233) );
  INV_X1 U5250 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5277) );
  INV_X1 U5251 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6452) );
  INV_X1 U5252 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6221) );
  INV_X1 U5253 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6423) );
  INV_X1 U5254 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6394) );
  INV_X1 U5255 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6212) );
  NOR3_X1 U5256 ( .A1(n6423), .A2(n6394), .A3(n6212), .ZN(n5345) );
  NAND3_X1 U5257 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        n5345), .ZN(n5297) );
  NAND3_X1 U5258 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5299) );
  NOR4_X1 U5259 ( .A1(n6452), .A2(n6221), .A3(n5297), .A4(n5299), .ZN(n5287)
         );
  NAND2_X1 U5260 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5287), .ZN(n5276) );
  NOR2_X1 U5261 ( .A1(n5277), .A2(n5276), .ZN(n5256) );
  NAND3_X1 U5262 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n5256), .ZN(n4236) );
  NAND2_X1 U5263 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5251), .ZN(n5241) );
  NOR2_X2 U5264 ( .A1(n4237), .A2(n5055), .ZN(n5032) );
  NAND4_X1 U5265 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5032), .ZN(n5014) );
  NOR2_X1 U5266 ( .A1(n4239), .A2(n5014), .ZN(n4240) );
  NAND2_X1 U5267 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4240), .ZN(n4241) );
  NOR2_X1 U5268 ( .A1(REIP_REG_30__SCAN_IN), .A2(n4241), .ZN(n4987) );
  INV_X1 U5269 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6397) );
  INV_X1 U5270 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6233) );
  OR2_X1 U5271 ( .A1(n4236), .A2(n5295), .ZN(n5248) );
  NOR4_X1 U5272 ( .A1(n6397), .A2(n6233), .A3(n6230), .A4(n5248), .ZN(n5074)
         );
  NAND4_X1 U5273 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5074), .A4(REIP_REG_18__SCAN_IN), .ZN(n5051) );
  NOR2_X1 U5274 ( .A1(n5051), .A2(n4237), .ZN(n5031) );
  INV_X1 U5275 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6364) );
  INV_X1 U5276 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5019) );
  INV_X1 U5277 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6246) );
  NOR3_X1 U5278 ( .A1(n6364), .A2(n5019), .A3(n6246), .ZN(n4238) );
  NAND2_X1 U5279 ( .A1(n4605), .A2(n5275), .ZN(n5368) );
  AOI21_X1 U5280 ( .B1(n5031), .B2(n4238), .A(n5330), .ZN(n5023) );
  AOI21_X1 U5281 ( .B1(n5346), .B2(n4239), .A(n5023), .ZN(n5006) );
  INV_X1 U5282 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U5283 ( .A1(n4240), .A2(n6254), .ZN(n4998) );
  NAND2_X1 U5284 ( .A1(n5006), .A2(n4998), .ZN(n4989) );
  OAI21_X1 U5285 ( .B1(n4987), .B2(n4989), .A(REIP_REG_31__SCAN_IN), .ZN(n4249) );
  INV_X1 U5286 ( .A(n4241), .ZN(n4242) );
  INV_X1 U5287 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6258) );
  NAND3_X1 U5288 ( .A1(REIP_REG_30__SCAN_IN), .A2(n4242), .A3(n6258), .ZN(
        n4248) );
  OR2_X1 U5289 ( .A1(n6198), .A2(n6168), .ZN(n4243) );
  NAND2_X1 U5290 ( .A1(n4244), .A2(n4243), .ZN(n4607) );
  INV_X1 U5291 ( .A(n4607), .ZN(n4246) );
  NAND2_X1 U5292 ( .A1(n4605), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5343) );
  AOI22_X1 U5293 ( .A1(n4246), .A2(n4245), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n5375), .ZN(n4247) );
  NAND3_X1 U5294 ( .A1(n4249), .A2(n4248), .A3(n4247), .ZN(n4250) );
  XNOR2_X1 U5295 ( .A(n3980), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5134)
         );
  NAND2_X1 U5296 ( .A1(n5135), .A2(n5134), .ZN(n4864) );
  XNOR2_X1 U5297 ( .A(n3980), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4877)
         );
  INV_X1 U5298 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4255) );
  XNOR2_X1 U5299 ( .A(n3980), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5126)
         );
  OR2_X2 U5300 ( .A1(n4873), .A2(n3033), .ZN(n4259) );
  NOR2_X1 U5301 ( .A1(n3980), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4871)
         );
  NAND2_X1 U5302 ( .A1(n4871), .A2(n6354), .ZN(n4257) );
  OAI21_X1 U5303 ( .B1(n4262), .B2(n4264), .A(n4263), .ZN(n4815) );
  INV_X1 U5304 ( .A(n4815), .ZN(n5092) );
  NOR2_X1 U5305 ( .A1(n5599), .A2(n6364), .ZN(n4924) );
  AOI21_X1 U5306 ( .B1(n5517), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4924), 
        .ZN(n4265) );
  OAI21_X1 U5307 ( .B1(n4266), .B2(n5525), .A(n4265), .ZN(n4267) );
  AOI21_X1 U5308 ( .B1(n5092), .B2(n5631), .A(n4267), .ZN(n4268) );
  OAI21_X1 U5309 ( .B1(n4926), .B2(n5503), .A(n4268), .ZN(U2962) );
  INV_X1 U5310 ( .A(n4850), .ZN(n4273) );
  NAND3_X1 U5311 ( .A1(n4273), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4269), .ZN(n4272) );
  INV_X1 U5312 ( .A(n4270), .ZN(n4271) );
  NAND2_X1 U5313 ( .A1(n4286), .A2(n5591), .ZN(n4285) );
  INV_X1 U5314 ( .A(n4885), .ZN(n4279) );
  INV_X1 U5315 ( .A(n4274), .ZN(n4275) );
  NAND2_X1 U5316 ( .A1(n4773), .A2(n4275), .ZN(n4276) );
  NAND2_X1 U5317 ( .A1(n4277), .A2(n4276), .ZN(n5000) );
  NAND2_X1 U5318 ( .A1(n5585), .A2(REIP_REG_29__SCAN_IN), .ZN(n4291) );
  OAI21_X1 U5319 ( .B1(n5000), .B2(n5540), .A(n4291), .ZN(n4278) );
  AOI21_X1 U5320 ( .B1(n4279), .B2(n4280), .A(n4278), .ZN(n4283) );
  OR2_X1 U5321 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  NAND2_X1 U5322 ( .A1(n4285), .A2(n4284), .ZN(U2989) );
  INV_X1 U5323 ( .A(n5082), .ZN(n4796) );
  NAND2_X1 U5324 ( .A1(n5517), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4290)
         );
  OAI211_X1 U5325 ( .C1(n5525), .C2(n4995), .A(n4291), .B(n4290), .ZN(n4292)
         );
  AOI21_X1 U5326 ( .B1(n5082), .B2(n5631), .A(n4292), .ZN(n4293) );
  NAND2_X1 U5327 ( .A1(n4294), .A2(n4293), .ZN(U2957) );
  INV_X1 U5328 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4296) );
  INV_X1 U5329 ( .A(n4385), .ZN(n4295) );
  OAI211_X1 U5330 ( .C1(n4297), .C2(n4296), .A(n4295), .B(n6316), .ZN(U2788)
         );
  INV_X1 U5331 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4301) );
  INV_X1 U5332 ( .A(n6136), .ZN(n4425) );
  NAND2_X1 U5333 ( .A1(n6169), .A2(n4425), .ZN(n4299) );
  NOR2_X1 U5334 ( .A1(n6395), .A2(n5766), .ZN(n6285) );
  NAND2_X1 U5335 ( .A1(n6180), .A2(n6285), .ZN(n5435) );
  AOI22_X1 U5336 ( .A1(n6170), .A2(UWORD_REG_1__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4300) );
  OAI21_X1 U5337 ( .B1(n4301), .B2(n5410), .A(n4300), .ZN(U2906) );
  INV_X1 U5338 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6348) );
  AOI22_X1 U5339 ( .A1(n6170), .A2(UWORD_REG_3__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4302) );
  OAI21_X1 U5340 ( .B1(n6348), .B2(n5410), .A(n4302), .ZN(U2904) );
  AOI22_X1 U5341 ( .A1(n6307), .A2(UWORD_REG_5__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4303) );
  OAI21_X1 U5342 ( .B1(n4304), .B2(n5410), .A(n4303), .ZN(U2902) );
  INV_X1 U5343 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U5344 ( .A1(n6170), .A2(UWORD_REG_6__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4305) );
  OAI21_X1 U5345 ( .B1(n4306), .B2(n5410), .A(n4305), .ZN(U2901) );
  INV_X1 U5346 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U5347 ( .A1(n6170), .A2(UWORD_REG_2__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4307) );
  OAI21_X1 U5348 ( .B1(n4308), .B2(n5410), .A(n4307), .ZN(U2905) );
  INV_X1 U5349 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5350 ( .A1(n6307), .A2(UWORD_REG_8__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4309) );
  OAI21_X1 U5351 ( .B1(n4310), .B2(n5410), .A(n4309), .ZN(U2899) );
  INV_X1 U5352 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U5353 ( .A1(n6170), .A2(UWORD_REG_4__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4311) );
  OAI21_X1 U5354 ( .B1(n4312), .B2(n5410), .A(n4311), .ZN(U2903) );
  INV_X1 U5355 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U5356 ( .A1(n6307), .A2(UWORD_REG_10__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4313) );
  OAI21_X1 U5357 ( .B1(n4314), .B2(n5410), .A(n4313), .ZN(U2897) );
  INV_X1 U5358 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U5359 ( .A1(n6307), .A2(UWORD_REG_9__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4315) );
  OAI21_X1 U5360 ( .B1(n4316), .B2(n5410), .A(n4315), .ZN(U2898) );
  INV_X1 U5361 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4318) );
  AOI22_X1 U5362 ( .A1(n6307), .A2(UWORD_REG_7__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4317) );
  OAI21_X1 U5363 ( .B1(n4318), .B2(n5410), .A(n4317), .ZN(U2900) );
  INV_X1 U5364 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U5365 ( .A1(n6170), .A2(UWORD_REG_0__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4319) );
  OAI21_X1 U5366 ( .B1(n4320), .B2(n5410), .A(n4319), .ZN(U2907) );
  AOI22_X1 U5367 ( .A1(n6307), .A2(UWORD_REG_14__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4321) );
  OAI21_X1 U5368 ( .B1(n3820), .B2(n5410), .A(n4321), .ZN(U2893) );
  INV_X1 U5369 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U5370 ( .A1(n6307), .A2(UWORD_REG_11__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4322) );
  OAI21_X1 U5371 ( .B1(n4323), .B2(n5410), .A(n4322), .ZN(U2896) );
  INV_X1 U5372 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5373 ( .A1(n6307), .A2(UWORD_REG_13__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4324) );
  OAI21_X1 U5374 ( .B1(n4325), .B2(n5410), .A(n4324), .ZN(U2894) );
  INV_X1 U5375 ( .A(n4326), .ZN(n4334) );
  AOI21_X1 U5376 ( .B1(n4425), .B2(n4041), .A(n4327), .ZN(n4328) );
  OAI211_X1 U5377 ( .C1(n3828), .C2(n4329), .A(n4328), .B(n6157), .ZN(n4332)
         );
  INV_X1 U5378 ( .A(n6157), .ZN(n4330) );
  OR2_X1 U5379 ( .A1(n6150), .A2(n4330), .ZN(n4331) );
  NAND2_X1 U5380 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6285), .ZN(n6189) );
  INV_X1 U5381 ( .A(n6189), .ZN(n6264) );
  AOI22_X1 U5382 ( .A1(n6181), .A2(n6138), .B1(FLUSH_REG_SCAN_IN), .B2(n6264), 
        .ZN(n5198) );
  INV_X1 U5383 ( .A(n5198), .ZN(n4337) );
  NOR2_X1 U5384 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6034), .ZN(n6265) );
  NOR2_X1 U5385 ( .A1(n4337), .A2(n6265), .ZN(n4792) );
  AOI21_X1 U5386 ( .B1(n6269), .B2(n4339), .A(n4338), .ZN(n4355) );
  OAI21_X1 U5387 ( .B1(n4340), .B2(n4785), .A(n6269), .ZN(n4782) );
  NAND2_X1 U5388 ( .A1(n4782), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4354) );
  INV_X1 U5389 ( .A(n4342), .ZN(n4346) );
  AND3_X1 U5390 ( .A1(n4344), .A2(n4343), .A3(n4041), .ZN(n4345) );
  NAND2_X1 U5391 ( .A1(n4346), .A2(n4345), .ZN(n6135) );
  NAND2_X1 U5392 ( .A1(n6029), .A2(n6135), .ZN(n4352) );
  NAND2_X1 U5393 ( .A1(n4347), .A2(n6150), .ZN(n4423) );
  INV_X1 U5394 ( .A(n4340), .ZN(n4783) );
  NAND2_X1 U5395 ( .A1(n4783), .A2(n3013), .ZN(n4421) );
  XNOR2_X1 U5396 ( .A(n4421), .B(n3037), .ZN(n4350) );
  XNOR2_X1 U5397 ( .A(n4348), .B(n3012), .ZN(n4349) );
  AOI22_X1 U5398 ( .A1(n4423), .A2(n4350), .B1(n6136), .B2(n4349), .ZN(n4351)
         );
  NAND2_X1 U5399 ( .A1(n4352), .A2(n4351), .ZN(n4429) );
  NAND3_X1 U5400 ( .A1(n6269), .A2(n6182), .A3(n4429), .ZN(n4353) );
  OAI211_X1 U5401 ( .C1(n4355), .C2(n4785), .A(n4354), .B(n4353), .ZN(U3456)
         );
  NAND2_X1 U5402 ( .A1(n5764), .A2(n6135), .ZN(n4359) );
  INV_X1 U5403 ( .A(n4357), .ZN(n4437) );
  NAND3_X1 U5404 ( .A1(n6134), .A2(n4783), .A3(n4437), .ZN(n4358) );
  OAI211_X1 U5405 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4425), .A(n4359), .B(n4358), .ZN(n6137) );
  NOR2_X1 U5406 ( .A1(n6395), .A2(n6461), .ZN(n4790) );
  INV_X1 U5407 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5408 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4360), .B2(n5587), .ZN(n4789)
         );
  INV_X1 U5409 ( .A(n4789), .ZN(n4362) );
  INV_X1 U5410 ( .A(n4785), .ZN(n6174) );
  AOI222_X1 U5411 ( .A1(n6137), .A2(n6182), .B1(n4790), .B2(n4362), .C1(n4361), 
        .C2(n6174), .ZN(n4365) );
  OAI21_X1 U5412 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4785), .A(n6269), 
        .ZN(n6270) );
  INV_X1 U5413 ( .A(n6270), .ZN(n4364) );
  OAI22_X1 U5414 ( .A1(n4792), .A2(n4365), .B1(n4363), .B2(n4364), .ZN(U3460)
         );
  OR2_X1 U5415 ( .A1(n4367), .A2(n4366), .ZN(n4368) );
  AND2_X1 U5416 ( .A1(n4369), .A2(n4368), .ZN(n5522) );
  INV_X1 U5417 ( .A(n5522), .ZN(n4734) );
  INV_X1 U5418 ( .A(n4370), .ZN(n4371) );
  INV_X1 U5419 ( .A(DATAI_1_), .ZN(n4499) );
  INV_X1 U5420 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6460) );
  OAI222_X1 U5421 ( .A1(n4734), .A2(n5403), .B1(n4457), .B2(n4499), .C1(n4839), 
        .C2(n6460), .ZN(U2890) );
  AOI21_X1 U5422 ( .B1(n4374), .B2(n4372), .A(n4373), .ZN(n4603) );
  INV_X1 U5423 ( .A(n4603), .ZN(n4572) );
  INV_X1 U5424 ( .A(DATAI_3_), .ZN(n5620) );
  INV_X1 U5425 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5432) );
  OAI222_X1 U5426 ( .A1(n4572), .A2(n5403), .B1(n4457), .B2(n5620), .C1(n4839), 
        .C2(n5432), .ZN(U2888) );
  AOI21_X1 U5427 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(n4378) );
  INV_X1 U5428 ( .A(n4378), .ZN(n5536) );
  INV_X1 U5429 ( .A(DATAI_0_), .ZN(n4496) );
  INV_X1 U5430 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5440) );
  OAI222_X1 U5431 ( .A1(n5536), .A2(n5403), .B1(n4457), .B2(n4496), .C1(n4839), 
        .C2(n5440), .ZN(U2891) );
  OAI21_X1 U5432 ( .B1(n4380), .B2(n4379), .A(n4372), .ZN(n4681) );
  INV_X1 U5433 ( .A(DATAI_2_), .ZN(n4493) );
  INV_X1 U5434 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5434) );
  OAI222_X1 U5435 ( .A1(n4681), .A2(n5403), .B1(n4457), .B2(n4493), .C1(n4839), 
        .C2(n5434), .ZN(U2889) );
  OAI21_X1 U5436 ( .B1(n4373), .B2(n4382), .A(n4381), .ZN(n5361) );
  INV_X1 U5437 ( .A(DATAI_4_), .ZN(n5623) );
  OAI222_X1 U5438 ( .A1(n5361), .A2(n5403), .B1(n4457), .B2(n5623), .C1(n4839), 
        .C2(n6441), .ZN(U2887) );
  INV_X1 U5439 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4387) );
  INV_X1 U5440 ( .A(DATAI_7_), .ZN(n4778) );
  NOR2_X1 U5441 ( .A1(n4403), .A2(n4778), .ZN(n4393) );
  AOI21_X1 U5442 ( .B1(n5459), .B2(EAX_REG_23__SCAN_IN), .A(n4393), .ZN(n4386)
         );
  OAI21_X1 U5443 ( .B1(n4522), .B2(n4387), .A(n4386), .ZN(U2931) );
  INV_X1 U5444 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n4389) );
  INV_X1 U5445 ( .A(DATAI_8_), .ZN(n6408) );
  NOR2_X1 U5446 ( .A1(n4403), .A2(n6408), .ZN(n4390) );
  AOI21_X1 U5447 ( .B1(n5459), .B2(EAX_REG_8__SCAN_IN), .A(n4390), .ZN(n4388)
         );
  OAI21_X1 U5448 ( .B1(n4522), .B2(n4389), .A(n4388), .ZN(U2947) );
  INV_X1 U5449 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4392) );
  AOI21_X1 U5450 ( .B1(n5459), .B2(EAX_REG_24__SCAN_IN), .A(n4390), .ZN(n4391)
         );
  OAI21_X1 U5451 ( .B1(n4522), .B2(n4392), .A(n4391), .ZN(U2932) );
  INV_X1 U5452 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4395) );
  AOI21_X1 U5453 ( .B1(n5459), .B2(EAX_REG_7__SCAN_IN), .A(n4393), .ZN(n4394)
         );
  OAI21_X1 U5454 ( .B1(n4522), .B2(n4395), .A(n4394), .ZN(U2946) );
  INV_X1 U5455 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5456 ( .A1(n6437), .A2(DATAI_1_), .ZN(n4530) );
  NAND2_X1 U5457 ( .A1(n5459), .A2(EAX_REG_1__SCAN_IN), .ZN(n4396) );
  OAI211_X1 U5458 ( .C1(n4522), .C2(n4397), .A(n4530), .B(n4396), .ZN(U2940)
         );
  XNOR2_X1 U5459 ( .A(n4399), .B(n4398), .ZN(n4417) );
  NAND2_X1 U5460 ( .A1(n4603), .A2(n5631), .ZN(n4402) );
  NOR2_X1 U5461 ( .A1(n5599), .A2(n6212), .ZN(n4414) );
  AND2_X1 U5462 ( .A1(n5517), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4400)
         );
  AOI211_X1 U5463 ( .C1(n5483), .C2(n4616), .A(n4414), .B(n4400), .ZN(n4401)
         );
  OAI211_X1 U5464 ( .C1(n4417), .C2(n5503), .A(n4402), .B(n4401), .ZN(U2983)
         );
  INV_X1 U5465 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4404) );
  OAI222_X1 U5466 ( .A1(n4404), .A2(n4522), .B1(n4403), .B2(n5623), .C1(n6440), 
        .C2(n4312), .ZN(U2928) );
  OAI21_X1 U5467 ( .B1(n2964), .B2(n4407), .A(n4406), .ZN(n5500) );
  AOI22_X1 U5468 ( .A1(n4654), .A2(DATAI_6_), .B1(n5406), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4408) );
  OAI21_X1 U5469 ( .B1(n5500), .B2(n5403), .A(n4408), .ZN(U2885) );
  INV_X1 U5470 ( .A(n4468), .ZN(n4409) );
  INV_X1 U5471 ( .A(n5574), .ZN(n4410) );
  AOI21_X1 U5472 ( .B1(n4409), .B2(n4410), .A(n5581), .ZN(n5569) );
  NAND2_X1 U5473 ( .A1(n5582), .A2(n4411), .ZN(n5576) );
  NAND2_X1 U5474 ( .A1(n5569), .A2(n5576), .ZN(n4981) );
  OAI21_X1 U5475 ( .B1(n4410), .B2(n5568), .A(n4662), .ZN(n4508) );
  INV_X1 U5476 ( .A(n4508), .ZN(n4470) );
  NOR2_X1 U5477 ( .A1(n4411), .A2(n4470), .ZN(n4977) );
  AOI22_X1 U5478 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4981), .B1(n4977), 
        .B2(n6463), .ZN(n4416) );
  AOI21_X1 U5479 ( .B1(n4413), .B2(n4412), .A(n4758), .ZN(n4571) );
  AOI21_X1 U5480 ( .B1(n5590), .B2(n4571), .A(n4414), .ZN(n4415) );
  OAI211_X1 U5481 ( .C1(n5541), .C2(n4417), .A(n4416), .B(n4415), .ZN(U3015)
         );
  INV_X1 U5482 ( .A(n6188), .ZN(n6310) );
  INV_X1 U5483 ( .A(n4419), .ZN(n5765) );
  XNOR2_X1 U5484 ( .A(n4784), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4426)
         );
  NAND2_X1 U5485 ( .A1(n4340), .A2(n4784), .ZN(n4420) );
  NAND2_X1 U5486 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  NAND2_X1 U5487 ( .A1(n4423), .A2(n4422), .ZN(n4424) );
  OAI21_X1 U5488 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4427) );
  AOI21_X1 U5489 ( .B1(n5765), .B2(n6135), .A(n4427), .ZN(n4786) );
  NOR2_X1 U5490 ( .A1(n6138), .A2(n4784), .ZN(n4428) );
  AOI21_X1 U5491 ( .B1(n4786), .B2(n6138), .A(n4428), .ZN(n6143) );
  NAND2_X1 U5492 ( .A1(n4429), .A2(n6138), .ZN(n4432) );
  INV_X1 U5493 ( .A(n6138), .ZN(n4430) );
  NAND2_X1 U5494 ( .A1(n4430), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5495 ( .A1(n4432), .A2(n4431), .ZN(n6146) );
  NAND3_X1 U5496 ( .A1(n6143), .A2(n6395), .A3(n6146), .ZN(n4436) );
  INV_X1 U5497 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5209) );
  NAND2_X1 U5498 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5209), .ZN(n4443) );
  INV_X1 U5499 ( .A(n4443), .ZN(n4433) );
  NAND2_X1 U5500 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  NAND2_X1 U5501 ( .A1(n4436), .A2(n4435), .ZN(n6164) );
  NAND2_X1 U5502 ( .A1(n6164), .A2(n4437), .ZN(n4445) );
  INV_X1 U5503 ( .A(n5966), .ZN(n5710) );
  NOR2_X1 U5504 ( .A1(n4438), .A2(n5710), .ZN(n4439) );
  XOR2_X1 U5505 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n4439), .Z(n5352) );
  NAND2_X1 U5506 ( .A1(n5352), .A2(n4440), .ZN(n5197) );
  OAI21_X1 U5507 ( .B1(n6138), .B2(n5200), .A(n5197), .ZN(n4441) );
  INV_X1 U5508 ( .A(n4441), .ZN(n4442) );
  OAI22_X1 U5509 ( .A1(n4443), .A2(n5200), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n4442), .ZN(n4444) );
  INV_X1 U5510 ( .A(n4444), .ZN(n6161) );
  NAND2_X1 U5511 ( .A1(n4445), .A2(n6161), .ZN(n6167) );
  OAI21_X1 U5512 ( .B1(n6167), .B2(FLUSH_REG_SCAN_IN), .A(n6264), .ZN(n4446)
         );
  NAND2_X1 U5513 ( .A1(n5630), .A2(n4446), .ZN(n6291) );
  INV_X1 U5514 ( .A(n5926), .ZN(n5606) );
  AOI21_X1 U5515 ( .B1(n5606), .B2(n6026), .A(n6275), .ZN(n4448) );
  NAND2_X1 U5516 ( .A1(n5926), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5919) );
  NOR2_X1 U5517 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6395), .ZN(n6278) );
  INV_X1 U5518 ( .A(n6278), .ZN(n6287) );
  AOI22_X1 U5519 ( .A1(n4448), .A2(n5919), .B1(n5764), .B2(n6287), .ZN(n4450)
         );
  NAND2_X1 U5520 ( .A1(n6294), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5521 ( .B1(n6294), .B2(n4450), .A(n4449), .ZN(U3464) );
  XNOR2_X1 U5522 ( .A(n4452), .B(n5919), .ZN(n4453) );
  AOI22_X1 U5523 ( .A1(n4453), .A2(n6289), .B1(n5765), .B2(n6287), .ZN(n4455)
         );
  NAND2_X1 U5524 ( .A1(n6294), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4454) );
  OAI21_X1 U5525 ( .B1(n6294), .B2(n4455), .A(n4454), .ZN(U3463) );
  AOI21_X1 U5526 ( .B1(n4456), .B2(n4381), .A(n2964), .ZN(n5506) );
  INV_X1 U5527 ( .A(n5506), .ZN(n4558) );
  INV_X1 U5528 ( .A(DATAI_5_), .ZN(n4485) );
  INV_X1 U5529 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4535) );
  OAI222_X1 U5530 ( .A1(n4558), .A2(n5403), .B1(n4457), .B2(n4485), .C1(n4839), 
        .C2(n4535), .ZN(U2886) );
  XOR2_X1 U5531 ( .A(n4459), .B(n4458), .Z(n4980) );
  INV_X1 U5532 ( .A(n4980), .ZN(n4462) );
  INV_X1 U5533 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6451) );
  NOR2_X1 U5534 ( .A1(n5599), .A2(n6451), .ZN(n4979) );
  OAI22_X1 U5535 ( .A1(n5525), .A2(n5360), .B1(n6076), .B2(n5361), .ZN(n4460)
         );
  AOI211_X1 U5536 ( .C1(n5517), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4979), 
        .B(n4460), .ZN(n4461) );
  OAI21_X1 U5537 ( .B1(n4462), .B2(n5503), .A(n4461), .ZN(U2982) );
  XNOR2_X1 U5538 ( .A(n4463), .B(n4465), .ZN(n5488) );
  AOI21_X1 U5539 ( .B1(n5582), .B2(n4471), .A(n5581), .ZN(n4466) );
  OAI21_X1 U5540 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n5548) );
  XNOR2_X1 U5541 ( .A(n4469), .B(n4506), .ZN(n5326) );
  NAND2_X1 U5542 ( .A1(n5585), .A2(REIP_REG_7__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U5543 ( .B1(n5540), .B2(n5326), .A(n5491), .ZN(n4473) );
  NOR2_X1 U5544 ( .A1(n5552), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4472)
         );
  AOI211_X1 U5545 ( .C1(n5548), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4473), 
        .B(n4472), .ZN(n4474) );
  OAI21_X1 U5546 ( .B1(n5541), .B2(n5488), .A(n4474), .ZN(U3011) );
  INV_X1 U5547 ( .A(n4475), .ZN(n5920) );
  NAND2_X1 U5548 ( .A1(n5920), .A2(n6284), .ZN(n4781) );
  NAND2_X1 U5549 ( .A1(n4777), .A2(n4477), .ZN(n5626) );
  NAND2_X1 U5550 ( .A1(n4419), .A2(n5764), .ZN(n5891) );
  INV_X1 U5551 ( .A(n5673), .ZN(n4478) );
  INV_X1 U5552 ( .A(n4781), .ZN(n5701) );
  AOI21_X1 U5553 ( .B1(n4478), .B2(n6288), .A(n5701), .ZN(n4487) );
  INV_X1 U5554 ( .A(n4487), .ZN(n4484) );
  NOR2_X1 U5555 ( .A1(n5926), .A2(n5797), .ZN(n4479) );
  NAND2_X1 U5556 ( .A1(n4452), .A2(n4479), .ZN(n5999) );
  INV_X1 U5557 ( .A(n5999), .ZN(n4480) );
  NAND2_X1 U5558 ( .A1(n4480), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5995) );
  AND2_X1 U5559 ( .A1(n5995), .A2(n5928), .ZN(n6277) );
  INV_X1 U5560 ( .A(n4452), .ZN(n4481) );
  INV_X1 U5561 ( .A(n5919), .ZN(n5796) );
  NAND3_X1 U5562 ( .A1(n6277), .A2(n4481), .A3(n5796), .ZN(n4482) );
  NAND2_X1 U5563 ( .A1(n4482), .A2(n6289), .ZN(n4486) );
  NAND3_X1 U5564 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6284), .A3(n6145), .ZN(n5670) );
  OAI21_X1 U5565 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6034), .A(n5831), 
        .ZN(n5736) );
  AOI21_X1 U5566 ( .B1(n6275), .B2(n5670), .A(n5736), .ZN(n4483) );
  OAI21_X1 U5567 ( .B1(n4484), .B2(n4486), .A(n4483), .ZN(n5703) );
  NOR2_X2 U5568 ( .A1(n4485), .A2(n5630), .ZN(n6111) );
  OAI22_X1 U5569 ( .A1(n4487), .A2(n4486), .B1(n5766), .B2(n5670), .ZN(n5702)
         );
  AOI22_X1 U5570 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5703), .B1(n6111), 
        .B2(n5702), .ZN(n4491) );
  NAND2_X1 U5571 ( .A1(n3933), .A2(n5926), .ZN(n4488) );
  AND2_X1 U5572 ( .A1(n5631), .A2(DATAI_21_), .ZN(n6113) );
  NOR2_X2 U5573 ( .A1(n4489), .A2(n6290), .ZN(n5700) );
  AND2_X1 U5574 ( .A1(n5631), .A2(DATAI_29_), .ZN(n6055) );
  AOI22_X1 U5575 ( .A1(n5726), .A2(n6113), .B1(n5700), .B2(n6055), .ZN(n4490)
         );
  OAI211_X1 U5576 ( .C1(n4781), .C2(n5626), .A(n4491), .B(n4490), .ZN(U3049)
         );
  NAND2_X1 U5577 ( .A1(n4777), .A2(n4492), .ZN(n5616) );
  NOR2_X2 U5578 ( .A1(n4493), .A2(n5630), .ZN(n6093) );
  AOI22_X1 U5579 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5703), .B1(n6093), 
        .B2(n5702), .ZN(n4495) );
  AND2_X1 U5580 ( .A1(n5631), .A2(DATAI_18_), .ZN(n6095) );
  AND2_X1 U5581 ( .A1(n5631), .A2(DATAI_26_), .ZN(n6043) );
  AOI22_X1 U5582 ( .A1(n5726), .A2(n6095), .B1(n5700), .B2(n6043), .ZN(n4494)
         );
  OAI211_X1 U5583 ( .C1(n4781), .C2(n5616), .A(n4495), .B(n4494), .ZN(U3046)
         );
  NAND2_X1 U5584 ( .A1(n4777), .A2(n3843), .ZN(n5601) );
  NOR2_X2 U5585 ( .A1(n4496), .A2(n5630), .ZN(n6074) );
  AOI22_X1 U5586 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5703), .B1(n6074), 
        .B2(n5702), .ZN(n4498) );
  AND2_X1 U5587 ( .A1(n5631), .A2(DATAI_16_), .ZN(n6083) );
  AND2_X1 U5588 ( .A1(n5631), .A2(DATAI_24_), .ZN(n6035) );
  AOI22_X1 U5589 ( .A1(n5726), .A2(n6083), .B1(n5700), .B2(n6035), .ZN(n4497)
         );
  OAI211_X1 U5590 ( .C1(n4781), .C2(n5601), .A(n4498), .B(n4497), .ZN(U3044)
         );
  NAND2_X1 U5591 ( .A1(n4777), .A2(n2980), .ZN(n5613) );
  NOR2_X2 U5592 ( .A1(n4499), .A2(n5630), .ZN(n6087) );
  AOI22_X1 U5593 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5703), .B1(n6087), 
        .B2(n5702), .ZN(n4501) );
  AND2_X1 U5594 ( .A1(n5631), .A2(DATAI_17_), .ZN(n6089) );
  AND2_X1 U5595 ( .A1(n5631), .A2(DATAI_25_), .ZN(n6039) );
  AOI22_X1 U5596 ( .A1(n5726), .A2(n6089), .B1(n5700), .B2(n6039), .ZN(n4500)
         );
  OAI211_X1 U5597 ( .C1(n4781), .C2(n5613), .A(n4501), .B(n4500), .ZN(U3045)
         );
  AND2_X1 U5598 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4972), .ZN(n4502)
         );
  OAI21_X1 U5599 ( .B1(n4949), .B2(n4502), .A(n5569), .ZN(n4971) );
  INV_X1 U5600 ( .A(n4971), .ZN(n4514) );
  XOR2_X1 U5601 ( .A(n4503), .B(n4504), .Z(n5494) );
  OR2_X1 U5602 ( .A1(n4505), .A2(n4555), .ZN(n4507) );
  NAND2_X1 U5603 ( .A1(n4507), .A2(n4506), .ZN(n4735) );
  NAND4_X1 U5604 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4972), .A3(n4508), 
        .A4(n4513), .ZN(n4510) );
  INV_X1 U5605 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6217) );
  NOR2_X1 U5606 ( .A1(n5599), .A2(n6217), .ZN(n5498) );
  INV_X1 U5607 ( .A(n5498), .ZN(n4509) );
  OAI211_X1 U5608 ( .C1(n5540), .C2(n4735), .A(n4510), .B(n4509), .ZN(n4511)
         );
  AOI21_X1 U5609 ( .B1(n5591), .B2(n5494), .A(n4511), .ZN(n4512) );
  OAI21_X1 U5610 ( .B1(n4514), .B2(n4513), .A(n4512), .ZN(U3012) );
  AOI21_X1 U5611 ( .B1(n4516), .B2(n4406), .A(n4515), .ZN(n5490) );
  INV_X1 U5612 ( .A(n5490), .ZN(n4521) );
  AOI22_X1 U5613 ( .A1(n4654), .A2(DATAI_7_), .B1(n5406), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4517) );
  OAI21_X1 U5614 ( .B1(n4521), .B2(n5403), .A(n4517), .ZN(U2884) );
  XOR2_X1 U5615 ( .A(n4515), .B(n4518), .Z(n5317) );
  INV_X1 U5616 ( .A(n5317), .ZN(n4581) );
  AOI22_X1 U5617 ( .A1(n4654), .A2(DATAI_8_), .B1(n5406), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4519) );
  OAI21_X1 U5618 ( .B1(n4581), .B2(n5403), .A(n4519), .ZN(U2883) );
  OAI222_X1 U5619 ( .A1(n4521), .A2(n4835), .B1(n4838), .B2(n5326), .C1(n4833), 
        .C2(n4520), .ZN(U2852) );
  NAND2_X1 U5620 ( .A1(n6438), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5621 ( .A1(n6437), .A2(DATAI_5_), .ZN(n4533) );
  OAI211_X1 U5622 ( .C1(n6440), .C2(n4304), .A(n4523), .B(n4533), .ZN(U2929)
         );
  INV_X1 U5623 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5624 ( .A1(n6438), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5625 ( .A1(n6437), .A2(DATAI_6_), .ZN(n4538) );
  OAI211_X1 U5626 ( .C1(n6440), .C2(n4525), .A(n4524), .B(n4538), .ZN(U2945)
         );
  NAND2_X1 U5627 ( .A1(n6438), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U5628 ( .A1(n6437), .A2(DATAI_3_), .ZN(n4536) );
  OAI211_X1 U5629 ( .C1(n6440), .C2(n6348), .A(n4526), .B(n4536), .ZN(U2927)
         );
  NAND2_X1 U5630 ( .A1(n6438), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4527) );
  NAND2_X1 U5631 ( .A1(n6437), .A2(DATAI_0_), .ZN(n4528) );
  OAI211_X1 U5632 ( .C1(n6440), .C2(n5440), .A(n4527), .B(n4528), .ZN(U2939)
         );
  NAND2_X1 U5633 ( .A1(n6438), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4529) );
  OAI211_X1 U5634 ( .C1(n6440), .C2(n4320), .A(n4529), .B(n4528), .ZN(U2924)
         );
  NAND2_X1 U5635 ( .A1(n6438), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4531) );
  OAI211_X1 U5636 ( .C1(n6440), .C2(n4301), .A(n4531), .B(n4530), .ZN(U2925)
         );
  NAND2_X1 U5637 ( .A1(n6438), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4532) );
  NAND2_X1 U5638 ( .A1(n6437), .A2(DATAI_2_), .ZN(n4540) );
  OAI211_X1 U5639 ( .C1(n6440), .C2(n4308), .A(n4532), .B(n4540), .ZN(U2926)
         );
  NAND2_X1 U5640 ( .A1(n6438), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4534) );
  OAI211_X1 U5641 ( .C1(n6440), .C2(n4535), .A(n4534), .B(n4533), .ZN(U2944)
         );
  NAND2_X1 U5642 ( .A1(n6438), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4537) );
  OAI211_X1 U5643 ( .C1(n6440), .C2(n5432), .A(n4537), .B(n4536), .ZN(U2942)
         );
  NAND2_X1 U5644 ( .A1(n6438), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4539) );
  OAI211_X1 U5645 ( .C1(n6440), .C2(n4306), .A(n4539), .B(n4538), .ZN(U2930)
         );
  NAND2_X1 U5646 ( .A1(n6438), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4541) );
  OAI211_X1 U5647 ( .C1(n6440), .C2(n5434), .A(n4541), .B(n4540), .ZN(U2941)
         );
  OAI21_X1 U5648 ( .B1(n4542), .B2(n4545), .A(n4544), .ZN(n5486) );
  AOI22_X1 U5649 ( .A1(n4654), .A2(DATAI_10_), .B1(n5406), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4546) );
  OAI21_X1 U5650 ( .B1(n5486), .B2(n5403), .A(n4546), .ZN(U2881) );
  AOI21_X1 U5651 ( .B1(n4548), .B2(n4547), .A(n4542), .ZN(n5307) );
  INV_X1 U5652 ( .A(n5307), .ZN(n4592) );
  AOI22_X1 U5653 ( .A1(n4654), .A2(DATAI_9_), .B1(n5406), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4549) );
  OAI21_X1 U5654 ( .B1(n4592), .B2(n5403), .A(n4549), .ZN(U2882) );
  AOI21_X1 U5655 ( .B1(n4551), .B2(n6461), .A(n4550), .ZN(n5589) );
  INV_X1 U5656 ( .A(n5589), .ZN(n4552) );
  OAI222_X1 U5657 ( .A1(n4552), .A2(n4838), .B1(n4833), .B2(n5371), .C1(n4835), 
        .C2(n5536), .ZN(U2859) );
  NAND2_X1 U5658 ( .A1(n4554), .A2(n4553), .ZN(n4557) );
  INV_X1 U5659 ( .A(n4555), .ZN(n4556) );
  NAND2_X1 U5660 ( .A1(n4557), .A2(n4556), .ZN(n5342) );
  OAI222_X1 U5661 ( .A1(n5342), .A2(n4838), .B1(n4559), .B2(n4833), .C1(n4835), 
        .C2(n4558), .ZN(U2854) );
  XNOR2_X1 U5662 ( .A(n3980), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4561)
         );
  XNOR2_X1 U5663 ( .A(n2953), .B(n4561), .ZN(n5560) );
  NAND2_X1 U5664 ( .A1(n5307), .A2(n5631), .ZN(n4564) );
  NAND2_X1 U5665 ( .A1(n5585), .A2(REIP_REG_9__SCAN_IN), .ZN(n5557) );
  OAI21_X1 U5666 ( .B1(n5530), .B2(n3454), .A(n5557), .ZN(n4562) );
  AOI21_X1 U5667 ( .B1(n5483), .B2(n5308), .A(n4562), .ZN(n4563) );
  OAI211_X1 U5668 ( .C1(n5560), .C2(n5503), .A(n4564), .B(n4563), .ZN(U2977)
         );
  OR2_X1 U5669 ( .A1(n4566), .A2(n4565), .ZN(n4568) );
  NAND2_X1 U5670 ( .A1(n4568), .A2(n4567), .ZN(n5314) );
  OAI22_X1 U5671 ( .A1(n4838), .A2(n5314), .B1(n5315), .B2(n4833), .ZN(n4569)
         );
  AOI21_X1 U5672 ( .B1(n5317), .B2(n5393), .A(n4569), .ZN(n4570) );
  INV_X1 U5673 ( .A(n4570), .ZN(U2851) );
  INV_X1 U5674 ( .A(n4571), .ZN(n4611) );
  OAI222_X1 U5675 ( .A1(n4611), .A2(n4838), .B1(n4573), .B2(n4833), .C1(n4572), 
        .C2(n4835), .ZN(U2856) );
  XOR2_X1 U5676 ( .A(n4575), .B(n2955), .Z(n4584) );
  INV_X1 U5677 ( .A(n5318), .ZN(n4578) );
  INV_X1 U5678 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4576) );
  NOR2_X1 U5679 ( .A1(n5599), .A2(n4576), .ZN(n4583) );
  AOI21_X1 U5680 ( .B1(n5517), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4583), 
        .ZN(n4577) );
  OAI21_X1 U5681 ( .B1(n5525), .B2(n4578), .A(n4577), .ZN(n4579) );
  AOI21_X1 U5682 ( .B1(n4584), .B2(n5533), .A(n4579), .ZN(n4580) );
  OAI21_X1 U5683 ( .B1(n4581), .B2(n6076), .A(n4580), .ZN(U2978) );
  OAI21_X1 U5684 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5553), .ZN(n4587) );
  NOR2_X1 U5685 ( .A1(n5540), .A2(n5314), .ZN(n4582) );
  AOI211_X1 U5686 ( .C1(n5548), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4583), 
        .B(n4582), .ZN(n4586) );
  NAND2_X1 U5687 ( .A1(n4584), .A2(n5591), .ZN(n4585) );
  OAI211_X1 U5688 ( .C1(n4587), .C2(n5552), .A(n4586), .B(n4585), .ZN(U3010)
         );
  OR2_X1 U5689 ( .A1(n4588), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U5690 ( .A1(n4589), .A2(n5284), .ZN(n5549) );
  OAI222_X1 U5691 ( .A1(n5549), .A2(n4838), .B1(n4833), .B2(n4083), .C1(n4835), 
        .C2(n5486), .ZN(U2849) );
  AOI21_X1 U5692 ( .B1(n4591), .B2(n4567), .A(n4590), .ZN(n5559) );
  INV_X1 U5693 ( .A(n5559), .ZN(n4594) );
  OAI222_X1 U5694 ( .A1(n4594), .A2(n4838), .B1(n4593), .B2(n4833), .C1(n4835), 
        .C2(n4592), .ZN(U2850) );
  AOI21_X1 U5695 ( .B1(n4544), .B2(n4596), .A(n4595), .ZN(n5473) );
  INV_X1 U5696 ( .A(n5473), .ZN(n4598) );
  AOI22_X1 U5697 ( .A1(n4654), .A2(DATAI_11_), .B1(n5406), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4597) );
  OAI21_X1 U5698 ( .B1(n4598), .B2(n5403), .A(n4597), .ZN(U2880) );
  OAI21_X1 U5699 ( .B1(n4595), .B2(n4600), .A(n4599), .ZN(n5468) );
  AOI22_X1 U5700 ( .A1(n4654), .A2(DATAI_12_), .B1(n5406), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4601) );
  OAI21_X1 U5701 ( .B1(n5468), .B2(n5403), .A(n4601), .ZN(U2879) );
  INV_X1 U5702 ( .A(n5351), .ZN(n5372) );
  NAND2_X1 U5703 ( .A1(n2977), .A2(n4608), .ZN(n4602) );
  NAND2_X1 U5704 ( .A1(n5336), .A2(n4602), .ZN(n5358) );
  NAND2_X1 U5705 ( .A1(n4603), .A2(n5358), .ZN(n4618) );
  INV_X1 U5706 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U5707 ( .A1(n4607), .A2(n4606), .ZN(n4609) );
  AOI22_X1 U5708 ( .A1(n5353), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n5375), .ZN(n4610) );
  OAI21_X1 U5709 ( .B1(n4611), .B2(n5367), .A(n4610), .ZN(n4615) );
  OAI21_X1 U5710 ( .B1(n5295), .B2(n6394), .A(n5368), .ZN(n4612) );
  NAND2_X1 U5711 ( .A1(n4612), .A2(REIP_REG_2__SCAN_IN), .ZN(n4686) );
  INV_X1 U5712 ( .A(n5345), .ZN(n4613) );
  OAI21_X1 U5713 ( .B1(n5295), .B2(n4613), .A(n5368), .ZN(n5356) );
  AOI21_X1 U5714 ( .B1(n6212), .B2(n4686), .A(n5356), .ZN(n4614) );
  AOI211_X1 U5715 ( .C1(n4616), .C2(n5374), .A(n4615), .B(n4614), .ZN(n4617)
         );
  OAI211_X1 U5716 ( .C1(n6279), .C2(n5372), .A(n4618), .B(n4617), .ZN(U2824)
         );
  OR2_X1 U5717 ( .A1(n4620), .A2(n4619), .ZN(n4621) );
  NAND2_X1 U5718 ( .A1(n4621), .A2(n4666), .ZN(n5280) );
  OAI222_X1 U5719 ( .A1(n5280), .A2(n4838), .B1(n4833), .B2(n4089), .C1(n4835), 
        .C2(n5468), .ZN(U2847) );
  AOI21_X1 U5720 ( .B1(n4599), .B2(n4623), .A(n4622), .ZN(n5386) );
  INV_X1 U5721 ( .A(n5386), .ZN(n4680) );
  AOI22_X1 U5722 ( .A1(n4654), .A2(DATAI_13_), .B1(n5406), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4624) );
  OAI21_X1 U5723 ( .B1(n4680), .B2(n5403), .A(n4624), .ZN(U2878) );
  OAI21_X1 U5724 ( .B1(n4622), .B2(n4627), .A(n4626), .ZN(n5260) );
  AOI22_X1 U5725 ( .A1(n4654), .A2(DATAI_14_), .B1(n5406), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U5726 ( .B1(n5260), .B2(n5403), .A(n4628), .ZN(U2877) );
  INV_X1 U5727 ( .A(n5764), .ZN(n5602) );
  INV_X1 U5728 ( .A(n4629), .ZN(n4732) );
  AOI22_X1 U5729 ( .A1(n4732), .A2(n5369), .B1(n5346), .B2(n6394), .ZN(n4630)
         );
  OAI21_X1 U5730 ( .B1(n5602), .B2(n5372), .A(n4630), .ZN(n4634) );
  INV_X1 U5731 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5732 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5353), .B1(n5295), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n4631) );
  OAI221_X1 U5733 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5359), .C1(n4632), 
        .C2(n5343), .A(n4631), .ZN(n4633) );
  AOI211_X1 U5734 ( .C1(n5522), .C2(n5358), .A(n4634), .B(n4633), .ZN(n4635)
         );
  INV_X1 U5735 ( .A(n4635), .ZN(U2826) );
  INV_X1 U5736 ( .A(n4637), .ZN(n4639) );
  NAND2_X1 U5737 ( .A1(n4639), .A2(n4638), .ZN(n4640) );
  XNOR2_X1 U5738 ( .A(n4636), .B(n4640), .ZN(n5465) );
  INV_X1 U5739 ( .A(n5465), .ZN(n4648) );
  INV_X1 U5740 ( .A(n4642), .ZN(n4959) );
  NOR3_X1 U5741 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n4959), .A3(n4643), 
        .ZN(n4646) );
  AOI21_X1 U5742 ( .B1(n4641), .B2(n5580), .A(n5548), .ZN(n5537) );
  NAND2_X1 U5743 ( .A1(n4643), .A2(n4642), .ZN(n5546) );
  AOI21_X1 U5744 ( .B1(n5537), .B2(n5546), .A(n3985), .ZN(n4645) );
  OAI22_X1 U5745 ( .A1(n5540), .A2(n5280), .B1(n5599), .B2(n5277), .ZN(n4644)
         );
  NOR3_X1 U5746 ( .A1(n4646), .A2(n4645), .A3(n4644), .ZN(n4647) );
  OAI21_X1 U5747 ( .B1(n4648), .B2(n5541), .A(n4647), .ZN(U3006) );
  OR2_X1 U5748 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  NAND2_X1 U5749 ( .A1(n4651), .A2(n4713), .ZN(n5257) );
  OAI222_X1 U5750 ( .A1(n5257), .A2(n4838), .B1(n4833), .B2(n4095), .C1(n4835), 
        .C2(n5260), .ZN(U2845) );
  AOI21_X1 U5751 ( .B1(n4626), .B2(n4653), .A(n4652), .ZN(n5383) );
  INV_X1 U5752 ( .A(n5383), .ZN(n4656) );
  AOI22_X1 U5753 ( .A1(n4654), .A2(DATAI_15_), .B1(n5406), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4655) );
  OAI21_X1 U5754 ( .B1(n4656), .B2(n5403), .A(n4655), .ZN(U2876) );
  OAI21_X1 U5755 ( .B1(n4659), .B2(n4658), .A(n4657), .ZN(n4677) );
  INV_X1 U5756 ( .A(n4677), .ZN(n4674) );
  NOR3_X1 U5757 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4660), .A3(n4669), 
        .ZN(n4665) );
  AND2_X1 U5758 ( .A1(n4662), .A2(n4661), .ZN(n5593) );
  INV_X1 U5759 ( .A(n5593), .ZN(n4663) );
  AOI21_X1 U5760 ( .B1(n4669), .B2(n4663), .A(n4665), .ZN(n4664) );
  OAI211_X1 U5761 ( .C1(n4701), .C2(n5595), .A(n5537), .B(n4664), .ZN(n4696)
         );
  OAI21_X1 U5762 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4665), .A(n4696), 
        .ZN(n4673) );
  AOI21_X1 U5763 ( .B1(n4667), .B2(n4666), .A(n4649), .ZN(n5385) );
  INV_X1 U5764 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6228) );
  NOR2_X1 U5765 ( .A1(n5599), .A2(n6228), .ZN(n4671) );
  NOR3_X1 U5766 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4669), .A3(n4668), 
        .ZN(n4670) );
  AOI211_X1 U5767 ( .C1(n5385), .C2(n5590), .A(n4671), .B(n4670), .ZN(n4672)
         );
  OAI211_X1 U5768 ( .C1(n4674), .C2(n5541), .A(n4673), .B(n4672), .ZN(U3005)
         );
  OAI22_X1 U5769 ( .A1(n5530), .A2(n4675), .B1(n5599), .B2(n6228), .ZN(n4676)
         );
  AOI21_X1 U5770 ( .B1(n5483), .B2(n5271), .A(n4676), .ZN(n4679) );
  NAND2_X1 U5771 ( .A1(n4677), .A2(n5533), .ZN(n4678) );
  OAI211_X1 U5772 ( .C1(n4680), .C2(n6076), .A(n4679), .B(n4678), .ZN(U2973)
         );
  INV_X1 U5773 ( .A(n4681), .ZN(n5513) );
  XNOR2_X1 U5774 ( .A(n4682), .B(n4683), .ZN(n5391) );
  OAI21_X1 U5775 ( .B1(n5275), .B2(n6394), .A(n6423), .ZN(n4685) );
  OAI22_X1 U5776 ( .A1(n5359), .A2(n5516), .B1(n4419), .B2(n5372), .ZN(n4684)
         );
  AOI21_X1 U5777 ( .B1(n4686), .B2(n4685), .A(n4684), .ZN(n4687) );
  OAI21_X1 U5778 ( .B1(n5391), .B2(n5367), .A(n4687), .ZN(n4689) );
  OAI22_X1 U5779 ( .A1(n5395), .A2(n5370), .B1(n3325), .B2(n5343), .ZN(n4688)
         );
  AOI211_X1 U5780 ( .C1(n5513), .C2(n5358), .A(n4689), .B(n4688), .ZN(n4690)
         );
  INV_X1 U5781 ( .A(n4690), .ZN(U2825) );
  OR2_X1 U5782 ( .A1(n4692), .A2(n4691), .ZN(n4693) );
  NAND2_X1 U5783 ( .A1(n4693), .A2(n5191), .ZN(n5247) );
  OAI21_X1 U5784 ( .B1(n4652), .B2(n4695), .A(n4694), .ZN(n5404) );
  OAI222_X1 U5785 ( .A1(n5247), .A2(n4838), .B1(n4833), .B2(n4101), .C1(n4835), 
        .C2(n5404), .ZN(U2843) );
  INV_X1 U5786 ( .A(n4696), .ZN(n4706) );
  XNOR2_X1 U5787 ( .A(n3980), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4698)
         );
  XNOR2_X1 U5788 ( .A(n4697), .B(n4698), .ZN(n5158) );
  NAND2_X1 U5789 ( .A1(n5158), .A2(n5591), .ZN(n4704) );
  NOR2_X1 U5790 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4959), .ZN(n4702)
         );
  INV_X1 U5791 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4699) );
  OAI22_X1 U5792 ( .A1(n5540), .A2(n5257), .B1(n5599), .B2(n4699), .ZN(n4700)
         );
  AOI21_X1 U5793 ( .B1(n4702), .B2(n4701), .A(n4700), .ZN(n4703) );
  OAI211_X1 U5794 ( .C1(n4706), .C2(n4705), .A(n4704), .B(n4703), .ZN(U3004)
         );
  INV_X1 U5795 ( .A(n4708), .ZN(n4710) );
  NAND2_X1 U5796 ( .A1(n4710), .A2(n4709), .ZN(n4711) );
  XNOR2_X1 U5797 ( .A(n4707), .B(n4711), .ZN(n4725) );
  INV_X1 U5798 ( .A(n4958), .ZN(n4712) );
  OAI21_X1 U5799 ( .B1(n4949), .B2(n4712), .A(n5537), .ZN(n4957) );
  AOI21_X1 U5800 ( .B1(n4714), .B2(n4713), .A(n4691), .ZN(n5382) );
  INV_X1 U5801 ( .A(n5382), .ZN(n4717) );
  NOR2_X1 U5802 ( .A1(n4959), .A2(n4958), .ZN(n4715) );
  NAND2_X1 U5803 ( .A1(n4715), .A2(n4960), .ZN(n4716) );
  NAND2_X1 U5804 ( .A1(n5585), .A2(REIP_REG_15__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5805 ( .C1(n5540), .C2(n4717), .A(n4716), .B(n4720), .ZN(n4718)
         );
  AOI21_X1 U5806 ( .B1(n4957), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n4718), 
        .ZN(n4719) );
  OAI21_X1 U5807 ( .B1(n4725), .B2(n5541), .A(n4719), .ZN(U3003) );
  NAND2_X1 U5808 ( .A1(n5250), .A2(n5483), .ZN(n4721) );
  OAI211_X1 U5809 ( .C1(n5530), .C2(n4722), .A(n4721), .B(n4720), .ZN(n4723)
         );
  AOI21_X1 U5810 ( .B1(n5383), .B2(n5631), .A(n4723), .ZN(n4724) );
  OAI21_X1 U5811 ( .B1(n5503), .B2(n4725), .A(n4724), .ZN(U2971) );
  OAI21_X1 U5812 ( .B1(n4726), .B2(n4729), .A(n4728), .ZN(n5230) );
  AOI22_X1 U5813 ( .A1(n5407), .A2(DATAI_2_), .B1(n5406), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5814 ( .A1(n5396), .A2(DATAI_18_), .ZN(n4730) );
  OAI211_X1 U5815 ( .C1(n5230), .C2(n5403), .A(n4731), .B(n4730), .ZN(U2873)
         );
  XNOR2_X1 U5816 ( .A(n4732), .B(n5207), .ZN(n5584) );
  AOI22_X1 U5817 ( .A1(n5392), .A2(n5584), .B1(n4774), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4733) );
  OAI21_X1 U5818 ( .B1(n4734), .B2(n4835), .A(n4733), .ZN(U2858) );
  INV_X1 U5819 ( .A(n4735), .ZN(n5339) );
  AOI22_X1 U5820 ( .A1(n5392), .A2(n5339), .B1(n4774), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4736) );
  OAI21_X1 U5821 ( .B1(n5500), .B2(n4835), .A(n4736), .ZN(U2853) );
  XOR2_X1 U5822 ( .A(n4737), .B(n4738), .Z(n5110) );
  INV_X1 U5823 ( .A(n5110), .ZN(n4744) );
  MUX2_X1 U5824 ( .A(n4740), .B(n4052), .S(n4739), .Z(n4742) );
  XNOR2_X1 U5825 ( .A(n4742), .B(n4741), .ZN(n5066) );
  AOI22_X1 U5826 ( .A1(n5392), .A2(n5066), .B1(n4774), .B2(EBX_REG_20__SCAN_IN), .ZN(n4743) );
  OAI21_X1 U5827 ( .B1(n4744), .B2(n4835), .A(n4743), .ZN(U2839) );
  INV_X1 U5828 ( .A(n4746), .ZN(n4747) );
  OAI21_X1 U5829 ( .B1(n4748), .B2(n4804), .A(n4747), .ZN(n5119) );
  OR2_X1 U5830 ( .A1(n4749), .A2(n4750), .ZN(n4751) );
  NAND2_X1 U5831 ( .A1(n4799), .A2(n4751), .ZN(n5020) );
  INV_X1 U5832 ( .A(n5020), .ZN(n4916) );
  AOI22_X1 U5833 ( .A1(n5392), .A2(n4916), .B1(n4774), .B2(EBX_REG_26__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5834 ( .B1(n5119), .B2(n4835), .A(n4752), .ZN(U2833) );
  INV_X1 U5835 ( .A(n4754), .ZN(n4755) );
  NAND2_X1 U5836 ( .A1(n4756), .A2(n4755), .ZN(n4829) );
  XOR2_X1 U5837 ( .A(n4753), .B(n4829), .Z(n5226) );
  AOI22_X1 U5838 ( .A1(n5226), .A2(n5392), .B1(n4774), .B2(EBX_REG_18__SCAN_IN), .ZN(n4757) );
  OAI21_X1 U5839 ( .B1(n5230), .B2(n4835), .A(n4757), .ZN(U2841) );
  OR2_X1 U5840 ( .A1(n4759), .A2(n4758), .ZN(n4760) );
  NAND2_X1 U5841 ( .A1(n4760), .A2(n4553), .ZN(n5366) );
  INV_X1 U5842 ( .A(n5366), .ZN(n4761) );
  AOI22_X1 U5843 ( .A1(n5392), .A2(n4761), .B1(n4774), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4762) );
  OAI21_X1 U5844 ( .B1(n5361), .B2(n4835), .A(n4762), .ZN(U2855) );
  NOR2_X1 U5845 ( .A1(n4763), .A2(n4764), .ZN(n4765) );
  OR2_X1 U5846 ( .A1(n4262), .A2(n4765), .ZN(n5096) );
  NOR2_X1 U5847 ( .A1(n4766), .A2(n4767), .ZN(n4768) );
  OR2_X1 U5848 ( .A1(n4811), .A2(n4768), .ZN(n5050) );
  OAI22_X1 U5849 ( .A1(n5050), .A2(n4838), .B1(n5043), .B2(n4833), .ZN(n4769)
         );
  INV_X1 U5850 ( .A(n4769), .ZN(n4770) );
  OAI21_X1 U5851 ( .B1(n5096), .B2(n4835), .A(n4770), .ZN(U2836) );
  NAND2_X1 U5852 ( .A1(n4801), .A2(n4771), .ZN(n4772) );
  NAND2_X1 U5853 ( .A1(n4773), .A2(n4772), .ZN(n5002) );
  INV_X1 U5854 ( .A(n5002), .ZN(n4775) );
  AOI22_X1 U5855 ( .A1(n5392), .A2(n4775), .B1(n4774), .B2(EBX_REG_28__SCAN_IN), .ZN(n4776) );
  OAI21_X1 U5856 ( .B1(n5003), .B2(n4835), .A(n4776), .ZN(U2831) );
  NAND2_X1 U5857 ( .A1(n4777), .A2(n3302), .ZN(n5634) );
  NOR2_X2 U5858 ( .A1(n4778), .A2(n5630), .ZN(n6124) );
  AOI22_X1 U5859 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5703), .B1(n6124), 
        .B2(n5702), .ZN(n4780) );
  AND2_X1 U5860 ( .A1(n5631), .A2(DATAI_23_), .ZN(n6128) );
  AND2_X1 U5861 ( .A1(n5631), .A2(DATAI_31_), .ZN(n6066) );
  AOI22_X1 U5862 ( .A1(n5726), .A2(n6128), .B1(n5700), .B2(n6066), .ZN(n4779)
         );
  OAI211_X1 U5863 ( .C1(n4781), .C2(n5634), .A(n4780), .B(n4779), .ZN(U3051)
         );
  INV_X1 U5864 ( .A(n4782), .ZN(n4793) );
  NOR3_X1 U5865 ( .A1(n4785), .A2(n4784), .A3(n4783), .ZN(n4788) );
  NOR2_X1 U5866 ( .A1(n4786), .A2(n6273), .ZN(n4787) );
  AOI211_X1 U5867 ( .C1(n4790), .C2(n4789), .A(n4788), .B(n4787), .ZN(n4791)
         );
  OAI22_X1 U5868 ( .A1(n4793), .A2(n3013), .B1(n4792), .B2(n4791), .ZN(U3459)
         );
  INV_X1 U5869 ( .A(n4888), .ZN(n4795) );
  OAI22_X1 U5870 ( .A1(n4795), .A2(n4838), .B1(n4833), .B2(n4794), .ZN(U2828)
         );
  INV_X1 U5871 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4797) );
  OAI222_X1 U5872 ( .A1(n5000), .A2(n4838), .B1(n4797), .B2(n4833), .C1(n4835), 
        .C2(n4796), .ZN(U2830) );
  NAND2_X1 U5873 ( .A1(n4799), .A2(n4798), .ZN(n4800) );
  NAND2_X1 U5874 ( .A1(n4801), .A2(n4800), .ZN(n5018) );
  OR2_X1 U5875 ( .A1(n4746), .A2(n4802), .ZN(n4803) );
  OAI222_X1 U5876 ( .A1(n5018), .A2(n4838), .B1(n4833), .B2(n4135), .C1(n4835), 
        .C2(n5086), .ZN(U2832) );
  AOI21_X1 U5877 ( .B1(n4805), .B2(n4263), .A(n4804), .ZN(n5121) );
  INV_X1 U5878 ( .A(n5121), .ZN(n4810) );
  AOI21_X1 U5879 ( .B1(n4807), .B2(n4806), .A(n4749), .ZN(n5163) );
  INV_X1 U5880 ( .A(n5163), .ZN(n4808) );
  OAI222_X1 U5881 ( .A1(n4810), .A2(n4835), .B1(n4809), .B2(n4833), .C1(n4838), 
        .C2(n4808), .ZN(U2834) );
  XOR2_X1 U5882 ( .A(n4812), .B(n4811), .Z(n5037) );
  INV_X1 U5883 ( .A(n5037), .ZN(n4814) );
  OAI222_X1 U5884 ( .A1(n4815), .A2(n4835), .B1(n4838), .B2(n4814), .C1(n4833), 
        .C2(n4813), .ZN(U2835) );
  NOR2_X1 U5885 ( .A1(n4816), .A2(n4817), .ZN(n4818) );
  OR2_X1 U5886 ( .A1(n4766), .A2(n4818), .ZN(n5053) );
  NOR2_X1 U5887 ( .A1(n4819), .A2(n4820), .ZN(n4821) );
  OR2_X1 U5888 ( .A1(n4763), .A2(n4821), .ZN(n5101) );
  OAI222_X1 U5889 ( .A1(n5053), .A2(n4838), .B1(n4833), .B2(n4118), .C1(n4835), 
        .C2(n5101), .ZN(U2837) );
  AND2_X1 U5890 ( .A1(n4823), .A2(n4822), .ZN(n4824) );
  OR2_X1 U5891 ( .A1(n4824), .A2(n4816), .ZN(n5169) );
  AND2_X1 U5892 ( .A1(n4826), .A2(n4825), .ZN(n4827) );
  OR2_X1 U5893 ( .A1(n4827), .A2(n4819), .ZN(n5106) );
  OAI222_X1 U5894 ( .A1(n5169), .A2(n4838), .B1(n4828), .B2(n4833), .C1(n4835), 
        .C2(n5106), .ZN(U2838) );
  NAND2_X1 U5895 ( .A1(n4753), .A2(n4829), .ZN(n4830) );
  XOR2_X1 U5896 ( .A(n4831), .B(n4830), .Z(n5176) );
  AOI21_X1 U5897 ( .B1(n4728), .B2(n4832), .A(n4737), .ZN(n5138) );
  INV_X1 U5898 ( .A(n5138), .ZN(n4834) );
  OAI22_X1 U5899 ( .A1(n4835), .A2(n4834), .B1(n5081), .B2(n4833), .ZN(n4836)
         );
  INV_X1 U5900 ( .A(n4836), .ZN(n4837) );
  OAI21_X1 U5901 ( .B1(n5176), .B2(n4838), .A(n4837), .ZN(U2840) );
  NAND3_X1 U5902 ( .A1(n4853), .A2(n4840), .A3(n4839), .ZN(n4842) );
  AOI22_X1 U5903 ( .A1(n5396), .A2(DATAI_31_), .B1(n5406), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U5904 ( .A1(n4842), .A2(n4841), .ZN(U2860) );
  AOI22_X1 U5905 ( .A1(n5407), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5406), .ZN(n4844) );
  NAND2_X1 U5906 ( .A1(n5396), .A2(DATAI_28_), .ZN(n4843) );
  OAI211_X1 U5907 ( .C1(n5003), .C2(n5403), .A(n4844), .B(n4843), .ZN(U2863)
         );
  AOI22_X1 U5908 ( .A1(n5407), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5406), .ZN(n4846) );
  NAND2_X1 U5909 ( .A1(n5396), .A2(DATAI_26_), .ZN(n4845) );
  OAI211_X1 U5910 ( .C1(n5119), .C2(n5403), .A(n4846), .B(n4845), .ZN(U2865)
         );
  NOR4_X1 U5911 ( .A1(n4847), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4848), .ZN(n4849) );
  AOI21_X1 U5912 ( .B1(n4850), .B2(n4883), .A(n4849), .ZN(n4851) );
  INV_X1 U5913 ( .A(n4851), .ZN(n4852) );
  XNOR2_X1 U5914 ( .A(n4852), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4892)
         );
  NAND2_X1 U5915 ( .A1(n4853), .A2(n5631), .ZN(n4857) );
  NOR2_X1 U5916 ( .A1(n5599), .A2(n6258), .ZN(n4887) );
  NOR2_X1 U5917 ( .A1(n5525), .A2(n4854), .ZN(n4855) );
  AOI211_X1 U5918 ( .C1(n5517), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4887), 
        .B(n4855), .ZN(n4856) );
  OAI211_X1 U5919 ( .C1(n4892), .C2(n5503), .A(n4857), .B(n4856), .ZN(U2955)
         );
  NAND2_X1 U5920 ( .A1(n4859), .A2(n4858), .ZN(n4860) );
  XOR2_X1 U5921 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n4860), .Z(n4902) );
  NAND2_X1 U5922 ( .A1(n5585), .A2(REIP_REG_27__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5923 ( .A1(n5517), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4861)
         );
  OAI211_X1 U5924 ( .C1(n5525), .C2(n5013), .A(n4905), .B(n4861), .ZN(n4862)
         );
  AOI21_X1 U5925 ( .B1(n4902), .B2(n5533), .A(n4862), .ZN(n4863) );
  OAI21_X1 U5926 ( .B1(n5086), .B2(n6076), .A(n4863), .ZN(U2959) );
  INV_X1 U5927 ( .A(n4871), .ZN(n4866) );
  INV_X1 U5928 ( .A(n4927), .ZN(n4865) );
  OAI22_X1 U5929 ( .A1(n5125), .A2(n4866), .B1(n4865), .B2(n4864), .ZN(n4867)
         );
  XNOR2_X1 U5930 ( .A(n4867), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4934)
         );
  INV_X1 U5931 ( .A(n5096), .ZN(n5047) );
  NAND2_X1 U5932 ( .A1(n5585), .A2(REIP_REG_23__SCAN_IN), .ZN(n4930) );
  NAND2_X1 U5933 ( .A1(n5517), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4868)
         );
  OAI211_X1 U5934 ( .C1(n5042), .C2(n5525), .A(n4930), .B(n4868), .ZN(n4869)
         );
  AOI21_X1 U5935 ( .B1(n5047), .B2(n5631), .A(n4869), .ZN(n4870) );
  OAI21_X1 U5936 ( .B1(n4934), .B2(n5503), .A(n4870), .ZN(U2963) );
  AOI21_X1 U5937 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3980), .A(n4871), 
        .ZN(n4872) );
  XNOR2_X1 U5938 ( .A(n4873), .B(n4872), .ZN(n4942) );
  NAND2_X1 U5939 ( .A1(n5585), .A2(REIP_REG_22__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U5940 ( .B1(n5530), .B2(n6412), .A(n4936), .ZN(n4875) );
  NOR2_X1 U5941 ( .A1(n5101), .A2(n6076), .ZN(n4874) );
  AOI211_X1 U5942 ( .C1(n5052), .C2(n5483), .A(n4875), .B(n4874), .ZN(n4876)
         );
  OAI21_X1 U5943 ( .B1(n4942), .B2(n5503), .A(n4876), .ZN(U2964) );
  XNOR2_X1 U5944 ( .A(n4878), .B(n4877), .ZN(n4952) );
  INV_X1 U5945 ( .A(n5069), .ZN(n4880) );
  NAND2_X1 U5946 ( .A1(n5585), .A2(REIP_REG_20__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U5947 ( .A1(n5517), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4879)
         );
  OAI211_X1 U5948 ( .C1(n4880), .C2(n5525), .A(n4943), .B(n4879), .ZN(n4881)
         );
  AOI21_X1 U5949 ( .B1(n5110), .B2(n5631), .A(n4881), .ZN(n4882) );
  OAI21_X1 U5950 ( .B1(n4952), .B2(n5503), .A(n4882), .ZN(U2966) );
  INV_X1 U5951 ( .A(n4883), .ZN(n4884) );
  NOR3_X1 U5952 ( .A1(n4885), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4884), 
        .ZN(n4886) );
  AOI211_X1 U5953 ( .C1(n5590), .C2(n4888), .A(n4887), .B(n4886), .ZN(n4891)
         );
  NAND2_X1 U5954 ( .A1(n4889), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4890) );
  OAI211_X1 U5955 ( .C1(n4892), .C2(n5541), .A(n4891), .B(n4890), .ZN(U2987)
         );
  INV_X1 U5956 ( .A(n4893), .ZN(n4901) );
  OAI21_X1 U5957 ( .B1(n5540), .B2(n5002), .A(n4894), .ZN(n4899) );
  INV_X1 U5958 ( .A(n4904), .ZN(n4897) );
  NOR3_X1 U5959 ( .A1(n4897), .A2(n4896), .A3(n4895), .ZN(n4898) );
  AOI211_X1 U5960 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n4908), .A(n4899), .B(n4898), .ZN(n4900) );
  OAI21_X1 U5961 ( .B1(n4901), .B2(n5541), .A(n4900), .ZN(U2990) );
  INV_X1 U5962 ( .A(n4902), .ZN(n4910) );
  INV_X1 U5963 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5964 ( .A1(n4904), .A2(n4903), .ZN(n4906) );
  OAI211_X1 U5965 ( .C1(n5018), .C2(n5540), .A(n4906), .B(n4905), .ZN(n4907)
         );
  AOI21_X1 U5966 ( .B1(n4908), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4907), 
        .ZN(n4909) );
  OAI21_X1 U5967 ( .B1(n4910), .B2(n5541), .A(n4909), .ZN(U2991) );
  NOR2_X1 U5968 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  XNOR2_X1 U5969 ( .A(n3999), .B(n4913), .ZN(n5116) );
  AOI211_X1 U5970 ( .C1(n4919), .C2(n5167), .A(n4914), .B(n5161), .ZN(n4915)
         );
  AOI21_X1 U5971 ( .B1(n5585), .B2(REIP_REG_26__SCAN_IN), .A(n4915), .ZN(n4918) );
  NAND2_X1 U5972 ( .A1(n5590), .A2(n4916), .ZN(n4917) );
  OAI211_X1 U5973 ( .C1(n5168), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4920)
         );
  AOI21_X1 U5974 ( .B1(n5116), .B2(n5591), .A(n4920), .ZN(n4921) );
  INV_X1 U5975 ( .A(n4921), .ZN(U2992) );
  INV_X1 U5976 ( .A(n5182), .ZN(n4928) );
  NAND3_X1 U5977 ( .A1(n4928), .A2(n4927), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4922) );
  AOI21_X1 U5978 ( .B1(n4260), .B2(n4922), .A(n5168), .ZN(n4923) );
  AOI211_X1 U5979 ( .C1(n5037), .C2(n5590), .A(n4924), .B(n4923), .ZN(n4925)
         );
  OAI21_X1 U5980 ( .B1(n4926), .B2(n5541), .A(n4925), .ZN(U2994) );
  INV_X1 U5981 ( .A(n5050), .ZN(n4932) );
  NAND3_X1 U5982 ( .A1(n4928), .A2(n4927), .A3(n6354), .ZN(n4929) );
  OAI211_X1 U5983 ( .C1(n4935), .C2(n6354), .A(n4930), .B(n4929), .ZN(n4931)
         );
  AOI21_X1 U5984 ( .B1(n4932), .B2(n5590), .A(n4931), .ZN(n4933) );
  OAI21_X1 U5985 ( .B1(n4934), .B2(n5541), .A(n4933), .ZN(U2995) );
  INV_X1 U5986 ( .A(n4935), .ZN(n4940) );
  OAI21_X1 U5987 ( .B1(n4937), .B2(n6455), .A(n4936), .ZN(n4939) );
  NOR2_X1 U5988 ( .A1(n5053), .A2(n5540), .ZN(n4938) );
  AOI211_X1 U5989 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n4940), .A(n4939), .B(n4938), .ZN(n4941) );
  OAI21_X1 U5990 ( .B1(n4942), .B2(n5541), .A(n4941), .ZN(U2996) );
  INV_X1 U5991 ( .A(n4943), .ZN(n4947) );
  NOR3_X1 U5992 ( .A1(n4945), .A2(n4944), .A3(n5182), .ZN(n4946) );
  AOI211_X1 U5993 ( .C1(n5590), .C2(n5066), .A(n4947), .B(n4946), .ZN(n4951)
         );
  AOI21_X1 U5994 ( .B1(n5183), .B2(n4948), .A(n5190), .ZN(n5189) );
  OAI21_X1 U5995 ( .B1(n4949), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5189), 
        .ZN(n5179) );
  NAND2_X1 U5996 ( .A1(n5179), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4950) );
  OAI211_X1 U5997 ( .C1(n4952), .C2(n5541), .A(n4951), .B(n4950), .ZN(U2998)
         );
  NOR2_X1 U5998 ( .A1(n3980), .A2(n3987), .ZN(n5149) );
  AOI21_X1 U5999 ( .B1(n3987), .B2(n3980), .A(n5149), .ZN(n4955) );
  BUF_X1 U6000 ( .A(n4953), .Z(n4954) );
  XOR2_X1 U6001 ( .A(n4955), .B(n4954), .Z(n5155) );
  INV_X1 U6002 ( .A(n5155), .ZN(n4965) );
  OAI22_X1 U6003 ( .A1(n5540), .A2(n5247), .B1(n5599), .B2(n6230), .ZN(n4956)
         );
  AOI21_X1 U6004 ( .B1(n4957), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n4956), 
        .ZN(n4964) );
  AOI211_X1 U6005 ( .C1(n4960), .C2(n3987), .A(n4959), .B(n4958), .ZN(n4962)
         );
  NAND2_X1 U6006 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  OAI211_X1 U6007 ( .C1(n4965), .C2(n5541), .A(n4964), .B(n4963), .ZN(U3002)
         );
  OR3_X1 U6008 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4966), .A3(n5568), 
        .ZN(n4975) );
  XOR2_X1 U6009 ( .A(n4967), .B(n4969), .Z(n5501) );
  NAND2_X1 U6010 ( .A1(n5585), .A2(REIP_REG_5__SCAN_IN), .ZN(n5507) );
  OAI21_X1 U6011 ( .B1(n5540), .B2(n5342), .A(n5507), .ZN(n4970) );
  AOI21_X1 U6012 ( .B1(n5501), .B2(n5591), .A(n4970), .ZN(n4974) );
  OAI221_X1 U6013 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5582), .C1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n4972), .A(n4971), .ZN(n4973) );
  NAND3_X1 U6014 ( .A1(n4975), .A2(n4974), .A3(n4973), .ZN(U3013) );
  OAI211_X1 U6015 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4977), .B(n4976), .ZN(n4984) );
  NOR2_X1 U6016 ( .A1(n5540), .A2(n5366), .ZN(n4978) );
  AOI211_X1 U6017 ( .C1(n4980), .C2(n5591), .A(n4979), .B(n4978), .ZN(n4983)
         );
  NAND2_X1 U6018 ( .A1(n4981), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4982)
         );
  NAND3_X1 U6019 ( .A1(n4984), .A2(n4983), .A3(n4982), .ZN(U3014) );
  AND2_X1 U6020 ( .A1(n5437), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI22_X1 U6021 ( .A1(n4985), .A2(n5370), .B1(n4011), .B2(n5343), .ZN(n4986)
         );
  AOI211_X1 U6022 ( .C1(n4988), .C2(n5374), .A(n4987), .B(n4986), .ZN(n4992)
         );
  OAI211_X1 U6023 ( .C1(n4993), .C2(n5336), .A(n4992), .B(n4991), .ZN(U2797)
         );
  AOI22_X1 U6024 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5375), .ZN(n4994) );
  INV_X1 U6025 ( .A(n4994), .ZN(n4997) );
  OAI22_X1 U6026 ( .A1(n5006), .A2(n6254), .B1(n4995), .B2(n5359), .ZN(n4996)
         );
  OAI211_X1 U6027 ( .C1(n5367), .C2(n5000), .A(n4999), .B(n4998), .ZN(U2798)
         );
  AOI22_X1 U6028 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5375), .B1(n5001), 
        .B2(n5374), .ZN(n5011) );
  OAI22_X1 U6029 ( .A1(n5003), .A2(n5336), .B1(n5002), .B2(n5367), .ZN(n5009)
         );
  INV_X1 U6030 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6249) );
  NOR3_X1 U6031 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6249), .A3(n5014), .ZN(n5008) );
  INV_X1 U6032 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5005) );
  OAI22_X1 U6033 ( .A1(n5006), .A2(n5005), .B1(n5004), .B2(n5370), .ZN(n5007)
         );
  NOR3_X1 U6034 ( .A1(n5009), .A2(n5008), .A3(n5007), .ZN(n5010) );
  NAND2_X1 U6035 ( .A1(n5011), .A2(n5010), .ZN(U2799) );
  AOI22_X1 U6036 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5375), .B1(
        REIP_REG_27__SCAN_IN), .B2(n5023), .ZN(n5012) );
  OAI21_X1 U6037 ( .B1(n5013), .B2(n5359), .A(n5012), .ZN(n5016) );
  OAI22_X1 U6038 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5014), .B1(n5086), .B2(
        n5336), .ZN(n5015) );
  OAI21_X1 U6039 ( .B1(n5018), .B2(n5367), .A(n5017), .ZN(U2800) );
  AOI22_X1 U6040 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5375), .B1(n5115), 
        .B2(n5374), .ZN(n5025) );
  NAND2_X1 U6041 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5032), .ZN(n5028) );
  OAI21_X1 U6042 ( .B1(n6246), .B2(n5028), .A(n5019), .ZN(n5022) );
  OAI22_X1 U6043 ( .A1(n5119), .A2(n5336), .B1(n5020), .B2(n5367), .ZN(n5021)
         );
  AOI21_X1 U6044 ( .B1(n5023), .B2(n5022), .A(n5021), .ZN(n5024) );
  OAI211_X1 U6045 ( .C1(n5026), .C2(n5370), .A(n5025), .B(n5024), .ZN(U2801)
         );
  AOI22_X1 U6046 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5375), .ZN(n5027) );
  INV_X1 U6047 ( .A(n5027), .ZN(n5030) );
  OAI22_X1 U6048 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5028), .B1(n5124), .B2(
        n5359), .ZN(n5029) );
  AOI211_X1 U6049 ( .C1(n5163), .C2(n5369), .A(n5030), .B(n5029), .ZN(n5035)
         );
  NOR2_X1 U6050 ( .A1(n5330), .A2(n5031), .ZN(n5046) );
  NAND2_X1 U6051 ( .A1(n6364), .A2(n5032), .ZN(n5038) );
  INV_X1 U6052 ( .A(n5038), .ZN(n5033) );
  OAI21_X1 U6053 ( .B1(n5046), .B2(n5033), .A(REIP_REG_25__SCAN_IN), .ZN(n5034) );
  OAI211_X1 U6054 ( .C1(n5336), .C2(n4810), .A(n5035), .B(n5034), .ZN(U2802)
         );
  AOI22_X1 U6055 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5375), .ZN(n5041) );
  AOI22_X1 U6056 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5046), .B1(n5036), .B2(
        n5374), .ZN(n5040) );
  AOI22_X1 U6057 ( .A1(n5037), .A2(n5369), .B1(n5092), .B2(n5328), .ZN(n5039)
         );
  NAND4_X1 U6058 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(U2803)
         );
  OAI22_X1 U6059 ( .A1(n5043), .A2(n5370), .B1(n5042), .B2(n5359), .ZN(n5044)
         );
  AOI21_X1 U6060 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5375), .A(n5044), 
        .ZN(n5049) );
  NAND2_X1 U6061 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5056) );
  INV_X1 U6062 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U6063 ( .B1(n5056), .B2(n5055), .A(n6243), .ZN(n5045) );
  AOI22_X1 U6064 ( .A1(n5047), .A2(n5328), .B1(n5046), .B2(n5045), .ZN(n5048)
         );
  OAI211_X1 U6065 ( .C1(n5050), .C2(n5367), .A(n5049), .B(n5048), .ZN(U2804)
         );
  AOI22_X1 U6066 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5375), .ZN(n5060) );
  AND2_X1 U6067 ( .A1(n5368), .A2(n5051), .ZN(n5067) );
  AOI22_X1 U6068 ( .A1(n5052), .A2(n5374), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5067), .ZN(n5059) );
  OAI22_X1 U6069 ( .A1(n5101), .A2(n5336), .B1(n5053), .B2(n5367), .ZN(n5054)
         );
  INV_X1 U6070 ( .A(n5054), .ZN(n5058) );
  INV_X1 U6071 ( .A(n5055), .ZN(n5063) );
  OAI211_X1 U6072 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5063), .B(n5056), .ZN(n5057) );
  NAND4_X1 U6073 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(U2805)
         );
  INV_X1 U6074 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6239) );
  AOI22_X1 U6075 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5375), .ZN(n5061) );
  OAI21_X1 U6076 ( .B1(n5129), .B2(n5359), .A(n5061), .ZN(n5062) );
  AOI221_X1 U6077 ( .B1(n5067), .B2(REIP_REG_21__SCAN_IN), .C1(n5063), .C2(
        n6239), .A(n5062), .ZN(n5065) );
  INV_X1 U6078 ( .A(n5106), .ZN(n5131) );
  NAND2_X1 U6079 ( .A1(n5131), .A2(n5328), .ZN(n5064) );
  OAI211_X1 U6080 ( .C1(n5367), .C2(n5169), .A(n5065), .B(n5064), .ZN(U2806)
         );
  AOI22_X1 U6081 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5353), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5375), .ZN(n5073) );
  AOI22_X1 U6082 ( .A1(n5110), .A2(n5328), .B1(n5066), .B2(n5369), .ZN(n5072)
         );
  OAI21_X1 U6083 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5068), .A(n5067), .ZN(n5071) );
  NAND2_X1 U6084 ( .A1(n5069), .A2(n5374), .ZN(n5070) );
  NAND4_X1 U6085 ( .A1(n5073), .A2(n5072), .A3(n5071), .A4(n5070), .ZN(U2807)
         );
  NOR2_X2 U6086 ( .A1(n5295), .A2(n6316), .ZN(n5354) );
  INV_X1 U6087 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6237) );
  OR2_X1 U6088 ( .A1(n5330), .A2(n5074), .ZN(n5233) );
  OAI21_X1 U6089 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5075), .ZN(n5076) );
  OAI22_X1 U6090 ( .A1(n6237), .A2(n5233), .B1(n5224), .B2(n5076), .ZN(n5077)
         );
  AOI211_X1 U6091 ( .C1(n5375), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5354), 
        .B(n5077), .ZN(n5080) );
  OAI22_X1 U6092 ( .A1(n5176), .A2(n5367), .B1(n5136), .B2(n5359), .ZN(n5078)
         );
  AOI21_X1 U6093 ( .B1(n5138), .B2(n5328), .A(n5078), .ZN(n5079) );
  OAI211_X1 U6094 ( .C1(n5081), .C2(n5370), .A(n5080), .B(n5079), .ZN(U2808)
         );
  AOI22_X1 U6095 ( .A1(n5082), .A2(n5397), .B1(n5396), .B2(DATAI_29_), .ZN(
        n5084) );
  AOI22_X1 U6096 ( .A1(n5407), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5406), .ZN(n5083) );
  NAND2_X1 U6097 ( .A1(n5084), .A2(n5083), .ZN(U2862) );
  INV_X1 U6098 ( .A(n5396), .ZN(n5402) );
  INV_X1 U6099 ( .A(DATAI_27_), .ZN(n5085) );
  OAI22_X1 U6100 ( .A1(n5086), .A2(n5403), .B1(n5402), .B2(n5085), .ZN(n5087)
         );
  INV_X1 U6101 ( .A(n5087), .ZN(n5089) );
  AOI22_X1 U6102 ( .A1(n5407), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5406), .ZN(n5088) );
  NAND2_X1 U6103 ( .A1(n5089), .A2(n5088), .ZN(U2864) );
  AOI22_X1 U6104 ( .A1(n5121), .A2(n5397), .B1(n5396), .B2(DATAI_25_), .ZN(
        n5091) );
  AOI22_X1 U6105 ( .A1(n5407), .A2(DATAI_9_), .B1(n5406), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6106 ( .A1(n5091), .A2(n5090), .ZN(U2866) );
  AOI22_X1 U6107 ( .A1(n5092), .A2(n5397), .B1(n5396), .B2(DATAI_24_), .ZN(
        n5094) );
  AOI22_X1 U6108 ( .A1(n5407), .A2(DATAI_8_), .B1(n5406), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6109 ( .A1(n5094), .A2(n5093), .ZN(U2867) );
  INV_X1 U6110 ( .A(DATAI_23_), .ZN(n5095) );
  OAI22_X1 U6111 ( .A1(n5096), .A2(n5403), .B1(n5402), .B2(n5095), .ZN(n5097)
         );
  INV_X1 U6112 ( .A(n5097), .ZN(n5099) );
  AOI22_X1 U6113 ( .A1(n5407), .A2(DATAI_7_), .B1(n5406), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6114 ( .A1(n5099), .A2(n5098), .ZN(U2868) );
  INV_X1 U6115 ( .A(DATAI_22_), .ZN(n5100) );
  OAI22_X1 U6116 ( .A1(n5101), .A2(n5403), .B1(n5402), .B2(n5100), .ZN(n5102)
         );
  INV_X1 U6117 ( .A(n5102), .ZN(n5104) );
  AOI22_X1 U6118 ( .A1(n5407), .A2(DATAI_6_), .B1(n5406), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6119 ( .A1(n5104), .A2(n5103), .ZN(U2869) );
  INV_X1 U6120 ( .A(DATAI_21_), .ZN(n5105) );
  OAI22_X1 U6121 ( .A1(n5106), .A2(n5403), .B1(n5402), .B2(n5105), .ZN(n5107)
         );
  INV_X1 U6122 ( .A(n5107), .ZN(n5109) );
  AOI22_X1 U6123 ( .A1(n5407), .A2(DATAI_5_), .B1(n5406), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6124 ( .A1(n5109), .A2(n5108), .ZN(U2870) );
  AOI22_X1 U6125 ( .A1(n5110), .A2(n5397), .B1(n5396), .B2(DATAI_20_), .ZN(
        n5112) );
  AOI22_X1 U6126 ( .A1(n5407), .A2(DATAI_4_), .B1(n5406), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6127 ( .A1(n5112), .A2(n5111), .ZN(U2871) );
  AOI22_X1 U6128 ( .A1(n5138), .A2(n5397), .B1(n5396), .B2(DATAI_19_), .ZN(
        n5114) );
  AOI22_X1 U6129 ( .A1(n5407), .A2(DATAI_3_), .B1(n5406), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6130 ( .A1(n5114), .A2(n5113), .ZN(U2872) );
  AOI22_X1 U6131 ( .A1(n5585), .A2(REIP_REG_26__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5118) );
  AOI22_X1 U6132 ( .A1(n5116), .A2(n5533), .B1(n5115), .B2(n5483), .ZN(n5117)
         );
  OAI211_X1 U6133 ( .C1(n6076), .C2(n5119), .A(n5118), .B(n5117), .ZN(U2960)
         );
  AOI22_X1 U6134 ( .A1(n5585), .A2(REIP_REG_25__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5123) );
  OAI21_X1 U6135 ( .B1(n5120), .B2(n4015), .A(n4847), .ZN(n5164) );
  AOI22_X1 U6136 ( .A1(n5121), .A2(n5631), .B1(n5533), .B2(n5164), .ZN(n5122)
         );
  OAI211_X1 U6137 ( .C1(n5525), .C2(n5124), .A(n5123), .B(n5122), .ZN(U2961)
         );
  INV_X1 U6138 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5133) );
  OAI21_X1 U6139 ( .B1(n5127), .B2(n5126), .A(n5125), .ZN(n5128) );
  INV_X1 U6140 ( .A(n5128), .ZN(n5170) );
  OAI22_X1 U6141 ( .A1(n5170), .A2(n5503), .B1(n5525), .B2(n5129), .ZN(n5130)
         );
  AOI21_X1 U6142 ( .B1(n5631), .B2(n5131), .A(n5130), .ZN(n5132) );
  NAND2_X1 U6143 ( .A1(n5585), .A2(REIP_REG_21__SCAN_IN), .ZN(n5173) );
  OAI211_X1 U6144 ( .C1(n5133), .C2(n5530), .A(n5132), .B(n5173), .ZN(U2965)
         );
  INV_X1 U6145 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5140) );
  OAI21_X1 U6146 ( .B1(n5135), .B2(n5134), .A(n4864), .ZN(n5177) );
  OAI22_X1 U6147 ( .A1(n5177), .A2(n5503), .B1(n5136), .B2(n5525), .ZN(n5137)
         );
  AOI21_X1 U6148 ( .B1(n5631), .B2(n5138), .A(n5137), .ZN(n5139) );
  NAND2_X1 U6149 ( .A1(n5585), .A2(REIP_REG_19__SCAN_IN), .ZN(n5180) );
  OAI211_X1 U6150 ( .C1(n5140), .C2(n5530), .A(n5139), .B(n5180), .ZN(U2967)
         );
  AOI22_X1 U6151 ( .A1(n5585), .A2(REIP_REG_18__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6152 ( .A1(n3981), .A2(n3987), .ZN(n5142) );
  OAI21_X1 U6153 ( .B1(n4954), .B2(n5142), .A(n5183), .ZN(n5143) );
  OAI21_X1 U6154 ( .B1(n5183), .B2(n3980), .A(n5143), .ZN(n5152) );
  AOI21_X1 U6155 ( .B1(n5141), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5152), 
        .ZN(n5144) );
  XOR2_X1 U6156 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5144), .Z(n5185) );
  AOI22_X1 U6157 ( .A1(n5533), .A2(n5185), .B1(n5483), .B2(n5227), .ZN(n5145)
         );
  OAI211_X1 U6158 ( .C1(n6076), .C2(n5230), .A(n5146), .B(n5145), .ZN(U2968)
         );
  AOI22_X1 U6159 ( .A1(n5585), .A2(REIP_REG_17__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5154) );
  AOI21_X1 U6160 ( .B1(n4694), .B2(n5147), .A(n4726), .ZN(n5398) );
  INV_X1 U6161 ( .A(n5141), .ZN(n5151) );
  MUX2_X1 U6162 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .B(n5183), .S(n3980), 
        .Z(n5148) );
  OAI21_X1 U6163 ( .B1(n5151), .B2(n5149), .A(n5148), .ZN(n5150) );
  OAI21_X1 U6164 ( .B1(n5152), .B2(n5151), .A(n5150), .ZN(n5193) );
  AOI22_X1 U6165 ( .A1(n5398), .A2(n5631), .B1(n5533), .B2(n5193), .ZN(n5153)
         );
  OAI211_X1 U6166 ( .C1(n5525), .C2(n5238), .A(n5154), .B(n5153), .ZN(U2969)
         );
  AOI22_X1 U6167 ( .A1(n5585), .A2(REIP_REG_16__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5157) );
  AOI22_X1 U6168 ( .A1(n5155), .A2(n5533), .B1(n5483), .B2(n5244), .ZN(n5156)
         );
  OAI211_X1 U6169 ( .C1(n6076), .C2(n5404), .A(n5157), .B(n5156), .ZN(U2970)
         );
  AOI22_X1 U6170 ( .A1(n5585), .A2(REIP_REG_14__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5160) );
  AOI22_X1 U6171 ( .A1(n5158), .A2(n5533), .B1(n5483), .B2(n5262), .ZN(n5159)
         );
  OAI211_X1 U6172 ( .C1(n6076), .C2(n5260), .A(n5160), .B(n5159), .ZN(U2972)
         );
  INV_X1 U6173 ( .A(n5161), .ZN(n5162) );
  AOI22_X1 U6174 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5585), .B1(n5162), .B2(
        n5167), .ZN(n5166) );
  AOI22_X1 U6175 ( .A1(n5164), .A2(n5591), .B1(n5590), .B2(n5163), .ZN(n5165)
         );
  OAI211_X1 U6176 ( .C1(n5168), .C2(n5167), .A(n5166), .B(n5165), .ZN(U2993)
         );
  OAI22_X1 U6177 ( .A1(n5170), .A2(n5541), .B1(n5540), .B2(n5169), .ZN(n5171)
         );
  AOI21_X1 U6178 ( .B1(n5172), .B2(n6455), .A(n5171), .ZN(n5174) );
  OAI211_X1 U6179 ( .C1(n5175), .C2(n6455), .A(n5174), .B(n5173), .ZN(U2997)
         );
  OAI22_X1 U6180 ( .A1(n5177), .A2(n5541), .B1(n5540), .B2(n5176), .ZN(n5178)
         );
  AOI21_X1 U6181 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5179), .A(n5178), 
        .ZN(n5181) );
  OAI211_X1 U6182 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5182), .A(n5181), .B(n5180), .ZN(U2999) );
  INV_X1 U6183 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5188) );
  NOR3_X1 U6184 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5183), .A3(n5196), 
        .ZN(n5184) );
  AOI21_X1 U6185 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5585), .A(n5184), .ZN(n5187) );
  AOI22_X1 U6186 ( .A1(n5185), .A2(n5591), .B1(n5590), .B2(n5226), .ZN(n5186)
         );
  OAI211_X1 U6187 ( .C1(n5189), .C2(n5188), .A(n5187), .B(n5186), .ZN(U3000)
         );
  AOI22_X1 U6188 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5190), .B1(n5585), .B2(REIP_REG_17__SCAN_IN), .ZN(n5195) );
  AOI21_X1 U6189 ( .B1(n5192), .B2(n5191), .A(n4753), .ZN(n5379) );
  AOI22_X1 U6190 ( .A1(n5193), .A2(n5591), .B1(n5590), .B2(n5379), .ZN(n5194)
         );
  OAI211_X1 U6191 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5196), .A(n5195), .B(n5194), .ZN(U3001) );
  OR3_X1 U6192 ( .A1(n5198), .A2(n5197), .A3(n6273), .ZN(n5199) );
  OAI21_X1 U6193 ( .B1(n6269), .B2(n5200), .A(n5199), .ZN(U3455) );
  AOI21_X1 U6194 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6209), .A(n6200), .ZN(n5205) );
  INV_X1 U6195 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5201) );
  NOR2_X2 U6196 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6199), .ZN(n6315) );
  AOI21_X1 U6197 ( .B1(n5205), .B2(n5201), .A(n6315), .ZN(U2789) );
  OAI22_X1 U6198 ( .A1(n3828), .A2(n5202), .B1(n2977), .B2(n6157), .ZN(n5208)
         );
  OAI21_X1 U6199 ( .B1(n5208), .B2(n6178), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5203) );
  OAI21_X1 U6200 ( .B1(n6316), .B2(n6180), .A(n5203), .ZN(U2790) );
  INV_X2 U6201 ( .A(n6315), .ZN(n6259) );
  NOR2_X1 U6202 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5206) );
  OAI21_X1 U6203 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5206), .A(n6259), .ZN(n5204)
         );
  OAI21_X1 U6204 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6259), .A(n5204), .ZN(
        U2791) );
  NOR2_X1 U6205 ( .A1(n6315), .A2(n5205), .ZN(n6263) );
  OAI21_X1 U6206 ( .B1(n5206), .B2(BS16_N), .A(n6263), .ZN(n6262) );
  OAI21_X1 U6207 ( .B1(n6263), .B2(n6026), .A(n6262), .ZN(U2792) );
  NOR2_X1 U6208 ( .A1(n5207), .A2(n2977), .ZN(n6320) );
  AOI21_X1 U6209 ( .B1(n6320), .B2(n6198), .A(READY_N), .ZN(n6308) );
  NOR2_X1 U6210 ( .A1(n5208), .A2(n6308), .ZN(n6159) );
  NOR2_X1 U6211 ( .A1(n6159), .A2(n6178), .ZN(n6305) );
  OAI21_X1 U6212 ( .B1(n6305), .B2(n5209), .A(n5503), .ZN(U2793) );
  INV_X1 U6213 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6363) );
  INV_X1 U6214 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U6215 ( .A1(n6363), .A2(n6353), .ZN(n6465) );
  OR4_X1 U6216 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5210) );
  AOI211_X1 U6217 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6465), .B(n5210), .ZN(n5218) );
  NOR4_X1 U6218 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5217) );
  NOR4_X1 U6219 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5216) );
  NOR4_X1 U6220 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5214) );
  NOR4_X1 U6221 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5213) );
  NOR4_X1 U6222 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5212) );
  NOR4_X1 U6223 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5211) );
  AND4_X1 U6224 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n5215)
         );
  NAND4_X1 U6225 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n6300)
         );
  NOR2_X1 U6226 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6300), .ZN(n6301) );
  INV_X1 U6227 ( .A(n6300), .ZN(n5219) );
  NOR2_X1 U6228 ( .A1(n5219), .A2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5220) );
  INV_X1 U6229 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6335) );
  INV_X1 U6230 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6383) );
  INV_X1 U6231 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6295) );
  NAND4_X1 U6232 ( .A1(n5219), .A2(n6335), .A3(n6383), .A4(n6295), .ZN(n5221)
         );
  OAI21_X1 U6233 ( .B1(n6301), .B2(n5220), .A(n5221), .ZN(U2794) );
  AOI22_X1 U6234 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6300), .B1(n6301), 
        .B2(n6383), .ZN(n5222) );
  NAND2_X1 U6235 ( .A1(n5222), .A2(n5221), .ZN(U2795) );
  INV_X1 U6236 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6235) );
  AOI21_X1 U6237 ( .B1(n5375), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5354), 
        .ZN(n5223) );
  OAI221_X1 U6238 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5224), .C1(n6235), .C2(
        n5233), .A(n5223), .ZN(n5225) );
  AOI21_X1 U6239 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5353), .A(n5225), .ZN(n5229)
         );
  AOI22_X1 U6240 ( .A1(n5227), .A2(n5374), .B1(n5369), .B2(n5226), .ZN(n5228)
         );
  OAI211_X1 U6241 ( .C1(n5336), .C2(n5230), .A(n5229), .B(n5228), .ZN(U2809)
         );
  NOR2_X1 U6242 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5231), .ZN(n5234) );
  INV_X1 U6243 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5232) );
  OAI22_X1 U6244 ( .A1(n5234), .A2(n5233), .B1(n5232), .B2(n5343), .ZN(n5235)
         );
  AOI211_X1 U6245 ( .C1(n5353), .C2(EBX_REG_17__SCAN_IN), .A(n5354), .B(n5235), 
        .ZN(n5237) );
  AOI22_X1 U6246 ( .A1(n5369), .A2(n5379), .B1(n5328), .B2(n5398), .ZN(n5236)
         );
  OAI211_X1 U6247 ( .C1(n5238), .C2(n5359), .A(n5237), .B(n5236), .ZN(U2810)
         );
  AOI22_X1 U6248 ( .A1(n5251), .A2(n6397), .B1(n5368), .B2(n5248), .ZN(n5240)
         );
  AOI21_X1 U6249 ( .B1(n5375), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5354), 
        .ZN(n5239) );
  OAI221_X1 U6250 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5241), .C1(n6230), .C2(
        n5240), .A(n5239), .ZN(n5242) );
  AOI21_X1 U6251 ( .B1(EBX_REG_16__SCAN_IN), .B2(n5353), .A(n5242), .ZN(n5246)
         );
  INV_X1 U6252 ( .A(n5404), .ZN(n5243) );
  AOI22_X1 U6253 ( .A1(n5244), .A2(n5374), .B1(n5328), .B2(n5243), .ZN(n5245)
         );
  OAI211_X1 U6254 ( .C1(n5367), .C2(n5247), .A(n5246), .B(n5245), .ZN(U2811)
         );
  NAND2_X1 U6255 ( .A1(n5368), .A2(n5248), .ZN(n5265) );
  OAI22_X1 U6256 ( .A1(n6378), .A2(n5370), .B1(n6397), .B2(n5265), .ZN(n5249)
         );
  AOI211_X1 U6257 ( .C1(n5375), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5354), 
        .B(n5249), .ZN(n5255) );
  AOI22_X1 U6258 ( .A1(n5250), .A2(n5374), .B1(n5328), .B2(n5383), .ZN(n5254)
         );
  NAND2_X1 U6259 ( .A1(n5251), .A2(n6397), .ZN(n5253) );
  NAND2_X1 U6260 ( .A1(n5369), .A2(n5382), .ZN(n5252) );
  NAND4_X1 U6261 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(U2812)
         );
  AND2_X1 U6262 ( .A1(n5346), .A2(n5256), .ZN(n5268) );
  AOI21_X1 U6263 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5268), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5266) );
  OAI22_X1 U6264 ( .A1(n5258), .A2(n5343), .B1(n5367), .B2(n5257), .ZN(n5259)
         );
  AOI211_X1 U6265 ( .C1(n5353), .C2(EBX_REG_14__SCAN_IN), .A(n5354), .B(n5259), 
        .ZN(n5264) );
  INV_X1 U6266 ( .A(n5260), .ZN(n5261) );
  AOI22_X1 U6267 ( .A1(n5262), .A2(n5374), .B1(n5328), .B2(n5261), .ZN(n5263)
         );
  OAI211_X1 U6268 ( .C1(n5266), .C2(n5265), .A(n5264), .B(n5263), .ZN(U2813)
         );
  OR3_X1 U6269 ( .A1(n5295), .A2(n5276), .A3(n5277), .ZN(n5267) );
  NAND2_X1 U6270 ( .A1(n5267), .A2(n5368), .ZN(n5274) );
  AOI22_X1 U6271 ( .A1(n5369), .A2(n5385), .B1(n5268), .B2(n6228), .ZN(n5269)
         );
  OAI21_X1 U6272 ( .B1(n5388), .B2(n5370), .A(n5269), .ZN(n5270) );
  AOI211_X1 U6273 ( .C1(n5375), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5354), 
        .B(n5270), .ZN(n5273) );
  AOI22_X1 U6274 ( .A1(n5271), .A2(n5374), .B1(n5328), .B2(n5386), .ZN(n5272)
         );
  OAI211_X1 U6275 ( .C1(n5274), .C2(n6228), .A(n5273), .B(n5272), .ZN(U2814)
         );
  NOR3_X1 U6276 ( .A1(n5275), .A2(n5276), .A3(REIP_REG_12__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6277 ( .A1(n5346), .A2(n5276), .ZN(n5286) );
  NOR2_X1 U6278 ( .A1(n5295), .A2(n5286), .ZN(n5288) );
  NOR2_X1 U6279 ( .A1(n5288), .A2(n5277), .ZN(n5278) );
  AOI211_X1 U6280 ( .C1(n5353), .C2(EBX_REG_12__SCAN_IN), .A(n5279), .B(n5278), 
        .ZN(n5283) );
  OAI22_X1 U6281 ( .A1(n6392), .A2(n5343), .B1(n5367), .B2(n5280), .ZN(n5281)
         );
  AOI211_X1 U6282 ( .C1(n5374), .C2(n5464), .A(n5354), .B(n5281), .ZN(n5282)
         );
  OAI211_X1 U6283 ( .C1(n5336), .C2(n5468), .A(n5283), .B(n5282), .ZN(U2815)
         );
  AOI21_X1 U6284 ( .B1(n5285), .B2(n5284), .A(n4619), .ZN(n5538) );
  AOI22_X1 U6285 ( .A1(n5369), .A2(n5538), .B1(n5287), .B2(n5286), .ZN(n5292)
         );
  INV_X1 U6286 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6225) );
  OAI22_X1 U6287 ( .A1(n5288), .A2(n6225), .B1(n3479), .B2(n5343), .ZN(n5289)
         );
  AOI211_X1 U6288 ( .C1(n5353), .C2(EBX_REG_11__SCAN_IN), .A(n5354), .B(n5289), 
        .ZN(n5291) );
  AOI22_X1 U6289 ( .A1(n5474), .A2(n5374), .B1(n5328), .B2(n5473), .ZN(n5290)
         );
  NAND3_X1 U6290 ( .A1(n5292), .A2(n5291), .A3(n5290), .ZN(U2816) );
  OAI22_X1 U6291 ( .A1(n4083), .A2(n5370), .B1(n5367), .B2(n5549), .ZN(n5293)
         );
  AOI211_X1 U6292 ( .C1(n5375), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5354), 
        .B(n5293), .ZN(n5305) );
  INV_X1 U6293 ( .A(n5486), .ZN(n5294) );
  AOI22_X1 U6294 ( .A1(n5482), .A2(n5374), .B1(n5328), .B2(n5294), .ZN(n5304)
         );
  INV_X1 U6295 ( .A(n5299), .ZN(n5296) );
  NOR2_X1 U6296 ( .A1(n5295), .A2(n5297), .ZN(n5329) );
  AOI21_X1 U6297 ( .B1(n5296), .B2(n5329), .A(n5330), .ZN(n5313) );
  INV_X1 U6298 ( .A(n5297), .ZN(n5298) );
  NAND2_X1 U6299 ( .A1(n5346), .A2(n5298), .ZN(n5331) );
  NOR2_X1 U6300 ( .A1(n5331), .A2(n5299), .ZN(n5301) );
  INV_X1 U6301 ( .A(n5301), .ZN(n5300) );
  NOR2_X1 U6302 ( .A1(n5300), .A2(REIP_REG_9__SCAN_IN), .ZN(n5306) );
  OAI21_X1 U6303 ( .B1(n5313), .B2(n5306), .A(REIP_REG_10__SCAN_IN), .ZN(n5303) );
  NAND3_X1 U6304 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5301), .A3(n6452), .ZN(n5302) );
  NAND4_X1 U6305 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(U2817)
         );
  AOI21_X1 U6306 ( .B1(n5313), .B2(REIP_REG_9__SCAN_IN), .A(n5306), .ZN(n5312)
         );
  AOI22_X1 U6307 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n5375), .B1(n5369), 
        .B2(n5559), .ZN(n5311) );
  AOI21_X1 U6308 ( .B1(n5353), .B2(EBX_REG_9__SCAN_IN), .A(n5354), .ZN(n5310)
         );
  AOI22_X1 U6309 ( .A1(n5308), .A2(n5374), .B1(n5328), .B2(n5307), .ZN(n5309)
         );
  NAND4_X1 U6310 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(U2818)
         );
  NOR2_X1 U6311 ( .A1(n5331), .A2(n6217), .ZN(n5323) );
  AOI21_X1 U6312 ( .B1(REIP_REG_7__SCAN_IN), .B2(n5323), .A(
        REIP_REG_8__SCAN_IN), .ZN(n5322) );
  INV_X1 U6313 ( .A(n5313), .ZN(n5321) );
  OAI22_X1 U6314 ( .A1(n5315), .A2(n5370), .B1(n5367), .B2(n5314), .ZN(n5316)
         );
  AOI211_X1 U6315 ( .C1(n5375), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5354), 
        .B(n5316), .ZN(n5320) );
  AOI22_X1 U6316 ( .A1(n5318), .A2(n5374), .B1(n5328), .B2(n5317), .ZN(n5319)
         );
  OAI211_X1 U6317 ( .C1(n5322), .C2(n5321), .A(n5320), .B(n5319), .ZN(U2819)
         );
  AOI21_X1 U6318 ( .B1(n5375), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5354), 
        .ZN(n5325) );
  INV_X1 U6319 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6220) );
  AOI22_X1 U6320 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5353), .B1(n5323), .B2(n6220), 
        .ZN(n5324) );
  OAI211_X1 U6321 ( .C1(n5367), .C2(n5326), .A(n5325), .B(n5324), .ZN(n5327)
         );
  AOI21_X1 U6322 ( .B1(n5328), .B2(n5490), .A(n5327), .ZN(n5333) );
  NOR2_X1 U6323 ( .A1(n5330), .A2(n5329), .ZN(n5348) );
  NOR2_X1 U6324 ( .A1(n5331), .A2(REIP_REG_6__SCAN_IN), .ZN(n5338) );
  OAI21_X1 U6325 ( .B1(n5348), .B2(n5338), .A(REIP_REG_7__SCAN_IN), .ZN(n5332)
         );
  OAI211_X1 U6326 ( .C1(n5359), .C2(n5487), .A(n5333), .B(n5332), .ZN(U2820)
         );
  AOI22_X1 U6327 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5375), .B1(
        REIP_REG_6__SCAN_IN), .B2(n5348), .ZN(n5335) );
  AOI21_X1 U6328 ( .B1(n5353), .B2(EBX_REG_6__SCAN_IN), .A(n5354), .ZN(n5334)
         );
  OAI211_X1 U6329 ( .C1(n5336), .C2(n5500), .A(n5335), .B(n5334), .ZN(n5337)
         );
  AOI211_X1 U6330 ( .C1(n5339), .C2(n5369), .A(n5338), .B(n5337), .ZN(n5340)
         );
  OAI21_X1 U6331 ( .B1(n5495), .B2(n5359), .A(n5340), .ZN(U2821) );
  INV_X1 U6332 ( .A(n5341), .ZN(n5502) );
  OAI22_X1 U6333 ( .A1(n5509), .A2(n5343), .B1(n5367), .B2(n5342), .ZN(n5344)
         );
  AOI211_X1 U6334 ( .C1(n5353), .C2(EBX_REG_5__SCAN_IN), .A(n5354), .B(n5344), 
        .ZN(n5350) );
  NAND2_X1 U6335 ( .A1(n5346), .A2(n5345), .ZN(n5357) );
  INV_X1 U6336 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6215) );
  OAI21_X1 U6337 ( .B1(n6451), .B2(n5357), .A(n6215), .ZN(n5347) );
  AOI22_X1 U6338 ( .A1(n5348), .A2(n5347), .B1(n5506), .B2(n5358), .ZN(n5349)
         );
  OAI211_X1 U6339 ( .C1(n5502), .C2(n5359), .A(n5350), .B(n5349), .ZN(U2822)
         );
  AOI22_X1 U6340 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5353), .B1(n5352), .B2(n5351), 
        .ZN(n5365) );
  INV_X1 U6341 ( .A(n5354), .ZN(n5355) );
  OAI221_X1 U6342 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5357), .C1(n6451), .C2(
        n5356), .A(n5355), .ZN(n5363) );
  INV_X1 U6343 ( .A(n5358), .ZN(n5378) );
  OAI22_X1 U6344 ( .A1(n5378), .A2(n5361), .B1(n5360), .B2(n5359), .ZN(n5362)
         );
  AOI211_X1 U6345 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n5375), .A(n5363), 
        .B(n5362), .ZN(n5364) );
  OAI211_X1 U6346 ( .C1(n5367), .C2(n5366), .A(n5365), .B(n5364), .ZN(U2823)
         );
  AOI22_X1 U6347 ( .A1(n5369), .A2(n5589), .B1(REIP_REG_0__SCAN_IN), .B2(n5368), .ZN(n5377) );
  OAI22_X1 U6348 ( .A1(n5921), .A2(n5372), .B1(n5371), .B2(n5370), .ZN(n5373)
         );
  AOI221_X1 U6349 ( .B1(n5375), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n5374), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n5373), .ZN(n5376) );
  OAI211_X1 U6350 ( .C1(n5378), .C2(n5536), .A(n5377), .B(n5376), .ZN(U2827)
         );
  AOI22_X1 U6351 ( .A1(n5398), .A2(n5393), .B1(n5392), .B2(n5379), .ZN(n5380)
         );
  OAI21_X1 U6352 ( .B1(n5381), .B2(n4833), .A(n5380), .ZN(U2842) );
  AOI22_X1 U6353 ( .A1(n5383), .A2(n5393), .B1(n5392), .B2(n5382), .ZN(n5384)
         );
  OAI21_X1 U6354 ( .B1(n6378), .B2(n4833), .A(n5384), .ZN(U2844) );
  AOI22_X1 U6355 ( .A1(n5386), .A2(n5393), .B1(n5392), .B2(n5385), .ZN(n5387)
         );
  OAI21_X1 U6356 ( .B1(n5388), .B2(n4833), .A(n5387), .ZN(U2846) );
  AOI22_X1 U6357 ( .A1(n5473), .A2(n5393), .B1(n5392), .B2(n5538), .ZN(n5389)
         );
  OAI21_X1 U6358 ( .B1(n5390), .B2(n4833), .A(n5389), .ZN(U2848) );
  INV_X1 U6359 ( .A(n5391), .ZN(n5567) );
  AOI22_X1 U6360 ( .A1(n5513), .A2(n5393), .B1(n5392), .B2(n5567), .ZN(n5394)
         );
  OAI21_X1 U6361 ( .B1(n5395), .B2(n4833), .A(n5394), .ZN(U2857) );
  AOI22_X1 U6362 ( .A1(n5398), .A2(n5397), .B1(n5396), .B2(DATAI_17_), .ZN(
        n5400) );
  AOI22_X1 U6363 ( .A1(n5407), .A2(DATAI_1_), .B1(n5406), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6364 ( .A1(n5400), .A2(n5399), .ZN(U2874) );
  INV_X1 U6365 ( .A(DATAI_16_), .ZN(n5401) );
  OAI22_X1 U6366 ( .A1(n5404), .A2(n5403), .B1(n5402), .B2(n5401), .ZN(n5405)
         );
  INV_X1 U6367 ( .A(n5405), .ZN(n5409) );
  AOI22_X1 U6368 ( .A1(n5407), .A2(DATAI_0_), .B1(n5406), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6369 ( .A1(n5409), .A2(n5408), .ZN(U2875) );
  INV_X1 U6370 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6420) );
  INV_X1 U6371 ( .A(n5410), .ZN(n5411) );
  AOI22_X1 U6372 ( .A1(n5411), .A2(EAX_REG_28__SCAN_IN), .B1(n6170), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5412) );
  OAI21_X1 U6373 ( .B1(n6420), .B2(n5436), .A(n5412), .ZN(U2895) );
  INV_X1 U6374 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5463) );
  AOI22_X1 U6375 ( .A1(n6170), .A2(LWORD_REG_15__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5413) );
  OAI21_X1 U6376 ( .B1(n5463), .B2(n5439), .A(n5413), .ZN(U2908) );
  INV_X1 U6377 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6366) );
  AOI22_X1 U6378 ( .A1(EAX_REG_14__SCAN_IN), .A2(n5426), .B1(n6307), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5414) );
  OAI21_X1 U6379 ( .B1(n6366), .B2(n5436), .A(n5414), .ZN(U2909) );
  INV_X1 U6380 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5416) );
  AOI22_X1 U6381 ( .A1(n6170), .A2(LWORD_REG_13__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U6382 ( .B1(n5416), .B2(n5439), .A(n5415), .ZN(U2910) );
  INV_X1 U6383 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n6384) );
  AOI22_X1 U6384 ( .A1(EAX_REG_12__SCAN_IN), .A2(n5426), .B1(n6307), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5417) );
  OAI21_X1 U6385 ( .B1(n6384), .B2(n5436), .A(n5417), .ZN(U2911) );
  INV_X1 U6386 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5419) );
  AOI22_X1 U6387 ( .A1(n6170), .A2(LWORD_REG_11__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5418) );
  OAI21_X1 U6388 ( .B1(n5419), .B2(n5439), .A(n5418), .ZN(U2912) );
  INV_X1 U6389 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5421) );
  AOI22_X1 U6390 ( .A1(n6170), .A2(LWORD_REG_10__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U6391 ( .B1(n5421), .B2(n5439), .A(n5420), .ZN(U2913) );
  INV_X1 U6392 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5423) );
  AOI22_X1 U6393 ( .A1(n6170), .A2(LWORD_REG_9__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5422) );
  OAI21_X1 U6394 ( .B1(n5423), .B2(n5439), .A(n5422), .ZN(U2914) );
  INV_X1 U6395 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5425) );
  AOI22_X1 U6396 ( .A1(n6170), .A2(LWORD_REG_8__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5424) );
  OAI21_X1 U6397 ( .B1(n5425), .B2(n5439), .A(n5424), .ZN(U2915) );
  AOI22_X1 U6398 ( .A1(EAX_REG_7__SCAN_IN), .A2(n5426), .B1(n5437), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5427) );
  OAI21_X1 U6399 ( .B1(n5435), .B2(n4395), .A(n5427), .ZN(U2916) );
  AOI22_X1 U6400 ( .A1(n6170), .A2(LWORD_REG_6__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5428) );
  OAI21_X1 U6401 ( .B1(n4525), .B2(n5439), .A(n5428), .ZN(U2917) );
  AOI22_X1 U6402 ( .A1(n6170), .A2(LWORD_REG_5__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5429) );
  OAI21_X1 U6403 ( .B1(n4535), .B2(n5439), .A(n5429), .ZN(U2918) );
  INV_X1 U6404 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n5430) );
  INV_X1 U6405 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6400) );
  OAI222_X1 U6406 ( .A1(n5435), .A2(n5430), .B1(n5439), .B2(n6441), .C1(n6400), 
        .C2(n5436), .ZN(U2919) );
  AOI22_X1 U6407 ( .A1(n6170), .A2(LWORD_REG_3__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5431) );
  OAI21_X1 U6408 ( .B1(n5432), .B2(n5439), .A(n5431), .ZN(U2920) );
  AOI22_X1 U6409 ( .A1(n6170), .A2(LWORD_REG_2__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5433) );
  OAI21_X1 U6410 ( .B1(n5434), .B2(n5439), .A(n5433), .ZN(U2921) );
  INV_X1 U6411 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6350) );
  OAI222_X1 U6412 ( .A1(n5436), .A2(n6350), .B1(n5439), .B2(n6460), .C1(n5435), 
        .C2(n4397), .ZN(U2922) );
  AOI22_X1 U6413 ( .A1(n6170), .A2(LWORD_REG_0__SCAN_IN), .B1(n5437), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5438) );
  OAI21_X1 U6414 ( .B1(n5440), .B2(n5439), .A(n5438), .ZN(U2923) );
  AOI22_X1 U6415 ( .A1(EAX_REG_25__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6416 ( .A1(n6437), .A2(DATAI_9_), .ZN(n5448) );
  NAND2_X1 U6417 ( .A1(n5441), .A2(n5448), .ZN(U2933) );
  AOI22_X1 U6418 ( .A1(EAX_REG_26__SCAN_IN), .A2(n5459), .B1(n6438), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6419 ( .A1(n6437), .A2(DATAI_10_), .ZN(n5450) );
  NAND2_X1 U6420 ( .A1(n5442), .A2(n5450), .ZN(U2934) );
  AOI22_X1 U6421 ( .A1(EAX_REG_27__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6422 ( .A1(n6437), .A2(DATAI_11_), .ZN(n5452) );
  NAND2_X1 U6423 ( .A1(n5443), .A2(n5452), .ZN(U2935) );
  AOI22_X1 U6424 ( .A1(EAX_REG_28__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6425 ( .A1(n6437), .A2(DATAI_12_), .ZN(n5454) );
  NAND2_X1 U6426 ( .A1(n5444), .A2(n5454), .ZN(U2936) );
  AOI22_X1 U6427 ( .A1(EAX_REG_29__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6428 ( .A1(n6437), .A2(DATAI_13_), .ZN(n5456) );
  NAND2_X1 U6429 ( .A1(n5445), .A2(n5456), .ZN(U2937) );
  NAND2_X1 U6430 ( .A1(n6437), .A2(DATAI_14_), .ZN(n5460) );
  INV_X1 U6431 ( .A(n5460), .ZN(n5446) );
  AOI21_X1 U6432 ( .B1(n6438), .B2(UWORD_REG_14__SCAN_IN), .A(n5446), .ZN(
        n5447) );
  OAI21_X1 U6433 ( .B1(n3820), .B2(n6440), .A(n5447), .ZN(U2938) );
  AOI22_X1 U6434 ( .A1(EAX_REG_9__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6435 ( .A1(n5449), .A2(n5448), .ZN(U2948) );
  AOI22_X1 U6436 ( .A1(EAX_REG_10__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6437 ( .A1(n5451), .A2(n5450), .ZN(U2949) );
  AOI22_X1 U6438 ( .A1(EAX_REG_11__SCAN_IN), .A2(n5459), .B1(n6438), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6439 ( .A1(n5453), .A2(n5452), .ZN(U2950) );
  AOI22_X1 U6440 ( .A1(EAX_REG_12__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6441 ( .A1(n5455), .A2(n5454), .ZN(U2951) );
  AOI22_X1 U6442 ( .A1(EAX_REG_13__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6443 ( .A1(n5457), .A2(n5456), .ZN(U2952) );
  AOI22_X1 U6444 ( .A1(EAX_REG_14__SCAN_IN), .A2(n5459), .B1(n5458), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6445 ( .A1(n5461), .A2(n5460), .ZN(U2953) );
  AOI22_X1 U6446 ( .A1(n6438), .A2(LWORD_REG_15__SCAN_IN), .B1(n6437), .B2(
        DATAI_15_), .ZN(n5462) );
  OAI21_X1 U6447 ( .B1(n5463), .B2(n6440), .A(n5462), .ZN(U2954) );
  AOI22_X1 U6448 ( .A1(n5585), .A2(REIP_REG_12__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5467) );
  AOI22_X1 U6449 ( .A1(n5465), .A2(n5533), .B1(n5483), .B2(n5464), .ZN(n5466)
         );
  OAI211_X1 U6450 ( .C1(n6076), .C2(n5468), .A(n5467), .B(n5466), .ZN(U2974)
         );
  AND2_X1 U6451 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  XNOR2_X1 U6452 ( .A(n2952), .B(n5472), .ZN(n5542) );
  AOI22_X1 U6453 ( .A1(n5585), .A2(REIP_REG_11__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5476) );
  AOI22_X1 U6454 ( .A1(n5483), .A2(n5474), .B1(n5631), .B2(n5473), .ZN(n5475)
         );
  OAI211_X1 U6455 ( .C1(n5542), .C2(n5503), .A(n5476), .B(n5475), .ZN(U2975)
         );
  AOI22_X1 U6456 ( .A1(n5585), .A2(REIP_REG_10__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5485) );
  INV_X1 U6457 ( .A(n5478), .ZN(n5480) );
  NOR2_X1 U6458 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  XNOR2_X1 U6459 ( .A(n5477), .B(n5481), .ZN(n5550) );
  AOI22_X1 U6460 ( .A1(n5550), .A2(n5533), .B1(n5483), .B2(n5482), .ZN(n5484)
         );
  OAI211_X1 U6461 ( .C1(n6076), .C2(n5486), .A(n5485), .B(n5484), .ZN(U2976)
         );
  OAI22_X1 U6462 ( .A1(n5488), .A2(n5503), .B1(n5487), .B2(n5525), .ZN(n5489)
         );
  AOI21_X1 U6463 ( .B1(n5631), .B2(n5490), .A(n5489), .ZN(n5492) );
  OAI211_X1 U6464 ( .C1(n5493), .C2(n5530), .A(n5492), .B(n5491), .ZN(U2979)
         );
  INV_X1 U6465 ( .A(n5494), .ZN(n5496) );
  OAI22_X1 U6466 ( .A1(n5496), .A2(n5503), .B1(n5495), .B2(n5525), .ZN(n5497)
         );
  AOI211_X1 U6467 ( .C1(PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n5517), .A(n5498), 
        .B(n5497), .ZN(n5499) );
  OAI21_X1 U6468 ( .B1(n6076), .B2(n5500), .A(n5499), .ZN(U2980) );
  INV_X1 U6469 ( .A(n5501), .ZN(n5504) );
  OAI22_X1 U6470 ( .A1(n5504), .A2(n5503), .B1(n5502), .B2(n5525), .ZN(n5505)
         );
  AOI21_X1 U6471 ( .B1(n5631), .B2(n5506), .A(n5505), .ZN(n5508) );
  OAI211_X1 U6472 ( .C1(n5509), .C2(n5530), .A(n5508), .B(n5507), .ZN(U2981)
         );
  AOI22_X1 U6473 ( .A1(n5585), .A2(REIP_REG_2__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5515) );
  XNOR2_X1 U6474 ( .A(n5511), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5512)
         );
  XNOR2_X1 U6475 ( .A(n5510), .B(n5512), .ZN(n5571) );
  AOI22_X1 U6476 ( .A1(n5533), .A2(n5571), .B1(n5631), .B2(n5513), .ZN(n5514)
         );
  OAI211_X1 U6477 ( .C1(n5525), .C2(n5516), .A(n5515), .B(n5514), .ZN(U2984)
         );
  AOI22_X1 U6478 ( .A1(n5585), .A2(REIP_REG_1__SCAN_IN), .B1(n5517), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5524) );
  OAI21_X1 U6479 ( .B1(n5520), .B2(n5519), .A(n5518), .ZN(n5521) );
  INV_X1 U6480 ( .A(n5521), .ZN(n5583) );
  AOI22_X1 U6481 ( .A1(n5533), .A2(n5583), .B1(n5631), .B2(n5522), .ZN(n5523)
         );
  OAI211_X1 U6482 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5525), .A(n5524), 
        .B(n5523), .ZN(U2985) );
  INV_X1 U6483 ( .A(n5526), .ZN(n5529) );
  INV_X1 U6484 ( .A(n5527), .ZN(n5528) );
  AOI21_X1 U6485 ( .B1(n5529), .B2(n6461), .A(n5528), .ZN(n5592) );
  NAND2_X1 U6486 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  AOI22_X1 U6487 ( .A1(n5533), .A2(n5592), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5532), .ZN(n5535) );
  NAND2_X1 U6488 ( .A1(n5585), .A2(REIP_REG_0__SCAN_IN), .ZN(n5534) );
  OAI211_X1 U6489 ( .C1(n5536), .C2(n6076), .A(n5535), .B(n5534), .ZN(U2986)
         );
  INV_X1 U6490 ( .A(n5537), .ZN(n5545) );
  INV_X1 U6491 ( .A(n5538), .ZN(n5539) );
  OAI22_X1 U6492 ( .A1(n5540), .A2(n5539), .B1(n6225), .B2(n5599), .ZN(n5544)
         );
  NOR2_X1 U6493 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  AOI211_X1 U6494 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n5545), .A(n5544), .B(n5543), .ZN(n5547) );
  NAND2_X1 U6495 ( .A1(n5547), .A2(n5546), .ZN(U3007) );
  AOI21_X1 U6496 ( .B1(n5553), .B2(n5580), .A(n5548), .ZN(n5566) );
  INV_X1 U6497 ( .A(n5549), .ZN(n5551) );
  AOI222_X1 U6498 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5585), .B1(n5590), .B2(
        n5551), .C1(n5591), .C2(n5550), .ZN(n5556) );
  NOR2_X1 U6499 ( .A1(n5553), .A2(n5552), .ZN(n5562) );
  OAI211_X1 U6500 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5562), .B(n5554), .ZN(n5555) );
  OAI211_X1 U6501 ( .C1(n5566), .C2(n6398), .A(n5556), .B(n5555), .ZN(U3008)
         );
  INV_X1 U6502 ( .A(n5557), .ZN(n5558) );
  AOI21_X1 U6503 ( .B1(n5590), .B2(n5559), .A(n5558), .ZN(n5564) );
  INV_X1 U6504 ( .A(n5560), .ZN(n5561) );
  AOI22_X1 U6505 ( .A1(n5562), .A2(n5565), .B1(n5591), .B2(n5561), .ZN(n5563)
         );
  OAI211_X1 U6506 ( .C1(n5566), .C2(n5565), .A(n5564), .B(n5563), .ZN(U3009)
         );
  AOI22_X1 U6507 ( .A1(n5567), .A2(n5590), .B1(n5585), .B2(REIP_REG_2__SCAN_IN), .ZN(n5578) );
  OAI33_X1 U6509 ( .A1(1'b0), .A2(n5569), .A3(n4059), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n5587), .B3(n5568), .ZN(n5573) );
  AND2_X1 U6510 ( .A1(n5571), .A2(n5591), .ZN(n5572) );
  NOR2_X1 U6511 ( .A1(n5573), .A2(n5572), .ZN(n5577) );
  NAND3_X1 U6512 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5582), .A3(n5574), 
        .ZN(n5575) );
  NAND4_X1 U6513 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(U3016)
         );
  NAND2_X1 U6514 ( .A1(n5580), .A2(n5579), .ZN(n5588) );
  AOI21_X1 U6515 ( .B1(n5582), .B2(n6461), .A(n5581), .ZN(n5594) );
  AOI222_X1 U6516 ( .A1(REIP_REG_1__SCAN_IN), .A2(n5585), .B1(n5590), .B2(
        n5584), .C1(n5591), .C2(n5583), .ZN(n5586) );
  OAI221_X1 U6517 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n5588), .C1(n5587), .C2(n5594), .A(n5586), .ZN(U3017) );
  AOI22_X1 U6518 ( .A1(n5592), .A2(n5591), .B1(n5590), .B2(n5589), .ZN(n5598)
         );
  AOI22_X1 U6519 ( .A1(n5595), .A2(n5594), .B1(n6461), .B2(n5593), .ZN(n5596)
         );
  INV_X1 U6520 ( .A(n5596), .ZN(n5597) );
  OAI211_X1 U6521 ( .C1(n6335), .C2(n5599), .A(n5598), .B(n5597), .ZN(U3018)
         );
  NOR2_X1 U6522 ( .A1(n6445), .A2(n6291), .ZN(U3019) );
  INV_X1 U6523 ( .A(n6035), .ZN(n6086) );
  AND2_X1 U6524 ( .A1(n5706), .A2(n5926), .ZN(n5600) );
  NAND2_X1 U6525 ( .A1(n4452), .A2(n5600), .ZN(n6021) );
  NAND3_X1 U6526 ( .A1(n6284), .A2(n6145), .A3(n6140), .ZN(n5646) );
  NOR2_X1 U6527 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5646), .ZN(n5636)
         );
  NAND2_X1 U6528 ( .A1(n5602), .A2(n4419), .ZN(n5827) );
  OR2_X1 U6529 ( .A1(n5827), .A2(n6029), .ZN(n5641) );
  NOR2_X1 U6530 ( .A1(n5767), .A2(n5766), .ZN(n5968) );
  INV_X1 U6531 ( .A(n5968), .ZN(n5830) );
  NOR2_X1 U6532 ( .A1(n6022), .A2(n5828), .ZN(n5604) );
  INV_X1 U6533 ( .A(n5604), .ZN(n5708) );
  OAI22_X1 U6534 ( .A1(n5641), .A2(n6275), .B1(n5830), .B2(n5708), .ZN(n5635)
         );
  AOI22_X1 U6535 ( .A1(n6075), .A2(n5636), .B1(n6074), .B2(n5635), .ZN(n5612)
         );
  INV_X1 U6536 ( .A(n5636), .ZN(n5605) );
  INV_X1 U6537 ( .A(n5767), .ZN(n5603) );
  NOR2_X1 U6538 ( .A1(n5603), .A2(n5766), .ZN(n6023) );
  OAI21_X1 U6539 ( .B1(n5604), .B2(n5766), .A(n5831), .ZN(n5712) );
  AOI211_X1 U6540 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5605), .A(n6023), .B(
        n5712), .ZN(n5610) );
  AND2_X1 U6541 ( .A1(n3933), .A2(n5606), .ZN(n5607) );
  NAND2_X1 U6542 ( .A1(n5643), .A2(n3920), .ZN(n5669) );
  OAI21_X1 U6543 ( .B1(n5657), .B2(n6127), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5608) );
  NAND3_X1 U6544 ( .A1(n5608), .A2(n6289), .A3(n5641), .ZN(n5609) );
  NAND2_X1 U6545 ( .A1(n5610), .A2(n5609), .ZN(n5637) );
  AOI22_X1 U6546 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5637), .B1(n6083), 
        .B2(n5657), .ZN(n5611) );
  OAI211_X1 U6547 ( .C1(n6086), .C2(n5640), .A(n5612), .B(n5611), .ZN(U3020)
         );
  INV_X1 U6548 ( .A(n6039), .ZN(n6092) );
  AOI22_X1 U6549 ( .A1(n6088), .A2(n5636), .B1(n6087), .B2(n5635), .ZN(n5615)
         );
  AOI22_X1 U6550 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5637), .B1(n6089), 
        .B2(n5657), .ZN(n5614) );
  OAI211_X1 U6551 ( .C1(n6092), .C2(n5640), .A(n5615), .B(n5614), .ZN(U3021)
         );
  INV_X1 U6552 ( .A(n6043), .ZN(n6098) );
  AOI22_X1 U6553 ( .A1(n6094), .A2(n5636), .B1(n6093), .B2(n5635), .ZN(n5618)
         );
  AOI22_X1 U6554 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5637), .B1(n6095), 
        .B2(n5657), .ZN(n5617) );
  OAI211_X1 U6555 ( .C1(n6098), .C2(n5640), .A(n5618), .B(n5617), .ZN(U3022)
         );
  AND2_X1 U6556 ( .A1(n5631), .A2(DATAI_27_), .ZN(n6047) );
  INV_X1 U6557 ( .A(n6047), .ZN(n6104) );
  NOR2_X2 U6558 ( .A1(n5629), .A2(n5619), .ZN(n6100) );
  NOR2_X2 U6559 ( .A1(n5620), .A2(n5630), .ZN(n6099) );
  AOI22_X1 U6560 ( .A1(n6100), .A2(n5636), .B1(n6099), .B2(n5635), .ZN(n5622)
         );
  AND2_X1 U6561 ( .A1(n5631), .A2(DATAI_19_), .ZN(n6101) );
  AOI22_X1 U6562 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5637), .B1(n6101), 
        .B2(n5657), .ZN(n5621) );
  OAI211_X1 U6563 ( .C1(n6104), .C2(n5640), .A(n5622), .B(n5621), .ZN(U3023)
         );
  AND2_X1 U6564 ( .A1(n5631), .A2(DATAI_28_), .ZN(n6051) );
  INV_X1 U6565 ( .A(n6051), .ZN(n6110) );
  NOR2_X2 U6566 ( .A1(n5629), .A2(n3216), .ZN(n6106) );
  NOR2_X2 U6567 ( .A1(n5623), .A2(n5630), .ZN(n6105) );
  AOI22_X1 U6568 ( .A1(n6106), .A2(n5636), .B1(n6105), .B2(n5635), .ZN(n5625)
         );
  AND2_X1 U6569 ( .A1(n5631), .A2(DATAI_20_), .ZN(n6107) );
  AOI22_X1 U6570 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5637), .B1(n6107), 
        .B2(n5657), .ZN(n5624) );
  OAI211_X1 U6571 ( .C1(n6110), .C2(n5640), .A(n5625), .B(n5624), .ZN(U3024)
         );
  INV_X1 U6572 ( .A(n6055), .ZN(n6116) );
  AOI22_X1 U6573 ( .A1(n6112), .A2(n5636), .B1(n6111), .B2(n5635), .ZN(n5628)
         );
  AOI22_X1 U6574 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5637), .B1(n6113), 
        .B2(n5657), .ZN(n5627) );
  OAI211_X1 U6575 ( .C1(n6116), .C2(n5640), .A(n5628), .B(n5627), .ZN(U3025)
         );
  AND2_X1 U6576 ( .A1(n5631), .A2(DATAI_30_), .ZN(n6059) );
  INV_X1 U6577 ( .A(n6059), .ZN(n6122) );
  NOR2_X2 U6578 ( .A1(n5629), .A2(n3320), .ZN(n6118) );
  INV_X1 U6579 ( .A(DATAI_6_), .ZN(n6381) );
  NOR2_X2 U6580 ( .A1(n6381), .A2(n5630), .ZN(n6117) );
  AOI22_X1 U6581 ( .A1(n6118), .A2(n5636), .B1(n6117), .B2(n5635), .ZN(n5633)
         );
  AND2_X1 U6582 ( .A1(n5631), .A2(DATAI_22_), .ZN(n6119) );
  AOI22_X1 U6583 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5637), .B1(n6119), 
        .B2(n5657), .ZN(n5632) );
  OAI211_X1 U6584 ( .C1(n6122), .C2(n5640), .A(n5633), .B(n5632), .ZN(U3026)
         );
  INV_X1 U6585 ( .A(n6066), .ZN(n6133) );
  AOI22_X1 U6586 ( .A1(n6126), .A2(n5636), .B1(n6124), .B2(n5635), .ZN(n5639)
         );
  AOI22_X1 U6587 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5637), .B1(n6128), 
        .B2(n5657), .ZN(n5638) );
  OAI211_X1 U6588 ( .C1(n6133), .C2(n5640), .A(n5639), .B(n5638), .ZN(U3027)
         );
  INV_X1 U6589 ( .A(n6083), .ZN(n6038) );
  NOR2_X1 U6590 ( .A1(n6293), .A2(n5646), .ZN(n5664) );
  AOI22_X1 U6591 ( .A1(n6075), .A2(n5664), .B1(n6035), .B2(n5657), .ZN(n5650)
         );
  INV_X1 U6592 ( .A(n5641), .ZN(n5642) );
  AOI21_X1 U6593 ( .B1(n5642), .B2(n6288), .A(n5664), .ZN(n5648) );
  AOI21_X1 U6594 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5643), .A(n6275), .ZN(
        n5645) );
  AOI22_X1 U6595 ( .A1(n5648), .A2(n5645), .B1(n6275), .B2(n5646), .ZN(n5644)
         );
  NAND2_X1 U6596 ( .A1(n6082), .A2(n5644), .ZN(n5666) );
  INV_X1 U6597 ( .A(n5645), .ZN(n5647) );
  OAI22_X1 U6598 ( .A1(n5648), .A2(n5647), .B1(n5766), .B2(n5646), .ZN(n5665)
         );
  AOI22_X1 U6599 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5666), .B1(n6074), 
        .B2(n5665), .ZN(n5649) );
  OAI211_X1 U6600 ( .C1(n5695), .C2(n6038), .A(n5650), .B(n5649), .ZN(U3028)
         );
  INV_X1 U6601 ( .A(n6089), .ZN(n6042) );
  AOI22_X1 U6602 ( .A1(n6088), .A2(n5664), .B1(n6039), .B2(n5657), .ZN(n5652)
         );
  AOI22_X1 U6603 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5666), .B1(n6087), 
        .B2(n5665), .ZN(n5651) );
  OAI211_X1 U6604 ( .C1(n5695), .C2(n6042), .A(n5652), .B(n5651), .ZN(U3029)
         );
  AOI22_X1 U6605 ( .A1(n6094), .A2(n5664), .B1(n6095), .B2(n5672), .ZN(n5654)
         );
  AOI22_X1 U6606 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5666), .B1(n6093), 
        .B2(n5665), .ZN(n5653) );
  OAI211_X1 U6607 ( .C1(n6098), .C2(n5669), .A(n5654), .B(n5653), .ZN(U3030)
         );
  INV_X1 U6608 ( .A(n6101), .ZN(n6050) );
  AOI22_X1 U6609 ( .A1(n6100), .A2(n5664), .B1(n5657), .B2(n6047), .ZN(n5656)
         );
  AOI22_X1 U6610 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5666), .B1(n6099), 
        .B2(n5665), .ZN(n5655) );
  OAI211_X1 U6611 ( .C1(n5695), .C2(n6050), .A(n5656), .B(n5655), .ZN(U3031)
         );
  INV_X1 U6612 ( .A(n6107), .ZN(n6054) );
  AOI22_X1 U6613 ( .A1(n6106), .A2(n5664), .B1(n5657), .B2(n6051), .ZN(n5659)
         );
  AOI22_X1 U6614 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5666), .B1(n6105), 
        .B2(n5665), .ZN(n5658) );
  OAI211_X1 U6615 ( .C1(n5695), .C2(n6054), .A(n5659), .B(n5658), .ZN(U3032)
         );
  AOI22_X1 U6616 ( .A1(n6112), .A2(n5664), .B1(n6113), .B2(n5672), .ZN(n5661)
         );
  AOI22_X1 U6617 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5666), .B1(n6111), 
        .B2(n5665), .ZN(n5660) );
  OAI211_X1 U6618 ( .C1(n6116), .C2(n5669), .A(n5661), .B(n5660), .ZN(U3033)
         );
  AOI22_X1 U6619 ( .A1(n6118), .A2(n5664), .B1(n5672), .B2(n6119), .ZN(n5663)
         );
  AOI22_X1 U6620 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5666), .B1(n6117), 
        .B2(n5665), .ZN(n5662) );
  OAI211_X1 U6621 ( .C1(n6122), .C2(n5669), .A(n5663), .B(n5662), .ZN(U3034)
         );
  AOI22_X1 U6622 ( .A1(n6126), .A2(n5664), .B1(n6128), .B2(n5672), .ZN(n5668)
         );
  AOI22_X1 U6623 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5666), .B1(n6124), 
        .B2(n5665), .ZN(n5667) );
  OAI211_X1 U6624 ( .C1(n6133), .C2(n5669), .A(n5668), .B(n5667), .ZN(U3035)
         );
  NOR2_X1 U6625 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5670), .ZN(n5691)
         );
  NAND3_X1 U6626 ( .A1(n5968), .A2(n6022), .A3(n6284), .ZN(n5671) );
  OAI21_X1 U6627 ( .B1(n5673), .B2(n6275), .A(n5671), .ZN(n5690) );
  AOI22_X1 U6628 ( .A1(n6075), .A2(n5691), .B1(n6074), .B2(n5690), .ZN(n5677)
         );
  NAND2_X1 U6629 ( .A1(n6289), .A2(n6026), .ZN(n6280) );
  OAI21_X1 U6630 ( .B1(n5672), .B2(n5700), .A(n6280), .ZN(n5674) );
  AOI21_X1 U6631 ( .B1(n5674), .B2(n5673), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5675) );
  OAI21_X1 U6632 ( .B1(n6022), .B2(n5766), .A(n5831), .ZN(n5773) );
  NOR2_X1 U6633 ( .A1(n6023), .A2(n5773), .ZN(n5895) );
  AOI22_X1 U6634 ( .A1(n5692), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5700), 
        .B2(n6083), .ZN(n5676) );
  OAI211_X1 U6635 ( .C1(n6086), .C2(n5695), .A(n5677), .B(n5676), .ZN(U3036)
         );
  AOI22_X1 U6636 ( .A1(n6088), .A2(n5691), .B1(n6087), .B2(n5690), .ZN(n5679)
         );
  AOI22_X1 U6637 ( .A1(n5692), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5700), 
        .B2(n6089), .ZN(n5678) );
  OAI211_X1 U6638 ( .C1(n5695), .C2(n6092), .A(n5679), .B(n5678), .ZN(U3037)
         );
  AOI22_X1 U6639 ( .A1(n6094), .A2(n5691), .B1(n6093), .B2(n5690), .ZN(n5681)
         );
  AOI22_X1 U6640 ( .A1(n5692), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5700), 
        .B2(n6095), .ZN(n5680) );
  OAI211_X1 U6641 ( .C1(n5695), .C2(n6098), .A(n5681), .B(n5680), .ZN(U3038)
         );
  AOI22_X1 U6642 ( .A1(n6100), .A2(n5691), .B1(n6099), .B2(n5690), .ZN(n5683)
         );
  AOI22_X1 U6643 ( .A1(n5692), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5700), 
        .B2(n6101), .ZN(n5682) );
  OAI211_X1 U6644 ( .C1(n5695), .C2(n6104), .A(n5683), .B(n5682), .ZN(U3039)
         );
  AOI22_X1 U6645 ( .A1(n6106), .A2(n5691), .B1(n6105), .B2(n5690), .ZN(n5685)
         );
  AOI22_X1 U6646 ( .A1(n5692), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5700), 
        .B2(n6107), .ZN(n5684) );
  OAI211_X1 U6647 ( .C1(n5695), .C2(n6110), .A(n5685), .B(n5684), .ZN(U3040)
         );
  AOI22_X1 U6648 ( .A1(n6112), .A2(n5691), .B1(n6111), .B2(n5690), .ZN(n5687)
         );
  AOI22_X1 U6649 ( .A1(n5692), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5700), 
        .B2(n6113), .ZN(n5686) );
  OAI211_X1 U6650 ( .C1(n5695), .C2(n6116), .A(n5687), .B(n5686), .ZN(U3041)
         );
  AOI22_X1 U6651 ( .A1(n6118), .A2(n5691), .B1(n6117), .B2(n5690), .ZN(n5689)
         );
  AOI22_X1 U6652 ( .A1(n5692), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5700), 
        .B2(n6119), .ZN(n5688) );
  OAI211_X1 U6653 ( .C1(n5695), .C2(n6122), .A(n5689), .B(n5688), .ZN(U3042)
         );
  AOI22_X1 U6654 ( .A1(n6126), .A2(n5691), .B1(n6124), .B2(n5690), .ZN(n5694)
         );
  AOI22_X1 U6655 ( .A1(n5692), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5700), 
        .B2(n6128), .ZN(n5693) );
  OAI211_X1 U6656 ( .C1(n5695), .C2(n6133), .A(n5694), .B(n5693), .ZN(U3043)
         );
  AOI22_X1 U6657 ( .A1(n6100), .A2(n5701), .B1(n5700), .B2(n6047), .ZN(n5697)
         );
  AOI22_X1 U6658 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5703), .B1(n6099), 
        .B2(n5702), .ZN(n5696) );
  OAI211_X1 U6659 ( .C1(n6050), .C2(n5734), .A(n5697), .B(n5696), .ZN(U3047)
         );
  AOI22_X1 U6660 ( .A1(n6106), .A2(n5701), .B1(n5700), .B2(n6051), .ZN(n5699)
         );
  AOI22_X1 U6661 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5703), .B1(n6105), 
        .B2(n5702), .ZN(n5698) );
  OAI211_X1 U6662 ( .C1(n6054), .C2(n5734), .A(n5699), .B(n5698), .ZN(U3048)
         );
  INV_X1 U6663 ( .A(n6119), .ZN(n6062) );
  AOI22_X1 U6664 ( .A1(n6118), .A2(n5701), .B1(n5700), .B2(n6059), .ZN(n5705)
         );
  AOI22_X1 U6665 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5703), .B1(n6117), 
        .B2(n5702), .ZN(n5704) );
  OAI211_X1 U6666 ( .C1(n6062), .C2(n5734), .A(n5705), .B(n5704), .ZN(U3050)
         );
  NOR2_X1 U6667 ( .A1(n5706), .A2(n5926), .ZN(n5707) );
  NAND2_X1 U6668 ( .A1(n4452), .A2(n5707), .ZN(n5735) );
  NAND2_X1 U6669 ( .A1(n6140), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5993) );
  OR2_X1 U6670 ( .A1(n5993), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5739)
         );
  NOR2_X1 U6671 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5739), .ZN(n5730)
         );
  NOR2_X1 U6672 ( .A1(n4419), .A2(n5764), .ZN(n5992) );
  NAND2_X1 U6673 ( .A1(n5992), .A2(n6289), .ZN(n5963) );
  INV_X1 U6674 ( .A(n6023), .ZN(n5962) );
  OAI22_X1 U6675 ( .A1(n5963), .A2(n6029), .B1(n5708), .B2(n5962), .ZN(n5729)
         );
  AOI22_X1 U6676 ( .A1(n6075), .A2(n5730), .B1(n6074), .B2(n5729), .ZN(n5715)
         );
  AOI21_X1 U6677 ( .B1(n5734), .B2(n5763), .A(n6026), .ZN(n5709) );
  AOI211_X1 U6678 ( .C1(n5710), .C2(n5992), .A(n6275), .B(n5709), .ZN(n5711)
         );
  NOR3_X1 U6679 ( .A1(n5712), .A2(n5968), .A3(n5711), .ZN(n5713) );
  AOI22_X1 U6680 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n5731), .B1(n6035), 
        .B2(n5726), .ZN(n5714) );
  OAI211_X1 U6681 ( .C1(n6038), .C2(n5763), .A(n5715), .B(n5714), .ZN(U3052)
         );
  AOI22_X1 U6682 ( .A1(n6088), .A2(n5730), .B1(n6087), .B2(n5729), .ZN(n5717)
         );
  AOI22_X1 U6683 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n5731), .B1(n6039), 
        .B2(n5726), .ZN(n5716) );
  OAI211_X1 U6684 ( .C1(n6042), .C2(n5763), .A(n5717), .B(n5716), .ZN(U3053)
         );
  AOI22_X1 U6685 ( .A1(n6094), .A2(n5730), .B1(n6093), .B2(n5729), .ZN(n5719)
         );
  AOI22_X1 U6686 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n5731), .B1(n6095), 
        .B2(n5748), .ZN(n5718) );
  OAI211_X1 U6687 ( .C1(n6098), .C2(n5734), .A(n5719), .B(n5718), .ZN(U3054)
         );
  AOI22_X1 U6688 ( .A1(n6100), .A2(n5730), .B1(n6099), .B2(n5729), .ZN(n5721)
         );
  AOI22_X1 U6689 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n5731), .B1(n6047), 
        .B2(n5726), .ZN(n5720) );
  OAI211_X1 U6690 ( .C1(n6050), .C2(n5763), .A(n5721), .B(n5720), .ZN(U3055)
         );
  AOI22_X1 U6691 ( .A1(n6106), .A2(n5730), .B1(n6105), .B2(n5729), .ZN(n5723)
         );
  AOI22_X1 U6692 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5731), .B1(n6051), 
        .B2(n5726), .ZN(n5722) );
  OAI211_X1 U6693 ( .C1(n6054), .C2(n5763), .A(n5723), .B(n5722), .ZN(U3056)
         );
  AOI22_X1 U6694 ( .A1(n6112), .A2(n5730), .B1(n6111), .B2(n5729), .ZN(n5725)
         );
  AOI22_X1 U6695 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n5731), .B1(n6113), 
        .B2(n5748), .ZN(n5724) );
  OAI211_X1 U6696 ( .C1(n6116), .C2(n5734), .A(n5725), .B(n5724), .ZN(U3057)
         );
  AOI22_X1 U6697 ( .A1(n6118), .A2(n5730), .B1(n6117), .B2(n5729), .ZN(n5728)
         );
  AOI22_X1 U6698 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n5731), .B1(n6059), 
        .B2(n5726), .ZN(n5727) );
  OAI211_X1 U6699 ( .C1(n6062), .C2(n5763), .A(n5728), .B(n5727), .ZN(U3058)
         );
  AOI22_X1 U6700 ( .A1(n6126), .A2(n5730), .B1(n6124), .B2(n5729), .ZN(n5733)
         );
  AOI22_X1 U6701 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n5731), .B1(n6128), 
        .B2(n5748), .ZN(n5732) );
  OAI211_X1 U6702 ( .C1(n6133), .C2(n5734), .A(n5733), .B(n5732), .ZN(U3059)
         );
  NOR2_X1 U6703 ( .A1(n6293), .A2(n5739), .ZN(n5758) );
  AOI22_X1 U6704 ( .A1(n6075), .A2(n5758), .B1(n6035), .B2(n5748), .ZN(n5743)
         );
  NOR2_X1 U6705 ( .A1(n5921), .A2(n5966), .ZN(n5798) );
  AOI21_X1 U6706 ( .B1(n5992), .B2(n5798), .A(n5758), .ZN(n5741) );
  INV_X1 U6707 ( .A(n5741), .ZN(n5738) );
  OAI21_X1 U6708 ( .B1(n6026), .B2(n5735), .A(n6289), .ZN(n5740) );
  AOI21_X1 U6709 ( .B1(n6275), .B2(n5739), .A(n5736), .ZN(n5737) );
  OAI21_X1 U6710 ( .B1(n5738), .B2(n5740), .A(n5737), .ZN(n5760) );
  OAI22_X1 U6711 ( .A1(n5741), .A2(n5740), .B1(n5766), .B2(n5739), .ZN(n5759)
         );
  AOI22_X1 U6712 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5760), .B1(n6074), 
        .B2(n5759), .ZN(n5742) );
  OAI211_X1 U6713 ( .C1(n6038), .C2(n5795), .A(n5743), .B(n5742), .ZN(U3060)
         );
  AOI22_X1 U6714 ( .A1(n6088), .A2(n5758), .B1(n6039), .B2(n5748), .ZN(n5745)
         );
  AOI22_X1 U6715 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5760), .B1(n6087), 
        .B2(n5759), .ZN(n5744) );
  OAI211_X1 U6716 ( .C1(n6042), .C2(n5795), .A(n5745), .B(n5744), .ZN(U3061)
         );
  INV_X1 U6717 ( .A(n6095), .ZN(n6046) );
  AOI22_X1 U6718 ( .A1(n6094), .A2(n5758), .B1(n6043), .B2(n5748), .ZN(n5747)
         );
  AOI22_X1 U6719 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5760), .B1(n6093), 
        .B2(n5759), .ZN(n5746) );
  OAI211_X1 U6720 ( .C1(n6046), .C2(n5795), .A(n5747), .B(n5746), .ZN(U3062)
         );
  AOI22_X1 U6721 ( .A1(n6100), .A2(n5758), .B1(n5748), .B2(n6047), .ZN(n5750)
         );
  AOI22_X1 U6722 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5760), .B1(n6099), 
        .B2(n5759), .ZN(n5749) );
  OAI211_X1 U6723 ( .C1(n6050), .C2(n5795), .A(n5750), .B(n5749), .ZN(U3063)
         );
  INV_X1 U6724 ( .A(n5795), .ZN(n5757) );
  AOI22_X1 U6725 ( .A1(n6106), .A2(n5758), .B1(n6107), .B2(n5757), .ZN(n5752)
         );
  AOI22_X1 U6726 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5760), .B1(n6105), 
        .B2(n5759), .ZN(n5751) );
  OAI211_X1 U6727 ( .C1(n6110), .C2(n5763), .A(n5752), .B(n5751), .ZN(U3064)
         );
  AOI22_X1 U6728 ( .A1(n6112), .A2(n5758), .B1(n6113), .B2(n5757), .ZN(n5754)
         );
  AOI22_X1 U6729 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5760), .B1(n6111), 
        .B2(n5759), .ZN(n5753) );
  OAI211_X1 U6730 ( .C1(n6116), .C2(n5763), .A(n5754), .B(n5753), .ZN(U3065)
         );
  AOI22_X1 U6731 ( .A1(n6118), .A2(n5758), .B1(n6119), .B2(n5757), .ZN(n5756)
         );
  AOI22_X1 U6732 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5760), .B1(n6117), 
        .B2(n5759), .ZN(n5755) );
  OAI211_X1 U6733 ( .C1(n6122), .C2(n5763), .A(n5756), .B(n5755), .ZN(U3066)
         );
  AOI22_X1 U6734 ( .A1(n6126), .A2(n5758), .B1(n6128), .B2(n5757), .ZN(n5762)
         );
  AOI22_X1 U6735 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5760), .B1(n6124), 
        .B2(n5759), .ZN(n5761) );
  OAI211_X1 U6736 ( .C1(n6133), .C2(n5763), .A(n5762), .B(n5761), .ZN(U3067)
         );
  NAND2_X1 U6737 ( .A1(n6293), .A2(n5805), .ZN(n5772) );
  INV_X1 U6738 ( .A(n5772), .ZN(n5791) );
  NAND2_X1 U6739 ( .A1(n6072), .A2(n6289), .ZN(n6025) );
  NOR2_X1 U6740 ( .A1(n5766), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6030)
         );
  NAND3_X1 U6741 ( .A1(n5767), .A2(n6022), .A3(n6030), .ZN(n5768) );
  OAI21_X1 U6742 ( .B1(n6025), .B2(n6029), .A(n5768), .ZN(n5790) );
  AOI22_X1 U6743 ( .A1(n6075), .A2(n5791), .B1(n6074), .B2(n5790), .ZN(n5777)
         );
  AND2_X1 U6744 ( .A1(n5926), .A2(n5797), .ZN(n5769) );
  NAND2_X1 U6745 ( .A1(n4452), .A2(n5769), .ZN(n5806) );
  OR2_X1 U6746 ( .A1(n5806), .A2(n6290), .ZN(n5775) );
  NAND3_X1 U6747 ( .A1(n5795), .A2(n5775), .A3(n6289), .ZN(n5770) );
  AOI21_X1 U6748 ( .B1(n6280), .B2(n5770), .A(n6072), .ZN(n5771) );
  AOI21_X1 U6749 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5772), .A(n5771), .ZN(
        n5774) );
  NOR2_X1 U6750 ( .A1(n5968), .A2(n5773), .ZN(n6033) );
  NAND3_X1 U6751 ( .A1(n6284), .A2(n5774), .A3(n6033), .ZN(n5792) );
  AOI22_X1 U6752 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n5792), .B1(n6083), 
        .B2(n5822), .ZN(n5776) );
  OAI211_X1 U6753 ( .C1(n6086), .C2(n5795), .A(n5777), .B(n5776), .ZN(U3068)
         );
  AOI22_X1 U6754 ( .A1(n6088), .A2(n5791), .B1(n6087), .B2(n5790), .ZN(n5779)
         );
  AOI22_X1 U6755 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n5792), .B1(n6089), 
        .B2(n5822), .ZN(n5778) );
  OAI211_X1 U6756 ( .C1(n6092), .C2(n5795), .A(n5779), .B(n5778), .ZN(U3069)
         );
  AOI22_X1 U6757 ( .A1(n6094), .A2(n5791), .B1(n6093), .B2(n5790), .ZN(n5781)
         );
  AOI22_X1 U6758 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n5792), .B1(n6095), 
        .B2(n5822), .ZN(n5780) );
  OAI211_X1 U6759 ( .C1(n6098), .C2(n5795), .A(n5781), .B(n5780), .ZN(U3070)
         );
  AOI22_X1 U6760 ( .A1(n6100), .A2(n5791), .B1(n6099), .B2(n5790), .ZN(n5783)
         );
  AOI22_X1 U6761 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n5792), .B1(n6101), 
        .B2(n5822), .ZN(n5782) );
  OAI211_X1 U6762 ( .C1(n6104), .C2(n5795), .A(n5783), .B(n5782), .ZN(U3071)
         );
  AOI22_X1 U6763 ( .A1(n6106), .A2(n5791), .B1(n6105), .B2(n5790), .ZN(n5785)
         );
  AOI22_X1 U6764 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5792), .B1(n6107), 
        .B2(n5822), .ZN(n5784) );
  OAI211_X1 U6765 ( .C1(n6110), .C2(n5795), .A(n5785), .B(n5784), .ZN(U3072)
         );
  AOI22_X1 U6766 ( .A1(n6112), .A2(n5791), .B1(n6111), .B2(n5790), .ZN(n5787)
         );
  AOI22_X1 U6767 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n5792), .B1(n6113), 
        .B2(n5822), .ZN(n5786) );
  OAI211_X1 U6768 ( .C1(n6116), .C2(n5795), .A(n5787), .B(n5786), .ZN(U3073)
         );
  AOI22_X1 U6769 ( .A1(n6118), .A2(n5791), .B1(n6117), .B2(n5790), .ZN(n5789)
         );
  AOI22_X1 U6770 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n5792), .B1(n6119), 
        .B2(n5822), .ZN(n5788) );
  OAI211_X1 U6771 ( .C1(n6122), .C2(n5795), .A(n5789), .B(n5788), .ZN(U3074)
         );
  AOI22_X1 U6772 ( .A1(n6126), .A2(n5791), .B1(n6124), .B2(n5790), .ZN(n5794)
         );
  AOI22_X1 U6773 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n5792), .B1(n6128), 
        .B2(n5822), .ZN(n5793) );
  OAI211_X1 U6774 ( .C1(n6133), .C2(n5795), .A(n5794), .B(n5793), .ZN(U3075)
         );
  NAND3_X1 U6775 ( .A1(n4452), .A2(n5797), .A3(n5796), .ZN(n6276) );
  AND2_X1 U6776 ( .A1(n6276), .A2(n6289), .ZN(n5803) );
  NAND2_X1 U6777 ( .A1(n6072), .A2(n5798), .ZN(n5799) );
  NAND2_X1 U6778 ( .A1(n5799), .A2(n5800), .ZN(n5801) );
  AOI22_X1 U6779 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5805), .B1(n5803), .B2(
        n5801), .ZN(n5826) );
  INV_X1 U6780 ( .A(n6074), .ZN(n5935) );
  INV_X1 U6781 ( .A(n5800), .ZN(n5821) );
  AOI22_X1 U6782 ( .A1(n6075), .A2(n5821), .B1(n6035), .B2(n5822), .ZN(n5808)
         );
  INV_X1 U6783 ( .A(n5801), .ZN(n5802) );
  NAND2_X1 U6784 ( .A1(n5803), .A2(n5802), .ZN(n5804) );
  OAI211_X1 U6785 ( .C1(n6289), .C2(n5805), .A(n6082), .B(n5804), .ZN(n5823)
         );
  AOI22_X1 U6786 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5823), .B1(n6083), 
        .B2(n5850), .ZN(n5807) );
  OAI211_X1 U6787 ( .C1(n5826), .C2(n5935), .A(n5808), .B(n5807), .ZN(U3076)
         );
  INV_X1 U6788 ( .A(n6087), .ZN(n5938) );
  AOI22_X1 U6789 ( .A1(n6088), .A2(n5821), .B1(n6039), .B2(n5822), .ZN(n5810)
         );
  AOI22_X1 U6790 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5823), .B1(n6089), 
        .B2(n5850), .ZN(n5809) );
  OAI211_X1 U6791 ( .C1(n5826), .C2(n5938), .A(n5810), .B(n5809), .ZN(U3077)
         );
  INV_X1 U6792 ( .A(n6093), .ZN(n5941) );
  AOI22_X1 U6793 ( .A1(n6094), .A2(n5821), .B1(n6043), .B2(n5822), .ZN(n5812)
         );
  AOI22_X1 U6794 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5823), .B1(n6095), 
        .B2(n5850), .ZN(n5811) );
  OAI211_X1 U6795 ( .C1(n5826), .C2(n5941), .A(n5812), .B(n5811), .ZN(U3078)
         );
  INV_X1 U6796 ( .A(n6099), .ZN(n5944) );
  AOI22_X1 U6797 ( .A1(n6100), .A2(n5821), .B1(n6101), .B2(n5850), .ZN(n5814)
         );
  AOI22_X1 U6798 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5823), .B1(n6047), 
        .B2(n5822), .ZN(n5813) );
  OAI211_X1 U6799 ( .C1(n5826), .C2(n5944), .A(n5814), .B(n5813), .ZN(U3079)
         );
  INV_X1 U6800 ( .A(n6105), .ZN(n5947) );
  AOI22_X1 U6801 ( .A1(n6106), .A2(n5821), .B1(n5822), .B2(n6051), .ZN(n5816)
         );
  AOI22_X1 U6802 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5823), .B1(n6107), 
        .B2(n5850), .ZN(n5815) );
  OAI211_X1 U6803 ( .C1(n5826), .C2(n5947), .A(n5816), .B(n5815), .ZN(U3080)
         );
  INV_X1 U6804 ( .A(n6111), .ZN(n5950) );
  AOI22_X1 U6805 ( .A1(n6112), .A2(n5821), .B1(n6055), .B2(n5822), .ZN(n5818)
         );
  AOI22_X1 U6806 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5823), .B1(n6113), 
        .B2(n5850), .ZN(n5817) );
  OAI211_X1 U6807 ( .C1(n5826), .C2(n5950), .A(n5818), .B(n5817), .ZN(U3081)
         );
  INV_X1 U6808 ( .A(n6117), .ZN(n5953) );
  AOI22_X1 U6809 ( .A1(n6118), .A2(n5821), .B1(n6119), .B2(n5850), .ZN(n5820)
         );
  AOI22_X1 U6810 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5823), .B1(n6059), 
        .B2(n5822), .ZN(n5819) );
  OAI211_X1 U6811 ( .C1(n5826), .C2(n5953), .A(n5820), .B(n5819), .ZN(U3082)
         );
  INV_X1 U6812 ( .A(n6124), .ZN(n5959) );
  AOI22_X1 U6813 ( .A1(n6126), .A2(n5821), .B1(n6128), .B2(n5850), .ZN(n5825)
         );
  AOI22_X1 U6814 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5823), .B1(n6066), 
        .B2(n5822), .ZN(n5824) );
  OAI211_X1 U6815 ( .C1(n5826), .C2(n5959), .A(n5825), .B(n5824), .ZN(U3083)
         );
  NAND2_X1 U6816 ( .A1(n5859), .A2(n3920), .ZN(n5875) );
  NAND3_X1 U6817 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6145), .A3(n6140), .ZN(n5863) );
  NOR2_X1 U6818 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5863), .ZN(n5854)
         );
  INV_X1 U6819 ( .A(n5827), .ZN(n5860) );
  NAND2_X1 U6820 ( .A1(n5860), .A2(n6029), .ZN(n5834) );
  INV_X1 U6821 ( .A(n5828), .ZN(n5829) );
  NOR2_X1 U6822 ( .A1(n5829), .A2(n6022), .ZN(n5832) );
  INV_X1 U6823 ( .A(n5832), .ZN(n5961) );
  OAI22_X1 U6824 ( .A1(n5834), .A2(n6275), .B1(n5830), .B2(n5961), .ZN(n5853)
         );
  AOI22_X1 U6825 ( .A1(n6075), .A2(n5854), .B1(n6074), .B2(n5853), .ZN(n5839)
         );
  INV_X1 U6826 ( .A(n5854), .ZN(n5833) );
  OAI21_X1 U6827 ( .B1(n5832), .B2(n5766), .A(n5831), .ZN(n5970) );
  AOI211_X1 U6828 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5833), .A(n6023), .B(
        n5970), .ZN(n5837) );
  OAI21_X1 U6829 ( .B1(n5882), .B2(n5850), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5835) );
  NAND3_X1 U6830 ( .A1(n5835), .A2(n6289), .A3(n5834), .ZN(n5836) );
  NAND2_X1 U6831 ( .A1(n5837), .A2(n5836), .ZN(n5855) );
  AOI22_X1 U6832 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5855), .B1(n6035), 
        .B2(n5850), .ZN(n5838) );
  OAI211_X1 U6833 ( .C1(n6038), .C2(n5875), .A(n5839), .B(n5838), .ZN(U3084)
         );
  AOI22_X1 U6834 ( .A1(n6088), .A2(n5854), .B1(n6087), .B2(n5853), .ZN(n5841)
         );
  AOI22_X1 U6835 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n5855), .B1(n6039), 
        .B2(n5850), .ZN(n5840) );
  OAI211_X1 U6836 ( .C1(n6042), .C2(n5875), .A(n5841), .B(n5840), .ZN(U3085)
         );
  AOI22_X1 U6837 ( .A1(n6094), .A2(n5854), .B1(n6093), .B2(n5853), .ZN(n5843)
         );
  AOI22_X1 U6838 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n5855), .B1(n6095), 
        .B2(n5882), .ZN(n5842) );
  OAI211_X1 U6839 ( .C1(n6098), .C2(n5858), .A(n5843), .B(n5842), .ZN(U3086)
         );
  AOI22_X1 U6840 ( .A1(n6100), .A2(n5854), .B1(n6099), .B2(n5853), .ZN(n5845)
         );
  AOI22_X1 U6841 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n5855), .B1(n6047), 
        .B2(n5850), .ZN(n5844) );
  OAI211_X1 U6842 ( .C1(n6050), .C2(n5875), .A(n5845), .B(n5844), .ZN(U3087)
         );
  AOI22_X1 U6843 ( .A1(n6106), .A2(n5854), .B1(n6105), .B2(n5853), .ZN(n5847)
         );
  AOI22_X1 U6844 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5855), .B1(n6051), 
        .B2(n5850), .ZN(n5846) );
  OAI211_X1 U6845 ( .C1(n6054), .C2(n5875), .A(n5847), .B(n5846), .ZN(U3088)
         );
  AOI22_X1 U6846 ( .A1(n6112), .A2(n5854), .B1(n6111), .B2(n5853), .ZN(n5849)
         );
  AOI22_X1 U6847 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n5855), .B1(n6113), 
        .B2(n5882), .ZN(n5848) );
  OAI211_X1 U6848 ( .C1(n6116), .C2(n5858), .A(n5849), .B(n5848), .ZN(U3089)
         );
  AOI22_X1 U6849 ( .A1(n6118), .A2(n5854), .B1(n6117), .B2(n5853), .ZN(n5852)
         );
  AOI22_X1 U6850 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n5855), .B1(n6059), 
        .B2(n5850), .ZN(n5851) );
  OAI211_X1 U6851 ( .C1(n6062), .C2(n5875), .A(n5852), .B(n5851), .ZN(U3090)
         );
  AOI22_X1 U6852 ( .A1(n6126), .A2(n5854), .B1(n6124), .B2(n5853), .ZN(n5857)
         );
  AOI22_X1 U6853 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n5855), .B1(n6128), 
        .B2(n5882), .ZN(n5856) );
  OAI211_X1 U6854 ( .C1(n6133), .C2(n5858), .A(n5857), .B(n5856), .ZN(U3091)
         );
  NOR2_X1 U6855 ( .A1(n6293), .A2(n5863), .ZN(n5883) );
  INV_X1 U6856 ( .A(n5918), .ZN(n5872) );
  AOI22_X1 U6857 ( .A1(n6075), .A2(n5883), .B1(n6083), .B2(n5872), .ZN(n5867)
         );
  AOI21_X1 U6858 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5859), .A(n6275), .ZN(
        n5862) );
  NOR2_X1 U6859 ( .A1(n6279), .A2(n5921), .ZN(n6073) );
  AOI21_X1 U6860 ( .B1(n6073), .B2(n5860), .A(n5883), .ZN(n5865) );
  AOI22_X1 U6861 ( .A1(n5862), .A2(n5865), .B1(n6275), .B2(n5863), .ZN(n5861)
         );
  NAND2_X1 U6862 ( .A1(n6082), .A2(n5861), .ZN(n5885) );
  INV_X1 U6863 ( .A(n5862), .ZN(n5864) );
  OAI22_X1 U6864 ( .A1(n5865), .A2(n5864), .B1(n5766), .B2(n5863), .ZN(n5884)
         );
  AOI22_X1 U6865 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5885), .B1(n6074), 
        .B2(n5884), .ZN(n5866) );
  OAI211_X1 U6866 ( .C1(n6086), .C2(n5875), .A(n5867), .B(n5866), .ZN(U3092)
         );
  AOI22_X1 U6867 ( .A1(n6088), .A2(n5883), .B1(n6039), .B2(n5882), .ZN(n5869)
         );
  AOI22_X1 U6868 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5885), .B1(n6087), 
        .B2(n5884), .ZN(n5868) );
  OAI211_X1 U6869 ( .C1(n6042), .C2(n5918), .A(n5869), .B(n5868), .ZN(U3093)
         );
  AOI22_X1 U6870 ( .A1(n6094), .A2(n5883), .B1(n6043), .B2(n5882), .ZN(n5871)
         );
  AOI22_X1 U6871 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5885), .B1(n6093), 
        .B2(n5884), .ZN(n5870) );
  OAI211_X1 U6872 ( .C1(n6046), .C2(n5918), .A(n5871), .B(n5870), .ZN(U3094)
         );
  AOI22_X1 U6873 ( .A1(n6100), .A2(n5883), .B1(n6101), .B2(n5872), .ZN(n5874)
         );
  AOI22_X1 U6874 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5885), .B1(n6099), 
        .B2(n5884), .ZN(n5873) );
  OAI211_X1 U6875 ( .C1(n6104), .C2(n5875), .A(n5874), .B(n5873), .ZN(U3095)
         );
  AOI22_X1 U6876 ( .A1(n6106), .A2(n5883), .B1(n5882), .B2(n6051), .ZN(n5877)
         );
  AOI22_X1 U6877 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5885), .B1(n6105), 
        .B2(n5884), .ZN(n5876) );
  OAI211_X1 U6878 ( .C1(n6054), .C2(n5918), .A(n5877), .B(n5876), .ZN(U3096)
         );
  INV_X1 U6879 ( .A(n6113), .ZN(n6058) );
  AOI22_X1 U6880 ( .A1(n6112), .A2(n5883), .B1(n6055), .B2(n5882), .ZN(n5879)
         );
  AOI22_X1 U6881 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5885), .B1(n6111), 
        .B2(n5884), .ZN(n5878) );
  OAI211_X1 U6882 ( .C1(n6058), .C2(n5918), .A(n5879), .B(n5878), .ZN(U3097)
         );
  AOI22_X1 U6883 ( .A1(n6118), .A2(n5883), .B1(n5882), .B2(n6059), .ZN(n5881)
         );
  AOI22_X1 U6884 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5885), .B1(n6117), 
        .B2(n5884), .ZN(n5880) );
  OAI211_X1 U6885 ( .C1(n6062), .C2(n5918), .A(n5881), .B(n5880), .ZN(U3098)
         );
  INV_X1 U6886 ( .A(n6128), .ZN(n6070) );
  AOI22_X1 U6887 ( .A1(n6126), .A2(n5883), .B1(n6066), .B2(n5882), .ZN(n5887)
         );
  AOI22_X1 U6888 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5885), .B1(n6124), 
        .B2(n5884), .ZN(n5886) );
  OAI211_X1 U6889 ( .C1(n6070), .C2(n5918), .A(n5887), .B(n5886), .ZN(U3099)
         );
  NAND3_X1 U6890 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6145), .ZN(n5929) );
  NOR2_X1 U6891 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5929), .ZN(n5913)
         );
  NAND2_X1 U6892 ( .A1(n5926), .A2(n3920), .ZN(n5888) );
  AOI22_X1 U6893 ( .A1(n6075), .A2(n5913), .B1(n6083), .B2(n5954), .ZN(n5900)
         );
  NAND3_X1 U6894 ( .A1(n5918), .A2(n6289), .A3(n5889), .ZN(n5890) );
  NAND2_X1 U6895 ( .A1(n5890), .A2(n6280), .ZN(n5896) );
  INV_X1 U6896 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U6897 ( .A1(n5892), .A2(n6029), .ZN(n5922) );
  INV_X1 U6898 ( .A(n5913), .ZN(n5893) );
  AOI22_X1 U6899 ( .A1(n5896), .A2(n5922), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5893), .ZN(n5894) );
  OAI211_X1 U6900 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5766), .A(n5895), .B(n5894), .ZN(n5915) );
  INV_X1 U6901 ( .A(n5896), .ZN(n5898) );
  NAND3_X1 U6902 ( .A1(n5968), .A2(n6022), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5897) );
  OAI21_X1 U6903 ( .B1(n5898), .B2(n5922), .A(n5897), .ZN(n5914) );
  AOI22_X1 U6904 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n5915), .B1(n6074), 
        .B2(n5914), .ZN(n5899) );
  OAI211_X1 U6905 ( .C1(n6086), .C2(n5918), .A(n5900), .B(n5899), .ZN(U3100)
         );
  AOI22_X1 U6906 ( .A1(n6088), .A2(n5913), .B1(n6089), .B2(n5954), .ZN(n5902)
         );
  AOI22_X1 U6907 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n5915), .B1(n6087), 
        .B2(n5914), .ZN(n5901) );
  OAI211_X1 U6908 ( .C1(n6092), .C2(n5918), .A(n5902), .B(n5901), .ZN(U3101)
         );
  AOI22_X1 U6909 ( .A1(n6094), .A2(n5913), .B1(n6095), .B2(n5954), .ZN(n5904)
         );
  AOI22_X1 U6910 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n5915), .B1(n6093), 
        .B2(n5914), .ZN(n5903) );
  OAI211_X1 U6911 ( .C1(n6098), .C2(n5918), .A(n5904), .B(n5903), .ZN(U3102)
         );
  AOI22_X1 U6912 ( .A1(n6100), .A2(n5913), .B1(n6101), .B2(n5954), .ZN(n5906)
         );
  AOI22_X1 U6913 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n5915), .B1(n6099), 
        .B2(n5914), .ZN(n5905) );
  OAI211_X1 U6914 ( .C1(n6104), .C2(n5918), .A(n5906), .B(n5905), .ZN(U3103)
         );
  AOI22_X1 U6915 ( .A1(n6106), .A2(n5913), .B1(n6107), .B2(n5954), .ZN(n5908)
         );
  AOI22_X1 U6916 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5915), .B1(n6105), 
        .B2(n5914), .ZN(n5907) );
  OAI211_X1 U6917 ( .C1(n6110), .C2(n5918), .A(n5908), .B(n5907), .ZN(U3104)
         );
  AOI22_X1 U6918 ( .A1(n6112), .A2(n5913), .B1(n6113), .B2(n5954), .ZN(n5910)
         );
  AOI22_X1 U6919 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n5915), .B1(n6111), 
        .B2(n5914), .ZN(n5909) );
  OAI211_X1 U6920 ( .C1(n6116), .C2(n5918), .A(n5910), .B(n5909), .ZN(U3105)
         );
  AOI22_X1 U6921 ( .A1(n6118), .A2(n5913), .B1(n6119), .B2(n5954), .ZN(n5912)
         );
  AOI22_X1 U6922 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n5915), .B1(n6117), 
        .B2(n5914), .ZN(n5911) );
  OAI211_X1 U6923 ( .C1(n6122), .C2(n5918), .A(n5912), .B(n5911), .ZN(U3106)
         );
  AOI22_X1 U6924 ( .A1(n6126), .A2(n5913), .B1(n6128), .B2(n5954), .ZN(n5917)
         );
  AOI22_X1 U6925 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n5915), .B1(n6124), 
        .B2(n5914), .ZN(n5916) );
  OAI211_X1 U6926 ( .C1(n6133), .C2(n5918), .A(n5917), .B(n5916), .ZN(U3107)
         );
  OAI21_X1 U6927 ( .B1(n5928), .B2(n5919), .A(n6289), .ZN(n5932) );
  INV_X1 U6928 ( .A(n5932), .ZN(n5924) );
  NAND2_X1 U6929 ( .A1(n5920), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U6930 ( .B1(n5922), .B2(n5921), .A(n5925), .ZN(n5931) );
  INV_X1 U6931 ( .A(n5929), .ZN(n5923) );
  AOI22_X1 U6932 ( .A1(n5924), .A2(n5931), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5923), .ZN(n5960) );
  INV_X1 U6933 ( .A(n5925), .ZN(n5955) );
  NAND2_X1 U6934 ( .A1(n5926), .A2(n6290), .ZN(n5927) );
  AOI22_X1 U6935 ( .A1(n6075), .A2(n5955), .B1(n6083), .B2(n5987), .ZN(n5934)
         );
  NAND2_X1 U6936 ( .A1(n6275), .A2(n5929), .ZN(n5930) );
  OAI211_X1 U6937 ( .C1(n5932), .C2(n5931), .A(n6082), .B(n5930), .ZN(n5956)
         );
  AOI22_X1 U6938 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n5956), .B1(n6035), 
        .B2(n5954), .ZN(n5933) );
  OAI211_X1 U6939 ( .C1(n5960), .C2(n5935), .A(n5934), .B(n5933), .ZN(U3108)
         );
  AOI22_X1 U6940 ( .A1(n6088), .A2(n5955), .B1(n6089), .B2(n5987), .ZN(n5937)
         );
  AOI22_X1 U6941 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n5956), .B1(n6039), 
        .B2(n5954), .ZN(n5936) );
  OAI211_X1 U6942 ( .C1(n5960), .C2(n5938), .A(n5937), .B(n5936), .ZN(U3109)
         );
  AOI22_X1 U6943 ( .A1(n6094), .A2(n5955), .B1(n6043), .B2(n5954), .ZN(n5940)
         );
  AOI22_X1 U6944 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n5956), .B1(n6095), 
        .B2(n5987), .ZN(n5939) );
  OAI211_X1 U6945 ( .C1(n5960), .C2(n5941), .A(n5940), .B(n5939), .ZN(U3110)
         );
  AOI22_X1 U6946 ( .A1(n6100), .A2(n5955), .B1(n6101), .B2(n5987), .ZN(n5943)
         );
  AOI22_X1 U6947 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n5956), .B1(n6047), 
        .B2(n5954), .ZN(n5942) );
  OAI211_X1 U6948 ( .C1(n5960), .C2(n5944), .A(n5943), .B(n5942), .ZN(U3111)
         );
  AOI22_X1 U6949 ( .A1(n6106), .A2(n5955), .B1(n6107), .B2(n5987), .ZN(n5946)
         );
  AOI22_X1 U6950 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5956), .B1(n6051), 
        .B2(n5954), .ZN(n5945) );
  OAI211_X1 U6951 ( .C1(n5960), .C2(n5947), .A(n5946), .B(n5945), .ZN(U3112)
         );
  AOI22_X1 U6952 ( .A1(n6112), .A2(n5955), .B1(n6113), .B2(n5987), .ZN(n5949)
         );
  AOI22_X1 U6953 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n5956), .B1(n6055), 
        .B2(n5954), .ZN(n5948) );
  OAI211_X1 U6954 ( .C1(n5960), .C2(n5950), .A(n5949), .B(n5948), .ZN(U3113)
         );
  AOI22_X1 U6955 ( .A1(n6118), .A2(n5955), .B1(n6059), .B2(n5954), .ZN(n5952)
         );
  AOI22_X1 U6956 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n5956), .B1(n6119), 
        .B2(n5987), .ZN(n5951) );
  OAI211_X1 U6957 ( .C1(n5960), .C2(n5953), .A(n5952), .B(n5951), .ZN(U3114)
         );
  AOI22_X1 U6958 ( .A1(n6126), .A2(n5955), .B1(n6066), .B2(n5954), .ZN(n5958)
         );
  AOI22_X1 U6959 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n5956), .B1(n6128), 
        .B2(n5987), .ZN(n5957) );
  OAI211_X1 U6960 ( .C1(n5960), .C2(n5959), .A(n5958), .B(n5957), .ZN(U3115)
         );
  NOR2_X1 U6961 ( .A1(n6284), .A2(n5993), .ZN(n5998) );
  INV_X1 U6962 ( .A(n5998), .ZN(n5991) );
  NOR2_X1 U6963 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5991), .ZN(n5986)
         );
  OAI22_X1 U6964 ( .A1(n5963), .A2(n6279), .B1(n5962), .B2(n5961), .ZN(n5985)
         );
  AOI22_X1 U6965 ( .A1(n6075), .A2(n5986), .B1(n6074), .B2(n5985), .ZN(n5972)
         );
  AOI21_X1 U6966 ( .B1(n5964), .B2(n6020), .A(n6026), .ZN(n5965) );
  AOI211_X1 U6967 ( .C1(n5992), .C2(n5966), .A(n6275), .B(n5965), .ZN(n5969)
         );
  NOR2_X1 U6968 ( .A1(n5986), .A2(n6034), .ZN(n5967) );
  AOI22_X1 U6969 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n5988), .B1(n6035), 
        .B2(n5987), .ZN(n5971) );
  OAI211_X1 U6970 ( .C1(n6038), .C2(n6020), .A(n5972), .B(n5971), .ZN(U3116)
         );
  AOI22_X1 U6971 ( .A1(n6088), .A2(n5986), .B1(n6087), .B2(n5985), .ZN(n5974)
         );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n5988), .B1(n6039), 
        .B2(n5987), .ZN(n5973) );
  OAI211_X1 U6973 ( .C1(n6042), .C2(n6020), .A(n5974), .B(n5973), .ZN(U3117)
         );
  AOI22_X1 U6974 ( .A1(n6094), .A2(n5986), .B1(n6093), .B2(n5985), .ZN(n5976)
         );
  AOI22_X1 U6975 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n5988), .B1(n6043), 
        .B2(n5987), .ZN(n5975) );
  OAI211_X1 U6976 ( .C1(n6046), .C2(n6020), .A(n5976), .B(n5975), .ZN(U3118)
         );
  AOI22_X1 U6977 ( .A1(n6100), .A2(n5986), .B1(n6099), .B2(n5985), .ZN(n5978)
         );
  AOI22_X1 U6978 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n5988), .B1(n6047), 
        .B2(n5987), .ZN(n5977) );
  OAI211_X1 U6979 ( .C1(n6050), .C2(n6020), .A(n5978), .B(n5977), .ZN(U3119)
         );
  AOI22_X1 U6980 ( .A1(n6106), .A2(n5986), .B1(n6105), .B2(n5985), .ZN(n5980)
         );
  AOI22_X1 U6981 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5988), .B1(n6051), 
        .B2(n5987), .ZN(n5979) );
  OAI211_X1 U6982 ( .C1(n6054), .C2(n6020), .A(n5980), .B(n5979), .ZN(U3120)
         );
  AOI22_X1 U6983 ( .A1(n6112), .A2(n5986), .B1(n6111), .B2(n5985), .ZN(n5982)
         );
  AOI22_X1 U6984 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n5988), .B1(n6055), 
        .B2(n5987), .ZN(n5981) );
  OAI211_X1 U6985 ( .C1(n6058), .C2(n6020), .A(n5982), .B(n5981), .ZN(U3121)
         );
  AOI22_X1 U6986 ( .A1(n6118), .A2(n5986), .B1(n6117), .B2(n5985), .ZN(n5984)
         );
  AOI22_X1 U6987 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n5988), .B1(n6059), 
        .B2(n5987), .ZN(n5983) );
  OAI211_X1 U6988 ( .C1(n6062), .C2(n6020), .A(n5984), .B(n5983), .ZN(U3122)
         );
  AOI22_X1 U6989 ( .A1(n6126), .A2(n5986), .B1(n6124), .B2(n5985), .ZN(n5990)
         );
  AOI22_X1 U6990 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n5988), .B1(n6066), 
        .B2(n5987), .ZN(n5989) );
  OAI211_X1 U6991 ( .C1(n6070), .C2(n6020), .A(n5990), .B(n5989), .ZN(U3123)
         );
  NOR2_X1 U6992 ( .A1(n6293), .A2(n5991), .ZN(n6016) );
  AOI21_X1 U6993 ( .B1(n6073), .B2(n5992), .A(n6016), .ZN(n5996) );
  NAND2_X1 U6994 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5994) );
  OAI22_X1 U6995 ( .A1(n5996), .A2(n6275), .B1(n5994), .B2(n5993), .ZN(n6015)
         );
  AOI22_X1 U6996 ( .A1(n6075), .A2(n6016), .B1(n6074), .B2(n6015), .ZN(n6001)
         );
  NAND2_X1 U6997 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  OAI221_X1 U6998 ( .B1(n6289), .B2(n5998), .C1(n6275), .C2(n5997), .A(n6082), 
        .ZN(n6017) );
  AOI22_X1 U6999 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6017), .B1(n6083), 
        .B2(n6065), .ZN(n6000) );
  OAI211_X1 U7000 ( .C1(n6086), .C2(n6020), .A(n6001), .B(n6000), .ZN(U3124)
         );
  AOI22_X1 U7001 ( .A1(n6088), .A2(n6016), .B1(n6087), .B2(n6015), .ZN(n6003)
         );
  INV_X1 U7002 ( .A(n6020), .ZN(n6006) );
  AOI22_X1 U7003 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6017), .B1(n6039), 
        .B2(n6006), .ZN(n6002) );
  OAI211_X1 U7004 ( .C1(n6042), .C2(n6027), .A(n6003), .B(n6002), .ZN(U3125)
         );
  AOI22_X1 U7005 ( .A1(n6094), .A2(n6016), .B1(n6093), .B2(n6015), .ZN(n6005)
         );
  AOI22_X1 U7006 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6017), .B1(n6043), 
        .B2(n6006), .ZN(n6004) );
  OAI211_X1 U7007 ( .C1(n6046), .C2(n6027), .A(n6005), .B(n6004), .ZN(U3126)
         );
  AOI22_X1 U7008 ( .A1(n6100), .A2(n6016), .B1(n6099), .B2(n6015), .ZN(n6008)
         );
  AOI22_X1 U7009 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6017), .B1(n6047), 
        .B2(n6006), .ZN(n6007) );
  OAI211_X1 U7010 ( .C1(n6050), .C2(n6027), .A(n6008), .B(n6007), .ZN(U3127)
         );
  AOI22_X1 U7011 ( .A1(n6106), .A2(n6016), .B1(n6105), .B2(n6015), .ZN(n6010)
         );
  AOI22_X1 U7012 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6017), .B1(n6107), 
        .B2(n6065), .ZN(n6009) );
  OAI211_X1 U7013 ( .C1(n6110), .C2(n6020), .A(n6010), .B(n6009), .ZN(U3128)
         );
  AOI22_X1 U7014 ( .A1(n6112), .A2(n6016), .B1(n6111), .B2(n6015), .ZN(n6012)
         );
  AOI22_X1 U7015 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6017), .B1(n6113), 
        .B2(n6065), .ZN(n6011) );
  OAI211_X1 U7016 ( .C1(n6116), .C2(n6020), .A(n6012), .B(n6011), .ZN(U3129)
         );
  AOI22_X1 U7017 ( .A1(n6118), .A2(n6016), .B1(n6117), .B2(n6015), .ZN(n6014)
         );
  AOI22_X1 U7018 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6017), .B1(n6119), 
        .B2(n6065), .ZN(n6013) );
  OAI211_X1 U7019 ( .C1(n6122), .C2(n6020), .A(n6014), .B(n6013), .ZN(U3130)
         );
  AOI22_X1 U7020 ( .A1(n6126), .A2(n6016), .B1(n6124), .B2(n6015), .ZN(n6019)
         );
  AOI22_X1 U7021 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6017), .B1(n6128), 
        .B2(n6065), .ZN(n6018) );
  OAI211_X1 U7022 ( .C1(n6133), .C2(n6020), .A(n6019), .B(n6018), .ZN(U3131)
         );
  INV_X1 U7023 ( .A(n6021), .ZN(n6077) );
  NOR2_X1 U7024 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6078), .ZN(n6064)
         );
  NAND3_X1 U7025 ( .A1(n6023), .A2(n6022), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7026 ( .B1(n6025), .B2(n6279), .A(n6024), .ZN(n6063) );
  AOI22_X1 U7027 ( .A1(n6075), .A2(n6064), .B1(n6074), .B2(n6063), .ZN(n6037)
         );
  AOI21_X1 U7028 ( .B1(n6132), .B2(n6027), .A(n6026), .ZN(n6028) );
  AOI211_X1 U7029 ( .C1(n6072), .C2(n6029), .A(n6275), .B(n6028), .ZN(n6031)
         );
  NOR2_X1 U7030 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  OAI211_X1 U7031 ( .C1(n6064), .C2(n6034), .A(n6033), .B(n6032), .ZN(n6067)
         );
  AOI22_X1 U7032 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6067), .B1(n6035), 
        .B2(n6065), .ZN(n6036) );
  OAI211_X1 U7033 ( .C1(n6038), .C2(n6132), .A(n6037), .B(n6036), .ZN(U3132)
         );
  AOI22_X1 U7034 ( .A1(n6088), .A2(n6064), .B1(n6087), .B2(n6063), .ZN(n6041)
         );
  AOI22_X1 U7035 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6067), .B1(n6039), 
        .B2(n6065), .ZN(n6040) );
  OAI211_X1 U7036 ( .C1(n6042), .C2(n6132), .A(n6041), .B(n6040), .ZN(U3133)
         );
  AOI22_X1 U7037 ( .A1(n6094), .A2(n6064), .B1(n6093), .B2(n6063), .ZN(n6045)
         );
  AOI22_X1 U7038 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6067), .B1(n6043), 
        .B2(n6065), .ZN(n6044) );
  OAI211_X1 U7039 ( .C1(n6046), .C2(n6132), .A(n6045), .B(n6044), .ZN(U3134)
         );
  AOI22_X1 U7040 ( .A1(n6100), .A2(n6064), .B1(n6099), .B2(n6063), .ZN(n6049)
         );
  AOI22_X1 U7041 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6067), .B1(n6047), 
        .B2(n6065), .ZN(n6048) );
  OAI211_X1 U7042 ( .C1(n6050), .C2(n6132), .A(n6049), .B(n6048), .ZN(U3135)
         );
  AOI22_X1 U7043 ( .A1(n6106), .A2(n6064), .B1(n6105), .B2(n6063), .ZN(n6053)
         );
  AOI22_X1 U7044 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6067), .B1(n6051), 
        .B2(n6065), .ZN(n6052) );
  OAI211_X1 U7045 ( .C1(n6054), .C2(n6132), .A(n6053), .B(n6052), .ZN(U3136)
         );
  AOI22_X1 U7046 ( .A1(n6112), .A2(n6064), .B1(n6111), .B2(n6063), .ZN(n6057)
         );
  AOI22_X1 U7047 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6067), .B1(n6055), 
        .B2(n6065), .ZN(n6056) );
  OAI211_X1 U7048 ( .C1(n6058), .C2(n6132), .A(n6057), .B(n6056), .ZN(U3137)
         );
  AOI22_X1 U7049 ( .A1(n6118), .A2(n6064), .B1(n6117), .B2(n6063), .ZN(n6061)
         );
  AOI22_X1 U7050 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6067), .B1(n6059), 
        .B2(n6065), .ZN(n6060) );
  OAI211_X1 U7051 ( .C1(n6062), .C2(n6132), .A(n6061), .B(n6060), .ZN(U3138)
         );
  AOI22_X1 U7052 ( .A1(n6126), .A2(n6064), .B1(n6124), .B2(n6063), .ZN(n6069)
         );
  AOI22_X1 U7053 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6067), .B1(n6066), 
        .B2(n6065), .ZN(n6068) );
  OAI211_X1 U7054 ( .C1(n6070), .C2(n6132), .A(n6069), .B(n6068), .ZN(U3139)
         );
  INV_X1 U7055 ( .A(n6071), .ZN(n6125) );
  AOI21_X1 U7056 ( .B1(n6073), .B2(n6072), .A(n6125), .ZN(n6080) );
  OAI22_X1 U7057 ( .A1(n6080), .A2(n6275), .B1(n5766), .B2(n6078), .ZN(n6123)
         );
  AOI22_X1 U7058 ( .A1(n6075), .A2(n6125), .B1(n6074), .B2(n6123), .ZN(n6085)
         );
  OAI21_X1 U7059 ( .B1(n6077), .B2(n6076), .A(n6280), .ZN(n6079) );
  AOI22_X1 U7060 ( .A1(n6080), .A2(n6079), .B1(n6275), .B2(n6078), .ZN(n6081)
         );
  NAND2_X1 U7061 ( .A1(n6082), .A2(n6081), .ZN(n6129) );
  AOI22_X1 U7062 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6129), .B1(n6083), 
        .B2(n6127), .ZN(n6084) );
  OAI211_X1 U7063 ( .C1(n6086), .C2(n6132), .A(n6085), .B(n6084), .ZN(U3140)
         );
  AOI22_X1 U7064 ( .A1(n6088), .A2(n6125), .B1(n6087), .B2(n6123), .ZN(n6091)
         );
  AOI22_X1 U7065 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6129), .B1(n6089), 
        .B2(n6127), .ZN(n6090) );
  OAI211_X1 U7066 ( .C1(n6092), .C2(n6132), .A(n6091), .B(n6090), .ZN(U3141)
         );
  AOI22_X1 U7067 ( .A1(n6094), .A2(n6125), .B1(n6093), .B2(n6123), .ZN(n6097)
         );
  AOI22_X1 U7068 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6129), .B1(n6095), 
        .B2(n6127), .ZN(n6096) );
  OAI211_X1 U7069 ( .C1(n6098), .C2(n6132), .A(n6097), .B(n6096), .ZN(U3142)
         );
  AOI22_X1 U7070 ( .A1(n6100), .A2(n6125), .B1(n6099), .B2(n6123), .ZN(n6103)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6129), .B1(n6101), 
        .B2(n6127), .ZN(n6102) );
  OAI211_X1 U7072 ( .C1(n6104), .C2(n6132), .A(n6103), .B(n6102), .ZN(U3143)
         );
  AOI22_X1 U7073 ( .A1(n6106), .A2(n6125), .B1(n6105), .B2(n6123), .ZN(n6109)
         );
  AOI22_X1 U7074 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6129), .B1(n6107), 
        .B2(n6127), .ZN(n6108) );
  OAI211_X1 U7075 ( .C1(n6110), .C2(n6132), .A(n6109), .B(n6108), .ZN(U3144)
         );
  AOI22_X1 U7076 ( .A1(n6112), .A2(n6125), .B1(n6111), .B2(n6123), .ZN(n6115)
         );
  AOI22_X1 U7077 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6129), .B1(n6113), 
        .B2(n6127), .ZN(n6114) );
  OAI211_X1 U7078 ( .C1(n6116), .C2(n6132), .A(n6115), .B(n6114), .ZN(U3145)
         );
  AOI22_X1 U7079 ( .A1(n6118), .A2(n6125), .B1(n6117), .B2(n6123), .ZN(n6121)
         );
  AOI22_X1 U7080 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6129), .B1(n6119), 
        .B2(n6127), .ZN(n6120) );
  OAI211_X1 U7081 ( .C1(n6122), .C2(n6132), .A(n6121), .B(n6120), .ZN(U3146)
         );
  AOI22_X1 U7082 ( .A1(n6126), .A2(n6125), .B1(n6124), .B2(n6123), .ZN(n6131)
         );
  AOI22_X1 U7083 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6129), .B1(n6128), 
        .B2(n6127), .ZN(n6130) );
  OAI211_X1 U7084 ( .C1(n6133), .C2(n6132), .A(n6131), .B(n6130), .ZN(U3147)
         );
  AOI22_X1 U7085 ( .A1(n6288), .A2(n6135), .B1(n6134), .B2(n3312), .ZN(n6268)
         );
  NAND2_X1 U7086 ( .A1(n6136), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6274) );
  NAND3_X1 U7087 ( .A1(n6268), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6274), .ZN(n6139) );
  OAI211_X1 U7088 ( .C1(n6140), .C2(n6139), .A(n6138), .B(n6137), .ZN(n6142)
         );
  NAND2_X1 U7089 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  NAND2_X1 U7090 ( .A1(n6142), .A2(n6141), .ZN(n6144) );
  AOI21_X1 U7091 ( .B1(n6144), .B2(n6145), .A(n6143), .ZN(n6148) );
  NOR2_X1 U7092 ( .A1(n6145), .A2(n6144), .ZN(n6147) );
  INV_X1 U7093 ( .A(n6146), .ZN(n6149) );
  OAI22_X1 U7094 ( .A1(n6148), .A2(n6147), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6149), .ZN(n6166) );
  AOI21_X1 U7095 ( .B1(n6149), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6165) );
  INV_X1 U7096 ( .A(n6150), .ZN(n6152) );
  NOR3_X1 U7097 ( .A1(n6152), .A2(n6151), .A3(n3828), .ZN(n6155) );
  INV_X1 U7098 ( .A(n6153), .ZN(n6154) );
  OAI22_X1 U7099 ( .A1(n6155), .A2(n6157), .B1(n4033), .B2(n6154), .ZN(n6156)
         );
  AOI21_X1 U7100 ( .B1(n6158), .B2(n6157), .A(n6156), .ZN(n6304) );
  OAI21_X1 U7101 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6159), 
        .ZN(n6160) );
  NAND4_X1 U7102 ( .A1(n6304), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n6163)
         );
  AOI211_X1 U7103 ( .C1(n6166), .C2(n6165), .A(n6164), .B(n6163), .ZN(n6179)
         );
  INV_X1 U7104 ( .A(n6167), .ZN(n6286) );
  NOR2_X1 U7105 ( .A1(n6198), .A2(n6168), .ZN(n6173) );
  INV_X1 U7106 ( .A(n6169), .ZN(n6172) );
  AOI22_X1 U7107 ( .A1(n6179), .A2(n6181), .B1(READY_N), .B2(n6170), .ZN(n6171) );
  AOI21_X1 U7108 ( .B1(n6173), .B2(n6172), .A(n6171), .ZN(n6266) );
  AOI211_X1 U7109 ( .C1(n6174), .C2(n6310), .A(STATE2_REG_0__SCAN_IN), .B(
        n6266), .ZN(n6175) );
  AOI211_X1 U7110 ( .C1(n6286), .C2(n6264), .A(n6176), .B(n6175), .ZN(n6177)
         );
  OAI221_X1 U7111 ( .B1(n6266), .B2(READY_N), .C1(n6266), .C2(n5766), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7112 ( .C1(n6179), .C2(n6178), .A(n6177), .B(n6187), .ZN(U3148)
         );
  NOR2_X1 U7113 ( .A1(READY_N), .A2(n6180), .ZN(n6190) );
  AOI21_X1 U7114 ( .B1(n6182), .B2(n6190), .A(n6181), .ZN(n6183) );
  NOR2_X1 U7115 ( .A1(n6183), .A2(n6266), .ZN(n6184) );
  AOI211_X1 U7116 ( .C1(n6266), .C2(n6285), .A(n6185), .B(n6184), .ZN(n6186)
         );
  OAI21_X1 U7117 ( .B1(n6395), .B2(n6187), .A(n6186), .ZN(U3149) );
  OAI211_X1 U7118 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6190), .A(n6189), .B(
        n6188), .ZN(n6191) );
  NAND2_X1 U7119 ( .A1(n6192), .A2(n6191), .ZN(U3150) );
  AND2_X1 U7120 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6261), .ZN(U3151) );
  AND2_X1 U7121 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6261), .ZN(U3152) );
  AND2_X1 U7122 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6261), .ZN(U3153) );
  AND2_X1 U7123 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6261), .ZN(U3154) );
  AND2_X1 U7124 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6261), .ZN(U3155) );
  AND2_X1 U7125 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6261), .ZN(U3156) );
  AND2_X1 U7126 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6261), .ZN(U3157) );
  AND2_X1 U7127 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6261), .ZN(U3158) );
  AND2_X1 U7128 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6261), .ZN(U3159) );
  AND2_X1 U7129 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6261), .ZN(U3160) );
  AND2_X1 U7130 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6261), .ZN(U3161) );
  AND2_X1 U7131 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6261), .ZN(U3162) );
  AND2_X1 U7132 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6261), .ZN(U3163) );
  AND2_X1 U7133 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6261), .ZN(U3164) );
  AND2_X1 U7134 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6261), .ZN(U3165) );
  AND2_X1 U7135 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6261), .ZN(U3166) );
  AND2_X1 U7136 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6261), .ZN(U3167) );
  AND2_X1 U7137 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6261), .ZN(U3168) );
  AND2_X1 U7138 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6261), .ZN(U3169) );
  NOR2_X1 U7139 ( .A1(n6263), .A2(n6353), .ZN(U3170) );
  AND2_X1 U7140 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6261), .ZN(U3171) );
  AND2_X1 U7141 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6261), .ZN(U3172) );
  AND2_X1 U7142 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6261), .ZN(U3173) );
  AND2_X1 U7143 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6261), .ZN(U3174) );
  AND2_X1 U7144 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6261), .ZN(U3175) );
  AND2_X1 U7145 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6261), .ZN(U3176) );
  AND2_X1 U7146 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6261), .ZN(U3177) );
  AND2_X1 U7147 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6261), .ZN(U3178) );
  NOR2_X1 U7148 ( .A1(n6263), .A2(n6363), .ZN(U3179) );
  AND2_X1 U7149 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6261), .ZN(U3180) );
  AOI22_X1 U7150 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6206) );
  INV_X1 U7151 ( .A(HOLD), .ZN(n6450) );
  NOR2_X1 U7152 ( .A1(n6199), .A2(n6450), .ZN(n6196) );
  INV_X1 U7153 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6194) );
  INV_X1 U7154 ( .A(NA_N), .ZN(n6203) );
  AOI211_X1 U7155 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6203), .A(
        STATE_REG_0__SCAN_IN), .B(n6202), .ZN(n6208) );
  AOI221_X1 U7156 ( .B1(n6196), .B2(n6259), .C1(n6194), .C2(n6259), .A(n6208), 
        .ZN(n6193) );
  OAI21_X1 U7157 ( .B1(n6202), .B2(n6206), .A(n6193), .ZN(U3181) );
  NOR2_X1 U7158 ( .A1(n6200), .A2(n6194), .ZN(n6204) );
  NAND2_X1 U7159 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6195) );
  OAI21_X1 U7160 ( .B1(n6204), .B2(n6196), .A(n6195), .ZN(n6197) );
  OAI211_X1 U7161 ( .C1(n6199), .C2(n4384), .A(n6198), .B(n6197), .ZN(U3182)
         );
  AOI221_X1 U7162 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4384), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6201) );
  AOI221_X1 U7163 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6201), .C2(HOLD), .A(n6200), .ZN(n6207) );
  AOI21_X1 U7164 ( .B1(n6204), .B2(n6203), .A(n6202), .ZN(n6205) );
  OAI22_X1 U7165 ( .A1(n6208), .A2(n6207), .B1(n6206), .B2(n6205), .ZN(U3183)
         );
  NAND2_X1 U7166 ( .A1(n6315), .A2(n6209), .ZN(n6257) );
  NOR2_X2 U7167 ( .A1(n6209), .A2(n6259), .ZN(n6255) );
  AOI22_X1 U7168 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6259), .ZN(n6210) );
  OAI21_X1 U7169 ( .B1(n6423), .B2(n6257), .A(n6210), .ZN(U3184) );
  AOI22_X1 U7170 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6259), .ZN(n6211) );
  OAI21_X1 U7171 ( .B1(n6212), .B2(n6257), .A(n6211), .ZN(U3185) );
  AOI22_X1 U7172 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6259), .ZN(n6213) );
  OAI21_X1 U7173 ( .B1(n6451), .B2(n6257), .A(n6213), .ZN(U3186) );
  AOI22_X1 U7174 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6259), .ZN(n6214) );
  OAI21_X1 U7175 ( .B1(n6215), .B2(n6257), .A(n6214), .ZN(U3187) );
  AOI22_X1 U7176 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6259), .ZN(n6216) );
  OAI21_X1 U7177 ( .B1(n6217), .B2(n6257), .A(n6216), .ZN(U3188) );
  AOI22_X1 U7178 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6259), .ZN(n6218) );
  OAI21_X1 U7179 ( .B1(n6220), .B2(n6257), .A(n6218), .ZN(U3189) );
  INV_X1 U7180 ( .A(n6257), .ZN(n6251) );
  AOI22_X1 U7181 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6259), .ZN(n6219) );
  OAI21_X1 U7182 ( .B1(n6220), .B2(n6253), .A(n6219), .ZN(U3190) );
  INV_X1 U7183 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6380) );
  OAI222_X1 U7184 ( .A1(n6253), .A2(n4576), .B1(n6380), .B2(n6315), .C1(n6221), 
        .C2(n6257), .ZN(U3191) );
  AOI22_X1 U7185 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6259), .ZN(n6222) );
  OAI21_X1 U7186 ( .B1(n6452), .B2(n6257), .A(n6222), .ZN(U3192) );
  AOI22_X1 U7187 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6259), .ZN(n6223) );
  OAI21_X1 U7188 ( .B1(n6452), .B2(n6253), .A(n6223), .ZN(U3193) );
  AOI22_X1 U7189 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6259), .ZN(n6224) );
  OAI21_X1 U7190 ( .B1(n6225), .B2(n6253), .A(n6224), .ZN(U3194) );
  AOI22_X1 U7191 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6259), .ZN(n6226) );
  OAI21_X1 U7192 ( .B1(n6228), .B2(n6257), .A(n6226), .ZN(U3195) );
  AOI22_X1 U7193 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6259), .ZN(n6227) );
  OAI21_X1 U7194 ( .B1(n6228), .B2(n6253), .A(n6227), .ZN(U3196) );
  AOI22_X1 U7195 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6259), .ZN(n6229) );
  OAI21_X1 U7196 ( .B1(n6397), .B2(n6257), .A(n6229), .ZN(U3197) );
  INV_X1 U7197 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6401) );
  OAI222_X1 U7198 ( .A1(n6257), .A2(n6230), .B1(n6401), .B2(n6315), .C1(n6397), 
        .C2(n6253), .ZN(U3198) );
  AOI22_X1 U7199 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6259), .ZN(n6231) );
  OAI21_X1 U7200 ( .B1(n6233), .B2(n6257), .A(n6231), .ZN(U3199) );
  AOI22_X1 U7201 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6259), .ZN(n6232) );
  OAI21_X1 U7202 ( .B1(n6233), .B2(n6253), .A(n6232), .ZN(U3200) );
  AOI22_X1 U7203 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6259), .ZN(n6234) );
  OAI21_X1 U7204 ( .B1(n6235), .B2(n6253), .A(n6234), .ZN(U3201) );
  AOI22_X1 U7205 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6259), .ZN(n6236) );
  OAI21_X1 U7206 ( .B1(n6237), .B2(n6253), .A(n6236), .ZN(U3202) );
  AOI22_X1 U7207 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6259), .ZN(n6238) );
  OAI21_X1 U7208 ( .B1(n6239), .B2(n6257), .A(n6238), .ZN(U3203) );
  INV_X1 U7209 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6351) );
  INV_X1 U7210 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6241) );
  OAI222_X1 U7211 ( .A1(n6253), .A2(n6239), .B1(n6351), .B2(n6315), .C1(n6241), 
        .C2(n6257), .ZN(U3204) );
  AOI22_X1 U7212 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6259), .ZN(n6240) );
  OAI21_X1 U7213 ( .B1(n6241), .B2(n6253), .A(n6240), .ZN(U3205) );
  AOI22_X1 U7214 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6259), .ZN(n6242) );
  OAI21_X1 U7215 ( .B1(n6243), .B2(n6253), .A(n6242), .ZN(U3206) );
  AOI22_X1 U7216 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6259), .ZN(n6244) );
  OAI21_X1 U7217 ( .B1(n6246), .B2(n6257), .A(n6244), .ZN(U3207) );
  AOI22_X1 U7218 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6259), .ZN(n6245) );
  OAI21_X1 U7219 ( .B1(n6246), .B2(n6253), .A(n6245), .ZN(U3208) );
  AOI22_X1 U7220 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6259), .ZN(n6247) );
  OAI21_X1 U7221 ( .B1(n6249), .B2(n6257), .A(n6247), .ZN(U3209) );
  AOI22_X1 U7222 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6259), .ZN(n6248) );
  OAI21_X1 U7223 ( .B1(n6249), .B2(n6253), .A(n6248), .ZN(U3210) );
  AOI22_X1 U7224 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6259), .ZN(n6250) );
  OAI21_X1 U7225 ( .B1(n6254), .B2(n6257), .A(n6250), .ZN(U3211) );
  AOI22_X1 U7226 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6251), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6259), .ZN(n6252) );
  OAI21_X1 U7227 ( .B1(n6254), .B2(n6253), .A(n6252), .ZN(U3212) );
  AOI22_X1 U7228 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6255), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6259), .ZN(n6256) );
  OAI21_X1 U7229 ( .B1(n6258), .B2(n6257), .A(n6256), .ZN(U3213) );
  MUX2_X1 U7230 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6315), .Z(U3445) );
  MUX2_X1 U7231 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6315), .Z(U3446) );
  MUX2_X1 U7232 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6315), .Z(U3447) );
  INV_X1 U7233 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6299) );
  INV_X1 U7234 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6361) );
  AOI22_X1 U7235 ( .A1(n6315), .A2(n6299), .B1(n6361), .B2(n6259), .ZN(U3448)
         );
  INV_X1 U7236 ( .A(n6262), .ZN(n6260) );
  AOI21_X1 U7237 ( .B1(n6295), .B2(n6261), .A(n6260), .ZN(U3451) );
  OAI21_X1 U7238 ( .B1(n6263), .B2(n6383), .A(n6262), .ZN(U3452) );
  AOI211_X1 U7239 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6266), .A(n6265), .B(
        n6264), .ZN(n6267) );
  INV_X1 U7240 ( .A(n6267), .ZN(U3453) );
  OAI22_X1 U7241 ( .A1(n6268), .A2(n6273), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6395), .ZN(n6271) );
  OAI22_X1 U7242 ( .A1(n6271), .A2(n6270), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6269), .ZN(n6272) );
  OAI21_X1 U7243 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(U3461) );
  AOI21_X1 U7244 ( .B1(n6277), .B2(n6276), .A(n6275), .ZN(n6282) );
  OAI22_X1 U7245 ( .A1(n3933), .A2(n6280), .B1(n6279), .B2(n6278), .ZN(n6281)
         );
  NOR2_X1 U7246 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  AOI22_X1 U7247 ( .A1(n6294), .A2(n6284), .B1(n6283), .B2(n6291), .ZN(U3462)
         );
  AOI222_X1 U7248 ( .A1(n6290), .A2(n6289), .B1(n6288), .B2(n6287), .C1(n6286), 
        .C2(n6285), .ZN(n6292) );
  AOI22_X1 U7249 ( .A1(n6294), .A2(n6293), .B1(n6292), .B2(n6291), .ZN(U3465)
         );
  OAI211_X1 U7250 ( .C1(n6295), .C2(n6335), .A(n6383), .B(n6301), .ZN(n6298)
         );
  NOR2_X1 U7251 ( .A1(n6300), .A2(n6335), .ZN(n6296) );
  AOI22_X1 U7252 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6300), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6296), .ZN(n6297) );
  NAND2_X1 U7253 ( .A1(n6298), .A2(n6297), .ZN(U3468) );
  AOI22_X1 U7254 ( .A1(n6301), .A2(n6335), .B1(n6300), .B2(n6299), .ZN(U3469)
         );
  INV_X1 U7255 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6338) );
  MUX2_X1 U7256 ( .A(W_R_N_REG_SCAN_IN), .B(n6338), .S(n6315), .Z(U3470) );
  INV_X1 U7257 ( .A(MORE_REG_SCAN_IN), .ZN(n6303) );
  INV_X1 U7258 ( .A(n6305), .ZN(n6302) );
  AOI22_X1 U7259 ( .A1(n6305), .A2(n6304), .B1(n6303), .B2(n6302), .ZN(U3471)
         );
  AOI211_X1 U7260 ( .C1(n6307), .C2(n4384), .A(n6306), .B(n6319), .ZN(n6314)
         );
  OAI211_X1 U7261 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6309), .A(n6308), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6311) );
  AOI21_X1 U7262 ( .B1(n6311), .B2(STATE2_REG_0__SCAN_IN), .A(n6310), .ZN(
        n6313) );
  NAND2_X1 U7263 ( .A1(n6314), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6312) );
  OAI21_X1 U7264 ( .B1(n6314), .B2(n6313), .A(n6312), .ZN(U3472) );
  MUX2_X1 U7265 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6315), .Z(U3473) );
  INV_X1 U7266 ( .A(n6316), .ZN(n6317) );
  NOR2_X1 U7267 ( .A1(n6319), .A2(n6317), .ZN(n6318) );
  AOI22_X1 U7268 ( .A1(n6320), .A2(n6319), .B1(n6338), .B2(n6318), .ZN(U3474)
         );
  INV_X1 U7269 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6322) );
  AOI22_X1 U7270 ( .A1(n6322), .A2(keyinput40), .B1(keyinput6), .B2(n6452), 
        .ZN(n6321) );
  OAI221_X1 U7271 ( .B1(n6322), .B2(keyinput40), .C1(n6452), .C2(keyinput6), 
        .A(n6321), .ZN(n6331) );
  AOI22_X1 U7272 ( .A1(n6453), .A2(keyinput49), .B1(keyinput21), .B2(n5105), 
        .ZN(n6323) );
  OAI221_X1 U7273 ( .B1(n6453), .B2(keyinput49), .C1(n5105), .C2(keyinput21), 
        .A(n6323), .ZN(n6330) );
  INV_X1 U7274 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6325) );
  AOI22_X1 U7275 ( .A1(n6325), .A2(keyinput61), .B1(keyinput42), .B2(n4011), 
        .ZN(n6324) );
  OAI221_X1 U7276 ( .B1(n6325), .B2(keyinput61), .C1(n4011), .C2(keyinput42), 
        .A(n6324), .ZN(n6329) );
  INV_X1 U7277 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6327) );
  AOI22_X1 U7278 ( .A1(n6455), .A2(keyinput25), .B1(n6327), .B2(keyinput10), 
        .ZN(n6326) );
  OAI221_X1 U7279 ( .B1(n6455), .B2(keyinput25), .C1(n6327), .C2(keyinput10), 
        .A(n6326), .ZN(n6328) );
  NOR4_X1 U7280 ( .A1(n6331), .A2(n6330), .A3(n6329), .A4(n6328), .ZN(n6376)
         );
  AOI22_X1 U7281 ( .A1(n6450), .A2(keyinput14), .B1(n6333), .B2(keyinput1), 
        .ZN(n6332) );
  OAI221_X1 U7282 ( .B1(n6450), .B2(keyinput14), .C1(n6333), .C2(keyinput1), 
        .A(n6332), .ZN(n6343) );
  AOI22_X1 U7283 ( .A1(n6335), .A2(keyinput11), .B1(n6460), .B2(keyinput50), 
        .ZN(n6334) );
  OAI221_X1 U7284 ( .B1(n6335), .B2(keyinput11), .C1(n6460), .C2(keyinput50), 
        .A(n6334), .ZN(n6342) );
  AOI22_X1 U7285 ( .A1(n6451), .A2(keyinput53), .B1(n6454), .B2(keyinput54), 
        .ZN(n6336) );
  OAI221_X1 U7286 ( .B1(n6451), .B2(keyinput53), .C1(n6454), .C2(keyinput54), 
        .A(n6336), .ZN(n6341) );
  NOR4_X1 U7287 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n6375)
         );
  INV_X1 U7288 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6345) );
  AOI22_X1 U7289 ( .A1(n6461), .A2(keyinput17), .B1(n6345), .B2(keyinput29), 
        .ZN(n6344) );
  OAI221_X1 U7290 ( .B1(n6461), .B2(keyinput17), .C1(n6345), .C2(keyinput29), 
        .A(n6344), .ZN(n6358) );
  INV_X1 U7291 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6347) );
  AOI22_X1 U7292 ( .A1(n6348), .A2(keyinput51), .B1(n6347), .B2(keyinput63), 
        .ZN(n6346) );
  OAI221_X1 U7293 ( .B1(n6348), .B2(keyinput51), .C1(n6347), .C2(keyinput63), 
        .A(n6346), .ZN(n6357) );
  AOI22_X1 U7294 ( .A1(n6351), .A2(keyinput44), .B1(keyinput59), .B2(n6350), 
        .ZN(n6349) );
  OAI221_X1 U7295 ( .B1(n6351), .B2(keyinput44), .C1(n6350), .C2(keyinput59), 
        .A(n6349), .ZN(n6356) );
  AOI22_X1 U7296 ( .A1(n6354), .A2(keyinput0), .B1(keyinput34), .B2(n6353), 
        .ZN(n6352) );
  OAI221_X1 U7297 ( .B1(n6354), .B2(keyinput0), .C1(n6353), .C2(keyinput34), 
        .A(n6352), .ZN(n6355) );
  NOR4_X1 U7298 ( .A1(n6358), .A2(n6357), .A3(n6356), .A4(n6355), .ZN(n6374)
         );
  INV_X1 U7299 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6360) );
  AOI22_X1 U7300 ( .A1(n6361), .A2(keyinput39), .B1(n6360), .B2(keyinput62), 
        .ZN(n6359) );
  OAI221_X1 U7301 ( .B1(n6361), .B2(keyinput39), .C1(n6360), .C2(keyinput62), 
        .A(n6359), .ZN(n6372) );
  AOI22_X1 U7302 ( .A1(n6364), .A2(keyinput56), .B1(keyinput28), .B2(n6363), 
        .ZN(n6362) );
  OAI221_X1 U7303 ( .B1(n6364), .B2(keyinput56), .C1(n6363), .C2(keyinput28), 
        .A(n6362), .ZN(n6371) );
  AOI22_X1 U7304 ( .A1(n6366), .A2(keyinput24), .B1(n6442), .B2(keyinput57), 
        .ZN(n6365) );
  OAI221_X1 U7305 ( .B1(n6366), .B2(keyinput24), .C1(n6442), .C2(keyinput57), 
        .A(n6365), .ZN(n6370) );
  INV_X1 U7306 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6368) );
  AOI22_X1 U7307 ( .A1(n6368), .A2(keyinput58), .B1(keyinput47), .B2(n6463), 
        .ZN(n6367) );
  OAI221_X1 U7308 ( .B1(n6368), .B2(keyinput58), .C1(n6463), .C2(keyinput47), 
        .A(n6367), .ZN(n6369) );
  NOR4_X1 U7309 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n6373)
         );
  NAND4_X1 U7310 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n6436)
         );
  AOI22_X1 U7311 ( .A1(n6446), .A2(keyinput16), .B1(keyinput5), .B2(n6378), 
        .ZN(n6377) );
  OAI221_X1 U7312 ( .B1(n6446), .B2(keyinput16), .C1(n6378), .C2(keyinput5), 
        .A(n6377), .ZN(n6390) );
  AOI22_X1 U7313 ( .A1(n6381), .A2(keyinput23), .B1(keyinput60), .B2(n6380), 
        .ZN(n6379) );
  OAI221_X1 U7314 ( .B1(n6381), .B2(keyinput23), .C1(n6380), .C2(keyinput60), 
        .A(n6379), .ZN(n6389) );
  AOI22_X1 U7315 ( .A1(n6384), .A2(keyinput55), .B1(n6383), .B2(keyinput37), 
        .ZN(n6382) );
  OAI221_X1 U7316 ( .B1(n6384), .B2(keyinput55), .C1(n6383), .C2(keyinput37), 
        .A(n6382), .ZN(n6388) );
  INV_X1 U7317 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U7318 ( .A1(n4397), .A2(keyinput41), .B1(n6386), .B2(keyinput26), 
        .ZN(n6385) );
  OAI221_X1 U7319 ( .B1(n4397), .B2(keyinput41), .C1(n6386), .C2(keyinput26), 
        .A(n6385), .ZN(n6387) );
  NOR4_X1 U7320 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n6434)
         );
  AOI22_X1 U7321 ( .A1(n6395), .A2(keyinput33), .B1(keyinput35), .B2(n6394), 
        .ZN(n6393) );
  OAI221_X1 U7322 ( .B1(n6395), .B2(keyinput33), .C1(n6394), .C2(keyinput35), 
        .A(n6393), .ZN(n6404) );
  AOI22_X1 U7323 ( .A1(n6398), .A2(keyinput30), .B1(keyinput22), .B2(n6397), 
        .ZN(n6396) );
  OAI221_X1 U7324 ( .B1(n6398), .B2(keyinput30), .C1(n6397), .C2(keyinput22), 
        .A(n6396), .ZN(n6403) );
  AOI22_X1 U7325 ( .A1(n6401), .A2(keyinput32), .B1(n6400), .B2(keyinput19), 
        .ZN(n6399) );
  OAI221_X1 U7326 ( .B1(n6401), .B2(keyinput32), .C1(n6400), .C2(keyinput19), 
        .A(n6399), .ZN(n6402) );
  NOR4_X1 U7327 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n6433)
         );
  INV_X1 U7328 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6407) );
  AOI22_X1 U7329 ( .A1(n6408), .A2(keyinput43), .B1(n6407), .B2(keyinput4), 
        .ZN(n6406) );
  OAI221_X1 U7330 ( .B1(n6408), .B2(keyinput43), .C1(n6407), .C2(keyinput4), 
        .A(n6406), .ZN(n6418) );
  INV_X1 U7331 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6444) );
  INV_X1 U7332 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6410) );
  AOI22_X1 U7333 ( .A1(n6444), .A2(keyinput46), .B1(n6410), .B2(keyinput13), 
        .ZN(n6409) );
  OAI221_X1 U7334 ( .B1(n6444), .B2(keyinput46), .C1(n6410), .C2(keyinput13), 
        .A(n6409), .ZN(n6417) );
  AOI22_X1 U7335 ( .A1(n6445), .A2(keyinput52), .B1(keyinput8), .B2(n6412), 
        .ZN(n6411) );
  OAI221_X1 U7336 ( .B1(n6445), .B2(keyinput52), .C1(n6412), .C2(keyinput8), 
        .A(n6411), .ZN(n6416) );
  INV_X1 U7337 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6414) );
  AOI22_X1 U7338 ( .A1(n6462), .A2(keyinput45), .B1(keyinput3), .B2(n6414), 
        .ZN(n6413) );
  OAI221_X1 U7339 ( .B1(n6462), .B2(keyinput45), .C1(n6414), .C2(keyinput3), 
        .A(n6413), .ZN(n6415) );
  NOR4_X1 U7340 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n6432)
         );
  AOI22_X1 U7341 ( .A1(n5401), .A2(keyinput27), .B1(keyinput15), .B2(n6420), 
        .ZN(n6419) );
  OAI221_X1 U7342 ( .B1(n5401), .B2(keyinput27), .C1(n6420), .C2(keyinput15), 
        .A(n6419), .ZN(n6430) );
  AOI22_X1 U7343 ( .A1(n4395), .A2(keyinput9), .B1(n3820), .B2(keyinput18), 
        .ZN(n6421) );
  OAI221_X1 U7344 ( .B1(n4395), .B2(keyinput9), .C1(n3820), .C2(keyinput18), 
        .A(n6421), .ZN(n6429) );
  INV_X1 U7345 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6424) );
  AOI22_X1 U7346 ( .A1(n6424), .A2(keyinput48), .B1(n6423), .B2(keyinput12), 
        .ZN(n6422) );
  OAI221_X1 U7347 ( .B1(n6424), .B2(keyinput48), .C1(n6423), .C2(keyinput12), 
        .A(n6422), .ZN(n6428) );
  INV_X1 U7348 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6443) );
  AOI22_X1 U7349 ( .A1(n6426), .A2(keyinput2), .B1(n6443), .B2(keyinput7), 
        .ZN(n6425) );
  OAI221_X1 U7350 ( .B1(n6426), .B2(keyinput2), .C1(n6443), .C2(keyinput7), 
        .A(n6425), .ZN(n6427) );
  NOR4_X1 U7351 ( .A1(n6430), .A2(n6429), .A3(n6428), .A4(n6427), .ZN(n6431)
         );
  NAND4_X1 U7352 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n6435)
         );
  NOR2_X1 U7353 ( .A1(n6436), .A2(n6435), .ZN(n6481) );
  AOI22_X1 U7354 ( .A1(n6438), .A2(LWORD_REG_4__SCAN_IN), .B1(n6437), .B2(
        DATAI_4_), .ZN(n6439) );
  OAI21_X1 U7355 ( .B1(n6441), .B2(n6440), .A(n6439), .ZN(n6479) );
  NAND4_X1 U7356 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(
        INSTQUEUE_REG_4__6__SCAN_IN), .A3(n6443), .A4(n6442), .ZN(n6477) );
  NOR3_X1 U7357 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(
        INSTQUEUE_REG_4__1__SCAN_IN), .A3(n6444), .ZN(n6449) );
  NOR4_X1 U7358 ( .A1(STATE2_REG_1__SCAN_IN), .A2(INSTQUEUE_REG_8__5__SCAN_IN), 
        .A3(INSTQUEUE_REG_10__5__SCAN_IN), .A4(n6445), .ZN(n6448) );
  NOR4_X1 U7359 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(
        INSTQUEUE_REG_5__6__SCAN_IN), .A3(INSTQUEUE_REG_13__6__SCAN_IN), .A4(
        n6446), .ZN(n6447) );
  NAND4_X1 U7360 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6449), .A3(n6448), 
        .A4(n6447), .ZN(n6476) );
  NOR4_X1 U7361 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        EBX_REG_15__SCAN_IN), .A3(PHYADDRPOINTER_REG_18__SCAN_IN), .A4(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6459) );
  NOR4_X1 U7362 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(EBX_REG_31__SCAN_IN), .A3(DATAI_8_), .A4(DATAI_21_), .ZN(n6458) );
  NOR4_X1 U7363 ( .A1(REIP_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n6451), .A4(n6450), .ZN(n6457) );
  NOR4_X1 U7364 ( .A1(n6455), .A2(n6454), .A3(n6453), .A4(n6452), .ZN(n6456)
         );
  NAND4_X1 U7365 ( .A1(n6459), .A2(n6458), .A3(n6457), .A4(n6456), .ZN(n6475)
         );
  NOR4_X1 U7366 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(
        ADDRESS_REG_20__SCAN_IN), .A3(ADDRESS_REG_7__SCAN_IN), .A4(
        READREQUEST_REG_SCAN_IN), .ZN(n6473) );
  NOR4_X1 U7367 ( .A1(REIP_REG_2__SCAN_IN), .A2(DATAI_16_), .A3(
        DATAO_REG_4__SCAN_IN), .A4(DATAO_REG_14__SCAN_IN), .ZN(n6472) );
  NAND4_X1 U7368 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n6464)
         );
  NOR4_X1 U7369 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6465), .A4(n6464), .ZN(n6471) );
  NAND4_X1 U7370 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .A3(EAX_REG_19__SCAN_IN), .A4(
        BE_N_REG_0__SCAN_IN), .ZN(n6469) );
  NAND4_X1 U7371 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        DATAO_REG_1__SCAN_IN), .A4(ADDRESS_REG_14__SCAN_IN), .ZN(n6468) );
  NAND4_X1 U7372 ( .A1(DATAI_6_), .A2(LWORD_REG_1__SCAN_IN), .A3(
        DATAO_REG_12__SCAN_IN), .A4(LWORD_REG_7__SCAN_IN), .ZN(n6467) );
  NAND4_X1 U7373 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        EAX_REG_30__SCAN_IN), .A3(DATAO_REG_28__SCAN_IN), .A4(
        BYTEENABLE_REG_3__SCAN_IN), .ZN(n6466) );
  NOR4_X1 U7374 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n6470)
         );
  NAND4_X1 U7375 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n6474)
         );
  NOR4_X1 U7376 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n6478)
         );
  XNOR2_X1 U7377 ( .A(n6479), .B(n6478), .ZN(n6480) );
  XNOR2_X1 U7378 ( .A(n6481), .B(n6480), .ZN(U2943) );
  CLKBUF_X2 U3524 ( .A(n3222), .Z(n3794) );
  AND2_X1 U3401 ( .A1(n3838), .A2(n3216), .ZN(n3211) );
  CLKBUF_X2 U3426 ( .A(n3082), .Z(n3203) );
  CLKBUF_X1 U3440 ( .A(n3185), .Z(n4046) );
  OR2_X1 U3554 ( .A1(n3094), .A2(n3093), .ZN(n3201) );
  CLKBUF_X2 U3851 ( .A(n4058), .Z(n4231) );
  OR2_X1 U4043 ( .A1(n2956), .A2(n2957), .ZN(n4823) );
endmodule

