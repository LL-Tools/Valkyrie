

module b22_C_gen_AntiSAT_k_128_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6469, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091;

  XNOR2_X1 U7217 ( .A(n8306), .B(n8305), .ZN(n13579) );
  AND2_X1 U7218 ( .A1(n8731), .A2(n8730), .ZN(n13532) );
  OAI21_X1 U7219 ( .B1(n8134), .B2(n6730), .A(n6727), .ZN(n7752) );
  AND2_X1 U7220 ( .A1(n12414), .A2(n12410), .ZN(n12565) );
  AND2_X1 U7222 ( .A1(n8402), .A2(n6511), .ZN(n10618) );
  INV_X1 U7223 ( .A(n9088), .ZN(n9089) );
  INV_X1 U7224 ( .A(n8518), .ZN(n8568) );
  AND4_X1 U7225 ( .A1(n7881), .A2(n7880), .A3(n7879), .A4(n7878), .ZN(n10732)
         );
  INV_X2 U7227 ( .A(n6485), .ZN(n8184) );
  CLKBUF_X1 U7228 ( .A(n8205), .Z(n6482) );
  NAND4_X2 U7231 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n13688)
         );
  NAND2_X1 U7232 ( .A1(n7855), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7832) );
  AND2_X1 U7233 ( .A1(n9896), .A2(n7798), .ZN(n7837) );
  AND2_X2 U7234 ( .A1(n14119), .A2(n7812), .ZN(n7855) );
  OAI21_X1 U7235 ( .B1(n8470), .B2(n8469), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8472) );
  INV_X1 U7236 ( .A(n8501), .ZN(n7798) );
  NOR2_X1 U7238 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7670) );
  INV_X1 U7239 ( .A(n12525), .ZN(n12514) );
  INV_X2 U7241 ( .A(n8375), .ZN(n8377) );
  AND3_X1 U7242 ( .A1(n7672), .A2(n7673), .A3(n7671), .ZN(n8427) );
  BUF_X1 U7243 ( .A(n8568), .Z(n6490) );
  NAND2_X1 U7245 ( .A1(n8485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8483) );
  AND2_X1 U7246 ( .A1(n9896), .A2(n8501), .ZN(n7862) );
  NAND3_X1 U7247 ( .A1(n7118), .A2(n7117), .A3(n7685), .ZN(n7801) );
  NAND2_X1 U7248 ( .A1(n6975), .A2(n15014), .ZN(n14995) );
  INV_X1 U7249 ( .A(n12538), .ZN(n9369) );
  CLKBUF_X3 U7250 ( .A(n9113), .Z(n9475) );
  INV_X1 U7251 ( .A(n9107), .ZN(n14992) );
  OR2_X1 U7252 ( .A1(n9131), .A2(n9098), .ZN(n9132) );
  NAND2_X2 U7254 ( .A1(n9770), .A2(n9727), .ZN(n8990) );
  AND2_X1 U7255 ( .A1(n7114), .A2(n7112), .ZN(n11693) );
  BUF_X2 U7256 ( .A(n7862), .Z(n8178) );
  INV_X1 U7257 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U7258 ( .A1(n9095), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9097) );
  INV_X1 U7259 ( .A(n8935), .ZN(n8580) );
  XNOR2_X1 U7260 ( .A(n8472), .B(n8471), .ZN(n11346) );
  AND4_X1 U7261 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n14357)
         );
  OR2_X1 U7262 ( .A1(n8205), .A2(n7829), .ZN(n7831) );
  OR2_X1 U7263 ( .A1(n7700), .A2(n9754), .ZN(n6469) );
  NOR2_X2 U7264 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9068) );
  NAND4_X2 U7265 ( .A1(n9068), .A2(n9067), .A3(n9275), .A4(n9343), .ZN(n9382)
         );
  AOI21_X2 U7266 ( .B1(n11780), .B2(n11779), .A(n6546), .ZN(n11781) );
  XNOR2_X2 U7267 ( .A(n7472), .B(n7471), .ZN(n14332) );
  OAI21_X1 U7268 ( .B1(n14036), .B2(n14095), .A(n14034), .ZN(n6618) );
  AOI21_X2 U7269 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n11714), .A(n11713), .ZN(
        n12613) );
  OAI21_X2 U7270 ( .B1(n7697), .B2(n6648), .A(n6647), .ZN(n7699) );
  NAND2_X2 U7271 ( .A1(n6792), .A2(n6793), .ZN(n7697) );
  NAND2_X2 U7272 ( .A1(n7697), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7273 ( .A1(n11331), .A2(n11272), .ZN(n11495) );
  NOR2_X2 U7274 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n9067) );
  NAND2_X2 U7275 ( .A1(n12010), .A2(n12009), .ZN(n13983) );
  OAI21_X2 U7277 ( .B1(n8260), .B2(n10917), .A(n7772), .ZN(n7774) );
  XNOR2_X1 U7278 ( .A(n7861), .B(n7867), .ZN(n9728) );
  AND2_X2 U7279 ( .A1(n9647), .A2(n9079), .ZN(n7383) );
  AND3_X2 U7280 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(n9647) );
  XNOR2_X2 U7281 ( .A(n8480), .B(n9039), .ZN(n8487) );
  NOR2_X2 U7282 ( .A1(n10996), .A2(n11052), .ZN(n11064) );
  NOR2_X2 U7283 ( .A1(n12004), .A2(n12006), .ZN(n13836) );
  NOR2_X2 U7284 ( .A1(n13877), .A2(n12003), .ZN(n12004) );
  XNOR2_X2 U7285 ( .A(n6941), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n7433) );
  INV_X2 U7286 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U7287 ( .A1(n10807), .A2(n14492), .ZN(n6473) );
  NAND2_X1 U7288 ( .A1(n10807), .A2(n14492), .ZN(n6474) );
  INV_X1 U7289 ( .A(n8972), .ZN(n6475) );
  INV_X4 U7290 ( .A(n6475), .ZN(n6476) );
  NAND2_X1 U7291 ( .A1(n8458), .A2(n8457), .ZN(n8972) );
  AND2_X2 U7292 ( .A1(n9131), .A2(n9074), .ZN(n9148) );
  NOR2_X4 U7293 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9131) );
  INV_X1 U7294 ( .A(n8332), .ZN(n6477) );
  XNOR2_X2 U7295 ( .A(n7708), .B(SI_4_), .ZN(n7896) );
  NOR2_X2 U7296 ( .A1(n14446), .A2(n14447), .ZN(n14451) );
  INV_X1 U7297 ( .A(n10794), .ZN(n14963) );
  XOR2_X2 U7298 ( .A(n7431), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15081) );
  XNOR2_X2 U7299 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n7430), .ZN(n7431) );
  OAI222_X1 U7300 ( .A1(P3_U3151), .A2(n9090), .B1(n13058), .B2(n12528), .C1(
        n13056), .C2(n12227), .ZN(P3_U3265) );
  AND2_X1 U7301 ( .A1(n8453), .A2(n8455), .ZN(n8935) );
  XNOR2_X2 U7302 ( .A(n7702), .B(SI_2_), .ZN(n7868) );
  INV_X2 U7303 ( .A(n8479), .ZN(n10181) );
  OAI211_X2 U7304 ( .C1(P2_IR_REG_21__SCAN_IN), .C2(P2_IR_REG_31__SCAN_IN), 
        .A(n8478), .B(n8477), .ZN(n8479) );
  NAND2_X2 U7305 ( .A1(n9118), .A2(n9107), .ZN(n12394) );
  AND4_X4 U7306 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n9118)
         );
  NAND2_X2 U7307 ( .A1(n13050), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9083) );
  CLKBUF_X1 U7308 ( .A(n9561), .Z(n6480) );
  CLKBUF_X2 U7309 ( .A(n9561), .Z(n6481) );
  NAND2_X1 U7310 ( .A1(n9103), .A2(n9733), .ZN(n9561) );
  OR2_X2 U7312 ( .A1(n7394), .A2(n6945), .ZN(n6944) );
  XNOR2_X2 U7313 ( .A(n8450), .B(n8449), .ZN(n8453) );
  XNOR2_X2 U7314 ( .A(n6936), .B(n9102), .ZN(n10028) );
  OR2_X2 U7315 ( .A1(n8435), .A2(n10256), .ZN(n10278) );
  INV_X4 U7316 ( .A(n12627), .ZN(n12729) );
  BUF_X4 U7317 ( .A(n7855), .Z(n6485) );
  XNOR2_X2 U7318 ( .A(n11748), .B(n13185), .ZN(n11742) );
  INV_X2 U7319 ( .A(n13523), .ZN(n11748) );
  NAND2_X1 U7320 ( .A1(n14447), .A2(n10732), .ZN(n10585) );
  NAND2_X2 U7321 ( .A1(n7875), .A2(n7874), .ZN(n14447) );
  XNOR2_X2 U7322 ( .A(n7678), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7813) );
  OR2_X2 U7323 ( .A1(n14111), .A2(n8135), .ZN(n7678) );
  XNOR2_X2 U7324 ( .A(n9132), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U7325 ( .A1(n6760), .A2(n11842), .ZN(n7329) );
  OAI21_X1 U7326 ( .B1(n8033), .B2(n8032), .A(n7737), .ZN(n8055) );
  NAND2_X1 U7327 ( .A1(n7733), .A2(n7732), .ZN(n8033) );
  OAI211_X1 U7328 ( .C1(n8990), .C2(n9752), .A(n7234), .B(n7233), .ZN(n11356)
         );
  INV_X1 U7329 ( .A(n10690), .ZN(n12610) );
  NAND2_X1 U7330 ( .A1(n7865), .A2(n7019), .ZN(n10637) );
  CLKBUF_X3 U7331 ( .A(n10426), .Z(n12213) );
  AND4_X1 U7332 ( .A1(n9162), .A2(n9161), .A3(n9160), .A4(n9159), .ZN(n10794)
         );
  INV_X1 U7333 ( .A(n14983), .ZN(n12611) );
  NAND2_X2 U7334 ( .A1(n10807), .A2(n14492), .ZN(n10373) );
  CLKBUF_X2 U7335 ( .A(n9139), .Z(n12540) );
  INV_X4 U7337 ( .A(n6512), .ZN(n8490) );
  CLKBUF_X2 U7338 ( .A(n6512), .Z(n8996) );
  NAND4_X1 U7339 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n13197)
         );
  INV_X1 U7340 ( .A(n10230), .ZN(n6486) );
  NAND2_X4 U7341 ( .A1(n11925), .A2(n9616), .ZN(n9103) );
  CLKBUF_X2 U7342 ( .A(n8501), .Z(n6627) );
  NOR2_X1 U7343 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7667) );
  NOR2_X1 U7344 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n7665) );
  NOR2_X1 U7345 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7666) );
  NOR2_X1 U7346 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n9076) );
  INV_X1 U7347 ( .A(n6618), .ZN(n6617) );
  OR2_X1 U7348 ( .A1(n14036), .A2(n14497), .ZN(n12024) );
  NOR2_X1 U7349 ( .A1(n12025), .A2(n13586), .ZN(n6652) );
  AND2_X1 U7350 ( .A1(n6852), .A2(n11975), .ZN(n13433) );
  OAI21_X1 U7351 ( .B1(n13278), .B2(n6889), .A(n6888), .ZN(n13243) );
  OR2_X1 U7352 ( .A1(n6828), .A2(n13231), .ZN(n6827) );
  NAND2_X1 U7353 ( .A1(n9488), .A2(n9487), .ZN(n12843) );
  NAND2_X1 U7354 ( .A1(n12248), .A2(n12247), .ZN(n12335) );
  NOR2_X1 U7355 ( .A1(n14134), .A2(n6753), .ZN(n14137) );
  AND2_X1 U7356 ( .A1(n14135), .A2(n14136), .ZN(n6753) );
  NAND2_X1 U7357 ( .A1(n12840), .A2(n12839), .ZN(n12961) );
  INV_X1 U7358 ( .A(n12246), .ZN(n12248) );
  NOR2_X1 U7359 ( .A1(n14135), .A2(n14136), .ZN(n14134) );
  NAND2_X1 U7360 ( .A1(n6616), .A2(n6513), .ZN(n6926) );
  NAND2_X1 U7361 ( .A1(n14253), .A2(n12064), .ZN(n14266) );
  NAND2_X1 U7362 ( .A1(n11864), .A2(n11863), .ZN(n12007) );
  NAND2_X1 U7363 ( .A1(n8946), .A2(n8945), .ZN(n13442) );
  NAND2_X1 U7364 ( .A1(n7329), .A2(n7328), .ZN(n14234) );
  NAND2_X1 U7365 ( .A1(n8293), .A2(n8292), .ZN(n14045) );
  NAND2_X1 U7366 ( .A1(n8896), .A2(n8895), .ZN(n13462) );
  NAND2_X1 U7367 ( .A1(n6651), .A2(n11376), .ZN(n11604) );
  NAND2_X1 U7368 ( .A1(n11768), .A2(n11769), .ZN(n9334) );
  NAND2_X1 U7369 ( .A1(n8114), .A2(n8113), .ZN(n14298) );
  NAND2_X1 U7370 ( .A1(n7346), .A2(n6507), .ZN(n11768) );
  OAI21_X1 U7371 ( .B1(n14192), .B2(n12453), .A(n12446), .ZN(n11831) );
  NAND2_X1 U7372 ( .A1(n6896), .A2(n6897), .ZN(n11234) );
  AND2_X1 U7373 ( .A1(n11662), .A2(n8123), .ZN(n11615) );
  NAND2_X1 U7374 ( .A1(n11245), .A2(n12433), .ZN(n14934) );
  NAND2_X1 U7375 ( .A1(n14948), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U7376 ( .A1(n10593), .A2(n10592), .ZN(n10767) );
  NAND2_X1 U7377 ( .A1(n8684), .A2(n8683), .ZN(n11302) );
  NAND2_X1 U7378 ( .A1(n10922), .A2(n12406), .ZN(n10921) );
  NAND2_X1 U7379 ( .A1(n8017), .A2(n8016), .ZN(n11591) );
  NAND2_X1 U7380 ( .A1(n10565), .A2(n10564), .ZN(n10589) );
  NAND2_X1 U7381 ( .A1(n6509), .A2(n9154), .ZN(n14966) );
  INV_X1 U7382 ( .A(n10581), .ZN(n14437) );
  AOI21_X1 U7383 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14876), .A(n14868), .ZN(
        n11147) );
  AOI21_X1 U7384 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14838) );
  AND2_X1 U7385 ( .A1(n7886), .A2(n10585), .ZN(n10581) );
  INV_X1 U7386 ( .A(n10751), .ZN(n14516) );
  NAND2_X2 U7387 ( .A1(n9621), .A2(n12394), .ZN(n10119) );
  NAND2_X1 U7388 ( .A1(n8550), .A2(n8549), .ZN(n10994) );
  AND4_X1 U7389 ( .A1(n9199), .A2(n9198), .A3(n9197), .A4(n9196), .ZN(n10838)
         );
  AND4_X1 U7390 ( .A1(n9143), .A2(n9142), .A3(n9141), .A4(n9140), .ZN(n14983)
         );
  AND3_X1 U7391 ( .A1(n9135), .A2(n9134), .A3(n9133), .ZN(n10093) );
  NAND2_X2 U7392 ( .A1(n8506), .A2(n8505), .ZN(n10654) );
  AND2_X2 U7393 ( .A1(n10278), .A2(n10281), .ZN(n10807) );
  CLKBUF_X1 U7394 ( .A(n9387), .Z(n12543) );
  INV_X1 U7395 ( .A(n14354), .ZN(n10374) );
  NAND4_X2 U7396 ( .A1(n8500), .A2(n8499), .A3(n8498), .A4(n8497), .ZN(n13200)
         );
  NAND4_X1 U7397 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(n9020)
         );
  NAND2_X1 U7398 ( .A1(n9607), .A2(n9661), .ZN(n12393) );
  OR2_X1 U7399 ( .A1(n6477), .A2(n13703), .ZN(n7879) );
  OAI21_X1 U7400 ( .B1(n7835), .B2(n7834), .A(n6469), .ZN(n6806) );
  NOR2_X1 U7401 ( .A1(n7709), .A2(n7710), .ZN(n7711) );
  NAND2_X1 U7402 ( .A1(n9652), .A2(n9651), .ZN(n11632) );
  OR2_X2 U7403 ( .A1(n10470), .A2(n10284), .ZN(n14492) );
  NAND2_X2 U7404 ( .A1(n9733), .A2(P3_U3151), .ZN(n13058) );
  NAND2_X2 U7405 ( .A1(n9733), .A2(P1_U3086), .ZN(n14125) );
  NAND2_X2 U7406 ( .A1(n8455), .A2(n8458), .ZN(n8966) );
  XNOR2_X1 U7407 ( .A(n8426), .B(P1_IR_REG_24__SCAN_IN), .ZN(n10257) );
  XNOR2_X1 U7408 ( .A(n9609), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U7409 ( .A1(n8486), .A2(n8485), .ZN(n13576) );
  OAI21_X1 U7410 ( .B1(n8432), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8434) );
  NAND2_X2 U7411 ( .A1(n11928), .A2(n14122), .ZN(n9896) );
  NAND2_X1 U7412 ( .A1(n14119), .A2(n14120), .ZN(n8205) );
  AND2_X1 U7413 ( .A1(n8431), .A2(n7795), .ZN(n10262) );
  NAND2_X2 U7414 ( .A1(n9727), .A2(P1_U3086), .ZN(n14128) );
  OR2_X1 U7415 ( .A1(n9605), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n9661) );
  XNOR2_X1 U7416 ( .A(n7699), .B(SI_1_), .ZN(n7835) );
  MUX2_X1 U7417 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8484), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8486) );
  XNOR2_X1 U7418 ( .A(n7800), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U7419 ( .A(n7686), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10284) );
  INV_X1 U7420 ( .A(n7842), .ZN(n6487) );
  OR2_X1 U7421 ( .A1(n7796), .A2(n7212), .ZN(n6615) );
  OR2_X1 U7422 ( .A1(n8420), .A2(n8135), .ZN(n7800) );
  NAND2_X1 U7423 ( .A1(n7803), .A2(n8429), .ZN(n13897) );
  OR2_X1 U7424 ( .A1(n8451), .A2(n8728), .ZN(n7287) );
  NOR2_X2 U7425 ( .A1(n8713), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U7426 ( .A1(n7797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7794) );
  AOI21_X1 U7427 ( .B1(n6745), .B2(n6520), .A(n7432), .ZN(n7394) );
  AND3_X2 U7428 ( .A1(n6776), .A2(n6775), .A3(n8468), .ZN(n8473) );
  NAND2_X1 U7429 ( .A1(n6744), .A2(n7435), .ZN(n6745) );
  AND2_X1 U7430 ( .A1(n6514), .A2(n9148), .ZN(n9243) );
  AND2_X1 U7431 ( .A1(n7338), .A2(n7339), .ZN(n6776) );
  AND2_X1 U7432 ( .A1(n8547), .A2(n8443), .ZN(n6775) );
  AND3_X1 U7433 ( .A1(n8440), .A2(n6761), .A3(n8503), .ZN(n8547) );
  AND3_X1 U7434 ( .A1(n8465), .A2(n8442), .A3(n8441), .ZN(n8468) );
  AND2_X1 U7435 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n6940), .ZN(n7435) );
  AND2_X1 U7436 ( .A1(n7675), .A2(n7674), .ZN(n7685) );
  AND3_X1 U7437 ( .A1(n7341), .A2(n8587), .A3(n7340), .ZN(n7339) );
  AND3_X1 U7438 ( .A1(n7256), .A2(n7255), .A3(n7254), .ZN(n7338) );
  INV_X1 U7439 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8440) );
  NOR2_X1 U7440 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n9073) );
  NOR2_X1 U7441 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7674) );
  NOR2_X1 U7442 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n7675) );
  INV_X4 U7443 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7444 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9275) );
  INV_X1 U7445 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9256) );
  NOR2_X1 U7446 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8465) );
  INV_X1 U7447 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9168) );
  INV_X1 U7448 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9343) );
  INV_X4 U7449 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7450 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9082) );
  NOR3_X1 U7451 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .A3(
        P3_IR_REG_25__SCAN_IN), .ZN(n9079) );
  INV_X1 U7452 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7696) );
  NOR2_X1 U7453 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n9078) );
  NOR2_X1 U7454 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n9077) );
  INV_X4 U7455 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7456 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7256) );
  NOR2_X1 U7457 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7255) );
  NOR2_X1 U7458 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7254) );
  INV_X1 U7459 ( .A(n10201), .ZN(n10203) );
  AND2_X2 U7460 ( .A1(n9137), .A2(n9136), .ZN(n6509) );
  NAND2_X1 U7461 ( .A1(n9087), .A2(n9089), .ZN(n9139) );
  INV_X1 U7462 ( .A(n9896), .ZN(n6488) );
  NAND2_X2 U7463 ( .A1(n12771), .A2(n9573), .ZN(n12770) );
  AOI21_X2 U7464 ( .B1(n11007), .B2(n7195), .A(n7194), .ZN(n7193) );
  NOR2_X2 U7465 ( .A1(n11237), .A2(n11701), .ZN(n6820) );
  AND2_X1 U7466 ( .A1(n7813), .A2(n7812), .ZN(n7842) );
  XNOR2_X2 U7467 ( .A(n9085), .B(P3_IR_REG_29__SCAN_IN), .ZN(n9088) );
  NOR2_X2 U7468 ( .A1(n8476), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n9040) );
  XNOR2_X2 U7469 ( .A(n14276), .B(n13679), .ZN(n11227) );
  NAND2_X4 U7470 ( .A1(n8039), .A2(n8038), .ZN(n14276) );
  NOR2_X2 U7471 ( .A1(n13341), .A2(n13474), .ZN(n13325) );
  NOR2_X2 U7472 ( .A1(n11798), .A2(n14256), .ZN(n11873) );
  AOI21_X2 U7473 ( .B1(n7482), .B2(n7481), .A(n14335), .ZN(n14341) );
  OR2_X1 U7474 ( .A1(n12976), .A2(n12885), .ZN(n12488) );
  NAND2_X1 U7475 ( .A1(n7738), .A2(n9760), .ZN(n7741) );
  NAND2_X1 U7476 ( .A1(n7176), .A2(n12517), .ZN(n7175) );
  OR2_X1 U7477 ( .A1(n12268), .A2(n12773), .ZN(n12521) );
  NOR2_X1 U7478 ( .A1(n12873), .A2(n7361), .ZN(n7360) );
  INV_X1 U7479 ( .A(n9451), .ZN(n7361) );
  NOR2_X1 U7480 ( .A1(n6990), .A2(n6986), .ZN(n9099) );
  INV_X1 U7481 ( .A(n8455), .ZN(n8457) );
  INV_X1 U7482 ( .A(n11945), .ZN(n13432) );
  NAND2_X1 U7483 ( .A1(n7791), .A2(n7790), .ZN(n8368) );
  NAND2_X1 U7484 ( .A1(n7824), .A2(n7823), .ZN(n7791) );
  NAND2_X1 U7485 ( .A1(n9693), .A2(n12560), .ZN(n15001) );
  OR2_X1 U7486 ( .A1(n13376), .A2(n11954), .ZN(n11956) );
  INV_X1 U7487 ( .A(n8190), .ZN(n7043) );
  INV_X1 U7488 ( .A(n7071), .ZN(n7070) );
  INV_X1 U7489 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9100) );
  INV_X1 U7490 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U7491 ( .A1(n6890), .A2(n6808), .ZN(n6810) );
  INV_X1 U7492 ( .A(n6892), .ZN(n6808) );
  AND2_X1 U7493 ( .A1(n8445), .A2(n8444), .ZN(n9048) );
  NAND2_X1 U7494 ( .A1(n7771), .A2(n7770), .ZN(n7772) );
  AND2_X1 U7495 ( .A1(n7392), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7393) );
  INV_X1 U7496 ( .A(n9157), .ZN(n9312) );
  NAND2_X1 U7497 ( .A1(n14807), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U7498 ( .A1(n9090), .A2(n9089), .ZN(n9387) );
  NAND2_X1 U7499 ( .A1(n9629), .A2(n12448), .ZN(n14192) );
  NAND2_X1 U7500 ( .A1(n7373), .A2(n9100), .ZN(n6989) );
  OAI21_X1 U7501 ( .B1(n9504), .B2(n7172), .A(n7170), .ZN(n9519) );
  INV_X1 U7502 ( .A(n7173), .ZN(n7172) );
  AOI21_X1 U7503 ( .B1(n7173), .B2(n7171), .A(n6609), .ZN(n7170) );
  AOI21_X1 U7504 ( .B1(n9503), .B2(n9505), .A(n7174), .ZN(n7173) );
  NOR2_X1 U7505 ( .A1(n9646), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n9603) );
  AND2_X1 U7506 ( .A1(n7152), .A2(n6678), .ZN(n6677) );
  NAND2_X1 U7507 ( .A1(n9359), .A2(n9376), .ZN(n6678) );
  INV_X1 U7508 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9070) );
  INV_X1 U7509 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9074) );
  NOR2_X1 U7510 ( .A1(n11416), .A2(n7303), .ZN(n7302) );
  INV_X1 U7511 ( .A(n11102), .ZN(n7303) );
  INV_X1 U7512 ( .A(n8453), .ZN(n8458) );
  INV_X1 U7513 ( .A(n11279), .ZN(n6871) );
  NAND2_X1 U7514 ( .A1(n7235), .A2(n11356), .ZN(n10662) );
  AND2_X1 U7515 ( .A1(n8473), .A2(n9048), .ZN(n9051) );
  NOR2_X1 U7516 ( .A1(n14282), .A2(n7111), .ZN(n7110) );
  NOR2_X1 U7517 ( .A1(n14264), .A2(n14262), .ZN(n7111) );
  INV_X1 U7518 ( .A(n10373), .ZN(n12135) );
  OR2_X1 U7519 ( .A1(n14298), .A2(n12055), .ZN(n11795) );
  OR2_X1 U7520 ( .A1(n14247), .A2(n12041), .ZN(n11662) );
  AND2_X1 U7521 ( .A1(n10599), .A2(n8401), .ZN(n10595) );
  AND2_X1 U7522 ( .A1(n10284), .A2(n11297), .ZN(n10468) );
  OAI21_X1 U7523 ( .B1(n8339), .B2(n8338), .A(n7787), .ZN(n7824) );
  XNOR2_X1 U7524 ( .A(n7774), .B(n11295), .ZN(n7773) );
  INV_X1 U7525 ( .A(n7077), .ZN(n7076) );
  NOR2_X2 U7526 ( .A1(n7801), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n7687) );
  NAND2_X1 U7527 ( .A1(n6796), .A2(n6794), .ZN(n8134) );
  AOI21_X1 U7528 ( .B1(n6798), .B2(n6801), .A(n6795), .ZN(n6794) );
  INV_X1 U7529 ( .A(n7741), .ZN(n6801) );
  XNOR2_X1 U7530 ( .A(n7705), .B(SI_3_), .ZN(n7871) );
  XNOR2_X1 U7531 ( .A(n7007), .B(n12723), .ZN(n7006) );
  OAI22_X1 U7532 ( .A1(n12559), .A2(n12558), .B1(n12749), .B2(n12557), .ZN(
        n7007) );
  NAND2_X1 U7533 ( .A1(n7177), .A2(n12553), .ZN(n12549) );
  OAI211_X1 U7534 ( .C1(n12526), .C2(n12514), .A(n7178), .B(n12550), .ZN(n7177) );
  BUF_X1 U7535 ( .A(n9312), .Z(n9594) );
  INV_X1 U7536 ( .A(n9574), .ZN(n7354) );
  OR2_X1 U7537 ( .A1(n9537), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9566) );
  OR2_X1 U7538 ( .A1(n12963), .A2(n12845), .ZN(n12812) );
  NAND2_X1 U7539 ( .A1(n7011), .A2(n7009), .ZN(n12876) );
  AND2_X1 U7540 ( .A1(n12873), .A2(n7010), .ZN(n7009) );
  NAND2_X1 U7541 ( .A1(n7013), .A2(n7012), .ZN(n7010) );
  NAND2_X1 U7542 ( .A1(n12883), .A2(n9450), .ZN(n9452) );
  OR2_X1 U7543 ( .A1(n12367), .A2(n12886), .ZN(n12474) );
  AND2_X1 U7544 ( .A1(n14193), .A2(n6506), .ZN(n7358) );
  AND2_X1 U7545 ( .A1(n12525), .A2(n10114), .ZN(n14962) );
  NAND2_X1 U7546 ( .A1(n9645), .A2(n7368), .ZN(n7365) );
  INV_X1 U7547 ( .A(n9475), .ZN(n12537) );
  OAI21_X1 U7548 ( .B1(n9576), .B2(n9575), .A(n9577), .ZN(n9588) );
  XNOR2_X1 U7549 ( .A(n9654), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U7550 ( .A1(n7163), .A2(n7165), .ZN(n9456) );
  NAND2_X1 U7551 ( .A1(n6653), .A2(n6654), .ZN(n9183) );
  AOI21_X1 U7552 ( .B1(n7119), .B2(n9163), .A(n7120), .ZN(n6654) );
  INV_X1 U7553 ( .A(n9165), .ZN(n7120) );
  NOR2_X1 U7554 ( .A1(n13074), .A2(n7322), .ZN(n7321) );
  INV_X1 U7555 ( .A(n12174), .ZN(n7322) );
  NAND2_X2 U7556 ( .A1(n13576), .A2(n10209), .ZN(n9770) );
  AOI21_X1 U7557 ( .B1(n7321), .B2(n7319), .A(n7318), .ZN(n7317) );
  INV_X1 U7558 ( .A(n12180), .ZN(n7318) );
  INV_X1 U7559 ( .A(n7324), .ZN(n7319) );
  NOR2_X1 U7560 ( .A1(n7320), .A2(n6767), .ZN(n6766) );
  INV_X1 U7561 ( .A(n13111), .ZN(n6767) );
  INV_X1 U7562 ( .A(n7321), .ZN(n7320) );
  AND2_X1 U7563 ( .A1(n7062), .A2(n11971), .ZN(n7061) );
  NOR2_X1 U7564 ( .A1(n13244), .A2(n7063), .ZN(n7062) );
  NAND2_X1 U7565 ( .A1(n6890), .A2(n7064), .ZN(n7063) );
  NOR2_X1 U7566 ( .A1(n9032), .A2(n13280), .ZN(n7064) );
  AND4_X1 U7567 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n13061)
         );
  INV_X1 U7568 ( .A(n6829), .ZN(n6828) );
  AOI21_X1 U7569 ( .B1(n13238), .B2(n13432), .A(n10230), .ZN(n6829) );
  NAND2_X1 U7570 ( .A1(n13307), .A2(n11934), .ZN(n11937) );
  NAND2_X1 U7571 ( .A1(n6873), .A2(n6875), .ZN(n13293) );
  INV_X1 U7572 ( .A(n6876), .ZN(n6875) );
  NAND2_X1 U7573 ( .A1(n13337), .A2(n6874), .ZN(n6873) );
  OAI21_X1 U7574 ( .B1(n6878), .B2(n6877), .A(n7380), .ZN(n6876) );
  OAI21_X1 U7575 ( .B1(n7244), .B2(n7243), .A(n6557), .ZN(n11933) );
  INV_X1 U7576 ( .A(n7249), .ZN(n7243) );
  AOI21_X1 U7577 ( .B1(n13363), .B2(n6844), .A(n6531), .ZN(n6843) );
  INV_X1 U7578 ( .A(n11955), .ZN(n6844) );
  AND2_X1 U7579 ( .A1(n6855), .A2(n11951), .ZN(n6854) );
  NAND2_X1 U7580 ( .A1(n6860), .A2(n6859), .ZN(n6858) );
  NOR2_X1 U7581 ( .A1(n11782), .A2(n6863), .ZN(n6862) );
  INV_X1 U7582 ( .A(n11738), .ZN(n6863) );
  OAI22_X1 U7583 ( .A1(n11658), .A2(n11657), .B1(n13539), .B2(n13187), .ZN(
        n11740) );
  NOR2_X1 U7584 ( .A1(n6530), .A2(n6791), .ZN(n6790) );
  INV_X1 U7585 ( .A(n11515), .ZN(n6791) );
  OAI22_X1 U7586 ( .A1(n11495), .A2(n7237), .B1(n7236), .B2(n7238), .ZN(n11514) );
  INV_X1 U7587 ( .A(n7241), .ZN(n7236) );
  NAND2_X1 U7588 ( .A1(n11273), .A2(n7241), .ZN(n7237) );
  AND2_X1 U7589 ( .A1(n7239), .A2(n11298), .ZN(n7238) );
  INV_X2 U7590 ( .A(n9770), .ZN(n8815) );
  AND2_X1 U7591 ( .A1(n6521), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U7592 ( .A1(n14266), .A2(n7110), .ZN(n7108) );
  OR2_X1 U7593 ( .A1(n8414), .A2(n8379), .ZN(n6634) );
  NAND2_X1 U7594 ( .A1(n6813), .A2(n6812), .ZN(n6811) );
  NOR2_X1 U7595 ( .A1(n14071), .A2(n13947), .ZN(n6812) );
  INV_X1 U7596 ( .A(n6814), .ZN(n6813) );
  OR2_X1 U7597 ( .A1(n14131), .A2(n10284), .ZN(n10570) );
  NOR2_X1 U7598 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7213) );
  INV_X1 U7599 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6940) );
  OAI22_X1 U7600 ( .A1(n7427), .A2(n7415), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n11724), .ZN(n7425) );
  OAI21_X1 U7601 ( .B1(n12771), .B2(n7357), .A(n7353), .ZN(n9601) );
  AOI21_X1 U7602 ( .B1(n7356), .B2(n12769), .A(n6594), .ZN(n7353) );
  NAND2_X1 U7603 ( .A1(n14503), .A2(n14354), .ZN(n7883) );
  OR2_X1 U7604 ( .A1(n8524), .A2(n8523), .ZN(n7379) );
  NAND2_X1 U7605 ( .A1(n8537), .A2(n7283), .ZN(n7281) );
  NAND2_X1 U7606 ( .A1(n7016), .A2(n7015), .ZN(n7923) );
  NOR2_X1 U7607 ( .A1(n7030), .A2(n8001), .ZN(n7031) );
  NAND2_X1 U7608 ( .A1(n7030), .A2(n8001), .ZN(n7029) );
  NAND2_X1 U7609 ( .A1(n6640), .A2(n6639), .ZN(n8084) );
  NAND2_X1 U7610 ( .A1(n8060), .A2(n8062), .ZN(n6639) );
  NOR2_X1 U7611 ( .A1(n8803), .A2(n7294), .ZN(n7293) );
  INV_X1 U7612 ( .A(n8198), .ZN(n7038) );
  AND2_X1 U7613 ( .A1(n7039), .A2(n8147), .ZN(n7035) );
  OAI21_X1 U7614 ( .B1(n8264), .B2(n7024), .A(n7023), .ZN(n8279) );
  INV_X1 U7615 ( .A(n8947), .ZN(n7266) );
  INV_X1 U7616 ( .A(n8948), .ZN(n7262) );
  INV_X1 U7617 ( .A(n7750), .ZN(n6731) );
  INV_X1 U7618 ( .A(n8133), .ZN(n6728) );
  INV_X1 U7619 ( .A(n7069), .ZN(n7068) );
  OAI21_X1 U7620 ( .B1(n7072), .B2(n7070), .A(n7744), .ZN(n7069) );
  NAND2_X1 U7621 ( .A1(n7266), .A2(n7262), .ZN(n7260) );
  NOR2_X1 U7622 ( .A1(n7266), .A2(n7262), .ZN(n7261) );
  INV_X1 U7623 ( .A(n8980), .ZN(n7264) );
  INV_X1 U7624 ( .A(n8979), .ZN(n7265) );
  AND2_X1 U7625 ( .A1(n9035), .A2(n8981), .ZN(n8982) );
  AND2_X1 U7626 ( .A1(n13982), .A2(n14000), .ZN(n8398) );
  NAND2_X1 U7627 ( .A1(n7781), .A2(n11645), .ZN(n7056) );
  AND2_X1 U7628 ( .A1(n7058), .A2(n6508), .ZN(n7053) );
  AOI21_X1 U7629 ( .B1(n7077), .B2(n7074), .A(n6596), .ZN(n6802) );
  NAND2_X1 U7630 ( .A1(n8862), .A2(SI_22_), .ZN(n7079) );
  NAND2_X1 U7631 ( .A1(n7753), .A2(n7078), .ZN(n7077) );
  INV_X1 U7632 ( .A(n8164), .ZN(n7078) );
  NAND2_X1 U7633 ( .A1(n7734), .A2(n9745), .ZN(n7737) );
  AND2_X1 U7634 ( .A1(n6535), .A2(n6942), .ZN(n7398) );
  INV_X1 U7635 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7397) );
  INV_X1 U7636 ( .A(n12296), .ZN(n6703) );
  OR2_X1 U7637 ( .A1(n11075), .A2(n7124), .ZN(n7123) );
  OAI21_X1 U7638 ( .B1(n12243), .B2(n6523), .A(n6722), .ZN(n12246) );
  OR2_X1 U7639 ( .A1(n12242), .A2(n12857), .ZN(n6722) );
  NOR2_X1 U7640 ( .A1(n10948), .A2(n6707), .ZN(n6706) );
  INV_X1 U7641 ( .A(n10950), .ZN(n6707) );
  INV_X1 U7642 ( .A(n12289), .ZN(n6720) );
  NAND2_X1 U7643 ( .A1(n12520), .A2(n12514), .ZN(n7178) );
  NAND2_X1 U7644 ( .A1(n14810), .A2(n11155), .ZN(n11156) );
  OR2_X1 U7645 ( .A1(n12849), .A2(n12857), .ZN(n12500) );
  NOR2_X1 U7646 ( .A1(n6996), .A2(n12575), .ZN(n6992) );
  INV_X1 U7647 ( .A(n12923), .ZN(n6996) );
  AND2_X1 U7648 ( .A1(n9192), .A2(n9174), .ZN(n7370) );
  INV_X1 U7649 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U7650 ( .A1(n9454), .A2(n6510), .ZN(n7163) );
  INV_X1 U7651 ( .A(n7158), .ZN(n7157) );
  OAI21_X1 U7652 ( .B1(n9272), .B2(n7159), .A(n9298), .ZN(n7158) );
  INV_X1 U7653 ( .A(n9293), .ZN(n7159) );
  CLKBUF_X1 U7654 ( .A(n9243), .Z(n9244) );
  AND2_X1 U7655 ( .A1(n7139), .A2(n9222), .ZN(n7138) );
  INV_X1 U7656 ( .A(n9225), .ZN(n7139) );
  NOR2_X1 U7657 ( .A1(n13457), .A2(n6834), .ZN(n6833) );
  INV_X1 U7658 ( .A(n6835), .ZN(n6834) );
  INV_X1 U7659 ( .A(n11949), .ZN(n6859) );
  NOR2_X1 U7660 ( .A1(n11302), .A2(n6825), .ZN(n6824) );
  INV_X1 U7661 ( .A(n6826), .ZN(n6825) );
  INV_X1 U7662 ( .A(n6870), .ZN(n6869) );
  OAI21_X1 U7663 ( .B1(n11472), .B2(n6871), .A(n11280), .ZN(n6870) );
  OAI21_X1 U7664 ( .B1(n10981), .B2(n6780), .A(n11053), .ZN(n6777) );
  NAND2_X1 U7665 ( .A1(n6565), .A2(n6494), .ZN(n6878) );
  NAND2_X1 U7666 ( .A1(n11962), .A2(n11961), .ZN(n6881) );
  NAND2_X1 U7667 ( .A1(n10656), .A2(n10655), .ZN(n11349) );
  NAND2_X1 U7668 ( .A1(n10662), .A2(n9023), .ZN(n11348) );
  AND2_X1 U7669 ( .A1(n8479), .A2(n8487), .ZN(n10236) );
  INV_X1 U7670 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7333) );
  AND2_X1 U7671 ( .A1(n8465), .A2(n8464), .ZN(n7334) );
  NAND2_X1 U7672 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  INV_X1 U7673 ( .A(n8356), .ZN(n8361) );
  INV_X1 U7674 ( .A(n14022), .ZN(n13841) );
  NAND2_X1 U7675 ( .A1(n13893), .A2(n7207), .ZN(n7206) );
  INV_X1 U7676 ( .A(n12001), .ZN(n7207) );
  NAND2_X1 U7677 ( .A1(n13994), .A2(n11993), .ZN(n7199) );
  AOI21_X1 U7678 ( .B1(n7191), .B2(n7189), .A(n11374), .ZN(n7188) );
  NOR2_X2 U7679 ( .A1(n13915), .A2(n14045), .ZN(n13881) );
  OAI21_X1 U7680 ( .B1(n13942), .B2(n13944), .A(n11998), .ZN(n13929) );
  NAND2_X1 U7681 ( .A1(n13929), .A2(n13928), .ZN(n13927) );
  OAI21_X1 U7682 ( .B1(n8326), .B2(n7784), .A(n7783), .ZN(n8339) );
  AND2_X1 U7683 ( .A1(n7775), .A2(n7059), .ZN(n7058) );
  INV_X1 U7684 ( .A(n8290), .ZN(n7059) );
  AND2_X1 U7685 ( .A1(n7106), .A2(n7105), .ZN(n7104) );
  INV_X1 U7686 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U7687 ( .A1(n7067), .A2(n7071), .ZN(n8105) );
  XNOR2_X1 U7688 ( .A(n8105), .B(n9822), .ZN(n8102) );
  NAND2_X1 U7689 ( .A1(n7704), .A2(n7051), .ZN(n7050) );
  AND2_X1 U7690 ( .A1(n7703), .A2(n7712), .ZN(n7051) );
  NAND2_X1 U7691 ( .A1(n6806), .A2(SI_2_), .ZN(n7869) );
  NOR2_X1 U7692 ( .A1(n7405), .A2(n7404), .ZN(n7461) );
  INV_X1 U7693 ( .A(n6756), .ZN(n7408) );
  OAI21_X1 U7694 ( .B1(n7466), .B2(n7465), .A(n6757), .ZN(n6756) );
  NAND2_X1 U7695 ( .A1(n7407), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U7696 ( .A1(n6694), .A2(n6695), .ZN(n10941) );
  AOI21_X1 U7697 ( .B1(n6699), .B2(n10508), .A(n6552), .ZN(n6695) );
  OAI21_X1 U7698 ( .B1(n7148), .B2(n7149), .A(n7145), .ZN(n7143) );
  NAND2_X1 U7699 ( .A1(n6567), .A2(n12910), .ZN(n7145) );
  AOI21_X1 U7700 ( .B1(n12276), .B2(n12260), .A(n12264), .ZN(n7133) );
  INV_X1 U7701 ( .A(n7133), .ZN(n7129) );
  NAND2_X1 U7702 ( .A1(n6713), .A2(n12347), .ZN(n6712) );
  NAND2_X1 U7703 ( .A1(n6717), .A2(n6719), .ZN(n6713) );
  NAND2_X1 U7704 ( .A1(n12283), .A2(n12335), .ZN(n12253) );
  NOR2_X1 U7705 ( .A1(n7168), .A2(n10399), .ZN(n7167) );
  INV_X1 U7706 ( .A(n10396), .ZN(n7168) );
  AND2_X1 U7707 ( .A1(n9261), .A2(n9260), .ZN(n12432) );
  NAND2_X1 U7708 ( .A1(n12297), .A2(n12296), .ZN(n6708) );
  NAND2_X1 U7709 ( .A1(n6708), .A2(n6706), .ZN(n11076) );
  NAND2_X1 U7710 ( .A1(n15014), .A2(n14999), .ZN(n14993) );
  AOI21_X1 U7711 ( .B1(n7143), .B2(n6720), .A(n6718), .ZN(n6717) );
  NOR2_X1 U7712 ( .A1(n12236), .A2(n12899), .ZN(n6718) );
  NOR2_X1 U7713 ( .A1(n12230), .A2(n12229), .ZN(n12232) );
  NOR2_X1 U7714 ( .A1(n10059), .A2(n10060), .ZN(n11151) );
  NAND2_X1 U7715 ( .A1(n14812), .A2(n14811), .ZN(n14810) );
  XNOR2_X1 U7716 ( .A(n11156), .B(n11181), .ZN(n14828) );
  NAND2_X1 U7717 ( .A1(n14799), .A2(n6920), .ZN(n6917) );
  AOI21_X1 U7718 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n14842), .A(n14833), .ZN(
        n11144) );
  NOR2_X1 U7719 ( .A1(n11193), .A2(n11144), .ZN(n11145) );
  OR2_X1 U7720 ( .A1(n14853), .A2(n14958), .ZN(n6908) );
  OR2_X1 U7721 ( .A1(n14920), .A2(n14919), .ZN(n6916) );
  NAND2_X1 U7722 ( .A1(n6916), .A2(n6915), .ZN(n6914) );
  NAND2_X1 U7723 ( .A1(n11213), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U7724 ( .A1(n12639), .A2(n6642), .ZN(n12660) );
  AND2_X1 U7725 ( .A1(n12644), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U7726 ( .A1(n12642), .A2(n12645), .ZN(n12666) );
  NAND2_X1 U7727 ( .A1(n9633), .A2(n12510), .ZN(n12783) );
  AOI21_X1 U7728 ( .B1(n12800), .B2(n7345), .A(n6556), .ZN(n7344) );
  NAND2_X1 U7729 ( .A1(n12815), .A2(n9531), .ZN(n12801) );
  NAND2_X1 U7730 ( .A1(n12817), .A2(n12816), .ZN(n12815) );
  AND2_X1 U7731 ( .A1(n12812), .A2(n12501), .ZN(n12839) );
  NAND2_X1 U7732 ( .A1(n12897), .A2(n7014), .ZN(n7013) );
  NAND2_X1 U7733 ( .A1(n6503), .A2(n7014), .ZN(n7012) );
  NAND2_X1 U7734 ( .A1(n9632), .A2(n12472), .ZN(n12902) );
  OR2_X1 U7735 ( .A1(n12902), .A2(n9429), .ZN(n12900) );
  AND3_X1 U7736 ( .A1(n9408), .A2(n9407), .A3(n9406), .ZN(n12922) );
  INV_X1 U7737 ( .A(n11831), .ZN(n6966) );
  NAND2_X1 U7738 ( .A1(n11888), .A2(n12460), .ZN(n11887) );
  AOI21_X1 U7739 ( .B1(n7001), .B2(n6999), .A(n6998), .ZN(n6997) );
  INV_X1 U7740 ( .A(n7001), .ZN(n7000) );
  INV_X1 U7741 ( .A(n12437), .ZN(n6999) );
  NOR2_X1 U7742 ( .A1(n7352), .A2(n7351), .ZN(n7350) );
  AND4_X1 U7743 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), .ZN(n14202)
         );
  AND2_X1 U7744 ( .A1(n12442), .A2(n12443), .ZN(n14205) );
  NAND2_X1 U7745 ( .A1(n14934), .A2(n14933), .ZN(n14932) );
  INV_X1 U7746 ( .A(n14962), .ZN(n14996) );
  NAND2_X1 U7747 ( .A1(n9441), .A2(n9440), .ZN(n12561) );
  NAND2_X1 U7748 ( .A1(n9402), .A2(n9401), .ZN(n12988) );
  AND2_X1 U7749 ( .A1(n13046), .A2(n10080), .ZN(n10337) );
  AND2_X1 U7750 ( .A1(n9075), .A2(n6988), .ZN(n6983) );
  NOR2_X1 U7751 ( .A1(n6989), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n6988) );
  OR2_X1 U7752 ( .A1(n9588), .A2(n9587), .ZN(n9591) );
  NAND2_X1 U7753 ( .A1(n6684), .A2(n9559), .ZN(n9576) );
  OR2_X1 U7754 ( .A1(n9558), .A2(n9557), .ZN(n6684) );
  OR2_X1 U7755 ( .A1(n7372), .A2(n9398), .ZN(n9651) );
  INV_X1 U7756 ( .A(n7383), .ZN(n7372) );
  OR2_X1 U7757 ( .A1(n9519), .A2(n11839), .ZN(n9532) );
  INV_X1 U7758 ( .A(n9532), .ZN(n6670) );
  NAND2_X1 U7759 ( .A1(n9520), .A2(n6672), .ZN(n6671) );
  AND2_X1 U7760 ( .A1(n9647), .A2(n6693), .ZN(n6691) );
  NAND2_X1 U7761 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6692) );
  OAI21_X1 U7762 ( .B1(n9647), .B2(n6692), .A(n6690), .ZN(n6689) );
  NAND2_X1 U7763 ( .A1(n6693), .A2(n9098), .ZN(n6690) );
  NAND2_X1 U7764 ( .A1(n9490), .A2(n9489), .ZN(n9504) );
  NAND2_X1 U7765 ( .A1(n9473), .A2(n9472), .ZN(n9490) );
  NAND2_X1 U7766 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U7767 ( .A1(n9455), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7165) );
  INV_X1 U7768 ( .A(n6677), .ZN(n6676) );
  AND2_X1 U7769 ( .A1(n6674), .A2(n7150), .ZN(n6673) );
  AOI21_X1 U7770 ( .B1(n7152), .B2(n7154), .A(n7151), .ZN(n7150) );
  NOR2_X1 U7771 ( .A1(n9071), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U7772 ( .A1(n9377), .A2(n9376), .ZN(n9380) );
  AND2_X1 U7773 ( .A1(n9395), .A2(n9378), .ZN(n9379) );
  NAND2_X1 U7774 ( .A1(n9380), .A2(n9379), .ZN(n9396) );
  NAND2_X1 U7775 ( .A1(n9339), .A2(n9338), .ZN(n9356) );
  NAND2_X1 U7776 ( .A1(n9335), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9339) );
  XNOR2_X1 U7777 ( .A(n9337), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U7778 ( .A1(n9270), .A2(n9269), .ZN(n9273) );
  NAND2_X1 U7779 ( .A1(n9273), .A2(n9272), .ZN(n9294) );
  AND2_X1 U7780 ( .A1(n9250), .A2(n9239), .ZN(n9240) );
  OAI21_X1 U7781 ( .B1(n9223), .B2(n7137), .A(n7135), .ZN(n9251) );
  INV_X1 U7782 ( .A(n7136), .ZN(n7135) );
  OAI21_X1 U7783 ( .B1(n7138), .B2(n7137), .A(n9240), .ZN(n7136) );
  INV_X1 U7784 ( .A(n9237), .ZN(n7137) );
  NAND2_X1 U7785 ( .A1(n9223), .A2(n7138), .ZN(n9238) );
  AND2_X1 U7786 ( .A1(n9184), .A2(n9166), .ZN(n9182) );
  AND2_X1 U7787 ( .A1(n9147), .A2(n9165), .ZN(n9163) );
  NAND2_X1 U7788 ( .A1(n9129), .A2(n9128), .ZN(n9145) );
  AND2_X1 U7789 ( .A1(n9146), .A2(n9130), .ZN(n9144) );
  NAND2_X1 U7790 ( .A1(n7305), .A2(n7308), .ZN(n7304) );
  INV_X1 U7791 ( .A(n7306), .ZN(n7305) );
  AOI21_X1 U7792 ( .B1(n11103), .B2(n11102), .A(n7307), .ZN(n7306) );
  NAND2_X1 U7793 ( .A1(n11104), .A2(n7302), .ZN(n7299) );
  INV_X1 U7794 ( .A(n6763), .ZN(n6762) );
  INV_X1 U7795 ( .A(n7317), .ZN(n6765) );
  NOR2_X1 U7796 ( .A1(n7304), .A2(n7301), .ZN(n7300) );
  INV_X1 U7797 ( .A(n11420), .ZN(n7301) );
  NAND2_X1 U7798 ( .A1(n11104), .A2(n6532), .ZN(n7298) );
  NOR2_X1 U7799 ( .A1(n12204), .A2(n12203), .ZN(n7313) );
  AND4_X1 U7800 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n11648)
         );
  OR2_X1 U7801 ( .A1(n8526), .A2(n8456), .ZN(n8460) );
  AND2_X1 U7802 ( .A1(n8463), .A2(n8440), .ZN(n7336) );
  INV_X1 U7803 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8463) );
  XOR2_X1 U7804 ( .A(n14653), .B(n11117), .Z(n14656) );
  NAND2_X1 U7805 ( .A1(n8963), .A2(n8962), .ZN(n13227) );
  AOI21_X1 U7806 ( .B1(n13569), .B2(n6489), .A(n8978), .ZN(n11945) );
  AND2_X1 U7807 ( .A1(n9017), .A2(n11940), .ZN(n13244) );
  AOI21_X1 U7808 ( .B1(n11969), .B2(n11965), .A(n11968), .ZN(n6892) );
  NAND2_X1 U7809 ( .A1(n6894), .A2(n11969), .ZN(n6893) );
  AND2_X1 U7810 ( .A1(n11969), .A2(n11967), .ZN(n13266) );
  AOI21_X1 U7811 ( .B1(n7220), .B2(n7223), .A(n6559), .ZN(n7218) );
  NOR2_X1 U7812 ( .A1(n6495), .A2(n11935), .ZN(n7224) );
  AOI21_X1 U7813 ( .B1(n7222), .B2(n7221), .A(n6894), .ZN(n7220) );
  INV_X1 U7814 ( .A(n7224), .ZN(n7221) );
  AOI22_X1 U7815 ( .A1(n13293), .A2(n13292), .B1(n13094), .B2(n13462), .ZN(
        n13278) );
  NAND2_X1 U7816 ( .A1(n13331), .A2(n6537), .ZN(n13307) );
  AOI21_X1 U7817 ( .B1(n13339), .B2(n13338), .A(n6562), .ZN(n13333) );
  NAND2_X1 U7818 ( .A1(n13333), .A2(n13332), .ZN(n13331) );
  INV_X1 U7819 ( .A(n6840), .ZN(n11959) );
  INV_X1 U7820 ( .A(n13363), .ZN(n6845) );
  AND2_X1 U7821 ( .A1(n11932), .A2(n7250), .ZN(n7249) );
  INV_X1 U7822 ( .A(n7253), .ZN(n7250) );
  INV_X1 U7823 ( .A(n11957), .ZN(n13358) );
  NAND2_X1 U7824 ( .A1(n7244), .A2(n7251), .ZN(n7247) );
  NAND2_X1 U7825 ( .A1(n8750), .A2(n8749), .ZN(n13400) );
  NAND2_X1 U7826 ( .A1(n8762), .A2(n8761), .ZN(n12157) );
  AOI21_X1 U7827 ( .B1(n6862), .B2(n11739), .A(n6501), .ZN(n6860) );
  INV_X1 U7828 ( .A(n11740), .ZN(n6865) );
  OAI21_X1 U7829 ( .B1(n11301), .B2(n6884), .A(n6882), .ZN(n11658) );
  INV_X1 U7830 ( .A(n6885), .ZN(n6884) );
  AOI21_X1 U7831 ( .B1(n6885), .B2(n6883), .A(n6549), .ZN(n6882) );
  NOR2_X1 U7832 ( .A1(n11517), .A2(n6886), .ZN(n6885) );
  NAND2_X1 U7833 ( .A1(n8700), .A2(n8699), .ZN(n11520) );
  NAND2_X1 U7834 ( .A1(n11495), .A2(n11494), .ZN(n11497) );
  NAND2_X1 U7835 ( .A1(n11473), .A2(n11472), .ZN(n11471) );
  INV_X1 U7836 ( .A(n7226), .ZN(n7228) );
  OAI21_X1 U7837 ( .B1(n11466), .B2(n7229), .A(n11477), .ZN(n7226) );
  INV_X1 U7838 ( .A(n11271), .ZN(n7229) );
  NAND2_X1 U7839 ( .A1(n11467), .A2(n11466), .ZN(n11465) );
  OAI21_X1 U7840 ( .B1(n10701), .B2(n6850), .A(n11059), .ZN(n6846) );
  INV_X1 U7841 ( .A(n11057), .ZN(n6850) );
  NAND2_X1 U7842 ( .A1(n10702), .A2(n10701), .ZN(n11058) );
  AND2_X1 U7843 ( .A1(n8718), .A2(n8717), .ZN(n13539) );
  NAND2_X1 U7844 ( .A1(n10207), .A2(n10206), .ZN(n13541) );
  NAND2_X1 U7845 ( .A1(n8534), .A2(n8535), .ZN(n10694) );
  AOI21_X1 U7846 ( .B1(n10182), .B2(n11881), .A(n13582), .ZN(n14679) );
  AND2_X1 U7847 ( .A1(n8447), .A2(n6577), .ZN(n6872) );
  INV_X1 U7848 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9050) );
  OR2_X1 U7849 ( .A1(n9042), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n9046) );
  INV_X1 U7850 ( .A(n9051), .ZN(n9055) );
  INV_X1 U7851 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9039) );
  INV_X1 U7852 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8474) );
  INV_X1 U7853 ( .A(n8473), .ZN(n8476) );
  NAND2_X1 U7854 ( .A1(n8467), .A2(n6521), .ZN(n8799) );
  AND2_X1 U7855 ( .A1(n13657), .A2(n7093), .ZN(n7092) );
  OR2_X1 U7856 ( .A1(n13620), .A2(n7094), .ZN(n7093) );
  INV_X1 U7857 ( .A(n12123), .ZN(n7094) );
  AOI21_X1 U7858 ( .B1(n7110), .B2(n14264), .A(n6560), .ZN(n7109) );
  NAND2_X1 U7859 ( .A1(n13635), .A2(n7102), .ZN(n13609) );
  NOR2_X1 U7860 ( .A1(n13612), .A2(n7103), .ZN(n7102) );
  INV_X1 U7861 ( .A(n12093), .ZN(n7103) );
  INV_X1 U7862 ( .A(n7100), .ZN(n7099) );
  OAI21_X1 U7863 ( .B1(n13646), .B2(n7101), .A(n13593), .ZN(n7100) );
  INV_X1 U7864 ( .A(n12102), .ZN(n7101) );
  AND3_X1 U7865 ( .A1(n10288), .A2(n10287), .A3(n10286), .ZN(n10318) );
  AND2_X1 U7866 ( .A1(n7115), .A2(n7113), .ZN(n7112) );
  NOR2_X1 U7867 ( .A1(n11592), .A2(n11593), .ZN(n7113) );
  OR2_X1 U7868 ( .A1(n8116), .A2(n8115), .ZN(n8129) );
  INV_X1 U7869 ( .A(n10278), .ZN(n10289) );
  INV_X1 U7870 ( .A(n10727), .ZN(n7084) );
  NOR2_X1 U7871 ( .A1(n13861), .A2(n12006), .ZN(n6736) );
  INV_X1 U7872 ( .A(n13944), .ZN(n6739) );
  NOR2_X1 U7873 ( .A1(n13972), .A2(n6741), .ZN(n6740) );
  OR2_X1 U7874 ( .A1(n8205), .A2(n7843), .ZN(n7844) );
  NAND2_X1 U7875 ( .A1(n8374), .A2(n8373), .ZN(n8378) );
  AOI211_X1 U7876 ( .C1(n13868), .C2(n13841), .A(n13840), .B(n14492), .ZN(
        n14024) );
  OAI21_X1 U7877 ( .B1(n13836), .B2(n13854), .A(n13855), .ZN(n13853) );
  INV_X1 U7878 ( .A(n6931), .ZN(n6930) );
  OAI21_X1 U7879 ( .B1(n13873), .B2(n12018), .A(n6561), .ZN(n6931) );
  AOI21_X1 U7880 ( .B1(n6935), .B2(n13928), .A(n6558), .ZN(n6933) );
  INV_X1 U7881 ( .A(n6935), .ZN(n6934) );
  NOR2_X1 U7882 ( .A1(n13920), .A2(n13622), .ZN(n12001) );
  AND2_X1 U7883 ( .A1(n13905), .A2(n12016), .ZN(n6935) );
  NOR2_X1 U7884 ( .A1(n13906), .A2(n13905), .ZN(n13912) );
  NAND2_X1 U7885 ( .A1(n7389), .A2(n13926), .ZN(n13925) );
  AND2_X1 U7886 ( .A1(n14130), .A2(n9896), .ZN(n13947) );
  NAND2_X1 U7887 ( .A1(n8159), .A2(n8158), .ZN(n12068) );
  NAND2_X1 U7888 ( .A1(n11868), .A2(n11867), .ZN(n11870) );
  AND2_X1 U7889 ( .A1(n11796), .A2(n11795), .ZN(n7387) );
  NAND2_X1 U7890 ( .A1(n7387), .A2(n11797), .ZN(n11868) );
  NAND2_X1 U7891 ( .A1(n6818), .A2(n6817), .ZN(n11798) );
  AOI21_X1 U7892 ( .B1(n11007), .B2(n6898), .A(n6548), .ZN(n6897) );
  INV_X1 U7893 ( .A(n10906), .ZN(n6898) );
  NAND2_X1 U7894 ( .A1(n10897), .A2(n7215), .ZN(n10900) );
  NAND2_X1 U7895 ( .A1(n14402), .A2(n7214), .ZN(n10897) );
  NOR2_X1 U7896 ( .A1(n10902), .A2(n7216), .ZN(n7214) );
  INV_X1 U7897 ( .A(n10757), .ZN(n7216) );
  NAND2_X1 U7898 ( .A1(n7920), .A2(n7919), .ZN(n14431) );
  NAND2_X1 U7899 ( .A1(n10751), .A2(n14357), .ZN(n14420) );
  OR2_X1 U7900 ( .A1(n13690), .A2(n10622), .ZN(n10576) );
  INV_X1 U7901 ( .A(n14024), .ZN(n6816) );
  INV_X1 U7902 ( .A(n14023), .ZN(n6630) );
  NAND2_X1 U7903 ( .A1(n8180), .A2(n8179), .ZN(n14092) );
  AND2_X1 U7904 ( .A1(n14497), .A2(n14095), .ZN(n14517) );
  XNOR2_X1 U7905 ( .A(n8368), .B(n7792), .ZN(n12273) );
  XNOR2_X1 U7906 ( .A(n7680), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7812) );
  XNOR2_X1 U7907 ( .A(n7824), .B(n7823), .ZN(n13569) );
  NAND3_X1 U7908 ( .A1(n7677), .A2(n7212), .A3(n7384), .ZN(n7797) );
  XNOR2_X1 U7909 ( .A(n8339), .B(n8338), .ZN(n11927) );
  INV_X1 U7910 ( .A(n7797), .ZN(n6614) );
  NOR2_X1 U7911 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6613) );
  INV_X1 U7912 ( .A(n7773), .ZN(n8274) );
  XNOR2_X1 U7913 ( .A(n8244), .B(SI_22_), .ZN(n8863) );
  NAND2_X1 U7914 ( .A1(n7075), .A2(n7074), .ZN(n8243) );
  NAND2_X1 U7915 ( .A1(n7687), .A2(n7688), .ZN(n7799) );
  INV_X1 U7916 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7688) );
  AND2_X1 U7917 ( .A1(n8014), .A2(n7998), .ZN(n9968) );
  INV_X1 U7918 ( .A(n7435), .ZN(n7434) );
  NAND2_X1 U7919 ( .A1(n6944), .A2(n6947), .ZN(n7441) );
  NOR2_X1 U7920 ( .A1(n7450), .A2(n7451), .ZN(n7452) );
  NOR2_X1 U7921 ( .A1(n7400), .A2(n7401), .ZN(n7454) );
  NOR2_X1 U7922 ( .A1(n7458), .A2(n7459), .ZN(n7462) );
  AOI21_X1 U7923 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n7417), .A(n7416), .ZN(
        n7483) );
  NOR2_X1 U7924 ( .A1(n7426), .A2(n7425), .ZN(n7416) );
  AOI21_X1 U7925 ( .B1(n12761), .B2(n9594), .A(n9585), .ZN(n12773) );
  AND2_X1 U7926 ( .A1(n9468), .A2(n9467), .ZN(n12885) );
  AND3_X1 U7927 ( .A1(n9191), .A2(n9190), .A3(n9189), .ZN(n10511) );
  AND2_X1 U7928 ( .A1(n9428), .A2(n9427), .ZN(n12886) );
  NAND2_X1 U7929 ( .A1(n7182), .A2(n7180), .ZN(n12346) );
  NOR2_X1 U7930 ( .A1(n10013), .A2(n7181), .ZN(n7180) );
  NAND2_X1 U7931 ( .A1(n11294), .A2(n9727), .ZN(n7182) );
  NOR2_X1 U7932 ( .A1(n9727), .A2(SI_24_), .ZN(n7181) );
  INV_X1 U7933 ( .A(n12866), .ZN(n12899) );
  XNOR2_X1 U7934 ( .A(n6664), .B(n12740), .ZN(n12589) );
  NOR2_X1 U7935 ( .A1(n12585), .A2(n6666), .ZN(n6665) );
  NAND2_X1 U7936 ( .A1(n6683), .A2(n7004), .ZN(n6682) );
  NAND2_X1 U7937 ( .A1(n7006), .A2(n7005), .ZN(n6683) );
  NAND2_X1 U7938 ( .A1(n12591), .A2(n14979), .ZN(n7004) );
  INV_X1 U7939 ( .A(n12560), .ZN(n7005) );
  NAND2_X1 U7940 ( .A1(n9555), .A2(n9554), .ZN(n12802) );
  NAND2_X1 U7941 ( .A1(n9485), .A2(n9484), .ZN(n12872) );
  INV_X1 U7942 ( .A(n14202), .ZN(n12607) );
  OAI21_X1 U7943 ( .B1(n10009), .B2(n10028), .A(n10010), .ZN(n10011) );
  NOR2_X1 U7944 ( .A1(n10011), .A2(n10020), .ZN(n10042) );
  XNOR2_X1 U7945 ( .A(n11144), .B(n11193), .ZN(n14853) );
  XNOR2_X1 U7946 ( .A(n6914), .B(n11435), .ZN(n11150) );
  NAND2_X1 U7947 ( .A1(n11438), .A2(n11439), .ZN(n11716) );
  XNOR2_X1 U7948 ( .A(n12613), .B(n12625), .ZN(n11715) );
  XNOR2_X1 U7949 ( .A(n12666), .B(n12674), .ZN(n12643) );
  NAND2_X1 U7950 ( .A1(n12643), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12668) );
  AOI21_X1 U7951 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n12722) );
  XNOR2_X1 U7952 ( .A(n6773), .B(n12736), .ZN(n6772) );
  INV_X1 U7953 ( .A(n12737), .ZN(n6773) );
  AOI21_X1 U7954 ( .B1(n13049), .B2(n12537), .A(n12536), .ZN(n12749) );
  NAND2_X1 U7955 ( .A1(n12770), .A2(n7356), .ZN(n12755) );
  NAND2_X1 U7956 ( .A1(n9507), .A2(n9506), .ZN(n12963) );
  NAND2_X1 U7957 ( .A1(n9459), .A2(n9458), .ZN(n12976) );
  NOR2_X1 U7958 ( .A1(n7365), .A2(n15077), .ZN(n7364) );
  INV_X1 U7959 ( .A(n7365), .ZN(n7362) );
  AND2_X1 U7960 ( .A1(n7140), .A2(n9656), .ZN(n13047) );
  AND2_X1 U7961 ( .A1(n9664), .A2(n7142), .ZN(n7141) );
  XNOR2_X1 U7962 ( .A(n9604), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12595) );
  NAND2_X2 U7963 ( .A1(n10888), .A2(n10887), .ZN(n11104) );
  NAND2_X1 U7964 ( .A1(n8664), .A2(n8663), .ZN(n14736) );
  NAND2_X1 U7965 ( .A1(n8817), .A2(n8816), .ZN(n13498) );
  NAND2_X1 U7966 ( .A1(n8628), .A2(n8627), .ZN(n11484) );
  INV_X1 U7967 ( .A(n13539), .ZN(n11649) );
  NAND2_X1 U7968 ( .A1(n8802), .A2(n8801), .ZN(n13503) );
  NAND2_X1 U7969 ( .A1(n7316), .A2(n7315), .ZN(n7314) );
  NAND2_X1 U7970 ( .A1(n7314), .A2(n7311), .ZN(n13160) );
  INV_X1 U7971 ( .A(n7313), .ZN(n7311) );
  NOR2_X1 U7972 ( .A1(n13159), .A2(n7313), .ZN(n7312) );
  NAND2_X1 U7973 ( .A1(n10240), .A2(n13414), .ZN(n14240) );
  INV_X1 U7974 ( .A(n8487), .ZN(n10205) );
  NAND2_X1 U7975 ( .A1(n11121), .A2(n11120), .ZN(n11324) );
  XNOR2_X1 U7976 ( .A(n13206), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13214) );
  INV_X1 U7977 ( .A(n13411), .ZN(n13365) );
  INV_X1 U7978 ( .A(n10238), .ZN(n10239) );
  NAND2_X1 U7979 ( .A1(n6788), .A2(n6543), .ZN(n13548) );
  NAND2_X1 U7980 ( .A1(n8328), .A2(n8327), .ZN(n14033) );
  NAND2_X1 U7981 ( .A1(n8262), .A2(n8261), .ZN(n14058) );
  NAND2_X1 U7982 ( .A1(n10883), .A2(n8372), .ZN(n6725) );
  OR2_X1 U7983 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  INV_X1 U7984 ( .A(n7827), .ZN(n13665) );
  OR2_X1 U7985 ( .A1(n14441), .A2(n10559), .ZN(n13923) );
  XNOR2_X1 U7986 ( .A(n7436), .B(n6621), .ZN(n15090) );
  INV_X1 U7987 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U7988 ( .A1(n7443), .A2(n7442), .ZN(n15087) );
  XNOR2_X1 U7989 ( .A(n7462), .B(n6951), .ZN(n14146) );
  INV_X1 U7990 ( .A(n7463), .ZN(n6951) );
  AND2_X1 U7991 ( .A1(n6962), .A2(n14344), .ZN(n6958) );
  NAND2_X1 U7992 ( .A1(n6749), .A2(n6748), .ZN(n6963) );
  INV_X1 U7993 ( .A(n14340), .ZN(n6748) );
  INV_X1 U7994 ( .A(n14341), .ZN(n6749) );
  NAND2_X1 U7995 ( .A1(n6754), .A2(n14164), .ZN(n14135) );
  OAI21_X1 U7996 ( .B1(n14166), .B2(n14165), .A(n6755), .ZN(n6754) );
  INV_X1 U7997 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n6755) );
  AOI21_X1 U7998 ( .B1(n14135), .B2(n14136), .A(n14678), .ZN(n6954) );
  XNOR2_X1 U7999 ( .A(n7663), .B(n7662), .ZN(n7664) );
  NAND2_X1 U8000 ( .A1(n8536), .A2(n8538), .ZN(n7282) );
  NAND2_X1 U8001 ( .A1(n8573), .A2(n8575), .ZN(n7277) );
  NAND2_X1 U8002 ( .A1(n7290), .A2(n8615), .ZN(n7289) );
  AOI21_X1 U8003 ( .B1(n7031), .B2(n7029), .A(n7028), .ZN(n7027) );
  NAND2_X1 U8004 ( .A1(n8649), .A2(n8653), .ZN(n7285) );
  NAND2_X1 U8005 ( .A1(n8685), .A2(n8687), .ZN(n7279) );
  INV_X1 U8006 ( .A(n8803), .ZN(n7292) );
  OR2_X1 U8007 ( .A1(n7293), .A2(n8792), .ZN(n7291) );
  NOR2_X1 U8008 ( .A1(n7038), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U8009 ( .A1(n6566), .A2(n8142), .ZN(n7037) );
  NAND2_X1 U8010 ( .A1(n7040), .A2(n8198), .ZN(n7039) );
  NAND2_X1 U8011 ( .A1(n8398), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U8012 ( .A1(n7043), .A2(n6513), .ZN(n7041) );
  NAND2_X1 U8013 ( .A1(n8233), .A2(n8235), .ZN(n6637) );
  NAND2_X1 U8014 ( .A1(n7274), .A2(n7273), .ZN(n8868) );
  OR2_X1 U8015 ( .A1(n7275), .A2(n8854), .ZN(n7273) );
  NAND2_X1 U8016 ( .A1(n7024), .A2(n7023), .ZN(n7021) );
  NOR2_X1 U8017 ( .A1(n8266), .A2(n8263), .ZN(n7024) );
  NAND2_X1 U8018 ( .A1(n8263), .A2(n8266), .ZN(n7023) );
  NAND2_X1 U8019 ( .A1(n7268), .A2(n7267), .ZN(n8899) );
  NAND2_X1 U8020 ( .A1(n8886), .A2(n8888), .ZN(n7267) );
  NAND2_X1 U8021 ( .A1(n8294), .A2(n8296), .ZN(n7025) );
  NAND2_X1 U8022 ( .A1(n7271), .A2(n7270), .ZN(n8929) );
  NAND2_X1 U8023 ( .A1(n8916), .A2(n8918), .ZN(n7270) );
  NAND2_X1 U8024 ( .A1(n14687), .A2(n6526), .ZN(n9024) );
  INV_X1 U8025 ( .A(n9517), .ZN(n7174) );
  INV_X1 U8026 ( .A(n9505), .ZN(n7171) );
  INV_X1 U8027 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9324) );
  NOR2_X1 U8028 ( .A1(n13462), .A2(n13468), .ZN(n6835) );
  NAND2_X1 U8029 ( .A1(n8329), .A2(n7049), .ZN(n7048) );
  NOR2_X1 U8030 ( .A1(n8228), .A2(SI_21_), .ZN(n7761) );
  AND2_X1 U8031 ( .A1(n7688), .A2(n7107), .ZN(n7106) );
  INV_X1 U8032 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7107) );
  AOI21_X1 U8033 ( .B1(n6729), .B2(n6728), .A(n6555), .ZN(n6727) );
  INV_X1 U8034 ( .A(n7065), .ZN(n6795) );
  AOI21_X1 U8035 ( .B1(n7068), .B2(n7070), .A(n7066), .ZN(n7065) );
  INV_X1 U8036 ( .A(n7748), .ZN(n7066) );
  AND2_X1 U8037 ( .A1(n7068), .A2(n6799), .ZN(n6798) );
  NAND2_X1 U8038 ( .A1(n6800), .A2(n7741), .ZN(n6799) );
  INV_X1 U8039 ( .A(n7386), .ZN(n6800) );
  NAND2_X1 U8040 ( .A1(n7742), .A2(n9798), .ZN(n7071) );
  NAND2_X1 U8041 ( .A1(n8071), .A2(SI_13_), .ZN(n7072) );
  INV_X1 U8042 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7693) );
  OR2_X1 U8043 ( .A1(n12362), .A2(n6527), .ZN(n7148) );
  NAND2_X1 U8044 ( .A1(n14845), .A2(n11158), .ZN(n11159) );
  NAND2_X1 U8045 ( .A1(n12707), .A2(n12708), .ZN(n12710) );
  NOR2_X1 U8046 ( .A1(n12797), .A2(n12811), .ZN(n7343) );
  INV_X1 U8047 ( .A(n9531), .ZN(n7345) );
  AND2_X1 U8048 ( .A1(n12811), .A2(n12812), .ZN(n12508) );
  NAND2_X1 U8049 ( .A1(n9479), .A2(n9478), .ZN(n9494) );
  INV_X1 U8050 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9460) );
  AND2_X1 U8051 ( .A1(n9461), .A2(n9460), .ZN(n9479) );
  NOR2_X1 U8052 ( .A1(n9367), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9388) );
  NOR2_X1 U8053 ( .A1(n7003), .A2(n7002), .ZN(n7001) );
  AND2_X1 U8054 ( .A1(n9628), .A2(n12437), .ZN(n7002) );
  INV_X1 U8055 ( .A(n14205), .ZN(n7003) );
  INV_X1 U8056 ( .A(n12442), .ZN(n6998) );
  NOR2_X1 U8057 ( .A1(n11261), .A2(n14936), .ZN(n7349) );
  INV_X1 U8058 ( .A(n9285), .ZN(n7352) );
  AND2_X1 U8059 ( .A1(n11261), .A2(n14936), .ZN(n7351) );
  NOR2_X1 U8060 ( .A1(n7348), .A2(n7349), .ZN(n7347) );
  AND2_X1 U8061 ( .A1(n9248), .A2(n9230), .ZN(n7371) );
  INV_X1 U8062 ( .A(n12569), .ZN(n9248) );
  NOR2_X1 U8063 ( .A1(n12565), .A2(n6982), .ZN(n6981) );
  INV_X1 U8064 ( .A(n12414), .ZN(n6982) );
  INV_X1 U8065 ( .A(n12422), .ZN(n6978) );
  OR2_X1 U8066 ( .A1(n9369), .A2(n11173), .ZN(n9160) );
  NAND2_X1 U8067 ( .A1(n12392), .A2(n12399), .ZN(n6969) );
  NAND2_X1 U8068 ( .A1(n12399), .A2(n12391), .ZN(n12392) );
  INV_X1 U8069 ( .A(n12393), .ZN(n10791) );
  AND2_X1 U8070 ( .A1(n10725), .A2(n12740), .ZN(n9694) );
  OR2_X1 U8071 ( .A1(n9658), .A2(n9678), .ZN(n9698) );
  INV_X1 U8072 ( .A(n7153), .ZN(n7152) );
  OAI21_X1 U8073 ( .B1(n9379), .B2(n7154), .A(n9412), .ZN(n7153) );
  INV_X1 U8074 ( .A(n9395), .ZN(n7154) );
  INV_X1 U8075 ( .A(n9414), .ZN(n7151) );
  NAND2_X1 U8076 ( .A1(n6677), .A2(n6675), .ZN(n6674) );
  INV_X1 U8077 ( .A(n9376), .ZN(n6675) );
  INV_X1 U8078 ( .A(n11417), .ZN(n7307) );
  NOR2_X1 U8079 ( .A1(n13151), .A2(n7325), .ZN(n7324) );
  INV_X1 U8080 ( .A(n12169), .ZN(n7325) );
  AND2_X1 U8081 ( .A1(n8688), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8704) );
  AND2_X1 U8082 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n8856), .ZN(n8874) );
  NOR2_X1 U8083 ( .A1(n8674), .A2(n11107), .ZN(n8688) );
  NOR2_X1 U8084 ( .A1(n8768), .A2(n8751), .ZN(n8740) );
  NAND2_X1 U8085 ( .A1(n8982), .A2(n6554), .ZN(n7258) );
  NAND2_X1 U8086 ( .A1(n7265), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U8087 ( .A1(n7261), .A2(n7260), .ZN(n7259) );
  INV_X1 U8088 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7340) );
  OR2_X1 U8089 ( .A1(n13311), .A2(n13177), .ZN(n7380) );
  AND2_X1 U8090 ( .A1(n6496), .A2(n11964), .ZN(n6874) );
  NOR2_X1 U8091 ( .A1(n6547), .A2(n7248), .ZN(n7245) );
  NAND2_X1 U8092 ( .A1(n13387), .A2(n7249), .ZN(n7242) );
  NAND2_X1 U8093 ( .A1(n13358), .A2(n6842), .ZN(n6841) );
  NAND2_X1 U8094 ( .A1(n6843), .A2(n6845), .ZN(n6842) );
  NAND2_X1 U8095 ( .A1(n6838), .A2(n13371), .ZN(n13351) );
  INV_X1 U8096 ( .A(n11303), .ZN(n6886) );
  INV_X1 U8097 ( .A(n11300), .ZN(n6883) );
  OR2_X1 U8098 ( .A1(n11494), .A2(n7240), .ZN(n7239) );
  NAND2_X1 U8099 ( .A1(n11302), .A2(n13189), .ZN(n7241) );
  NOR2_X1 U8100 ( .A1(n14736), .A2(n14727), .ZN(n6826) );
  NOR2_X1 U8101 ( .A1(n8618), .A2(n8617), .ZN(n8635) );
  AND2_X1 U8102 ( .A1(n8576), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U8103 ( .A1(n6809), .A2(n6890), .ZN(n6889) );
  AND2_X1 U8104 ( .A1(n6810), .A2(n6568), .ZN(n6888) );
  NOR2_X1 U8105 ( .A1(n13174), .A2(n13274), .ZN(n11938) );
  NAND2_X1 U8106 ( .A1(n13325), .A2(n6835), .ZN(n13301) );
  NAND2_X1 U8107 ( .A1(n13325), .A2(n13311), .ZN(n13310) );
  NAND2_X1 U8108 ( .A1(n11339), .A2(n11340), .ZN(n11498) );
  NAND2_X1 U8109 ( .A1(n11349), .A2(n11348), .ZN(n11347) );
  INV_X1 U8110 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8448) );
  INV_X1 U8111 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7332) );
  OR2_X1 U8112 ( .A1(n8661), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8681) );
  OR2_X1 U8113 ( .A1(n8569), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8586) );
  OAI22_X1 U8114 ( .A1(n14443), .A2(n10731), .B1(n10732), .B2(n12139), .ZN(
        n10734) );
  OR2_X1 U8115 ( .A1(n13926), .A2(n6742), .ZN(n6741) );
  NAND2_X1 U8116 ( .A1(n8398), .A2(n6743), .ZN(n6742) );
  NOR2_X1 U8117 ( .A1(n8411), .A2(n11667), .ZN(n6743) );
  INV_X1 U8118 ( .A(n10468), .ZN(n10281) );
  NAND2_X1 U8119 ( .A1(n14077), .A2(n6815), .ZN(n6814) );
  INV_X1 U8120 ( .A(n7193), .ZN(n7189) );
  AOI21_X1 U8121 ( .B1(n7193), .B2(n7192), .A(n6550), .ZN(n7191) );
  INV_X1 U8122 ( .A(n7195), .ZN(n7192) );
  AND2_X1 U8123 ( .A1(n14388), .A2(n10896), .ZN(n7215) );
  OR2_X1 U8124 ( .A1(n7988), .A2(n7814), .ZN(n8004) );
  AND2_X1 U8125 ( .A1(n10755), .A2(n8399), .ZN(n10596) );
  INV_X1 U8126 ( .A(n10631), .ZN(n10579) );
  INV_X1 U8127 ( .A(n13666), .ZN(n13621) );
  CLKBUF_X1 U8128 ( .A(n10285), .Z(n6620) );
  AOI21_X1 U8129 ( .B1(n10327), .B2(n10264), .A(n10263), .ZN(n10555) );
  NAND2_X1 U8130 ( .A1(n7055), .A2(n7054), .ZN(n8326) );
  NAND2_X1 U8131 ( .A1(n6602), .A2(n6508), .ZN(n7054) );
  NAND2_X1 U8132 ( .A1(n7766), .A2(n7765), .ZN(n7768) );
  OAI21_X1 U8133 ( .B1(n7754), .B2(n7073), .A(n6802), .ZN(n7766) );
  OR2_X1 U8134 ( .A1(n8174), .A2(n6803), .ZN(n7754) );
  INV_X1 U8135 ( .A(n8173), .ZN(n6803) );
  XNOR2_X1 U8136 ( .A(n7752), .B(SI_18_), .ZN(n8174) );
  NAND2_X1 U8137 ( .A1(n6797), .A2(n7741), .ZN(n8073) );
  OR2_X1 U8138 ( .A1(n7972), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7996) );
  OR2_X1 U8139 ( .A1(n7953), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U8140 ( .A1(n6738), .A2(n7050), .ZN(n7936) );
  NAND2_X1 U8141 ( .A1(n6946), .A2(n7395), .ZN(n6945) );
  INV_X1 U8142 ( .A(n7393), .ZN(n6946) );
  INV_X1 U8143 ( .A(n6746), .ZN(n7399) );
  OAI21_X1 U8144 ( .B1(n7430), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6502), .ZN(
        n6746) );
  XNOR2_X1 U8145 ( .A(n7399), .B(n6938), .ZN(n7447) );
  INV_X1 U8146 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7402) );
  AND2_X1 U8147 ( .A1(n6752), .A2(n6751), .ZN(n7403) );
  NAND2_X1 U8148 ( .A1(n7402), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6751) );
  OR2_X1 U8149 ( .A1(n7454), .A2(n7453), .ZN(n6752) );
  NOR2_X1 U8150 ( .A1(n7410), .A2(n7409), .ZN(n7470) );
  AOI21_X1 U8151 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n7412), .A(n7411), .ZN(
        n7476) );
  NOR2_X1 U8152 ( .A1(n7470), .A2(n7469), .ZN(n7411) );
  OR2_X1 U8153 ( .A1(n9347), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U8154 ( .A1(n7148), .A2(n7146), .ZN(n7144) );
  NAND2_X1 U8155 ( .A1(n7147), .A2(n12910), .ZN(n7146) );
  INV_X1 U8156 ( .A(n12329), .ZN(n7147) );
  CLKBUF_X1 U8157 ( .A(n9621), .Z(n10094) );
  AND2_X1 U8158 ( .A1(n6709), .A2(n6702), .ZN(n6701) );
  NAND2_X1 U8159 ( .A1(n7122), .A2(n6491), .ZN(n6709) );
  NAND2_X1 U8160 ( .A1(n6704), .A2(n6703), .ZN(n6702) );
  AND2_X1 U8161 ( .A1(n12258), .A2(n12256), .ZN(n12318) );
  AND2_X1 U8162 ( .A1(n10310), .A2(n10307), .ZN(n10308) );
  AND2_X1 U8163 ( .A1(n12317), .A2(n12252), .ZN(n12336) );
  NOR2_X1 U8164 ( .A1(n9508), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U8165 ( .A1(n9523), .A2(n12341), .ZN(n9537) );
  INV_X1 U8166 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U8167 ( .A1(n6975), .A2(n10344), .ZN(n12389) );
  NAND2_X1 U8168 ( .A1(n7144), .A2(n6720), .ZN(n6719) );
  NAND2_X1 U8169 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  OR2_X1 U8170 ( .A1(n12243), .A2(n12242), .ZN(n7169) );
  NOR2_X1 U8171 ( .A1(n7134), .A2(n12612), .ZN(n10100) );
  NOR2_X1 U8172 ( .A1(n12328), .A2(n12329), .ZN(n12327) );
  OR2_X1 U8173 ( .A1(n9422), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9442) );
  INV_X1 U8174 ( .A(n7374), .ZN(n6700) );
  NAND2_X1 U8175 ( .A1(n6696), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8176 ( .A1(n12584), .A2(n6667), .ZN(n6666) );
  AND2_X1 U8177 ( .A1(n12753), .A2(n6668), .ZN(n6667) );
  AND2_X1 U8178 ( .A1(n12583), .A2(n12769), .ZN(n6668) );
  NAND2_X1 U8179 ( .A1(n12997), .A2(n12746), .ZN(n6669) );
  NOR2_X1 U8180 ( .A1(n10030), .A2(n10031), .ZN(n10057) );
  NOR2_X1 U8181 ( .A1(n10057), .A2(n10058), .ZN(n10059) );
  NAND2_X1 U8182 ( .A1(n11153), .A2(n6515), .ZN(n14812) );
  NAND2_X1 U8183 ( .A1(n14827), .A2(n11157), .ZN(n14847) );
  NAND2_X1 U8184 ( .A1(n14847), .A2(n14846), .ZN(n14845) );
  XNOR2_X1 U8185 ( .A(n11159), .B(n11193), .ZN(n14863) );
  INV_X1 U8186 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12299) );
  NAND2_X1 U8187 ( .A1(n11716), .A2(n6599), .ZN(n12616) );
  NOR2_X1 U8188 ( .A1(n12695), .A2(n6903), .ZN(n12696) );
  NOR2_X1 U8189 ( .A1(n12682), .A2(n6904), .ZN(n6903) );
  XNOR2_X1 U8190 ( .A(n12710), .B(n14173), .ZN(n14172) );
  OR2_X1 U8191 ( .A1(n14169), .A2(n14170), .ZN(n12701) );
  NAND2_X1 U8192 ( .A1(n14172), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14171) );
  AOI21_X1 U8193 ( .B1(n14171), .B2(n12712), .A(n12711), .ZN(n12733) );
  AND2_X1 U8194 ( .A1(n12531), .A2(n12550), .ZN(n12584) );
  OR2_X1 U8195 ( .A1(n9582), .A2(n12744), .ZN(n12761) );
  AND2_X1 U8196 ( .A1(n12521), .A2(n12387), .ZN(n12753) );
  AND2_X1 U8197 ( .A1(n9572), .A2(n9571), .ZN(n12786) );
  NAND2_X1 U8198 ( .A1(n12810), .A2(n12388), .ZN(n12798) );
  NAND2_X1 U8199 ( .A1(n12961), .A2(n12508), .ZN(n12810) );
  AND2_X1 U8200 ( .A1(n9388), .A2(n11760), .ZN(n9404) );
  INV_X1 U8201 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9403) );
  AOI21_X1 U8202 ( .B1(n12923), .B2(n6995), .A(n6994), .ZN(n6993) );
  INV_X1 U8203 ( .A(n12467), .ZN(n6995) );
  INV_X1 U8204 ( .A(n9631), .ZN(n12912) );
  OR2_X1 U8205 ( .A1(n9279), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9286) );
  OR2_X1 U8206 ( .A1(n9286), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9306) );
  OAI21_X1 U8207 ( .B1(n11244), .B2(n9626), .A(n9627), .ZN(n14931) );
  NAND2_X1 U8208 ( .A1(n9262), .A2(n10952), .ZN(n9279) );
  AND2_X1 U8209 ( .A1(n9231), .A2(n12299), .ZN(n9262) );
  AND2_X1 U8210 ( .A1(n12429), .A2(n12428), .ZN(n12569) );
  NAND2_X1 U8211 ( .A1(n14946), .A2(n9230), .ZN(n11089) );
  NOR2_X1 U8212 ( .A1(n9211), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9231) );
  INV_X1 U8213 ( .A(n14947), .ZN(n14944) );
  AND2_X1 U8214 ( .A1(n10933), .A2(n9193), .ZN(n7369) );
  AND2_X1 U8215 ( .A1(n10793), .A2(n9193), .ZN(n10934) );
  OR2_X1 U8216 ( .A1(n9194), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9211) );
  CLKBUF_X1 U8217 ( .A(n10792), .Z(n10793) );
  NOR2_X1 U8218 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9175) );
  NAND2_X1 U8219 ( .A1(n14976), .A2(n12399), .ZN(n14961) );
  NAND2_X1 U8220 ( .A1(n6970), .A2(n14982), .ZN(n14976) );
  AOI21_X1 U8221 ( .B1(n12538), .B2(P3_REG1_REG_0__SCAN_IN), .A(n9108), .ZN(
        n9112) );
  NOR2_X1 U8222 ( .A1(n9139), .A2(n10342), .ZN(n9108) );
  NAND2_X1 U8223 ( .A1(n9563), .A2(n9562), .ZN(n12778) );
  NAND2_X1 U8224 ( .A1(n9550), .A2(n9549), .ZN(n12791) );
  NAND2_X1 U8225 ( .A1(n9536), .A2(n9535), .ZN(n12315) );
  INV_X1 U8226 ( .A(n15047), .ZN(n15015) );
  NAND2_X1 U8227 ( .A1(n6659), .A2(n6610), .ZN(n6658) );
  OAI22_X1 U8228 ( .A1(n6661), .A2(n6658), .B1(n14117), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8229 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n6660), .ZN(n6659) );
  NOR2_X1 U8230 ( .A1(n12224), .A2(n6662), .ZN(n6661) );
  INV_X1 U8231 ( .A(n9590), .ZN(n6662) );
  INV_X1 U8232 ( .A(n6989), .ZN(n6987) );
  NAND2_X1 U8233 ( .A1(n9547), .A2(n9546), .ZN(n9558) );
  NAND2_X1 U8234 ( .A1(n9545), .A2(n9544), .ZN(n9547) );
  XNOR2_X1 U8235 ( .A(n9663), .B(n9662), .ZN(n10079) );
  INV_X1 U8236 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9662) );
  OAI21_X1 U8237 ( .B1(n9661), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9663) );
  NOR2_X1 U8238 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n6721) );
  NAND2_X1 U8239 ( .A1(n7161), .A2(n7165), .ZN(n9473) );
  AND2_X1 U8240 ( .A1(n9489), .A2(n9471), .ZN(n9472) );
  NAND2_X1 U8241 ( .A1(n9603), .A2(n9602), .ZN(n9608) );
  NAND2_X1 U8242 ( .A1(n9432), .A2(n9431), .ZN(n9435) );
  AND2_X1 U8243 ( .A1(n9453), .A2(n9433), .ZN(n9434) );
  NAND2_X1 U8244 ( .A1(n9435), .A2(n9434), .ZN(n9454) );
  OAI21_X1 U8245 ( .B1(n9356), .B2(n9355), .A(n9357), .ZN(n9360) );
  AND2_X1 U8246 ( .A1(n10614), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U8247 ( .A1(n6680), .A2(n6679), .ZN(n9377) );
  INV_X1 U8248 ( .A(n9359), .ZN(n6679) );
  INV_X1 U8249 ( .A(n9360), .ZN(n6680) );
  NAND2_X1 U8250 ( .A1(n7156), .A2(n7155), .ZN(n9323) );
  AOI21_X1 U8251 ( .B1(n7157), .B2(n7159), .A(n6595), .ZN(n7155) );
  NAND2_X1 U8252 ( .A1(n9251), .A2(n9250), .ZN(n9254) );
  AND2_X1 U8253 ( .A1(n9269), .A2(n9252), .ZN(n9253) );
  NAND2_X1 U8254 ( .A1(n9254), .A2(n9253), .ZN(n9270) );
  OR2_X1 U8255 ( .A1(n9258), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9383) );
  INV_X1 U8256 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9200) );
  AND2_X1 U8257 ( .A1(n9205), .A2(n9186), .ZN(n9203) );
  XNOR2_X1 U8258 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9127) );
  NAND2_X1 U8259 ( .A1(n13109), .A2(n7324), .ZN(n7323) );
  INV_X1 U8260 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8617) );
  AND2_X1 U8261 ( .A1(n8874), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U8262 ( .A1(n8889), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U8263 ( .A1(n7327), .A2(n7326), .ZN(n10888) );
  AND2_X1 U8264 ( .A1(n10874), .A2(n10873), .ZN(n7326) );
  NAND2_X1 U8265 ( .A1(n10872), .A2(n10871), .ZN(n7327) );
  NOR2_X1 U8266 ( .A1(n8805), .A2(n13078), .ZN(n8826) );
  NAND2_X1 U8267 ( .A1(n8704), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8722) );
  OR2_X1 U8268 ( .A1(n8795), .A2(n8794), .ZN(n8805) );
  NAND2_X1 U8269 ( .A1(n13110), .A2(n13111), .ZN(n13109) );
  AND2_X1 U8270 ( .A1(n10205), .A2(n10181), .ZN(n10228) );
  OR2_X1 U8271 ( .A1(n8766), .A2(n11855), .ZN(n8768) );
  NAND2_X1 U8272 ( .A1(n9043), .A2(n9046), .ZN(n9768) );
  INV_X1 U8273 ( .A(n8526), .ZN(n8986) );
  NOR2_X1 U8274 ( .A1(n14604), .A2(n14603), .ZN(n14602) );
  NOR2_X1 U8275 ( .A1(n14621), .A2(n14620), .ZN(n14619) );
  AOI21_X1 U8276 ( .B1(n9859), .B2(n9812), .A(n9811), .ZN(n9833) );
  AOI21_X1 U8277 ( .B1(n14632), .B2(n9852), .A(n9851), .ZN(n9875) );
  AND2_X1 U8278 ( .A1(n8467), .A2(n8464), .ZN(n8775) );
  NAND2_X1 U8279 ( .A1(n11116), .A2(n14647), .ZN(n11117) );
  INV_X1 U8280 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13078) );
  NAND2_X1 U8281 ( .A1(n8992), .A2(n8991), .ZN(n9033) );
  NOR2_X1 U8282 ( .A1(n13442), .A2(n13268), .ZN(n13255) );
  NAND2_X1 U8283 ( .A1(n13325), .A2(n6831), .ZN(n13268) );
  NOR2_X1 U8284 ( .A1(n13274), .A2(n6832), .ZN(n6831) );
  INV_X1 U8285 ( .A(n6833), .ZN(n6832) );
  NAND2_X1 U8286 ( .A1(n8865), .A2(n8864), .ZN(n13474) );
  NAND2_X1 U8287 ( .A1(n6837), .A2(n6836), .ZN(n13341) );
  INV_X1 U8288 ( .A(n6837), .ZN(n13352) );
  NAND2_X1 U8289 ( .A1(n8834), .A2(n8833), .ZN(n12181) );
  NOR2_X1 U8290 ( .A1(n13503), .A2(n13182), .ZN(n7253) );
  INV_X1 U8291 ( .A(n7247), .ZN(n13385) );
  OR2_X1 U8292 ( .A1(n13395), .A2(n13400), .ZN(n13396) );
  OR2_X1 U8293 ( .A1(n11784), .A2(n12157), .ZN(n13395) );
  AND2_X1 U8294 ( .A1(n11653), .A2(n13532), .ZN(n11743) );
  NAND2_X1 U8295 ( .A1(n11743), .A2(n13523), .ZN(n11784) );
  NAND2_X1 U8296 ( .A1(n7231), .A2(n7230), .ZN(n11780) );
  NAND2_X1 U8297 ( .A1(n13532), .A2(n11846), .ZN(n7230) );
  NAND2_X1 U8298 ( .A1(n6789), .A2(n6499), .ZN(n7231) );
  AND2_X1 U8299 ( .A1(n11523), .A2(n13539), .ZN(n11653) );
  NOR2_X1 U8300 ( .A1(n6822), .A2(n11520), .ZN(n6821) );
  INV_X1 U8301 ( .A(n6824), .ZN(n6822) );
  NAND2_X1 U8302 ( .A1(n11339), .A2(n6824), .ZN(n11307) );
  AOI21_X1 U8303 ( .B1(n6869), .B2(n6871), .A(n6538), .ZN(n6868) );
  NAND2_X1 U8304 ( .A1(n7225), .A2(n7227), .ZN(n11332) );
  AOI21_X1 U8305 ( .B1(n11477), .B2(n7229), .A(n6539), .ZN(n7227) );
  NAND2_X1 U8306 ( .A1(n11332), .A2(n11333), .ZN(n11331) );
  OR2_X1 U8307 ( .A1(n11484), .A2(n11459), .ZN(n11479) );
  AOI21_X1 U8308 ( .B1(n6849), .B2(n6850), .A(n6524), .ZN(n6847) );
  NAND2_X1 U8309 ( .A1(n10702), .A2(n6849), .ZN(n6848) );
  NAND2_X1 U8310 ( .A1(n6492), .A2(n10697), .ZN(n6779) );
  NAND2_X1 U8311 ( .A1(n10984), .A2(n10697), .ZN(n11054) );
  NAND2_X1 U8312 ( .A1(n10982), .A2(n10981), .ZN(n10984) );
  NAND2_X1 U8313 ( .A1(n11357), .A2(n11358), .ZN(n6839) );
  OR2_X1 U8314 ( .A1(n10198), .A2(n6774), .ZN(n10656) );
  OR2_X1 U8315 ( .A1(n10222), .A2(n14685), .ZN(n10822) );
  NAND2_X1 U8316 ( .A1(n11976), .A2(n13541), .ZN(n6852) );
  NAND2_X1 U8317 ( .A1(n13432), .A2(n14735), .ZN(n6830) );
  NAND2_X1 U8318 ( .A1(n6879), .A2(n6878), .ZN(n13315) );
  NAND2_X1 U8319 ( .A1(n13337), .A2(n6496), .ZN(n6879) );
  NAND2_X1 U8320 ( .A1(n6887), .A2(n11303), .ZN(n11518) );
  NAND2_X1 U8321 ( .A1(n11301), .A2(n11300), .ZN(n6887) );
  INV_X1 U8322 ( .A(n14735), .ZN(n14749) );
  AND2_X1 U8323 ( .A1(n8504), .A2(n7381), .ZN(n8505) );
  AND2_X1 U8324 ( .A1(n8447), .A2(n7286), .ZN(n7232) );
  NAND2_X1 U8325 ( .A1(n8467), .A2(n7334), .ZN(n8746) );
  OR2_X1 U8326 ( .A1(n8625), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8644) );
  INV_X1 U8327 ( .A(n8236), .ZN(n8255) );
  NAND2_X1 U8328 ( .A1(n8255), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U8329 ( .A1(n6646), .A2(n6645), .ZN(n6644) );
  INV_X1 U8330 ( .A(n11384), .ZN(n6645) );
  INV_X1 U8331 ( .A(n11383), .ZN(n6646) );
  OR2_X1 U8332 ( .A1(n7945), .A2(n7944), .ZN(n7988) );
  NAND2_X1 U8333 ( .A1(n10282), .A2(n10281), .ZN(n10733) );
  INV_X1 U8334 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8048) );
  NOR2_X1 U8335 ( .A1(n8129), .A2(n8128), .ZN(n8160) );
  INV_X1 U8336 ( .A(n8254), .ZN(n8268) );
  INV_X1 U8337 ( .A(n10807), .ZN(n10731) );
  OR2_X1 U8338 ( .A1(n11398), .A2(n11394), .ZN(n7115) );
  OR2_X1 U8339 ( .A1(n11558), .A2(n11557), .ZN(n7116) );
  NOR2_X1 U8340 ( .A1(n8199), .A2(n13639), .ZN(n8217) );
  NAND2_X1 U8341 ( .A1(n7108), .A2(n6529), .ZN(n13602) );
  OR2_X1 U8342 ( .A1(n8049), .A2(n8048), .ZN(n8064) );
  INV_X1 U8343 ( .A(n8216), .ZN(n8237) );
  NAND2_X1 U8344 ( .A1(n8237), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U8345 ( .A1(n13645), .A2(n13646), .ZN(n13644) );
  NOR2_X1 U8346 ( .A1(n8004), .A2(n9980), .ZN(n8025) );
  INV_X1 U8347 ( .A(n13678), .ZN(n11699) );
  OAI22_X1 U8348 ( .A1(n6474), .A2(n10623), .B1(n10285), .B2(n12139), .ZN(
        n10367) );
  OR2_X1 U8349 ( .A1(n10852), .A2(n10851), .ZN(n7085) );
  NAND2_X1 U8350 ( .A1(n12051), .A2(n12050), .ZN(n12054) );
  NAND2_X1 U8351 ( .A1(n8361), .A2(n8360), .ZN(n6635) );
  AND3_X1 U8352 ( .A1(n8122), .A2(n8121), .A3(n8120), .ZN(n12055) );
  INV_X1 U8353 ( .A(n13846), .ZN(n13831) );
  AOI21_X1 U8354 ( .B1(n13890), .B2(n6493), .A(n6927), .ZN(n13862) );
  INV_X1 U8355 ( .A(n6928), .ZN(n6927) );
  AOI21_X1 U8356 ( .B1(n6493), .B2(n13873), .A(n6932), .ZN(n6928) );
  NOR2_X1 U8357 ( .A1(n14033), .A2(n13834), .ZN(n6932) );
  NAND2_X1 U8358 ( .A1(n13881), .A2(n12019), .ZN(n13882) );
  NAND2_X1 U8359 ( .A1(n6518), .A2(n7205), .ZN(n7204) );
  NAND2_X1 U8360 ( .A1(n7206), .A2(n6518), .ZN(n7203) );
  NAND2_X1 U8361 ( .A1(n13946), .A2(n13938), .ZN(n13932) );
  INV_X1 U8362 ( .A(n7197), .ZN(n7196) );
  NOR2_X1 U8363 ( .A1(n13985), .A2(n14085), .ZN(n13984) );
  AOI21_X1 U8364 ( .B1(n7209), .B2(n11861), .A(n6551), .ZN(n7208) );
  NOR2_X1 U8365 ( .A1(n11615), .A2(n6923), .ZN(n6922) );
  INV_X1 U8366 ( .A(n11605), .ZN(n6923) );
  NAND2_X1 U8367 ( .A1(n8059), .A2(n8058), .ZN(n11701) );
  OR2_X1 U8368 ( .A1(n11591), .A2(n11589), .ZN(n7195) );
  NOR2_X1 U8369 ( .A1(n7185), .A2(n7186), .ZN(n7184) );
  INV_X1 U8370 ( .A(n10585), .ZN(n7186) );
  INV_X1 U8371 ( .A(n14356), .ZN(n14003) );
  NAND2_X1 U8372 ( .A1(n10584), .A2(n10585), .ZN(n7187) );
  OR2_X1 U8373 ( .A1(n10295), .A2(n10294), .ZN(n14356) );
  INV_X1 U8374 ( .A(n13658), .ZN(n14353) );
  AOI22_X1 U8375 ( .A1(n7862), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n10357), .B2(
        n8177), .ZN(n7019) );
  NOR2_X2 U8376 ( .A1(n10570), .A2(n10275), .ZN(n14549) );
  INV_X1 U8377 ( .A(n14517), .ZN(n14574) );
  NAND2_X1 U8378 ( .A1(n7057), .A2(n7780), .ZN(n8306) );
  NAND2_X1 U8379 ( .A1(n7776), .A2(n7058), .ZN(n7057) );
  XNOR2_X1 U8380 ( .A(n7768), .B(n7769), .ZN(n8260) );
  XNOR2_X1 U8381 ( .A(n8422), .B(n8421), .ZN(n9894) );
  INV_X1 U8382 ( .A(n8362), .ZN(n8363) );
  XNOR2_X1 U8383 ( .A(n8230), .B(n8229), .ZN(n11509) );
  XNOR2_X1 U8384 ( .A(n6726), .B(n8164), .ZN(n10883) );
  NAND2_X1 U8385 ( .A1(n7754), .A2(n7753), .ZN(n6726) );
  NAND2_X1 U8386 ( .A1(n6732), .A2(n7750), .ZN(n8150) );
  NAND2_X1 U8387 ( .A1(n8134), .A2(n8133), .ZN(n6732) );
  OR2_X1 U8388 ( .A1(n8056), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8057) );
  OR2_X1 U8389 ( .A1(n7913), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7915) );
  XNOR2_X1 U8390 ( .A(n7912), .B(n7911), .ZN(n9755) );
  AND2_X1 U8391 ( .A1(n7052), .A2(n7050), .ZN(n7912) );
  XNOR2_X1 U8392 ( .A(n7872), .B(n7871), .ZN(n9737) );
  NOR2_X2 U8393 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7863) );
  INV_X4 U8394 ( .A(n7798), .ZN(n9733) );
  XNOR2_X1 U8395 ( .A(n7447), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U8396 ( .A1(n6948), .A2(n7455), .ZN(n7457) );
  NAND2_X1 U8397 ( .A1(n14145), .A2(n14144), .ZN(n6948) );
  XNOR2_X1 U8398 ( .A(n7403), .B(n6750), .ZN(n7456) );
  AND2_X1 U8399 ( .A1(n6759), .A2(n6758), .ZN(n7466) );
  NAND2_X1 U8400 ( .A1(n7406), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n6758) );
  OR2_X1 U8401 ( .A1(n7461), .A2(n7460), .ZN(n6759) );
  AOI21_X1 U8402 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n7414), .A(n7413), .ZN(
        n7427) );
  NOR2_X1 U8403 ( .A1(n7476), .A2(n7475), .ZN(n7413) );
  NAND2_X1 U8404 ( .A1(n6961), .A2(n14345), .ZN(n6960) );
  INV_X1 U8405 ( .A(n14344), .ZN(n6961) );
  NAND2_X1 U8406 ( .A1(n14344), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6959) );
  AND4_X1 U8407 ( .A1(n9236), .A2(n9235), .A3(n9234), .A4(n9233), .ZN(n10946)
         );
  NAND2_X1 U8408 ( .A1(n12275), .A2(n12276), .ZN(n12274) );
  NAND2_X1 U8409 ( .A1(n12374), .A2(n12261), .ZN(n12275) );
  INV_X1 U8410 ( .A(n12283), .ZN(n12338) );
  NAND2_X1 U8411 ( .A1(n11076), .A2(n11075), .ZN(n11257) );
  NAND2_X1 U8412 ( .A1(n10308), .A2(n10309), .ZN(n10397) );
  INV_X1 U8413 ( .A(n6714), .ZN(n12290) );
  OAI21_X1 U8414 ( .B1(n12328), .B2(n6716), .A(n6715), .ZN(n6714) );
  INV_X1 U8415 ( .A(n7144), .ZN(n6716) );
  INV_X1 U8416 ( .A(n7143), .ZN(n6715) );
  NAND2_X1 U8417 ( .A1(n7131), .A2(n7128), .ZN(n7127) );
  NAND2_X1 U8418 ( .A1(n7130), .A2(n7129), .ZN(n7128) );
  AND2_X1 U8419 ( .A1(n12355), .A2(n6975), .ZN(n6974) );
  OR2_X1 U8420 ( .A1(n12237), .A2(n12885), .ZN(n12238) );
  NAND2_X1 U8421 ( .A1(n9477), .A2(n9476), .ZN(n12860) );
  NAND2_X1 U8422 ( .A1(n9386), .A2(n9385), .ZN(n12925) );
  INV_X1 U8423 ( .A(n6698), .ZN(n10684) );
  AND3_X1 U8424 ( .A1(n9172), .A2(n9171), .A3(n9170), .ZN(n10919) );
  AND2_X1 U8425 ( .A1(n10397), .A2(n7167), .ZN(n10507) );
  NAND2_X1 U8426 ( .A1(n10397), .A2(n10396), .ZN(n10400) );
  AND2_X1 U8427 ( .A1(n6708), .A2(n6710), .ZN(n10949) );
  OAI21_X1 U8428 ( .B1(n12328), .B2(n6719), .A(n6717), .ZN(n12348) );
  NAND2_X1 U8429 ( .A1(n9331), .A2(n9330), .ZN(n14193) );
  NAND2_X1 U8430 ( .A1(n7169), .A2(n12244), .ZN(n12354) );
  NAND2_X1 U8431 ( .A1(n9493), .A2(n9492), .ZN(n12849) );
  NAND2_X1 U8432 ( .A1(n11257), .A2(n11256), .ZN(n11534) );
  NOR2_X1 U8433 ( .A1(n10684), .A2(n7374), .ZN(n10687) );
  NAND2_X1 U8434 ( .A1(n6698), .A2(n6699), .ZN(n10835) );
  AND2_X1 U8435 ( .A1(n9543), .A2(n9542), .ZN(n12821) );
  INV_X1 U8436 ( .A(n12371), .ZN(n12376) );
  NAND2_X1 U8437 ( .A1(n10088), .A2(n10087), .ZN(n12383) );
  INV_X1 U8438 ( .A(n12786), .ZN(n12758) );
  INV_X1 U8439 ( .A(n12885), .ZN(n12601) );
  INV_X1 U8440 ( .A(n12921), .ZN(n12604) );
  INV_X1 U8441 ( .A(n10946), .ZN(n14950) );
  CLKBUF_X1 U8442 ( .A(n10096), .Z(n12612) );
  INV_X1 U8443 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14780) );
  CLKBUF_X1 U8444 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n14772) );
  OR2_X1 U8445 ( .A1(n10042), .A2(n10041), .ZN(n10043) );
  AND2_X1 U8446 ( .A1(n14784), .A2(n11139), .ZN(n14800) );
  INV_X1 U8447 ( .A(n14799), .ZN(n6918) );
  INV_X1 U8448 ( .A(n14800), .ZN(n6919) );
  NOR2_X1 U8449 ( .A1(n14817), .A2(n11142), .ZN(n14835) );
  INV_X1 U8450 ( .A(n6908), .ZN(n14852) );
  OAI21_X1 U8451 ( .B1(n14853), .B2(n6906), .A(n6905), .ZN(n14868) );
  NAND2_X1 U8452 ( .A1(n6909), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U8453 ( .A1(n11145), .A2(n6909), .ZN(n6905) );
  INV_X1 U8454 ( .A(n14869), .ZN(n6909) );
  INV_X1 U8455 ( .A(n11145), .ZN(n6907) );
  INV_X1 U8456 ( .A(n6916), .ZN(n14918) );
  NOR2_X1 U8457 ( .A1(n11431), .A2(n11430), .ZN(n11433) );
  INV_X1 U8458 ( .A(n6914), .ZN(n11429) );
  NAND2_X1 U8459 ( .A1(n11436), .A2(n11437), .ZN(n11438) );
  XNOR2_X1 U8460 ( .A(n12616), .B(n12625), .ZN(n11717) );
  INV_X1 U8461 ( .A(n6913), .ZN(n12614) );
  OR2_X1 U8462 ( .A1(n11715), .A2(n14190), .ZN(n6913) );
  INV_X1 U8463 ( .A(n12615), .ZN(n6912) );
  OAI21_X1 U8464 ( .B1(n11715), .B2(n6911), .A(n6910), .ZN(n12639) );
  NAND2_X1 U8465 ( .A1(n12628), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U8466 ( .A1(n12665), .A2(n12664), .ZN(n12695) );
  NAND2_X1 U8467 ( .A1(n12668), .A2(n12669), .ZN(n12670) );
  INV_X1 U8468 ( .A(n12701), .ZN(n14168) );
  INV_X1 U8469 ( .A(n9619), .ZN(n7368) );
  AND2_X1 U8470 ( .A1(n12768), .A2(n12767), .ZN(n12943) );
  NAND2_X1 U8471 ( .A1(n12801), .A2(n12800), .ZN(n12799) );
  INV_X1 U8472 ( .A(n12346), .ZN(n12958) );
  AND2_X1 U8473 ( .A1(n12834), .A2(n12833), .ZN(n12967) );
  NAND2_X1 U8474 ( .A1(n7008), .A2(n7012), .ZN(n12874) );
  OR2_X1 U8475 ( .A1(n12902), .A2(n7013), .ZN(n7008) );
  NAND2_X1 U8476 ( .A1(n9452), .A2(n9451), .ZN(n12869) );
  AND2_X1 U8477 ( .A1(n12900), .A2(n12474), .ZN(n12888) );
  NAND2_X1 U8478 ( .A1(n9410), .A2(n9409), .ZN(n12896) );
  NAND2_X1 U8479 ( .A1(n11887), .A2(n12467), .ZN(n12924) );
  NAND2_X1 U8480 ( .A1(n9334), .A2(n9332), .ZN(n14185) );
  NAND2_X1 U8481 ( .A1(n14932), .A2(n9285), .ZN(n14199) );
  INV_X1 U8482 ( .A(n12928), .ZN(n12878) );
  NAND2_X1 U8483 ( .A1(n6979), .A2(n12414), .ZN(n10929) );
  NAND2_X1 U8484 ( .A1(n10790), .A2(n12565), .ZN(n6979) );
  OR2_X1 U8485 ( .A1(n10340), .A2(n14979), .ZN(n14939) );
  NAND2_X1 U8486 ( .A1(n10337), .A2(n10336), .ZN(n14978) );
  INV_X1 U8487 ( .A(n12778), .ZN(n13011) );
  INV_X1 U8488 ( .A(n12791), .ZN(n13015) );
  INV_X1 U8489 ( .A(n12315), .ZN(n13019) );
  NAND2_X1 U8490 ( .A1(n9346), .A2(n9345), .ZN(n11912) );
  AND2_X1 U8491 ( .A1(n9660), .A2(n9659), .ZN(n13045) );
  OR2_X1 U8492 ( .A1(n9658), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9660) );
  AND2_X1 U8493 ( .A1(n10079), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13046) );
  INV_X1 U8494 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9080) );
  XNOR2_X1 U8495 ( .A(n6663), .B(n12535), .ZN(n13049) );
  OAI21_X1 U8496 ( .B1(n9591), .B2(n6658), .A(n6656), .ZN(n6663) );
  INV_X1 U8497 ( .A(n6657), .ZN(n6656) );
  NAND2_X1 U8498 ( .A1(n6655), .A2(n6659), .ZN(n12534) );
  INV_X1 U8499 ( .A(SI_29_), .ZN(n13057) );
  INV_X1 U8500 ( .A(SI_26_), .ZN(n11645) );
  OR2_X1 U8501 ( .A1(n6670), .A2(n6671), .ZN(n9533) );
  INV_X1 U8502 ( .A(n6689), .ZN(n6688) );
  OR2_X1 U8503 ( .A1(n9648), .A2(n6692), .ZN(n6687) );
  OAI21_X1 U8504 ( .B1(n9504), .B2(n9503), .A(n9505), .ZN(n9518) );
  INV_X1 U8505 ( .A(n9692), .ZN(n10725) );
  NAND2_X1 U8506 ( .A1(n7160), .A2(n7165), .ZN(n9470) );
  INV_X1 U8507 ( .A(n7161), .ZN(n7160) );
  INV_X1 U8508 ( .A(SI_19_), .ZN(n10465) );
  NAND2_X1 U8509 ( .A1(n9396), .A2(n9395), .ZN(n9413) );
  NAND2_X1 U8510 ( .A1(n9398), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9399) );
  INV_X1 U8511 ( .A(SI_16_), .ZN(n9991) );
  INV_X1 U8512 ( .A(SI_14_), .ZN(n9822) );
  INV_X1 U8513 ( .A(SI_12_), .ZN(n9760) );
  INV_X1 U8514 ( .A(n11721), .ZN(n11714) );
  NAND2_X1 U8515 ( .A1(n9294), .A2(n9293), .ZN(n9299) );
  INV_X1 U8516 ( .A(SI_11_), .ZN(n9745) );
  INV_X1 U8517 ( .A(n11200), .ZN(n14876) );
  NAND2_X1 U8518 ( .A1(n9238), .A2(n9237), .ZN(n9241) );
  NAND2_X1 U8519 ( .A1(n9223), .A2(n9222), .ZN(n9226) );
  INV_X1 U8520 ( .A(n11188), .ZN(n14842) );
  XNOR2_X1 U8521 ( .A(n9169), .B(n9168), .ZN(n14807) );
  NAND2_X1 U8522 ( .A1(n7121), .A2(n9146), .ZN(n9164) );
  NAND2_X1 U8523 ( .A1(n9145), .A2(n9144), .ZN(n7121) );
  INV_X1 U8524 ( .A(n12208), .ZN(n7310) );
  NAND2_X1 U8525 ( .A1(n7329), .A2(n11845), .ZN(n14232) );
  AND2_X1 U8526 ( .A1(n11852), .A2(n11845), .ZN(n7328) );
  NAND2_X1 U8527 ( .A1(n10413), .A2(n10412), .ZN(n10417) );
  AND2_X1 U8528 ( .A1(n10419), .A2(n10412), .ZN(n7309) );
  NAND2_X1 U8529 ( .A1(n7323), .A2(n12174), .ZN(n13075) );
  NAND2_X1 U8530 ( .A1(n7081), .A2(n8960), .ZN(n13436) );
  NAND2_X1 U8531 ( .A1(n11927), .A2(n6490), .ZN(n7081) );
  AND2_X1 U8532 ( .A1(n7298), .A2(n7295), .ZN(n11546) );
  NAND2_X1 U8533 ( .A1(n7299), .A2(n7304), .ZN(n11419) );
  INV_X1 U8534 ( .A(n7300), .ZN(n7295) );
  NAND2_X1 U8535 ( .A1(n6807), .A2(n8915), .ZN(n13457) );
  NAND2_X1 U8536 ( .A1(n11880), .A2(n6489), .ZN(n6807) );
  NAND2_X1 U8537 ( .A1(n7327), .A2(n10873), .ZN(n10876) );
  NAND2_X1 U8538 ( .A1(n6764), .A2(n7317), .ZN(n13127) );
  NAND2_X1 U8539 ( .A1(n13110), .A2(n6766), .ZN(n6764) );
  NAND2_X1 U8540 ( .A1(n7298), .A2(n7296), .ZN(n11840) );
  NOR2_X1 U8541 ( .A1(n7300), .A2(n7297), .ZN(n7296) );
  INV_X1 U8542 ( .A(n11545), .ZN(n7297) );
  OAI21_X1 U8543 ( .B1(n11104), .B2(n11103), .A(n11102), .ZN(n11418) );
  NAND2_X1 U8544 ( .A1(n13109), .A2(n12169), .ZN(n13152) );
  NAND2_X1 U8545 ( .A1(n10539), .A2(n7335), .ZN(n10717) );
  AND2_X1 U8546 ( .A1(n10545), .A2(n10538), .ZN(n7335) );
  AND2_X1 U8547 ( .A1(n10539), .A2(n10538), .ZN(n10546) );
  XNOR2_X1 U8548 ( .A(n7060), .B(n13217), .ZN(n9036) );
  INV_X1 U8549 ( .A(n13061), .ZN(n13172) );
  OR2_X1 U8550 ( .A1(n8580), .A2(n8528), .ZN(n8529) );
  NAND2_X1 U8551 ( .A1(n6478), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8500) );
  OR2_X1 U8552 ( .A1(n8966), .A2(n13412), .ZN(n8498) );
  OR2_X1 U8553 ( .A1(n6476), .A2(n13415), .ZN(n8499) );
  OR2_X2 U8554 ( .A1(n9772), .A2(P2_U3088), .ZN(n13199) );
  OR2_X1 U8555 ( .A1(n6476), .A2(n10829), .ZN(n8459) );
  NOR2_X1 U8556 ( .A1(n10129), .A2(n10128), .ZN(n10162) );
  AOI21_X1 U8557 ( .B1(n10524), .B2(n11309), .A(n10523), .ZN(n10528) );
  NAND2_X1 U8558 ( .A1(n11324), .A2(n6606), .ZN(n11327) );
  INV_X1 U8559 ( .A(n13214), .ZN(n13216) );
  NAND2_X1 U8560 ( .A1(n13224), .A2(n6486), .ZN(n13427) );
  INV_X1 U8561 ( .A(n9033), .ZN(n13430) );
  OR2_X1 U8562 ( .A1(n13236), .A2(n6787), .ZN(n6782) );
  NAND2_X1 U8563 ( .A1(n11971), .A2(n11940), .ZN(n6787) );
  OAI21_X1 U8564 ( .B1(n11941), .B2(n6785), .A(n6784), .ZN(n6783) );
  NOR2_X1 U8565 ( .A1(n13244), .A2(n6786), .ZN(n6785) );
  NAND2_X1 U8566 ( .A1(n11941), .A2(n11940), .ZN(n6784) );
  INV_X1 U8567 ( .A(n11940), .ZN(n6786) );
  INV_X1 U8568 ( .A(n6827), .ZN(n13431) );
  INV_X1 U8569 ( .A(n13436), .ZN(n13240) );
  INV_X1 U8570 ( .A(n6891), .ZN(n13251) );
  OAI21_X1 U8571 ( .B1(n13278), .B2(n6893), .A(n6892), .ZN(n6891) );
  OAI21_X1 U8572 ( .B1(n13278), .B2(n13280), .A(n11966), .ZN(n13267) );
  NAND2_X1 U8573 ( .A1(n7219), .A2(n7222), .ZN(n13281) );
  OAI21_X1 U8574 ( .B1(n11937), .B2(n7223), .A(n7220), .ZN(n13279) );
  NAND2_X1 U8575 ( .A1(n11937), .A2(n7224), .ZN(n7219) );
  NAND2_X1 U8576 ( .A1(n11937), .A2(n11936), .ZN(n13297) );
  NAND2_X1 U8577 ( .A1(n6880), .A2(n11961), .ZN(n13322) );
  OR2_X1 U8578 ( .A1(n13337), .A2(n11962), .ZN(n6880) );
  OAI21_X1 U8579 ( .B1(n11956), .B2(n6845), .A(n6843), .ZN(n13359) );
  AND2_X1 U8580 ( .A1(n7246), .A2(n7252), .ZN(n13350) );
  NAND2_X1 U8581 ( .A1(n7247), .A2(n7249), .ZN(n7246) );
  NAND2_X1 U8582 ( .A1(n11956), .A2(n11955), .ZN(n13362) );
  OAI21_X1 U8583 ( .B1(n11740), .B2(n6858), .A(n6522), .ZN(n13394) );
  NAND2_X1 U8584 ( .A1(n6856), .A2(n6860), .ZN(n11950) );
  NAND2_X1 U8585 ( .A1(n11740), .A2(n6862), .ZN(n6856) );
  NAND2_X1 U8586 ( .A1(n6864), .A2(n11738), .ZN(n11783) );
  NAND2_X1 U8587 ( .A1(n6865), .A2(n6866), .ZN(n6864) );
  AND2_X1 U8588 ( .A1(n6789), .A2(n6497), .ZN(n11741) );
  NAND2_X1 U8589 ( .A1(n11516), .A2(n11515), .ZN(n11647) );
  NAND2_X1 U8590 ( .A1(n11497), .A2(n11273), .ZN(n11299) );
  NAND2_X1 U8591 ( .A1(n11471), .A2(n11279), .ZN(n11334) );
  INV_X1 U8592 ( .A(n13422), .ZN(n13398) );
  OAI21_X1 U8593 ( .B1(n11467), .B2(n7229), .A(n7228), .ZN(n11476) );
  NAND2_X1 U8594 ( .A1(n11465), .A2(n11271), .ZN(n11478) );
  OAI21_X1 U8595 ( .B1(n10702), .B2(n6850), .A(n6849), .ZN(n11275) );
  NAND2_X1 U8596 ( .A1(n11058), .A2(n11057), .ZN(n11060) );
  NAND2_X1 U8597 ( .A1(n13406), .A2(n11051), .ZN(n13411) );
  INV_X1 U8598 ( .A(n10694), .ZN(n11044) );
  NAND2_X1 U8599 ( .A1(n8815), .A2(n9779), .ZN(n7233) );
  NAND2_X1 U8600 ( .A1(n8568), .A2(n9728), .ZN(n7234) );
  INV_X1 U8601 ( .A(n13417), .ZN(n13399) );
  INV_X2 U8602 ( .A(n14766), .ZN(n14768) );
  INV_X2 U8603 ( .A(n14755), .ZN(n14756) );
  AND2_X1 U8604 ( .A1(n10224), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14686) );
  INV_X1 U8605 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U8606 ( .A1(n13566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8450) );
  INV_X1 U8607 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11882) );
  NAND2_X1 U8608 ( .A1(n9058), .A2(n9057), .ZN(n11881) );
  NAND2_X1 U8609 ( .A1(n9049), .A2(n9055), .ZN(n11837) );
  OR2_X1 U8610 ( .A1(n9040), .A2(n8728), .ZN(n8480) );
  NAND2_X1 U8611 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  INV_X1 U8612 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8471) );
  INV_X1 U8613 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10886) );
  INV_X1 U8614 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10532) );
  INV_X1 U8615 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10680) );
  INV_X1 U8616 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10616) );
  INV_X1 U8617 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9901) );
  INV_X1 U8618 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9893) );
  INV_X1 U8619 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9819) );
  INV_X1 U8620 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9802) );
  INV_X1 U8621 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9795) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9765) );
  INV_X1 U8623 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9758) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9750) );
  INV_X1 U8625 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9748) );
  INV_X1 U8626 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9752) );
  AOI21_X1 U8627 ( .B1(n7092), .B2(n7094), .A(n6545), .ZN(n7090) );
  AOI22_X1 U8628 ( .A1(n12036), .A2(n12035), .B1(n12034), .B2(n12033), .ZN(
        n14245) );
  NAND2_X1 U8629 ( .A1(n13644), .A2(n12102), .ZN(n13592) );
  NAND2_X1 U8630 ( .A1(n7108), .A2(n7109), .ZN(n13604) );
  NAND2_X1 U8631 ( .A1(n13635), .A2(n12093), .ZN(n13611) );
  NAND2_X1 U8632 ( .A1(n7087), .A2(n7088), .ZN(n7086) );
  INV_X1 U8633 ( .A(n12068), .ZN(n14305) );
  NAND2_X1 U8634 ( .A1(n7097), .A2(n7098), .ZN(n13627) );
  AOI21_X1 U8635 ( .B1(n7099), .B2(n7101), .A(n6544), .ZN(n7098) );
  NAND2_X1 U8636 ( .A1(n7901), .A2(n7900), .ZN(n10751) );
  NAND2_X1 U8637 ( .A1(n7114), .A2(n7115), .ZN(n11594) );
  AND2_X1 U8638 ( .A1(n7116), .A2(n11394), .ZN(n11399) );
  AND2_X1 U8639 ( .A1(n11694), .A2(n11695), .ZN(n6619) );
  AOI21_X1 U8640 ( .B1(n14266), .B2(n14262), .A(n14264), .ZN(n14283) );
  NAND2_X1 U8641 ( .A1(n7091), .A2(n12123), .ZN(n13656) );
  NAND2_X1 U8642 ( .A1(n13619), .A2(n13620), .ZN(n7091) );
  OR2_X1 U8643 ( .A1(n10292), .A2(n10276), .ZN(n13663) );
  NAND2_X1 U8644 ( .A1(n7095), .A2(n12057), .ZN(n14296) );
  INV_X1 U8645 ( .A(n7096), .ZN(n7095) );
  INV_X1 U8646 ( .A(n14284), .ZN(n14364) );
  INV_X1 U8647 ( .A(n13663), .ZN(n14359) );
  NAND2_X1 U8648 ( .A1(n10728), .A2(n7083), .ZN(n10729) );
  NOR2_X1 U8649 ( .A1(n7084), .A2(n10289), .ZN(n7083) );
  AND2_X1 U8650 ( .A1(n6733), .A2(n8417), .ZN(n6633) );
  XNOR2_X1 U8651 ( .A(n6734), .B(n13897), .ZN(n6733) );
  NOR3_X1 U8652 ( .A1(n8413), .A2(n8414), .A3(n6735), .ZN(n6734) );
  OR2_X1 U8653 ( .A1(n8205), .A2(n7856), .ZN(n7857) );
  NAND2_X1 U8654 ( .A1(n6485), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7845) );
  OR2_X1 U8655 ( .A1(n10494), .A2(n10493), .ZN(n10969) );
  INV_X1 U8656 ( .A(n8378), .ZN(n14016) );
  AOI21_X1 U8657 ( .B1(n12273), .B2(n8372), .A(n7382), .ZN(n14019) );
  AND2_X1 U8658 ( .A1(n7826), .A2(n7825), .ZN(n14022) );
  NAND2_X1 U8659 ( .A1(n8341), .A2(n8340), .ZN(n14028) );
  AND2_X1 U8660 ( .A1(n13859), .A2(n13858), .ZN(n14030) );
  AND2_X1 U8661 ( .A1(n6929), .A2(n6493), .ZN(n13829) );
  AND2_X1 U8662 ( .A1(n13890), .A2(n12018), .ZN(n13874) );
  NOR2_X1 U8663 ( .A1(n13912), .A2(n12001), .ZN(n13889) );
  NAND2_X1 U8664 ( .A1(n13925), .A2(n6935), .ZN(n13904) );
  NAND2_X1 U8665 ( .A1(n13925), .A2(n12016), .ZN(n13902) );
  NAND2_X1 U8666 ( .A1(n8276), .A2(n8275), .ZN(n13920) );
  INV_X1 U8667 ( .A(n13947), .ZN(n14063) );
  NAND2_X1 U8668 ( .A1(n7202), .A2(n11993), .ZN(n13971) );
  OR2_X1 U8669 ( .A1(n13993), .A2(n13994), .ZN(n7202) );
  NAND2_X1 U8670 ( .A1(n6926), .A2(n12008), .ZN(n13999) );
  NAND2_X1 U8671 ( .A1(n11868), .A2(n7209), .ZN(n11989) );
  NAND2_X1 U8672 ( .A1(n8138), .A2(n8137), .ZN(n14256) );
  NAND2_X2 U8673 ( .A1(n8094), .A2(n8093), .ZN(n14247) );
  NAND2_X1 U8674 ( .A1(n6899), .A2(n10906), .ZN(n11008) );
  NAND2_X1 U8675 ( .A1(n14387), .A2(n14386), .ZN(n6899) );
  NAND2_X1 U8676 ( .A1(n10897), .A2(n10896), .ZN(n14389) );
  NAND2_X1 U8677 ( .A1(n8000), .A2(n7999), .ZN(n14557) );
  INV_X1 U8678 ( .A(n13897), .ZN(n13964) );
  INV_X1 U8679 ( .A(n13917), .ZN(n14452) );
  INV_X1 U8680 ( .A(n10637), .ZN(n14503) );
  OR2_X1 U8681 ( .A1(n13987), .A2(n10573), .ZN(n14444) );
  AND2_X1 U8682 ( .A1(n13923), .A2(n10560), .ZN(n13998) );
  INV_X1 U8683 ( .A(n14594), .ZN(n14591) );
  NAND2_X1 U8684 ( .A1(n14015), .A2(n6625), .ZN(n14097) );
  INV_X1 U8685 ( .A(n6626), .ZN(n6625) );
  OAI21_X1 U8686 ( .B1(n14016), .B2(n14570), .A(n14017), .ZN(n6626) );
  AND2_X1 U8687 ( .A1(n6816), .A2(n6630), .ZN(n6629) );
  NAND2_X1 U8688 ( .A1(n14025), .A2(n14522), .ZN(n6631) );
  OR2_X1 U8689 ( .A1(n14026), .A2(n14517), .ZN(n6628) );
  INV_X1 U8690 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7211) );
  INV_X1 U8691 ( .A(n7813), .ZN(n14119) );
  INV_X1 U8692 ( .A(n7812), .ZN(n14120) );
  NOR2_X1 U8693 ( .A1(n6614), .A2(n6613), .ZN(n6612) );
  NAND2_X1 U8694 ( .A1(n8432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8426) );
  OR2_X1 U8695 ( .A1(n8863), .A2(n8501), .ZN(n8245) );
  XNOR2_X1 U8696 ( .A(n7689), .B(n7688), .ZN(n11297) );
  INV_X1 U8697 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10884) );
  INV_X1 U8698 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10847) );
  INV_X1 U8699 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10534) );
  INV_X1 U8700 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10682) );
  INV_X1 U8701 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10614) );
  AND2_X1 U8702 ( .A1(n8091), .A2(n8079), .ZN(n10497) );
  INV_X1 U8703 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9891) );
  INV_X1 U8704 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9821) );
  INV_X1 U8705 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9804) );
  INV_X1 U8706 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9797) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9763) );
  INV_X1 U8708 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9756) );
  NAND2_X1 U8709 ( .A1(n15090), .A2(n15091), .ZN(n7437) );
  NOR2_X1 U8710 ( .A1(n15088), .A2(n7444), .ZN(n15080) );
  XNOR2_X1 U8711 ( .A(n7452), .B(n6949), .ZN(n14145) );
  NAND2_X1 U8712 ( .A1(n6950), .A2(n7464), .ZN(n14149) );
  NAND2_X1 U8713 ( .A1(n14146), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6950) );
  AND2_X1 U8714 ( .A1(n6957), .A2(n6955), .ZN(n14348) );
  NOR2_X1 U8715 ( .A1(n7487), .A2(n6956), .ZN(n6955) );
  INV_X1 U8716 ( .A(n6959), .ZN(n6956) );
  NAND2_X1 U8717 ( .A1(n14350), .A2(n14351), .ZN(n14347) );
  NAND2_X1 U8718 ( .A1(n6681), .A2(n12596), .ZN(P3_U3296) );
  OAI21_X1 U8719 ( .B1(n12590), .B2(n6682), .A(n10012), .ZN(n6681) );
  NAND2_X1 U8720 ( .A1(n6972), .A2(n6971), .ZN(P3_U3491) );
  NAND2_X1 U8721 ( .A1(P3_U3897), .A2(n6975), .ZN(n6971) );
  OR2_X1 U8722 ( .A1(P3_U3897), .A2(n6973), .ZN(n6972) );
  INV_X1 U8723 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U8724 ( .A1(n6772), .A2(n14910), .ZN(n6771) );
  AOI21_X1 U8725 ( .B1(n12742), .B2(n14892), .A(n12741), .ZN(n6770) );
  OR2_X1 U8726 ( .A1(n15079), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U8727 ( .A1(n12268), .A2(n9689), .ZN(n6650) );
  OAI21_X1 U8728 ( .B1(n9702), .B2(n15064), .A(n6622), .ZN(n9704) );
  NAND2_X1 U8729 ( .A1(n15064), .A2(n9597), .ZN(n6622) );
  NAND2_X1 U8730 ( .A1(n12268), .A2(n13000), .ZN(n6649) );
  AOI22_X1 U8731 ( .A1(n13160), .A2(n13159), .B1(n7312), .B2(n7314), .ZN(
        n13169) );
  NAND2_X1 U8732 ( .A1(n6851), .A2(n6607), .ZN(P2_U3496) );
  NAND2_X1 U8733 ( .A1(n13548), .A2(n14756), .ZN(n6851) );
  NAND2_X1 U8734 ( .A1(n6624), .A2(n6623), .ZN(P1_U3527) );
  NAND2_X1 U8735 ( .A1(n14576), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8736 ( .A1(n14097), .A2(n14578), .ZN(n6624) );
  INV_X1 U8737 ( .A(n6963), .ZN(n14339) );
  NAND2_X1 U8738 ( .A1(n6958), .A2(n6963), .ZN(n14343) );
  XNOR2_X1 U8739 ( .A(n6953), .B(n6952), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8740 ( .A(n7664), .B(n7490), .ZN(n6952) );
  NOR2_X1 U8741 ( .A1(n14134), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8742 ( .A1(n11532), .A2(n14936), .ZN(n6491) );
  AND2_X2 U8743 ( .A1(n10202), .A2(n8481), .ZN(n6512) );
  INV_X1 U8744 ( .A(n10097), .ZN(n12262) );
  NAND2_X2 U8745 ( .A1(n8453), .A2(n8457), .ZN(n8526) );
  INV_X1 U8746 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8135) );
  INV_X1 U8747 ( .A(n13905), .ZN(n7205) );
  OR2_X1 U8748 ( .A1(n11052), .A2(n13195), .ZN(n6492) );
  AND2_X1 U8749 ( .A1(n6930), .A2(n12006), .ZN(n6493) );
  OR2_X1 U8750 ( .A1(n13474), .A2(n11963), .ZN(n6494) );
  INV_X1 U8751 ( .A(n7223), .ZN(n7222) );
  NOR2_X1 U8752 ( .A1(n13296), .A2(n6495), .ZN(n7223) );
  AND2_X1 U8753 ( .A1(n13462), .A2(n13176), .ZN(n6495) );
  AND2_X1 U8754 ( .A1(n10947), .A2(n14950), .ZN(n10948) );
  INV_X1 U8755 ( .A(n6937), .ZN(n10583) );
  OAI21_X1 U8756 ( .B1(n14357), .B2(n10751), .A(n14420), .ZN(n6937) );
  INV_X1 U8757 ( .A(n12800), .ZN(n12797) );
  AND2_X1 U8758 ( .A1(n11961), .A2(n6494), .ZN(n6496) );
  NAND2_X1 U8759 ( .A1(n11649), .A2(n13187), .ZN(n6497) );
  INV_X1 U8760 ( .A(n12008), .ZN(n7042) );
  INV_X1 U8761 ( .A(n14298), .ZN(n6817) );
  AND2_X1 U8762 ( .A1(n12474), .A2(n12479), .ZN(n12897) );
  NAND2_X1 U8763 ( .A1(n12249), .A2(n12335), .ZN(n12282) );
  INV_X1 U8764 ( .A(n10508), .ZN(n6697) );
  AND2_X1 U8765 ( .A1(n12518), .A2(n12752), .ZN(n12769) );
  INV_X1 U8766 ( .A(n13274), .ZN(n13449) );
  NAND2_X1 U8767 ( .A1(n8926), .A2(n8925), .ZN(n13274) );
  AND2_X1 U8768 ( .A1(n7358), .A2(n7359), .ZN(n6498) );
  AND2_X1 U8769 ( .A1(n6563), .A2(n6497), .ZN(n6499) );
  OR2_X1 U8770 ( .A1(n7312), .A2(n7310), .ZN(n6500) );
  INV_X1 U8771 ( .A(n13532), .ZN(n14239) );
  AND2_X1 U8772 ( .A1(n11748), .A2(n11854), .ZN(n6501) );
  OR2_X1 U8773 ( .A1(n7398), .A2(n7397), .ZN(n6502) );
  NAND2_X1 U8774 ( .A1(n12485), .A2(n12474), .ZN(n6503) );
  AND2_X1 U8775 ( .A1(n9429), .A2(n9409), .ZN(n6504) );
  AND2_X1 U8776 ( .A1(n6783), .A2(n13525), .ZN(n6505) );
  INV_X1 U8777 ( .A(n7942), .ZN(n7046) );
  OR2_X1 U8778 ( .A1(n9332), .A2(n7359), .ZN(n6506) );
  OR2_X1 U8779 ( .A1(n7350), .A2(n7349), .ZN(n6507) );
  INV_X1 U8780 ( .A(n13387), .ZN(n7251) );
  INV_X1 U8781 ( .A(n7074), .ZN(n7073) );
  AND2_X1 U8782 ( .A1(n7080), .A2(n7758), .ZN(n7074) );
  INV_X1 U8783 ( .A(n12268), .ZN(n13007) );
  NAND2_X1 U8784 ( .A1(n9580), .A2(n9579), .ZN(n12268) );
  INV_X1 U8785 ( .A(n8862), .ZN(n7764) );
  NAND2_X1 U8786 ( .A1(n8081), .A2(n8080), .ZN(n11824) );
  INV_X1 U8787 ( .A(n11824), .ZN(n6819) );
  OR2_X1 U8788 ( .A1(n7781), .A2(n11645), .ZN(n6508) );
  AND2_X1 U8789 ( .A1(n7164), .A2(n9453), .ZN(n6510) );
  INV_X1 U8790 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U8791 ( .A1(n13688), .A2(n10285), .ZN(n6511) );
  XNOR2_X1 U8792 ( .A(n6921), .B(n7896), .ZN(n8545) );
  OR2_X1 U8793 ( .A1(n12068), .A2(n14002), .ZN(n6513) );
  AND4_X1 U8794 ( .A1(n9073), .A2(n9072), .A3(n9167), .A4(n9168), .ZN(n6514)
         );
  OR2_X1 U8795 ( .A1(n11154), .A2(n11168), .ZN(n6515) );
  AND2_X1 U8796 ( .A1(n13325), .A2(n6833), .ZN(n6516) );
  AND3_X1 U8797 ( .A1(n8350), .A2(n8349), .A3(n8348), .ZN(n6517) );
  NAND2_X1 U8798 ( .A1(n14045), .A2(n13659), .ZN(n6518) );
  XOR2_X1 U8799 ( .A(n13173), .B(n13442), .Z(n13256) );
  INV_X1 U8800 ( .A(n13256), .ZN(n6890) );
  INV_X1 U8801 ( .A(n12832), .ZN(n7179) );
  INV_X1 U8802 ( .A(n14933), .ZN(n7348) );
  OR2_X1 U8803 ( .A1(n14397), .A2(n14557), .ZN(n6519) );
  NAND2_X1 U8804 ( .A1(n6941), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6520) );
  AND2_X1 U8805 ( .A1(n7334), .A2(n7333), .ZN(n6521) );
  INV_X1 U8806 ( .A(n11227), .ZN(n7194) );
  NAND2_X1 U8807 ( .A1(n11997), .A2(n11996), .ZN(n13942) );
  AND2_X1 U8808 ( .A1(n6857), .A2(n11948), .ZN(n6522) );
  AND2_X1 U8809 ( .A1(n8210), .A2(n8209), .ZN(n14077) );
  INV_X1 U8810 ( .A(n14077), .ZN(n8395) );
  INV_X1 U8811 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7897) );
  AND2_X1 U8812 ( .A1(n12242), .A2(n12857), .ZN(n6523) );
  INV_X1 U8813 ( .A(n7697), .ZN(n7706) );
  XOR2_X1 U8814 ( .A(n13665), .B(n13841), .Z(n13838) );
  INV_X1 U8815 ( .A(n13838), .ZN(n6737) );
  AND2_X1 U8816 ( .A1(n14706), .A2(n11274), .ZN(n6524) );
  NAND2_X1 U8817 ( .A1(n8852), .A2(n8851), .ZN(n13346) );
  INV_X1 U8818 ( .A(n13346), .ZN(n6836) );
  NAND2_X1 U8819 ( .A1(n8885), .A2(n8884), .ZN(n13468) );
  INV_X1 U8820 ( .A(n12468), .ZN(n6994) );
  OR3_X1 U8821 ( .A1(n13985), .A2(n6814), .A3(n14071), .ZN(n6525) );
  AND2_X1 U8822 ( .A1(n10198), .A2(n9022), .ZN(n6526) );
  AND2_X1 U8823 ( .A1(n12329), .A2(n7149), .ZN(n6527) );
  NAND2_X1 U8824 ( .A1(n12054), .A2(n12057), .ZN(n14293) );
  INV_X1 U8825 ( .A(n8330), .ZN(n7049) );
  NAND3_X1 U8826 ( .A1(n12249), .A2(n12335), .A3(n12845), .ZN(n12283) );
  INV_X1 U8827 ( .A(n13091), .ZN(n7315) );
  AND3_X1 U8828 ( .A1(n7169), .A2(n12857), .A3(n12244), .ZN(n6528) );
  AND2_X1 U8829 ( .A1(n7109), .A2(n12083), .ZN(n6529) );
  AND2_X1 U8830 ( .A1(n13539), .A2(n11648), .ZN(n6530) );
  INV_X1 U8831 ( .A(n12811), .ZN(n12816) );
  XNOR2_X1 U8832 ( .A(n12346), .B(n7179), .ZN(n12811) );
  AND2_X1 U8833 ( .A1(n13498), .A2(n13154), .ZN(n6531) );
  INV_X1 U8834 ( .A(n7377), .ZN(n7149) );
  NAND2_X1 U8835 ( .A1(n8648), .A2(n8647), .ZN(n14727) );
  NOR2_X1 U8836 ( .A1(n13289), .A2(n13175), .ZN(n11965) );
  AND2_X1 U8837 ( .A1(n11420), .A2(n7302), .ZN(n6532) );
  AND2_X1 U8838 ( .A1(n12138), .A2(n12137), .ZN(n6533) );
  OR2_X1 U8839 ( .A1(n11970), .A2(n13162), .ZN(n6534) );
  OR2_X1 U8840 ( .A1(n7396), .A2(n7395), .ZN(n6535) );
  INV_X1 U8841 ( .A(n8021), .ZN(n7028) );
  OR2_X1 U8842 ( .A1(n6823), .A2(n11519), .ZN(n6536) );
  OR2_X1 U8843 ( .A1(n13150), .A2(n11963), .ZN(n6537) );
  INV_X1 U8844 ( .A(n8003), .ZN(n7030) );
  INV_X1 U8845 ( .A(n10697), .ZN(n6780) );
  INV_X1 U8846 ( .A(n8616), .ZN(n7290) );
  INV_X1 U8847 ( .A(n11256), .ZN(n7124) );
  INV_X1 U8848 ( .A(n11993), .ZN(n7201) );
  AND2_X1 U8849 ( .A1(n14727), .A2(n11281), .ZN(n6538) );
  AND2_X1 U8850 ( .A1(n11484), .A2(n13192), .ZN(n6539) );
  OR2_X1 U8851 ( .A1(n8235), .A2(n8233), .ZN(n6540) );
  INV_X1 U8852 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7395) );
  AND2_X1 U8853 ( .A1(n6827), .A2(n6830), .ZN(n6541) );
  AND2_X1 U8854 ( .A1(n6491), .A2(n11256), .ZN(n6542) );
  INV_X1 U8855 ( .A(n6894), .ZN(n13280) );
  XNOR2_X1 U8856 ( .A(n13457), .B(n13175), .ZN(n6894) );
  INV_X1 U8857 ( .A(n11520), .ZN(n6823) );
  AND2_X1 U8858 ( .A1(n13433), .A2(n6541), .ZN(n6543) );
  AND2_X1 U8859 ( .A1(n12108), .A2(n12107), .ZN(n6544) );
  AND2_X1 U8860 ( .A1(n12129), .A2(n12128), .ZN(n6545) );
  AND2_X1 U8861 ( .A1(n13523), .A2(n11854), .ZN(n6546) );
  AND2_X1 U8862 ( .A1(n12488), .A2(n12489), .ZN(n12873) );
  NOR2_X1 U8863 ( .A1(n13490), .A2(n13077), .ZN(n6547) );
  NOR2_X1 U8864 ( .A1(n11591), .A2(n13680), .ZN(n6548) );
  NOR2_X1 U8865 ( .A1(n11520), .A2(n11519), .ZN(n6549) );
  NOR2_X1 U8866 ( .A1(n14276), .A2(n11229), .ZN(n6550) );
  NOR2_X1 U8867 ( .A1(n12068), .A2(n11988), .ZN(n6551) );
  NOR2_X1 U8868 ( .A1(n10834), .A2(n10838), .ZN(n6552) );
  INV_X1 U8869 ( .A(n11416), .ZN(n7308) );
  NAND2_X1 U8870 ( .A1(n7383), .A2(n9243), .ZN(n6990) );
  AND2_X1 U8871 ( .A1(n14092), .A2(n13673), .ZN(n6553) );
  NAND2_X1 U8872 ( .A1(n7259), .A2(n7263), .ZN(n6554) );
  AND2_X1 U8873 ( .A1(n8148), .A2(SI_17_), .ZN(n6555) );
  AND2_X1 U8874 ( .A1(n12315), .A2(n12600), .ZN(n6556) );
  INV_X1 U8875 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7793) );
  AND2_X1 U8876 ( .A1(n7245), .A2(n7242), .ZN(n6557) );
  NOR2_X1 U8877 ( .A1(n13920), .A2(n13668), .ZN(n6558) );
  NOR2_X1 U8878 ( .A1(n13457), .A2(n13175), .ZN(n6559) );
  NOR2_X1 U8879 ( .A1(n12078), .A2(n12077), .ZN(n6560) );
  OR2_X1 U8880 ( .A1(n12019), .A2(n13621), .ZN(n6561) );
  AND2_X1 U8881 ( .A1(n6836), .A2(n11960), .ZN(n6562) );
  INV_X1 U8882 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9096) );
  INV_X1 U8883 ( .A(n7210), .ZN(n7209) );
  NAND2_X1 U8884 ( .A1(n11865), .A2(n11867), .ZN(n7210) );
  INV_X1 U8885 ( .A(n7357), .ZN(n7356) );
  NAND2_X1 U8886 ( .A1(n9586), .A2(n9574), .ZN(n7357) );
  OR2_X1 U8887 ( .A1(n13532), .A2(n11846), .ZN(n6563) );
  OR2_X1 U8888 ( .A1(n13091), .A2(n7310), .ZN(n6564) );
  INV_X1 U8889 ( .A(n6730), .ZN(n6729) );
  OR2_X1 U8890 ( .A1(n7751), .A2(n6731), .ZN(n6730) );
  INV_X1 U8891 ( .A(n11273), .ZN(n7240) );
  INV_X1 U8892 ( .A(n8536), .ZN(n7283) );
  NAND2_X1 U8893 ( .A1(n13321), .A2(n6881), .ZN(n6565) );
  OR2_X1 U8894 ( .A1(n7043), .A2(n7042), .ZN(n6566) );
  NAND2_X1 U8895 ( .A1(n12362), .A2(n7149), .ZN(n6567) );
  NAND2_X1 U8896 ( .A1(n7123), .A2(n11533), .ZN(n7122) );
  INV_X1 U8897 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n6693) );
  INV_X1 U8898 ( .A(n10901), .ZN(n11007) );
  OR2_X1 U8899 ( .A1(n11970), .A2(n13173), .ZN(n6568) );
  INV_X1 U8900 ( .A(n12484), .ZN(n7014) );
  AND2_X1 U8901 ( .A1(n6745), .A2(n6520), .ZN(n6569) );
  AND2_X1 U8902 ( .A1(n11941), .A2(n13244), .ZN(n6570) );
  NOR2_X1 U8903 ( .A1(n11398), .A2(n11557), .ZN(n6571) );
  AND2_X1 U8904 ( .A1(n7213), .A2(n7211), .ZN(n6572) );
  AND2_X1 U8905 ( .A1(n6963), .A2(n6962), .ZN(n6573) );
  AND2_X1 U8906 ( .A1(n11139), .A2(n6920), .ZN(n6574) );
  OR2_X1 U8907 ( .A1(n8296), .A2(n8294), .ZN(n6575) );
  OR2_X1 U8908 ( .A1(n8062), .A2(n8060), .ZN(n6576) );
  AND2_X1 U8909 ( .A1(n7286), .A2(n8448), .ZN(n6577) );
  OR2_X1 U8910 ( .A1(n8649), .A2(n8653), .ZN(n6578) );
  OR2_X1 U8911 ( .A1(n8575), .A2(n8573), .ZN(n6579) );
  OR2_X1 U8912 ( .A1(n8687), .A2(n8685), .ZN(n6580) );
  OR2_X1 U8913 ( .A1(n8329), .A2(n7049), .ZN(n6581) );
  AND2_X1 U8914 ( .A1(n6669), .A2(n12555), .ZN(n6582) );
  OR2_X1 U8915 ( .A1(n7046), .A2(n7943), .ZN(n6583) );
  OR2_X1 U8916 ( .A1(n8615), .A2(n7290), .ZN(n6584) );
  INV_X1 U8917 ( .A(n12456), .ZN(n9353) );
  AND2_X1 U8918 ( .A1(n12459), .A2(n12463), .ZN(n12456) );
  NAND2_X1 U8919 ( .A1(n8887), .A2(n7269), .ZN(n6585) );
  NAND2_X1 U8920 ( .A1(n8917), .A2(n7272), .ZN(n6586) );
  INV_X1 U8921 ( .A(n11964), .ZN(n6877) );
  OR2_X1 U8922 ( .A1(n13468), .A2(n13121), .ZN(n11964) );
  INV_X1 U8923 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7286) );
  AND2_X1 U8924 ( .A1(n10686), .A2(n6700), .ZN(n6699) );
  INV_X1 U8925 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7212) );
  OR2_X1 U8926 ( .A1(n8395), .A2(n13614), .ZN(n11994) );
  INV_X1 U8927 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U8928 ( .A1(n8854), .A2(n7275), .ZN(n6587) );
  INV_X1 U8929 ( .A(n6705), .ZN(n6704) );
  NAND2_X1 U8930 ( .A1(n6706), .A2(n6542), .ZN(n6705) );
  INV_X1 U8931 ( .A(n12606), .ZN(n7359) );
  INV_X1 U8932 ( .A(n14859), .ZN(n11193) );
  XOR2_X1 U8933 ( .A(n13468), .B(n12213), .Z(n6588) );
  INV_X1 U8934 ( .A(n7677), .ZN(n8111) );
  NOR2_X1 U8935 ( .A1(n14247), .A2(n11607), .ZN(n6818) );
  INV_X1 U8936 ( .A(n13174), .ZN(n13093) );
  AND4_X1 U8937 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n11854)
         );
  INV_X1 U8938 ( .A(n11846), .ZN(n13186) );
  NAND2_X1 U8939 ( .A1(n6776), .A2(n8547), .ZN(n8697) );
  INV_X1 U8940 ( .A(n6838), .ZN(n13379) );
  NOR2_X1 U8941 ( .A1(n13396), .A2(n13503), .ZN(n6838) );
  AND2_X1 U8942 ( .A1(n9593), .A2(n9592), .ZN(n11982) );
  INV_X1 U8943 ( .A(n6862), .ZN(n6861) );
  AND2_X1 U8944 ( .A1(n7202), .A2(n7200), .ZN(n6589) );
  AND2_X1 U8945 ( .A1(n7323), .A2(n7321), .ZN(n6590) );
  INV_X1 U8946 ( .A(SI_13_), .ZN(n9798) );
  INV_X1 U8947 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6938) );
  AND2_X1 U8948 ( .A1(n6913), .A2(n6912), .ZN(n6591) );
  OR2_X1 U8949 ( .A1(n12306), .A2(n12309), .ZN(n12307) );
  OR2_X1 U8950 ( .A1(n13011), .A2(n13043), .ZN(n6592) );
  OR2_X1 U8951 ( .A1(n13011), .A2(n12996), .ZN(n6593) );
  AND2_X1 U8952 ( .A1(n12268), .A2(n12599), .ZN(n6594) );
  AND2_X1 U8953 ( .A1(n9903), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8954 ( .A1(n8242), .A2(n7079), .ZN(n6596) );
  OR2_X1 U8955 ( .A1(n13985), .A2(n6814), .ZN(n6597) );
  AOI21_X1 U8956 ( .B1(n13172), .B2(n13141), .A(n11974), .ZN(n11975) );
  INV_X1 U8957 ( .A(n7252), .ZN(n7248) );
  NAND2_X1 U8958 ( .A1(n13498), .A2(n13181), .ZN(n7252) );
  NAND2_X1 U8959 ( .A1(n13845), .A2(n14439), .ZN(n14010) );
  NAND2_X1 U8960 ( .A1(n10905), .A2(n10904), .ZN(n14387) );
  INV_X2 U8961 ( .A(n15064), .ZN(n15066) );
  AND2_X2 U8962 ( .A1(n10335), .A2(n9688), .ZN(n15079) );
  AND2_X1 U8963 ( .A1(n11339), .A2(n6826), .ZN(n6598) );
  OR2_X1 U8964 ( .A1(n11721), .A2(n9305), .ZN(n6599) );
  INV_X1 U8965 ( .A(n14085), .ZN(n6815) );
  AND2_X1 U8966 ( .A1(n14402), .A2(n10757), .ZN(n6600) );
  INV_X1 U8967 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n6750) );
  INV_X1 U8968 ( .A(SI_22_), .ZN(n9491) );
  AND2_X1 U8969 ( .A1(n6924), .A2(n11605), .ZN(n6601) );
  INV_X1 U8970 ( .A(n6820), .ZN(n11377) );
  NAND2_X1 U8971 ( .A1(n7056), .A2(n7780), .ZN(n6602) );
  NAND3_X1 U8972 ( .A1(n6687), .A2(n6686), .A3(n6688), .ZN(n9655) );
  NOR2_X1 U8973 ( .A1(n10124), .A2(n6974), .ZN(n6603) );
  AND2_X1 U8974 ( .A1(n10921), .A2(n9174), .ZN(n6604) );
  INV_X1 U8975 ( .A(n14578), .ZN(n14576) );
  INV_X1 U8976 ( .A(n7082), .ZN(n10558) );
  NAND2_X1 U8977 ( .A1(n10278), .A2(n10328), .ZN(n7082) );
  NAND4_X1 U8978 ( .A1(n8517), .A2(n8516), .A3(n8515), .A4(n8514), .ZN(n13198)
         );
  INV_X1 U8979 ( .A(n13198), .ZN(n7235) );
  AND2_X2 U8980 ( .A1(n12595), .A2(n10791), .ZN(n12525) );
  INV_X1 U8981 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7164) );
  INV_X1 U8982 ( .A(n14769), .ZN(n14910) );
  INV_X1 U8983 ( .A(n10199), .ZN(n6774) );
  AND2_X1 U8984 ( .A1(n14739), .A2(n10245), .ZN(n14718) );
  INV_X1 U8985 ( .A(n14718), .ZN(n13525) );
  XOR2_X1 U8986 ( .A(n10852), .B(n10851), .Z(n6605) );
  OR2_X1 U8987 ( .A1(n11326), .A2(n11325), .ZN(n6606) );
  OR2_X1 U8988 ( .A1(n14756), .A2(n8973), .ZN(n6607) );
  AND2_X1 U8989 ( .A1(n6908), .A2(n6907), .ZN(n6608) );
  INV_X1 U8990 ( .A(n14975), .ZN(n6970) );
  AND2_X1 U8991 ( .A1(n11628), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6609) );
  INV_X1 U8992 ( .A(n10948), .ZN(n6710) );
  XNOR2_X1 U8993 ( .A(n9438), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12723) );
  INV_X1 U8994 ( .A(n12723), .ZN(n12740) );
  INV_X1 U8995 ( .A(n10202), .ZN(n13217) );
  OR2_X1 U8996 ( .A1(n12533), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6610) );
  AND2_X1 U8997 ( .A1(n6919), .A2(n6918), .ZN(n6611) );
  INV_X1 U8998 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n6904) );
  INV_X1 U8999 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7694) );
  INV_X1 U9000 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6901) );
  INV_X1 U9001 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7392) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6648) );
  INV_X1 U9003 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7162) );
  INV_X1 U9004 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6660) );
  INV_X1 U9005 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6949) );
  INV_X1 U9006 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U9007 ( .A1(n14254), .A2(n14255), .ZN(n14253) );
  NAND2_X1 U9008 ( .A1(n6643), .A2(n6571), .ZN(n7114) );
  OAI21_X1 U9009 ( .B1(n10855), .B2(n10854), .A(n10853), .ZN(n11024) );
  OAI21_X1 U9010 ( .B1(n10743), .B2(n10742), .A(n14358), .ZN(n10745) );
  AOI21_X1 U9011 ( .B1(n13584), .B2(n13585), .A(n6533), .ZN(n12145) );
  NAND2_X1 U9012 ( .A1(n14274), .A2(n14275), .ZN(n14273) );
  NAND2_X2 U9013 ( .A1(n6615), .A2(n6612), .ZN(n14122) );
  XNOR2_X1 U9014 ( .A(n10694), .B(n10426), .ZN(n10416) );
  NAND2_X1 U9015 ( .A1(n10783), .A2(n10782), .ZN(n10872) );
  NAND2_X2 U9016 ( .A1(n13100), .A2(n13101), .ZN(n13099) );
  NAND2_X2 U9017 ( .A1(n13099), .A2(n12163), .ZN(n13110) );
  INV_X1 U9018 ( .A(n11840), .ZN(n6760) );
  NAND2_X1 U9019 ( .A1(n13126), .A2(n12187), .ZN(n13084) );
  NAND2_X1 U9020 ( .A1(n10428), .A2(n10427), .ZN(n10432) );
  NAND2_X1 U9021 ( .A1(n11604), .A2(n11603), .ZN(n6924) );
  AOI21_X1 U9022 ( .B1(n13983), .B2(n13994), .A(n12011), .ZN(n13970) );
  INV_X1 U9023 ( .A(n12007), .ZN(n6616) );
  NAND2_X2 U9024 ( .A1(n12017), .A2(n13888), .ZN(n13890) );
  OAI21_X2 U9025 ( .B1(n13956), .B2(n12013), .A(n12014), .ZN(n13945) );
  OAI21_X2 U9026 ( .B1(n11792), .B2(n11793), .A(n11791), .ZN(n11862) );
  NAND2_X1 U9027 ( .A1(n10563), .A2(n10562), .ZN(n14435) );
  NAND2_X1 U9028 ( .A1(n13891), .A2(n13878), .ZN(n6929) );
  NAND2_X1 U9029 ( .A1(n11666), .A2(n11665), .ZN(n11792) );
  NAND2_X1 U9030 ( .A1(n14035), .A2(n6617), .ZN(n14101) );
  NAND3_X1 U9031 ( .A1(n6631), .A2(n6628), .A3(n6629), .ZN(n14099) );
  NAND2_X1 U9032 ( .A1(n6924), .A2(n6922), .ZN(n11666) );
  XNOR2_X1 U9033 ( .A(n13833), .B(n13838), .ZN(n14026) );
  NAND2_X1 U9034 ( .A1(n12908), .A2(n9631), .ZN(n9410) );
  NAND2_X1 U9035 ( .A1(n11884), .A2(n12575), .ZN(n11883) );
  AOI21_X1 U9036 ( .B1(n12940), .B2(n15063), .A(n12939), .ZN(n13004) );
  NAND2_X2 U9037 ( .A1(n7342), .A2(n7344), .ZN(n12784) );
  OAI22_X2 U9038 ( .A1(n9334), .A2(n6498), .B1(n7358), .B2(n9333), .ZN(n11828)
         );
  NAND2_X1 U9039 ( .A1(n11827), .A2(n9354), .ZN(n11884) );
  AND2_X1 U9040 ( .A1(n9109), .A2(n9110), .ZN(n9111) );
  NAND2_X1 U9041 ( .A1(n7370), .A2(n10921), .ZN(n10792) );
  NOR2_X1 U9042 ( .A1(n7355), .A2(n7354), .ZN(n12756) );
  INV_X2 U9043 ( .A(n14999), .ZN(n6975) );
  AND2_X2 U9044 ( .A1(n12024), .A2(n6652), .ZN(n14035) );
  INV_X1 U9045 ( .A(n13892), .ZN(n12017) );
  NAND2_X1 U9046 ( .A1(n13945), .A2(n13944), .ZN(n13943) );
  AND2_X2 U9047 ( .A1(n13943), .A2(n12015), .ZN(n7389) );
  OAI21_X2 U9048 ( .B1(n11386), .B2(n11385), .A(n6644), .ZN(n11558) );
  NOR2_X1 U9049 ( .A1(n11693), .A2(n6619), .ZN(n14274) );
  XNOR2_X1 U9050 ( .A(n10283), .B(n10733), .ZN(n10368) );
  NAND2_X1 U9051 ( .A1(n13602), .A2(n12087), .ZN(n13637) );
  NAND2_X1 U9052 ( .A1(n14245), .A2(n14246), .ZN(n14244) );
  NAND2_X1 U9053 ( .A1(n13969), .A2(n12012), .ZN(n13956) );
  INV_X1 U9054 ( .A(n11558), .ZN(n6643) );
  NAND2_X1 U9055 ( .A1(n13010), .A2(n6592), .ZN(P3_U3454) );
  NAND2_X1 U9056 ( .A1(n12947), .A2(n6593), .ZN(P3_U3486) );
  NAND2_X1 U9057 ( .A1(n8055), .A2(n7386), .ZN(n6797) );
  AOI21_X1 U9058 ( .B1(n15058), .B2(n12945), .A(n12944), .ZN(n13008) );
  INV_X1 U9059 ( .A(n7871), .ZN(n6805) );
  NOR2_X1 U9060 ( .A1(n14886), .A2(n11148), .ZN(n14920) );
  XNOR2_X1 U9061 ( .A(n12696), .B(n14173), .ZN(n14169) );
  XNOR2_X1 U9062 ( .A(n12660), .B(n12674), .ZN(n12640) );
  NOR2_X1 U9063 ( .A1(n14818), .A2(n11180), .ZN(n14817) );
  NAND2_X1 U9064 ( .A1(n14341), .A2(n14340), .ZN(n6747) );
  NAND2_X1 U9065 ( .A1(n6747), .A2(n14651), .ZN(n6962) );
  NAND2_X1 U9066 ( .A1(n6957), .A2(n6959), .ZN(n7488) );
  OAI21_X2 U9067 ( .B1(n7468), .B2(n14155), .A(n14152), .ZN(n7472) );
  NAND2_X1 U9068 ( .A1(n6929), .A2(n6930), .ZN(n12020) );
  OAI21_X2 U9069 ( .B1(n7389), .B2(n6934), .A(n6933), .ZN(n13892) );
  NAND2_X1 U9070 ( .A1(n10629), .A2(n10631), .ZN(n10563) );
  XNOR2_X2 U9071 ( .A(n10637), .B(n10374), .ZN(n10631) );
  NAND3_X1 U9072 ( .A1(n6967), .A2(n6969), .A3(n14960), .ZN(n6968) );
  NAND2_X1 U9073 ( .A1(n6966), .A2(n12456), .ZN(n9630) );
  NAND2_X1 U9074 ( .A1(n6965), .A2(n12493), .ZN(n12848) );
  NAND2_X1 U9075 ( .A1(n6964), .A2(n12500), .ZN(n12840) );
  NAND2_X1 U9076 ( .A1(n6985), .A2(n6984), .ZN(n9095) );
  OR2_X2 U9077 ( .A1(n13932), .A2(n13920), .ZN(n13915) );
  OR2_X2 U9078 ( .A1(n13882), .A2(n14033), .ZN(n13866) );
  NAND2_X1 U9079 ( .A1(n6820), .A2(n6819), .ZN(n11607) );
  NOR2_X2 U9080 ( .A1(n6519), .A2(n11591), .ZN(n11009) );
  NAND2_X1 U9081 ( .A1(n14451), .A2(n14516), .ZN(n14430) );
  NAND2_X1 U9082 ( .A1(n8055), .A2(n6798), .ZN(n6796) );
  NAND2_X1 U9083 ( .A1(n7075), .A2(n7758), .ZN(n8225) );
  NAND2_X1 U9084 ( .A1(n6636), .A2(n7025), .ZN(n8311) );
  NAND2_X1 U9085 ( .A1(n6638), .A2(n6637), .ZN(n8248) );
  NOR2_X1 U9086 ( .A1(n8390), .A2(n6634), .ZN(n8385) );
  AOI21_X1 U9087 ( .B1(n8419), .B2(n8418), .A(n6633), .ZN(n8439) );
  INV_X1 U9088 ( .A(n7868), .ZN(n7861) );
  NAND2_X1 U9089 ( .A1(n7701), .A2(n7868), .ZN(n7704) );
  NOR2_X1 U9090 ( .A1(n13879), .A2(n13878), .ZN(n13877) );
  NAND2_X1 U9091 ( .A1(n13993), .A2(n7200), .ZN(n7198) );
  AOI21_X2 U9092 ( .B1(n12784), .B2(n9556), .A(n7390), .ZN(n12771) );
  AND4_X2 U9093 ( .A1(n8034), .A2(n7665), .A3(n7666), .A4(n7669), .ZN(n7117)
         );
  NAND3_X1 U9094 ( .A1(n6632), .A2(n7866), .A3(n10579), .ZN(n7885) );
  NAND2_X1 U9095 ( .A1(n7854), .A2(n7853), .ZN(n6632) );
  OAI21_X1 U9096 ( .B1(n7017), .B2(n7903), .A(n7902), .ZN(n7016) );
  NAND2_X1 U9097 ( .A1(n7034), .A2(n7032), .ZN(n8213) );
  NOR2_X2 U9098 ( .A1(n6517), .A2(n6635), .ZN(n8390) );
  NAND3_X1 U9099 ( .A1(n8283), .A2(n8284), .A3(n6575), .ZN(n6636) );
  NAND3_X1 U9100 ( .A1(n8215), .A2(n8214), .A3(n6540), .ZN(n6638) );
  NAND3_X1 U9101 ( .A1(n8047), .A2(n8046), .A3(n6576), .ZN(n6640) );
  NOR2_X1 U9102 ( .A1(n12640), .A2(n12641), .ZN(n12662) );
  NAND2_X1 U9103 ( .A1(n12615), .A2(n12628), .ZN(n6910) );
  NOR2_X1 U9104 ( .A1(n14835), .A2(n14834), .ZN(n14833) );
  NOR2_X1 U9105 ( .A1(n14888), .A2(n14887), .ZN(n14886) );
  NAND2_X1 U9106 ( .A1(n6917), .A2(n6641), .ZN(n11141) );
  NAND2_X1 U9107 ( .A1(n6574), .A2(n14784), .ZN(n6641) );
  OAI211_X1 U9108 ( .C1(n12743), .C2(n14921), .A(n6771), .B(n6770), .ZN(
        P3_U3201) );
  NAND2_X1 U9109 ( .A1(n12054), .A2(n12056), .ZN(n7096) );
  NAND2_X2 U9110 ( .A1(n13609), .A2(n12097), .ZN(n13645) );
  NAND2_X2 U9111 ( .A1(n12116), .A2(n12115), .ZN(n13619) );
  INV_X1 U9112 ( .A(n6990), .ZN(n6985) );
  OR2_X4 U9113 ( .A1(n9090), .A2(n9089), .ZN(n9157) );
  NAND2_X1 U9114 ( .A1(n11883), .A2(n9375), .ZN(n12919) );
  NAND2_X1 U9115 ( .A1(n12867), .A2(n9469), .ZN(n12855) );
  NAND2_X1 U9116 ( .A1(n14966), .A2(n9155), .ZN(n10922) );
  NAND2_X1 U9117 ( .A1(n13006), .A2(n6649), .ZN(P3_U3455) );
  NAND2_X1 U9118 ( .A1(n12942), .A2(n6650), .ZN(P3_U3487) );
  NAND2_X1 U9119 ( .A1(n6985), .A2(n6983), .ZN(n9084) );
  NAND2_X2 U9120 ( .A1(n12828), .A2(n9516), .ZN(n12817) );
  NAND2_X1 U9121 ( .A1(n9452), .A2(n7360), .ZN(n12867) );
  NAND2_X1 U9122 ( .A1(n12894), .A2(n9430), .ZN(n12883) );
  INV_X1 U9123 ( .A(n12770), .ZN(n7355) );
  NAND2_X1 U9124 ( .A1(n10792), .A2(n7369), .ZN(n10932) );
  INV_X2 U9125 ( .A(n9387), .ZN(n9086) );
  INV_X1 U9126 ( .A(n9387), .ZN(n9156) );
  NAND2_X1 U9127 ( .A1(n11375), .A2(n11374), .ZN(n6651) );
  NOR2_X2 U9128 ( .A1(n13688), .A2(n10285), .ZN(n10578) );
  AND3_X2 U9129 ( .A1(n7839), .A2(n7841), .A3(n7840), .ZN(n10285) );
  NAND3_X1 U9130 ( .A1(n9145), .A2(n9163), .A3(n9144), .ZN(n6653) );
  NAND2_X1 U9131 ( .A1(n9183), .A2(n9182), .ZN(n9185) );
  NAND2_X1 U9132 ( .A1(n9591), .A2(n6661), .ZN(n6655) );
  NAND2_X1 U9133 ( .A1(n9591), .A2(n9590), .ZN(n12225) );
  NAND3_X1 U9134 ( .A1(n6582), .A2(n6665), .A3(n12554), .ZN(n6664) );
  NAND2_X1 U9135 ( .A1(n9532), .A2(n6671), .ZN(n9545) );
  NAND2_X1 U9136 ( .A1(n9532), .A2(n9520), .ZN(n9521) );
  INV_X1 U9137 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U9138 ( .B1(n9360), .B2(n6676), .A(n6673), .ZN(n9417) );
  NAND2_X1 U9139 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  NAND2_X1 U9140 ( .A1(n6685), .A2(n7141), .ZN(n7140) );
  NAND2_X1 U9141 ( .A1(n6685), .A2(n9664), .ZN(n9658) );
  NAND2_X1 U9142 ( .A1(n9653), .A2(n11632), .ZN(n6685) );
  NAND2_X1 U9143 ( .A1(n9648), .A2(n6691), .ZN(n6686) );
  NAND2_X1 U9144 ( .A1(n9648), .A2(n9647), .ZN(n9649) );
  INV_X1 U9145 ( .A(n9655), .ZN(n9665) );
  INV_X1 U9146 ( .A(n10509), .ZN(n6696) );
  NAND2_X1 U9147 ( .A1(n6699), .A2(n10509), .ZN(n6694) );
  OAI21_X1 U9148 ( .B1(n12297), .B2(n6705), .A(n6701), .ZN(n11535) );
  NAND2_X1 U9149 ( .A1(n11535), .A2(n11536), .ZN(n11575) );
  AOI21_X1 U9150 ( .B1(n12328), .B2(n6717), .A(n6712), .ZN(n6711) );
  INV_X1 U9151 ( .A(n6711), .ZN(n12239) );
  NAND2_X1 U9152 ( .A1(n9603), .A2(n6721), .ZN(n9605) );
  NAND4_X1 U9153 ( .A1(n6724), .A2(n9148), .A3(n6514), .A4(n6723), .ZN(n9646)
         );
  INV_X1 U9154 ( .A(n9382), .ZN(n6724) );
  NAND2_X1 U9155 ( .A1(n9244), .A2(n9075), .ZN(n9398) );
  NOR2_X2 U9156 ( .A1(n9382), .A2(n9071), .ZN(n9075) );
  XNOR2_X1 U9157 ( .A(n10395), .B(n12611), .ZN(n10310) );
  XNOR2_X1 U9158 ( .A(n10097), .B(n14970), .ZN(n10395) );
  NAND2_X2 U9159 ( .A1(n6725), .A2(n8165), .ZN(n14085) );
  NAND3_X1 U9160 ( .A1(n6737), .A2(n8415), .A3(n6736), .ZN(n6735) );
  NOR2_X1 U9161 ( .A1(n7711), .A2(n7911), .ZN(n6738) );
  NAND3_X1 U9162 ( .A1(n12013), .A2(n6740), .A3(n6739), .ZN(n8412) );
  INV_X1 U9163 ( .A(n7433), .ZN(n6744) );
  XNOR2_X2 U9164 ( .A(n7398), .B(n7397), .ZN(n7430) );
  NAND3_X1 U9165 ( .A1(n6963), .A2(n6960), .A3(n6962), .ZN(n6957) );
  NAND2_X2 U9166 ( .A1(n14234), .A2(n11853), .ZN(n12153) );
  INV_X1 U9167 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U9168 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8519) );
  OAI21_X2 U9169 ( .B1(n13110), .B2(n6765), .A(n6762), .ZN(n13126) );
  OAI21_X1 U9170 ( .B1(n6765), .B2(n6766), .A(n13128), .ZN(n6763) );
  NAND2_X2 U9171 ( .A1(n10236), .A2(n6472), .ZN(n10230) );
  NAND2_X1 U9172 ( .A1(n13197), .A2(n10230), .ZN(n6769) );
  INV_X1 U9173 ( .A(n6769), .ZN(n10415) );
  NAND2_X1 U9174 ( .A1(n10427), .A2(n6768), .ZN(n10418) );
  NAND2_X1 U9175 ( .A1(n10414), .A2(n6769), .ZN(n6768) );
  NAND2_X1 U9176 ( .A1(n8473), .A2(n8447), .ZN(n9053) );
  NAND2_X1 U9177 ( .A1(n6777), .A2(n6492), .ZN(n6778) );
  OAI21_X1 U9178 ( .B1(n10982), .B2(n6779), .A(n6778), .ZN(n11056) );
  NAND2_X1 U9179 ( .A1(n11056), .A2(n11055), .ZN(n11270) );
  NAND2_X1 U9180 ( .A1(n13236), .A2(n6570), .ZN(n6781) );
  NAND2_X1 U9181 ( .A1(n13236), .A2(n13244), .ZN(n13235) );
  NAND3_X1 U9182 ( .A1(n6782), .A2(n6781), .A3(n6783), .ZN(n13434) );
  NAND3_X1 U9183 ( .A1(n6782), .A2(n6781), .A3(n6505), .ZN(n6788) );
  NAND2_X1 U9184 ( .A1(n11516), .A2(n6790), .ZN(n6789) );
  NAND2_X1 U9185 ( .A1(n6900), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U9186 ( .A1(n6902), .A2(n6901), .ZN(n6793) );
  INV_X1 U9187 ( .A(n7869), .ZN(n6804) );
  NAND2_X1 U9188 ( .A1(n6804), .A2(n6805), .ZN(n7703) );
  INV_X1 U9189 ( .A(n6806), .ZN(n7702) );
  NAND2_X1 U9190 ( .A1(n6893), .A2(n6892), .ZN(n6809) );
  NOR2_X2 U9191 ( .A1(n14428), .A2(n14533), .ZN(n14415) );
  OR2_X2 U9192 ( .A1(n14430), .A2(n14431), .ZN(n14428) );
  NOR2_X2 U9193 ( .A1(n13985), .A2(n6811), .ZN(n13946) );
  NOR2_X4 U9194 ( .A1(n13841), .A2(n13868), .ZN(n13840) );
  INV_X2 U9195 ( .A(n8990), .ZN(n8814) );
  XNOR2_X2 U9196 ( .A(n8483), .B(n8448), .ZN(n10209) );
  NAND2_X1 U9197 ( .A1(n11339), .A2(n6821), .ZN(n11522) );
  NOR2_X2 U9198 ( .A1(n13351), .A2(n12181), .ZN(n6837) );
  NAND2_X1 U9199 ( .A1(n6839), .A2(n10662), .ZN(n10665) );
  OAI21_X1 U9200 ( .B1(n11357), .B2(n11358), .A(n6839), .ZN(n11359) );
  AOI21_X1 U9201 ( .B1(n11956), .B2(n6843), .A(n6841), .ZN(n6840) );
  INV_X1 U9202 ( .A(n6846), .ZN(n6849) );
  NAND2_X1 U9203 ( .A1(n6848), .A2(n6847), .ZN(n11456) );
  NAND2_X1 U9204 ( .A1(n10198), .A2(n6774), .ZN(n10200) );
  OAI21_X1 U9205 ( .B1(n10204), .B2(n10198), .A(n10661), .ZN(n10208) );
  NAND2_X1 U9206 ( .A1(n10204), .A2(n10198), .ZN(n10661) );
  NAND2_X1 U9207 ( .A1(n6854), .A2(n6853), .ZN(n11953) );
  NAND2_X1 U9208 ( .A1(n6522), .A2(n11740), .ZN(n6853) );
  NAND3_X1 U9209 ( .A1(n6857), .A2(n11948), .A3(n6858), .ZN(n6855) );
  NAND3_X1 U9210 ( .A1(n6860), .A2(n6861), .A3(n6859), .ZN(n6857) );
  INV_X1 U9211 ( .A(n11739), .ZN(n6866) );
  NAND2_X1 U9212 ( .A1(n11473), .A2(n6869), .ZN(n6867) );
  NAND2_X1 U9213 ( .A1(n6867), .A2(n6868), .ZN(n11490) );
  AND2_X1 U9214 ( .A1(n6872), .A2(n8473), .ZN(n8451) );
  NAND3_X1 U9215 ( .A1(n6872), .A2(n8452), .A3(n8473), .ZN(n13566) );
  NOR2_X1 U9216 ( .A1(n13243), .A2(n13244), .ZN(n13242) );
  NAND2_X1 U9217 ( .A1(n14387), .A2(n6895), .ZN(n6896) );
  NOR2_X1 U9218 ( .A1(n14388), .A2(n10901), .ZN(n6895) );
  NAND3_X1 U9219 ( .A1(n7696), .A2(n7695), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6900) );
  NAND3_X1 U9220 ( .A1(n7694), .A2(n7693), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n6902) );
  NAND2_X1 U9221 ( .A1(n14781), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14784) );
  NAND3_X1 U9222 ( .A1(n7704), .A2(n7895), .A3(n7703), .ZN(n6921) );
  NAND2_X1 U9223 ( .A1(n6926), .A2(n6925), .ZN(n12010) );
  NOR2_X1 U9224 ( .A1(n6553), .A2(n7042), .ZN(n6925) );
  NAND2_X1 U9225 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n6936) );
  NAND3_X1 U9226 ( .A1(n6944), .A2(n6947), .A3(n6943), .ZN(n6942) );
  NOR2_X1 U9227 ( .A1(n7394), .A2(n7393), .ZN(n7396) );
  INV_X1 U9228 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6943) );
  OAI21_X1 U9229 ( .B1(n7394), .B2(n7393), .A(P3_ADDR_REG_3__SCAN_IN), .ZN(
        n6947) );
  NAND2_X1 U9230 ( .A1(n12848), .A2(n12498), .ZN(n6964) );
  NAND2_X1 U9231 ( .A1(n12858), .A2(n12492), .ZN(n6965) );
  NAND2_X1 U9232 ( .A1(n14975), .A2(n12399), .ZN(n6967) );
  NAND2_X1 U9233 ( .A1(n6968), .A2(n12400), .ZN(n10918) );
  AND2_X2 U9234 ( .A1(n9112), .A2(n9111), .ZN(n14999) );
  NAND2_X1 U9235 ( .A1(n10790), .A2(n6980), .ZN(n6976) );
  NAND2_X1 U9236 ( .A1(n6976), .A2(n6977), .ZN(n14945) );
  AOI21_X1 U9237 ( .B1(n6980), .B2(n6982), .A(n6978), .ZN(n6977) );
  NOR2_X1 U9238 ( .A1(n6981), .A2(n10933), .ZN(n6980) );
  AND2_X1 U9239 ( .A1(n9075), .A2(n6987), .ZN(n6984) );
  NAND2_X1 U9240 ( .A1(n9075), .A2(n7373), .ZN(n6986) );
  NAND2_X1 U9241 ( .A1(n11888), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U9242 ( .A1(n6991), .A2(n6993), .ZN(n12913) );
  OAI21_X1 U9243 ( .B1(n14931), .B2(n7000), .A(n6997), .ZN(n11767) );
  OAI21_X1 U9244 ( .B1(n14931), .B2(n9628), .A(n12437), .ZN(n14206) );
  NAND2_X1 U9245 ( .A1(n12902), .A2(n7012), .ZN(n7011) );
  NAND2_X1 U9246 ( .A1(n12766), .A2(n12769), .ZN(n12768) );
  NAND2_X1 U9247 ( .A1(n9625), .A2(n12429), .ZN(n11244) );
  NOR2_X1 U9248 ( .A1(n12552), .A2(n12551), .ZN(n12559) );
  NAND2_X1 U9249 ( .A1(n9630), .A2(n12459), .ZN(n11888) );
  AOI21_X2 U9250 ( .B1(n12021), .B2(n12020), .A(n13829), .ZN(n14036) );
  NAND2_X1 U9251 ( .A1(n13970), .A2(n13972), .ZN(n13969) );
  AND2_X4 U9252 ( .A1(n7118), .A2(n7117), .ZN(n7677) );
  INV_X4 U9253 ( .A(n9896), .ZN(n8177) );
  OR2_X2 U9254 ( .A1(n14007), .A2(n14092), .ZN(n13985) );
  INV_X1 U9255 ( .A(n7711), .ZN(n7052) );
  NAND2_X1 U9256 ( .A1(n10987), .A2(n10986), .ZN(n10985) );
  NOR2_X1 U9257 ( .A1(n13242), .A2(n7385), .ZN(n11972) );
  XNOR2_X2 U9258 ( .A(n13200), .B(n10654), .ZN(n10198) );
  NAND2_X1 U9259 ( .A1(n11959), .A2(n11958), .ZN(n13337) );
  NAND2_X1 U9260 ( .A1(n9623), .A2(n12409), .ZN(n10790) );
  NAND2_X1 U9261 ( .A1(n7017), .A2(n7903), .ZN(n7015) );
  NAND2_X1 U9262 ( .A1(n7018), .A2(n7887), .ZN(n7017) );
  NAND3_X1 U9263 ( .A1(n7884), .A2(n7885), .A3(n10581), .ZN(n7018) );
  NAND2_X1 U9264 ( .A1(n7022), .A2(n7020), .ZN(n8278) );
  AND2_X1 U9265 ( .A1(n8280), .A2(n7021), .ZN(n7020) );
  NAND2_X1 U9266 ( .A1(n8264), .A2(n7023), .ZN(n7022) );
  INV_X1 U9267 ( .A(n8311), .ZN(n8314) );
  NAND2_X1 U9268 ( .A1(n8002), .A2(n7029), .ZN(n7026) );
  OAI21_X1 U9269 ( .B1(n8002), .B2(n7031), .A(n7029), .ZN(n8020) );
  NAND2_X1 U9270 ( .A1(n7026), .A2(n7027), .ZN(n8019) );
  NAND2_X1 U9271 ( .A1(n7033), .A2(n7039), .ZN(n7032) );
  NAND2_X1 U9272 ( .A1(n8143), .A2(n7036), .ZN(n7033) );
  NAND2_X1 U9273 ( .A1(n7388), .A2(n7035), .ZN(n7034) );
  NAND3_X1 U9274 ( .A1(n7928), .A2(n7927), .A3(n7044), .ZN(n7045) );
  NAND2_X1 U9275 ( .A1(n7943), .A2(n7046), .ZN(n7044) );
  NAND2_X1 U9276 ( .A1(n7045), .A2(n6583), .ZN(n7959) );
  NAND2_X1 U9277 ( .A1(n8084), .A2(n8085), .ZN(n8083) );
  NAND2_X1 U9278 ( .A1(n8248), .A2(n8249), .ZN(n8247) );
  AND3_X2 U9279 ( .A1(n8427), .A2(n7676), .A3(n7685), .ZN(n7384) );
  NAND2_X1 U9280 ( .A1(n7047), .A2(n7048), .ZN(n8344) );
  NAND3_X1 U9281 ( .A1(n8316), .A2(n8315), .A3(n6581), .ZN(n7047) );
  INV_X2 U9282 ( .A(n7706), .ZN(n8501) );
  MUX2_X1 U9283 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7706), .Z(n7705) );
  AOI21_X2 U9284 ( .B1(n7936), .B2(n7718), .A(n7375), .ZN(n7952) );
  NAND2_X1 U9285 ( .A1(n7776), .A2(n7053), .ZN(n7055) );
  NAND2_X1 U9286 ( .A1(n7776), .A2(n7775), .ZN(n8291) );
  NAND3_X1 U9287 ( .A1(n9035), .A2(n9034), .A3(n7061), .ZN(n7060) );
  NAND2_X1 U9288 ( .A1(n8073), .A2(n7072), .ZN(n7067) );
  NAND2_X1 U9289 ( .A1(n7754), .A2(n7076), .ZN(n7075) );
  NOR2_X1 U9290 ( .A1(n7759), .A2(n7761), .ZN(n7080) );
  NOR2_X1 U9291 ( .A1(n10278), .A2(n9705), .ZN(P1_U4016) );
  NAND3_X1 U9292 ( .A1(n7088), .A2(n7087), .A3(n7085), .ZN(n10853) );
  XNOR2_X1 U9293 ( .A(n7086), .B(n6605), .ZN(n10819) );
  INV_X1 U9294 ( .A(n10804), .ZN(n7087) );
  NAND2_X1 U9295 ( .A1(n10805), .A2(n10806), .ZN(n7088) );
  NAND2_X1 U9296 ( .A1(n13619), .A2(n7092), .ZN(n7089) );
  NAND2_X1 U9297 ( .A1(n7089), .A2(n7090), .ZN(n13584) );
  NAND2_X1 U9298 ( .A1(n7096), .A2(n12057), .ZN(n14254) );
  NAND2_X1 U9299 ( .A1(n13645), .A2(n7099), .ZN(n7097) );
  NAND2_X2 U9300 ( .A1(n13637), .A2(n13636), .ZN(n13635) );
  AND2_X1 U9301 ( .A1(n7687), .A2(n7106), .ZN(n8420) );
  NAND2_X1 U9302 ( .A1(n7687), .A2(n7104), .ZN(n8424) );
  INV_X1 U9303 ( .A(n8424), .ZN(n8425) );
  INV_X1 U9304 ( .A(n7116), .ZN(n11556) );
  AND2_X1 U9305 ( .A1(n7863), .A2(n7669), .ZN(n7898) );
  AND4_X2 U9306 ( .A1(n7863), .A2(n7668), .A3(n7670), .A4(n7667), .ZN(n7118)
         );
  INV_X1 U9307 ( .A(n9146), .ZN(n7119) );
  OAI211_X1 U9308 ( .C1(n12374), .C2(n7132), .A(n7127), .B(n7125), .ZN(n12272)
         );
  NAND2_X1 U9309 ( .A1(n12374), .A2(n7126), .ZN(n7125) );
  NOR2_X1 U9310 ( .A1(n12265), .A2(n7129), .ZN(n7126) );
  INV_X1 U9311 ( .A(n12265), .ZN(n7130) );
  OAI21_X1 U9312 ( .B1(n12265), .B2(n12276), .A(n7133), .ZN(n7131) );
  NAND2_X1 U9313 ( .A1(n12265), .A2(n12276), .ZN(n7132) );
  XNOR2_X1 U9314 ( .A(n14992), .B(n10097), .ZN(n7134) );
  NAND3_X1 U9315 ( .A1(n10122), .A2(n10099), .A3(n14995), .ZN(n10121) );
  NOR2_X1 U9316 ( .A1(n10100), .A2(n10098), .ZN(n10122) );
  NAND2_X1 U9317 ( .A1(n10089), .A2(n13047), .ZN(n10092) );
  INV_X1 U9318 ( .A(n13047), .ZN(n9657) );
  INV_X1 U9319 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7142) );
  NOR2_X1 U9320 ( .A1(n12327), .A2(n7377), .ZN(n12364) );
  NAND2_X1 U9321 ( .A1(n9273), .A2(n7157), .ZN(n7156) );
  OAI21_X1 U9322 ( .B1(n7167), .B2(n10506), .A(n7166), .ZN(n10509) );
  NAND3_X1 U9323 ( .A1(n10308), .A2(n10309), .A3(n10505), .ZN(n7166) );
  NAND3_X1 U9324 ( .A1(n7175), .A2(n12753), .A3(n12769), .ZN(n12522) );
  NAND3_X1 U9325 ( .A1(n12512), .A2(n12513), .A3(n12511), .ZN(n7176) );
  OAI211_X1 U9326 ( .C1(n10583), .C2(n7185), .A(n7183), .B(n10595), .ZN(n10598) );
  NAND2_X1 U9327 ( .A1(n10584), .A2(n7184), .ZN(n7183) );
  INV_X1 U9328 ( .A(n14420), .ZN(n7185) );
  NAND2_X1 U9329 ( .A1(n7187), .A2(n10583), .ZN(n10594) );
  OAI21_X1 U9330 ( .B1(n11004), .B2(n7189), .A(n7191), .ZN(n11367) );
  NAND2_X1 U9331 ( .A1(n7190), .A2(n7188), .ZN(n11369) );
  NAND2_X1 U9332 ( .A1(n11004), .A2(n7191), .ZN(n7190) );
  OAI21_X1 U9333 ( .B1(n11004), .B2(n11007), .A(n7195), .ZN(n11228) );
  NOR2_X1 U9334 ( .A1(n13972), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U9335 ( .A1(n7198), .A2(n7196), .ZN(n13960) );
  OAI21_X1 U9336 ( .B1(n13972), .B2(n7199), .A(n11994), .ZN(n7197) );
  OAI21_X2 U9337 ( .B1(n13906), .B2(n7204), .A(n7203), .ZN(n13879) );
  OAI21_X2 U9338 ( .B1(n7387), .B2(n7210), .A(n7208), .ZN(n14001) );
  NAND2_X1 U9339 ( .A1(n7677), .A2(n7384), .ZN(n7795) );
  NAND3_X1 U9340 ( .A1(n7677), .A2(n7384), .A3(n7213), .ZN(n7679) );
  AND3_X2 U9341 ( .A1(n7677), .A2(n7384), .A3(n6572), .ZN(n14111) );
  NAND2_X1 U9342 ( .A1(n11937), .A2(n7220), .ZN(n7217) );
  NAND2_X1 U9343 ( .A1(n7218), .A2(n7217), .ZN(n13265) );
  NAND2_X1 U9344 ( .A1(n7228), .A2(n11467), .ZN(n7225) );
  NAND2_X1 U9345 ( .A1(n8473), .A2(n7232), .ZN(n8485) );
  INV_X1 U9346 ( .A(n11356), .ZN(n14693) );
  NAND2_X1 U9347 ( .A1(n11514), .A2(n6536), .ZN(n11516) );
  INV_X1 U9348 ( .A(n13386), .ZN(n7244) );
  NOR2_X1 U9349 ( .A1(n13385), .A2(n7253), .ZN(n13364) );
  NAND3_X1 U9350 ( .A1(n7257), .A2(n9001), .A3(n7258), .ZN(n9009) );
  NAND3_X1 U9351 ( .A1(n8949), .A2(n7260), .A3(n8982), .ZN(n7257) );
  NAND3_X1 U9352 ( .A1(n8873), .A2(n8872), .A3(n6585), .ZN(n7268) );
  INV_X1 U9353 ( .A(n8886), .ZN(n7269) );
  NAND3_X1 U9354 ( .A1(n8904), .A2(n8903), .A3(n6586), .ZN(n7271) );
  INV_X1 U9355 ( .A(n8916), .ZN(n7272) );
  NAND3_X1 U9356 ( .A1(n8842), .A2(n8841), .A3(n6587), .ZN(n7274) );
  INV_X1 U9357 ( .A(n8853), .ZN(n7275) );
  NAND2_X1 U9358 ( .A1(n7276), .A2(n7277), .ZN(n8594) );
  NAND3_X1 U9359 ( .A1(n8558), .A2(n6579), .A3(n8557), .ZN(n7276) );
  NAND3_X1 U9360 ( .A1(n8672), .A2(n6580), .A3(n8671), .ZN(n7278) );
  NAND2_X1 U9361 ( .A1(n7278), .A2(n7279), .ZN(n8703) );
  NAND2_X1 U9362 ( .A1(n7280), .A2(n7282), .ZN(n8553) );
  NAND3_X1 U9363 ( .A1(n7379), .A2(n8525), .A3(n7281), .ZN(n7280) );
  NAND3_X1 U9364 ( .A1(n8651), .A2(n8650), .A3(n6578), .ZN(n7284) );
  NAND2_X1 U9365 ( .A1(n7284), .A2(n7285), .ZN(n8667) );
  XNOR2_X2 U9366 ( .A(n7287), .B(n8452), .ZN(n8455) );
  NAND3_X1 U9367 ( .A1(n8599), .A2(n6584), .A3(n8598), .ZN(n7288) );
  NAND2_X1 U9368 ( .A1(n7288), .A2(n7289), .ZN(n8631) );
  OAI22_X1 U9369 ( .A1(n8793), .A2(n7291), .B1(n8804), .B2(n7292), .ZN(n8820)
         );
  INV_X1 U9370 ( .A(n8804), .ZN(n7294) );
  XNOR2_X2 U9371 ( .A(n10426), .B(n10654), .ZN(n10248) );
  NAND2_X2 U9372 ( .A1(n10245), .A2(n10244), .ZN(n10426) );
  NAND2_X2 U9373 ( .A1(n13217), .A2(n10203), .ZN(n10245) );
  NAND2_X1 U9374 ( .A1(n7309), .A2(n10413), .ZN(n10428) );
  INV_X1 U9375 ( .A(n13092), .ZN(n7316) );
  OAI21_X2 U9376 ( .B1(n13092), .B2(n6564), .A(n6500), .ZN(n13060) );
  NAND2_X1 U9377 ( .A1(n7330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U9378 ( .A1(n8467), .A2(n7331), .ZN(n7330) );
  NAND2_X1 U9379 ( .A1(n10481), .A2(n10482), .ZN(n10539) );
  NAND2_X1 U9380 ( .A1(n10717), .A2(n10716), .ZN(n10719) );
  AND2_X1 U9381 ( .A1(n7336), .A2(n8519), .ZN(n7337) );
  NAND3_X1 U9382 ( .A1(n7338), .A2(n7339), .A3(n7337), .ZN(n8713) );
  INV_X1 U9383 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7341) );
  NAND2_X1 U9384 ( .A1(n12817), .A2(n7343), .ZN(n7342) );
  NAND2_X1 U9385 ( .A1(n14934), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U9386 ( .A1(n11828), .A2(n9353), .ZN(n11827) );
  NAND2_X1 U9387 ( .A1(n9410), .A2(n6504), .ZN(n12894) );
  NAND2_X1 U9388 ( .A1(n9620), .A2(n15001), .ZN(n7366) );
  NAND2_X1 U9389 ( .A1(n7366), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U9390 ( .A1(n7366), .A2(n7362), .ZN(n9702) );
  AND2_X1 U9391 ( .A1(n7366), .A2(n7368), .ZN(n11980) );
  NAND2_X1 U9392 ( .A1(n7363), .A2(n7367), .ZN(n9691) );
  AND2_X2 U9393 ( .A1(n11087), .A2(n9249), .ZN(n11246) );
  NAND2_X1 U9394 ( .A1(n14946), .A2(n7371), .ZN(n11087) );
  NAND2_X1 U9395 ( .A1(n11236), .A2(n11235), .ZN(n11375) );
  OR2_X2 U9396 ( .A1(n10637), .A2(n10636), .ZN(n14446) );
  NAND2_X1 U9397 ( .A1(n9417), .A2(n9416), .ZN(n9432) );
  NAND2_X1 U9398 ( .A1(n9326), .A2(n9325), .ZN(n9337) );
  NAND2_X1 U9399 ( .A1(n10277), .A2(n10807), .ZN(n10280) );
  NAND2_X1 U9400 ( .A1(n10811), .A2(n13688), .ZN(n10279) );
  NAND2_X1 U9401 ( .A1(n11757), .A2(n11756), .ZN(n12233) );
  NAND2_X1 U9402 ( .A1(n8332), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7846) );
  INV_X1 U9403 ( .A(n12233), .ZN(n11759) );
  NAND2_X1 U9404 ( .A1(n10280), .A2(n10279), .ZN(n10283) );
  INV_X1 U9405 ( .A(n7687), .ZN(n8429) );
  INV_X1 U9406 ( .A(n8343), .ZN(n8349) );
  NAND2_X1 U9407 ( .A1(n13440), .A2(n6534), .ZN(n13236) );
  NOR2_X1 U9408 ( .A1(n10319), .A2(n10318), .ZN(n10320) );
  NAND2_X1 U9409 ( .A1(n10696), .A2(n10695), .ZN(n10982) );
  OR2_X1 U9410 ( .A1(n13200), .A2(n10654), .ZN(n10655) );
  INV_X1 U9411 ( .A(n8631), .ZN(n8634) );
  AND2_X1 U9412 ( .A1(n8748), .A2(n8799), .ZN(n13201) );
  NAND2_X1 U9413 ( .A1(n9020), .A2(n8489), .ZN(n8492) );
  NAND2_X1 U9414 ( .A1(n10096), .A2(n14992), .ZN(n9621) );
  INV_X1 U9415 ( .A(n9118), .ZN(n10096) );
  NAND2_X1 U9416 ( .A1(n10202), .A2(n6472), .ZN(n10828) );
  NAND2_X1 U9417 ( .A1(n9084), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9085) );
  AND4_X2 U9418 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n14997)
         );
  OR2_X1 U9419 ( .A1(n9157), .A2(n7575), .ZN(n9123) );
  NAND2_X1 U9420 ( .A1(n9086), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9122) );
  OAI21_X2 U9421 ( .B1(n13084), .B2(n13083), .A(n12192), .ZN(n12194) );
  NAND2_X1 U9422 ( .A1(n13257), .A2(n13256), .ZN(n13440) );
  AND2_X1 U9423 ( .A1(n13406), .A2(n13217), .ZN(n13422) );
  NAND2_X1 U9424 ( .A1(n13217), .A2(n6472), .ZN(n10232) );
  AND2_X1 U9425 ( .A1(n10683), .A2(n10690), .ZN(n7374) );
  INV_X1 U9426 ( .A(n13881), .ZN(n13894) );
  INV_X2 U9427 ( .A(n15010), .ZN(n15012) );
  NAND2_X2 U9428 ( .A1(n10340), .A2(n14978), .ZN(n15010) );
  INV_X1 U9429 ( .A(n12996), .ZN(n9689) );
  NOR2_X1 U9430 ( .A1(n7717), .A2(n7716), .ZN(n7375) );
  AND3_X1 U9431 ( .A1(n14982), .A2(n12396), .A3(n12395), .ZN(n7376) );
  AND2_X1 U9432 ( .A1(n12235), .A2(n12602), .ZN(n7377) );
  NOR2_X1 U9433 ( .A1(n7724), .A2(n7723), .ZN(n7378) );
  XNOR2_X1 U9434 ( .A(n12197), .B(n6588), .ZN(n13066) );
  OR2_X1 U9435 ( .A1(n9770), .A2(n14600), .ZN(n7381) );
  AND2_X1 U9436 ( .A1(n8178), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7382) );
  INV_X1 U9437 ( .A(n10241), .ZN(n8489) );
  AND2_X1 U9438 ( .A1(n13240), .A2(n13172), .ZN(n7385) );
  AND2_X1 U9439 ( .A1(n7741), .A2(n7740), .ZN(n7386) );
  AND2_X1 U9440 ( .A1(n8145), .A2(n8144), .ZN(n7388) );
  XNOR2_X1 U9441 ( .A(n8466), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10202) );
  AND2_X2 U9442 ( .A1(n10823), .A2(n13414), .ZN(n13402) );
  INV_X2 U9443 ( .A(n13402), .ZN(n13406) );
  AND2_X1 U9444 ( .A1(n12791), .A2(n12802), .ZN(n7390) );
  INV_X1 U9445 ( .A(n12769), .ZN(n9573) );
  INV_X1 U9446 ( .A(n12845), .ZN(n12818) );
  NAND2_X1 U9447 ( .A1(n9500), .A2(n9499), .ZN(n12831) );
  INV_X1 U9448 ( .A(n12831), .ZN(n12857) );
  NAND2_X1 U9449 ( .A1(n10241), .A2(n8490), .ZN(n8491) );
  OR2_X1 U9450 ( .A1(n7852), .A2(n7882), .ZN(n7853) );
  NAND2_X1 U9451 ( .A1(n8512), .A2(n8511), .ZN(n8524) );
  INV_X1 U9452 ( .A(n8632), .ZN(n8633) );
  INV_X1 U9453 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9072) );
  INV_X1 U9454 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9069) );
  INV_X1 U9455 ( .A(n12897), .ZN(n9429) );
  INV_X1 U9456 ( .A(n12753), .ZN(n9586) );
  NOR3_X1 U9457 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_13__SCAN_IN), .ZN(n8443) );
  AOI22_X1 U9458 ( .A1(n10637), .A2(n10807), .B1(n10811), .B2(n14354), .ZN(
        n10371) );
  INV_X1 U9459 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7695) );
  INV_X1 U9460 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9478) );
  INV_X1 U9461 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n11760) );
  OAI21_X1 U9462 ( .B1(n12843), .B2(n9502), .A(n9501), .ZN(n12829) );
  INV_X1 U9463 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U9464 ( .A1(n11246), .A2(n12427), .ZN(n11245) );
  INV_X1 U9465 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8751) );
  OR2_X1 U9466 ( .A1(n13468), .A2(n13177), .ZN(n11934) );
  NOR2_X1 U9467 ( .A1(n8474), .A2(n8728), .ZN(n8475) );
  INV_X1 U9468 ( .A(n7828), .ZN(n8350) );
  INV_X1 U9469 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7944) );
  INV_X1 U9470 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U9471 ( .A1(n10943), .A2(n12609), .ZN(n10944) );
  NAND2_X1 U9472 ( .A1(n11755), .A2(n12604), .ZN(n11756) );
  OR2_X1 U9473 ( .A1(n9566), .A2(n9565), .ZN(n9581) );
  OR2_X1 U9474 ( .A1(n9494), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9508) );
  NAND2_X1 U9475 ( .A1(n9103), .A2(n9727), .ZN(n9113) );
  NOR2_X1 U9476 ( .A1(n9306), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9314) );
  INV_X1 U9477 ( .A(n13045), .ZN(n10332) );
  AND2_X1 U9478 ( .A1(n9301), .A2(n9300), .ZN(n9328) );
  INV_X1 U9479 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9167) );
  INV_X1 U9480 ( .A(n14231), .ZN(n11852) );
  INV_X1 U9481 ( .A(n10877), .ZN(n10874) );
  NOR2_X1 U9482 ( .A1(n8907), .A2(n8906), .ZN(n8919) );
  INV_X1 U9483 ( .A(n8855), .ZN(n8856) );
  OR2_X1 U9484 ( .A1(n8655), .A2(n8654), .ZN(n8674) );
  INV_X1 U9485 ( .A(n11965), .ZN(n11966) );
  INV_X1 U9486 ( .A(n13163), .ZN(n13141) );
  AND2_X1 U9487 ( .A1(n8446), .A2(n9048), .ZN(n8447) );
  INV_X1 U9488 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U9489 ( .A1(n12053), .A2(n12052), .ZN(n12057) );
  OAI21_X1 U9490 ( .B1(n6473), .B2(n10291), .A(n10290), .ZN(n10319) );
  INV_X1 U9491 ( .A(n13605), .ZN(n12083) );
  NAND2_X1 U9492 ( .A1(n14448), .A2(n13964), .ZN(n10466) );
  NAND2_X1 U9493 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  INV_X1 U9494 ( .A(n8267), .ZN(n8285) );
  OR2_X1 U9495 ( .A1(n8183), .A2(n8166), .ZN(n8199) );
  INV_X1 U9496 ( .A(n8332), .ZN(n7876) );
  AND2_X1 U9497 ( .A1(n10969), .A2(n10968), .ZN(n10971) );
  NAND2_X1 U9498 ( .A1(n10580), .A2(n10579), .ZN(n10630) );
  AND2_X1 U9499 ( .A1(n11297), .A2(n13897), .ZN(n10275) );
  INV_X1 U9500 ( .A(n10466), .ZN(n10557) );
  INV_X1 U9501 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8433) );
  INV_X1 U9502 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U9503 ( .A1(n7755), .A2(n10465), .ZN(n7758) );
  NAND2_X1 U9504 ( .A1(n7952), .A2(n7719), .ZN(n7969) );
  AND2_X1 U9505 ( .A1(n7429), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n7409) );
  INV_X1 U9506 ( .A(n11632), .ZN(n9667) );
  NOR2_X1 U9507 ( .A1(n9442), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U9508 ( .A1(n9404), .A2(n9403), .ZN(n9422) );
  OR2_X1 U9509 ( .A1(n10395), .A2(n14983), .ZN(n10396) );
  AND2_X1 U9510 ( .A1(n12593), .A2(n10110), .ZN(n10115) );
  NAND2_X1 U9511 ( .A1(n10115), .A2(n10114), .ZN(n12380) );
  NOR2_X1 U9512 ( .A1(n9581), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U9513 ( .A1(n11138), .A2(n14792), .ZN(n11139) );
  INV_X1 U9514 ( .A(n12872), .ZN(n12846) );
  AND2_X1 U9515 ( .A1(n12469), .A2(n12468), .ZN(n12923) );
  INV_X1 U9516 ( .A(n12595), .ZN(n9644) );
  AND2_X1 U9517 ( .A1(n13047), .A2(n13045), .ZN(n9696) );
  INV_X1 U9518 ( .A(n6480), .ZN(n9439) );
  INV_X1 U9519 ( .A(n14965), .ZN(n14998) );
  INV_X1 U9520 ( .A(n12432), .ZN(n11249) );
  INV_X1 U9521 ( .A(n15001), .ZN(n14988) );
  AND2_X1 U9522 ( .A1(n9643), .A2(n9683), .ZN(n15004) );
  AND2_X1 U9523 ( .A1(n9431), .A2(n9415), .ZN(n9416) );
  AND2_X1 U9524 ( .A1(n9293), .A2(n9271), .ZN(n9272) );
  INV_X1 U9525 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8721) );
  INV_X1 U9526 ( .A(n10418), .ZN(n10419) );
  AND2_X1 U9527 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  NAND2_X1 U9528 ( .A1(n8843), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8855) );
  AND2_X1 U9529 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  INV_X1 U9530 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11855) );
  AOI21_X1 U9531 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9038) );
  AND2_X1 U9532 ( .A1(n8826), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8843) );
  INV_X1 U9533 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11107) );
  OR2_X1 U9534 ( .A1(n9787), .A2(n11973), .ZN(n14668) );
  INV_X1 U9535 ( .A(n13227), .ZN(n13223) );
  OR2_X1 U9536 ( .A1(n11520), .A2(n13188), .ZN(n11515) );
  INV_X1 U9537 ( .A(n11059), .ZN(n11055) );
  NAND2_X1 U9538 ( .A1(n13406), .A2(n10993), .ZN(n13417) );
  INV_X1 U9539 ( .A(n13468), .ZN(n13311) );
  NAND2_X1 U9540 ( .A1(n14746), .A2(n8479), .ZN(n10238) );
  NOR2_X1 U9541 ( .A1(n8064), .A2(n8063), .ZN(n8096) );
  AND2_X1 U9542 ( .A1(n11705), .A2(n11703), .ZN(n11704) );
  INV_X1 U9543 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8128) );
  INV_X1 U9544 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13639) );
  NAND2_X1 U9545 ( .A1(n12084), .A2(n12086), .ZN(n12087) );
  INV_X1 U9546 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8115) );
  INV_X1 U9547 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9980) );
  INV_X1 U9548 ( .A(n14019), .ZN(n13824) );
  NAND2_X1 U9549 ( .A1(n14045), .A2(n13667), .ZN(n12018) );
  INV_X1 U9550 ( .A(n11865), .ZN(n11869) );
  INV_X1 U9551 ( .A(n10596), .ZN(n10766) );
  INV_X1 U9552 ( .A(n14388), .ZN(n14386) );
  AND2_X1 U9553 ( .A1(n10297), .A2(n10296), .ZN(n10556) );
  OR2_X1 U9554 ( .A1(n10337), .A2(n10012), .ZN(n10018) );
  AND3_X2 U9555 ( .A1(n9152), .A2(n9151), .A3(n9150), .ZN(n14970) );
  INV_X1 U9556 ( .A(n9103), .ZN(n10013) );
  AND2_X1 U9557 ( .A1(n10115), .A2(n10111), .ZN(n12355) );
  AND2_X1 U9558 ( .A1(n10725), .A2(n12723), .ZN(n14979) );
  AND2_X1 U9559 ( .A1(n9515), .A2(n9514), .ZN(n12845) );
  AND3_X1 U9560 ( .A1(n9374), .A2(n9373), .A3(n9372), .ZN(n12921) );
  INV_X1 U9561 ( .A(n14896), .ZN(n14926) );
  AND2_X1 U9562 ( .A1(n10018), .A2(n10016), .ZN(n10035) );
  AND2_X1 U9563 ( .A1(n12525), .A2(n10111), .ZN(n14965) );
  AND2_X1 U9564 ( .A1(n15010), .A2(n14953), .ZN(n12930) );
  AND2_X1 U9565 ( .A1(n12433), .A2(n9268), .ZN(n12427) );
  INV_X1 U9566 ( .A(n14978), .ZN(n15007) );
  NAND2_X1 U9567 ( .A1(n9644), .A2(n12393), .ZN(n15047) );
  NOR2_X1 U9568 ( .A1(n9680), .A2(n9696), .ZN(n10335) );
  NAND2_X1 U9569 ( .A1(n15004), .A2(n15049), .ZN(n15063) );
  INV_X1 U9570 ( .A(n15049), .ZN(n15058) );
  INV_X1 U9571 ( .A(n9616), .ZN(n12627) );
  INV_X1 U9572 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9300) );
  OR2_X1 U9573 ( .A1(n8722), .A2(n8721), .ZN(n8766) );
  AND2_X1 U9574 ( .A1(n10237), .A2(n10233), .ZN(n14237) );
  INV_X1 U9575 ( .A(n13168), .ZN(n14235) );
  AND2_X1 U9576 ( .A1(n10232), .A2(n10236), .ZN(n14735) );
  AND4_X1 U9577 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n12218)
         );
  OR2_X1 U9578 ( .A1(n8966), .A2(n11043), .ZN(n8532) );
  OR2_X1 U9579 ( .A1(n8526), .A2(n9777), .ZN(n8497) );
  INV_X1 U9580 ( .A(n14668), .ZN(n14658) );
  AND2_X1 U9581 ( .A1(n9773), .A2(n11973), .ZN(n14655) );
  XNOR2_X1 U9582 ( .A(n13230), .B(n13223), .ZN(n13224) );
  NAND2_X1 U9583 ( .A1(n13392), .A2(n13393), .ZN(n13391) );
  NAND2_X2 U9584 ( .A1(n10239), .A2(n14686), .ZN(n13414) );
  OR2_X1 U9585 ( .A1(n10828), .A2(n10205), .ZN(n14739) );
  INV_X1 U9586 ( .A(n13541), .ZN(n13529) );
  INV_X1 U9587 ( .A(n14739), .ZN(n14746) );
  AND2_X1 U9588 ( .A1(n9706), .A2(n9768), .ZN(n10224) );
  AND2_X1 U9589 ( .A1(n9894), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10328) );
  AND2_X1 U9590 ( .A1(n8160), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U9591 ( .A1(n8181), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8183) );
  AND2_X1 U9592 ( .A1(n14352), .A2(n14549), .ZN(n14297) );
  AND2_X1 U9593 ( .A1(n8208), .A2(n8207), .ZN(n13614) );
  OR2_X1 U9594 ( .A1(n10074), .A2(n10294), .ZN(n14380) );
  AND2_X1 U9595 ( .A1(n9920), .A2(n14122), .ZN(n14375) );
  INV_X1 U9596 ( .A(n14370), .ZN(n13811) );
  INV_X1 U9597 ( .A(n14492), .ZN(n14448) );
  INV_X1 U9598 ( .A(n13923), .ZN(n14453) );
  INV_X1 U9599 ( .A(n14444), .ZN(n14396) );
  AOI21_X1 U9600 ( .B1(n10327), .B2(n10261), .A(n10260), .ZN(n10554) );
  INV_X1 U9601 ( .A(n14549), .ZN(n14570) );
  INV_X1 U9602 ( .A(n14522), .ZN(n14566) );
  NAND2_X1 U9603 ( .A1(n10472), .A2(n10471), .ZN(n14522) );
  AND2_X1 U9604 ( .A1(n10467), .A2(n10556), .ZN(n11684) );
  AND2_X1 U9605 ( .A1(n8157), .A2(n8175), .ZN(n13789) );
  AND2_X1 U9606 ( .A1(n10018), .A2(n10017), .ZN(n14899) );
  INV_X1 U9607 ( .A(n12383), .ZN(n10956) );
  AND2_X1 U9608 ( .A1(n10108), .A2(n10107), .ZN(n12371) );
  NAND2_X1 U9609 ( .A1(n9530), .A2(n9529), .ZN(n12832) );
  INV_X1 U9610 ( .A(n12886), .ZN(n12910) );
  INV_X1 U9611 ( .A(n14899), .ZN(n14930) );
  INV_X1 U9612 ( .A(n14892), .ZN(n14915) );
  NAND2_X1 U9613 ( .A1(n10035), .A2(n10015), .ZN(n14921) );
  OR2_X1 U9614 ( .A1(n14939), .A2(n15047), .ZN(n12928) );
  NAND2_X1 U9615 ( .A1(n15079), .A2(n15015), .ZN(n12996) );
  INV_X1 U9616 ( .A(n15079), .ZN(n15077) );
  NAND2_X1 U9617 ( .A1(n9600), .A2(n13000), .ZN(n9703) );
  AND2_X1 U9618 ( .A1(n9701), .A2(n9700), .ZN(n15064) );
  NAND2_X1 U9619 ( .A1(n9658), .A2(n13046), .ZN(n9824) );
  INV_X1 U9620 ( .A(SI_25_), .ZN(n11631) );
  INV_X1 U9621 ( .A(SI_20_), .ZN(n10724) );
  INV_X1 U9622 ( .A(SI_15_), .ZN(n9898) );
  INV_X1 U9623 ( .A(SI_10_), .ZN(n9740) );
  NAND2_X1 U9624 ( .A1(n10421), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14243) );
  INV_X1 U9625 ( .A(n12157), .ZN(n13516) );
  INV_X1 U9626 ( .A(n12181), .ZN(n13490) );
  OR3_X1 U9627 ( .A1(n10229), .A2(n10228), .A3(n14735), .ZN(n13168) );
  INV_X1 U9628 ( .A(n11854), .ZN(n13185) );
  INV_X1 U9629 ( .A(n14655), .ZN(n14670) );
  INV_X1 U9630 ( .A(n14673), .ZN(n14644) );
  INV_X1 U9631 ( .A(n13409), .ZN(n13375) );
  OR3_X1 U9632 ( .A1(n10653), .A2(n10652), .A3(n14681), .ZN(n14766) );
  OR2_X1 U9633 ( .A1(n10653), .A2(n10821), .ZN(n14755) );
  OR2_X1 U9634 ( .A1(n14683), .A2(n14679), .ZN(n14680) );
  INV_X1 U9635 ( .A(n14686), .ZN(n14683) );
  INV_X1 U9636 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13580) );
  INV_X1 U9637 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10221) );
  INV_X1 U9638 ( .A(n14297), .ZN(n14286) );
  AND2_X1 U9639 ( .A1(n10730), .A2(n11622), .ZN(n14367) );
  OR2_X1 U9640 ( .A1(n8100), .A2(n8099), .ZN(n13676) );
  INV_X1 U9641 ( .A(n14375), .ZN(n13767) );
  OR2_X1 U9642 ( .A1(n13845), .A2(n13964), .ZN(n13917) );
  INV_X1 U9643 ( .A(n14010), .ZN(n14395) );
  OR2_X1 U9644 ( .A1(n14395), .A2(n14566), .ZN(n13955) );
  AND2_X2 U9645 ( .A1(n11684), .A2(n10554), .ZN(n14594) );
  AND4_X1 U9646 ( .A1(n14539), .A2(n14538), .A3(n14537), .A4(n14536), .ZN(
        n14587) );
  AND2_X2 U9647 ( .A1(n11684), .A2(n11683), .ZN(n14578) );
  NOR2_X2 U9648 ( .A1(n10327), .A2(n7082), .ZN(n14472) );
  CLKBUF_X1 U9649 ( .A(n14472), .Z(n14488) );
  INV_X1 U9650 ( .A(n8363), .ZN(n14131) );
  INV_X1 U9651 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10678) );
  INV_X1 U9652 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9903) );
  AND2_X2 U9653 ( .A1(n13046), .A2(n9708), .ZN(P3_U3897) );
  INV_X1 U9654 ( .A(n13199), .ZN(P2_U3947) );
  INV_X1 U9655 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12679) );
  NAND2_X1 U9656 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12679), .ZN(n7420) );
  INV_X1 U9657 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7391) );
  AOI22_X1 U9658 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n7391), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n12679), .ZN(n7485) );
  INV_X1 U9659 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n7417) );
  XOR2_X1 U9660 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n7426) );
  INV_X1 U9661 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7414) );
  INV_X1 U9662 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7412) );
  INV_X1 U9663 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7407) );
  INV_X1 U9664 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7406) );
  XNOR2_X1 U9665 ( .A(n7392), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n7432) );
  NOR2_X1 U9666 ( .A1(n7399), .A2(n6938), .ZN(n7401) );
  NOR2_X1 U9667 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7447), .ZN(n7400) );
  XNOR2_X1 U9668 ( .A(n7402), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n7453) );
  NOR2_X1 U9669 ( .A1(n7403), .A2(n6750), .ZN(n7405) );
  NOR2_X1 U9670 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7456), .ZN(n7404) );
  XNOR2_X1 U9671 ( .A(n7406), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n7460) );
  XNOR2_X1 U9672 ( .A(n7407), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n7465) );
  NOR2_X1 U9673 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n7408), .ZN(n7410) );
  XOR2_X1 U9674 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n7408), .Z(n7429) );
  XNOR2_X1 U9675 ( .A(n7412), .B(P3_ADDR_REG_11__SCAN_IN), .ZN(n7469) );
  XNOR2_X1 U9676 ( .A(n7414), .B(P3_ADDR_REG_12__SCAN_IN), .ZN(n7475) );
  INV_X1 U9677 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n11724) );
  AND2_X1 U9678 ( .A1(n11724), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7415) );
  INV_X1 U9679 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U9680 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12651), .ZN(n7418) );
  INV_X1 U9681 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U9682 ( .A1(n7483), .A2(n7418), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n14385), .ZN(n7486) );
  NAND2_X1 U9683 ( .A1(n7485), .A2(n7486), .ZN(n7419) );
  NAND2_X1 U9684 ( .A1(n7420), .A2(n7419), .ZN(n7421) );
  NOR2_X1 U9685 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n7421), .ZN(n7423) );
  INV_X1 U9686 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14176) );
  XNOR2_X1 U9687 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7421), .ZN(n7424) );
  NOR2_X1 U9688 ( .A1(n14176), .A2(n7424), .ZN(n7422) );
  NOR2_X1 U9689 ( .A1(n7423), .A2(n7422), .ZN(n7492) );
  XOR2_X1 U9690 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n7491) );
  XOR2_X1 U9691 ( .A(n7492), .B(n7491), .Z(n14136) );
  XOR2_X1 U9692 ( .A(n14176), .B(n7424), .Z(n14165) );
  INV_X1 U9693 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14651) );
  XOR2_X1 U9694 ( .A(n7426), .B(n7425), .Z(n14340) );
  INV_X1 U9695 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7482) );
  XOR2_X1 U9696 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(n11724), .Z(n7428) );
  XOR2_X1 U9697 ( .A(n7428), .B(n7427), .Z(n14336) );
  INV_X1 U9698 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14929) );
  XOR2_X1 U9699 ( .A(n7429), .B(n14929), .Z(n14154) );
  NAND2_X1 U9700 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n7431), .ZN(n7446) );
  XNOR2_X1 U9701 ( .A(n6569), .B(n7432), .ZN(n14141) );
  XNOR2_X1 U9702 ( .A(n7434), .B(n7433), .ZN(n7436) );
  NAND2_X1 U9703 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n7436), .ZN(n7438) );
  AOI21_X1 U9704 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14780), .A(n7435), .ZN(
        n15084) );
  INV_X1 U9705 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15083) );
  NOR2_X1 U9706 ( .A1(n15084), .A2(n15083), .ZN(n15091) );
  NAND2_X1 U9707 ( .A1(n7438), .A2(n7437), .ZN(n14142) );
  AND2_X1 U9708 ( .A1(n14141), .A2(n14142), .ZN(n7440) );
  NOR2_X1 U9709 ( .A1(n14141), .A2(n14142), .ZN(n14140) );
  INV_X1 U9710 ( .A(n14140), .ZN(n7439) );
  OAI21_X1 U9711 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n7440), .A(n7439), .ZN(
        n7442) );
  XOR2_X1 U9712 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n7441), .Z(n7443) );
  AND2_X1 U9713 ( .A1(n7442), .A2(n7443), .ZN(n15088) );
  NOR2_X1 U9714 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15087), .ZN(n7444) );
  NAND2_X1 U9715 ( .A1(n15081), .A2(n15080), .ZN(n7445) );
  NAND2_X1 U9716 ( .A1(n7446), .A2(n7445), .ZN(n7449) );
  NOR2_X1 U9717 ( .A1(n7449), .A2(n7448), .ZN(n7451) );
  XNOR2_X1 U9718 ( .A(n7449), .B(n7448), .ZN(n15082) );
  NOR2_X1 U9719 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15082), .ZN(n7450) );
  NAND2_X1 U9720 ( .A1(n7452), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7455) );
  XNOR2_X1 U9721 ( .A(n7454), .B(n7453), .ZN(n14144) );
  NOR2_X1 U9722 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n7457), .ZN(n7459) );
  XNOR2_X1 U9723 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7456), .ZN(n15086) );
  XNOR2_X1 U9724 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n7457), .ZN(n15085) );
  NOR2_X1 U9725 ( .A1(n15086), .A2(n15085), .ZN(n7458) );
  XNOR2_X1 U9726 ( .A(n7461), .B(n7460), .ZN(n7463) );
  NAND2_X1 U9727 ( .A1(n7462), .A2(n7463), .ZN(n7464) );
  XNOR2_X1 U9728 ( .A(n7466), .B(n7465), .ZN(n14148) );
  NOR2_X1 U9729 ( .A1(n14149), .A2(n14148), .ZN(n7467) );
  INV_X1 U9730 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U9731 ( .A1(n14149), .A2(n14148), .ZN(n14147) );
  OAI21_X2 U9732 ( .B1(n7467), .B2(n14150), .A(n14147), .ZN(n14153) );
  NOR2_X1 U9733 ( .A1(n14154), .A2(n14153), .ZN(n7468) );
  INV_X1 U9734 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U9735 ( .A1(n14154), .A2(n14153), .ZN(n14152) );
  XNOR2_X1 U9736 ( .A(n7470), .B(n7469), .ZN(n7471) );
  NOR2_X1 U9737 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n14332), .ZN(n7474) );
  NOR2_X1 U9738 ( .A1(n7472), .A2(n7471), .ZN(n7473) );
  NOR2_X2 U9739 ( .A1(n7474), .A2(n7473), .ZN(n7478) );
  XNOR2_X1 U9740 ( .A(n7476), .B(n7475), .ZN(n7477) );
  XNOR2_X1 U9741 ( .A(n7478), .B(n7477), .ZN(n14333) );
  NOR2_X1 U9742 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n14333), .ZN(n7480) );
  NOR2_X1 U9743 ( .A1(n7478), .A2(n7477), .ZN(n7479) );
  NOR2_X2 U9744 ( .A1(n7480), .A2(n7479), .ZN(n14337) );
  NAND2_X1 U9745 ( .A1(n14336), .A2(n14337), .ZN(n7481) );
  NOR2_X1 U9746 ( .A1(n14336), .A2(n14337), .ZN(n14335) );
  XOR2_X1 U9747 ( .A(n14385), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n7484) );
  XNOR2_X1 U9748 ( .A(n7484), .B(n7483), .ZN(n14344) );
  INV_X1 U9749 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14345) );
  XOR2_X1 U9750 ( .A(n7486), .B(n7485), .Z(n7487) );
  NAND2_X1 U9751 ( .A1(n7488), .A2(n7487), .ZN(n14350) );
  INV_X1 U9752 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14351) );
  INV_X1 U9753 ( .A(n14348), .ZN(n14349) );
  NAND2_X1 U9754 ( .A1(n14347), .A2(n14349), .ZN(n14166) );
  NAND2_X1 U9755 ( .A1(n14165), .A2(n14166), .ZN(n14164) );
  XNOR2_X1 U9756 ( .A(n7696), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7489) );
  XNOR2_X1 U9757 ( .A(n7489), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7490) );
  INV_X1 U9758 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7494) );
  NOR2_X1 U9759 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  AOI21_X1 U9760 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n7494), .A(n7493), .ZN(
        n7663) );
  INV_X1 U9761 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U9762 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(keyinput_f57), .ZN(n7495) );
  OAI221_X1 U9763 ( .B1(SI_2_), .B2(keyinput_f30), .C1(P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n7495), .ZN(n7502) );
  AOI22_X1 U9764 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n7496) );
  OAI221_X1 U9765 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_6_), .C2(
        keyinput_f26), .A(n7496), .ZN(n7501) );
  AOI22_X1 U9766 ( .A1(keyinput_f33), .A2(P3_RD_REG_SCAN_IN), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n7497) );
  OAI221_X1 U9767 ( .B1(keyinput_f33), .B2(P3_RD_REG_SCAN_IN), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n7497), .ZN(n7500) );
  AOI22_X1 U9768 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n7498) );
  OAI221_X1 U9769 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n7498), .ZN(n7499) );
  NOR4_X1 U9770 ( .A1(n7502), .A2(n7501), .A3(n7500), .A4(n7499), .ZN(n7530)
         );
  INV_X1 U9771 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n7575) );
  XOR2_X1 U9772 ( .A(n7575), .B(keyinput_f59), .Z(n7510) );
  INV_X1 U9773 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7504) );
  AOI22_X1 U9774 ( .A1(SI_23_), .A2(keyinput_f9), .B1(n7504), .B2(keyinput_f47), .ZN(n7503) );
  OAI221_X1 U9775 ( .B1(SI_23_), .B2(keyinput_f9), .C1(n7504), .C2(
        keyinput_f47), .A(n7503), .ZN(n7509) );
  AOI22_X1 U9776 ( .A1(SI_26_), .A2(keyinput_f6), .B1(SI_28_), .B2(keyinput_f4), .ZN(n7505) );
  OAI221_X1 U9777 ( .B1(SI_26_), .B2(keyinput_f6), .C1(SI_28_), .C2(
        keyinput_f4), .A(n7505), .ZN(n7508) );
  AOI22_X1 U9778 ( .A1(SI_9_), .A2(keyinput_f23), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n7506) );
  OAI221_X1 U9779 ( .B1(SI_9_), .B2(keyinput_f23), .C1(P3_REG3_REG_5__SCAN_IN), 
        .C2(keyinput_f49), .A(n7506), .ZN(n7507) );
  NOR4_X1 U9780 ( .A1(n7510), .A2(n7509), .A3(n7508), .A4(n7507), .ZN(n7529)
         );
  AOI22_X1 U9781 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_f56), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n7511) );
  OAI221_X1 U9782 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n7511), .ZN(n7518) );
  AOI22_X1 U9783 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n7512) );
  OAI221_X1 U9784 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n7512), .ZN(n7517) );
  AOI22_X1 U9785 ( .A1(n10724), .A2(keyinput_f12), .B1(n13057), .B2(
        keyinput_f3), .ZN(n7513) );
  OAI221_X1 U9786 ( .B1(n10724), .B2(keyinput_f12), .C1(n13057), .C2(
        keyinput_f3), .A(n7513), .ZN(n7516) );
  AOI22_X1 U9787 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n7514) );
  OAI221_X1 U9788 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_17_), .C2(
        keyinput_f15), .A(n7514), .ZN(n7515) );
  NOR4_X1 U9789 ( .A1(n7518), .A2(n7517), .A3(n7516), .A4(n7515), .ZN(n7528)
         );
  AOI22_X1 U9790 ( .A1(SI_27_), .A2(keyinput_f5), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(keyinput_f36), .ZN(n7519) );
  OAI221_X1 U9791 ( .B1(SI_27_), .B2(keyinput_f5), .C1(P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n7519), .ZN(n7526) );
  AOI22_X1 U9792 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n7520) );
  OAI221_X1 U9793 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n7520), .ZN(n7525) );
  AOI22_X1 U9794 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n7521) );
  OAI221_X1 U9795 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n7521), .ZN(n7524) );
  AOI22_X1 U9796 ( .A1(SI_19_), .A2(keyinput_f13), .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n7522) );
  OAI221_X1 U9797 ( .B1(SI_19_), .B2(keyinput_f13), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n7522), .ZN(n7523) );
  NOR4_X1 U9798 ( .A1(n7526), .A2(n7525), .A3(n7524), .A4(n7523), .ZN(n7527)
         );
  NAND4_X1 U9799 ( .A1(n7530), .A2(n7529), .A3(n7528), .A4(n7527), .ZN(n7572)
         );
  INV_X1 U9800 ( .A(P3_WR_REG_SCAN_IN), .ZN(n7595) );
  AOI22_X1 U9801 ( .A1(n12341), .A2(keyinput_f51), .B1(keyinput_f0), .B2(n7595), .ZN(n7531) );
  OAI221_X1 U9802 ( .B1(n12341), .B2(keyinput_f51), .C1(n7595), .C2(
        keyinput_f0), .A(n7531), .ZN(n7539) );
  INV_X1 U9803 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10837) );
  INV_X1 U9804 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U9805 ( .A1(n10837), .A2(keyinput_f35), .B1(keyinput_f52), .B2(
        n10401), .ZN(n7532) );
  OAI221_X1 U9806 ( .B1(n10837), .B2(keyinput_f35), .C1(n10401), .C2(
        keyinput_f52), .A(n7532), .ZN(n7538) );
  INV_X1 U9807 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U9808 ( .A1(n11220), .A2(keyinput_f58), .B1(keyinput_f18), .B2(
        n9822), .ZN(n7533) );
  OAI221_X1 U9809 ( .B1(n11220), .B2(keyinput_f58), .C1(n9822), .C2(
        keyinput_f18), .A(n7533), .ZN(n7537) );
  XNOR2_X1 U9810 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_f50), .ZN(n7535)
         );
  XNOR2_X1 U9811 ( .A(SI_4_), .B(keyinput_f28), .ZN(n7534) );
  NAND2_X1 U9812 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NOR4_X1 U9813 ( .A1(n7539), .A2(n7538), .A3(n7537), .A4(n7536), .ZN(n7570)
         );
  INV_X1 U9814 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11447) );
  INV_X1 U9815 ( .A(SI_0_), .ZN(n7628) );
  AOI22_X1 U9816 ( .A1(n11447), .A2(keyinput_f46), .B1(keyinput_f32), .B2(
        n7628), .ZN(n7540) );
  OAI221_X1 U9817 ( .B1(n11447), .B2(keyinput_f46), .C1(n7628), .C2(
        keyinput_f32), .A(n7540), .ZN(n7548) );
  AOI22_X1 U9818 ( .A1(n9798), .A2(keyinput_f19), .B1(keyinput_f17), .B2(n9898), .ZN(n7541) );
  OAI221_X1 U9819 ( .B1(n9798), .B2(keyinput_f19), .C1(n9898), .C2(
        keyinput_f17), .A(n7541), .ZN(n7547) );
  INV_X1 U9820 ( .A(SI_24_), .ZN(n11295) );
  AOI22_X1 U9821 ( .A1(n11295), .A2(keyinput_f8), .B1(n11631), .B2(keyinput_f7), .ZN(n7542) );
  OAI221_X1 U9822 ( .B1(n11295), .B2(keyinput_f8), .C1(n11631), .C2(
        keyinput_f7), .A(n7542), .ZN(n7546) );
  XNOR2_X1 U9823 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_f41), .ZN(n7544)
         );
  XNOR2_X1 U9824 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7543) );
  NAND2_X1 U9825 ( .A1(n7544), .A2(n7543), .ZN(n7545) );
  NOR4_X1 U9826 ( .A1(n7548), .A2(n7547), .A3(n7546), .A4(n7545), .ZN(n7569)
         );
  INV_X1 U9827 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U9828 ( .A1(n10952), .A2(keyinput_f53), .B1(keyinput_f54), .B2(
        n14775), .ZN(n7549) );
  OAI221_X1 U9829 ( .B1(n10952), .B2(keyinput_f53), .C1(n14775), .C2(
        keyinput_f54), .A(n7549), .ZN(n7557) );
  INV_X1 U9830 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U9831 ( .A1(n10688), .A2(keyinput_f61), .B1(n11760), .B2(
        keyinput_f48), .ZN(n7550) );
  OAI221_X1 U9832 ( .B1(n10688), .B2(keyinput_f61), .C1(n11760), .C2(
        keyinput_f48), .A(n7550), .ZN(n7556) );
  XNOR2_X1 U9833 ( .A(SI_22_), .B(keyinput_f10), .ZN(n7554) );
  XNOR2_X1 U9834 ( .A(SI_7_), .B(keyinput_f25), .ZN(n7553) );
  XNOR2_X1 U9835 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_f40), .ZN(n7552) );
  XNOR2_X1 U9836 ( .A(SI_8_), .B(keyinput_f24), .ZN(n7551) );
  NAND4_X1 U9837 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n7555)
         );
  NOR3_X1 U9838 ( .A1(n7557), .A2(n7556), .A3(n7555), .ZN(n7568) );
  INV_X1 U9839 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7597) );
  AOI22_X1 U9840 ( .A1(n7597), .A2(keyinput_f60), .B1(keyinput_f22), .B2(n9740), .ZN(n7558) );
  OAI221_X1 U9841 ( .B1(n7597), .B2(keyinput_f60), .C1(n9740), .C2(
        keyinput_f22), .A(n7558), .ZN(n7566) );
  AOI22_X1 U9842 ( .A1(n9991), .A2(keyinput_f16), .B1(keyinput_f21), .B2(n9745), .ZN(n7559) );
  OAI221_X1 U9843 ( .B1(n9991), .B2(keyinput_f16), .C1(n9745), .C2(
        keyinput_f21), .A(n7559), .ZN(n7565) );
  INV_X1 U9844 ( .A(SI_18_), .ZN(n10325) );
  INV_X1 U9845 ( .A(SI_21_), .ZN(n11922) );
  AOI22_X1 U9846 ( .A1(n10325), .A2(keyinput_f14), .B1(n11922), .B2(
        keyinput_f11), .ZN(n7560) );
  OAI221_X1 U9847 ( .B1(n10325), .B2(keyinput_f14), .C1(n11922), .C2(
        keyinput_f11), .A(n7560), .ZN(n7564) );
  XNOR2_X1 U9848 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_f45), .ZN(n7562)
         );
  XNOR2_X1 U9849 ( .A(SI_3_), .B(keyinput_f29), .ZN(n7561) );
  NAND2_X1 U9850 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  NOR4_X1 U9851 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n7567)
         );
  NAND4_X1 U9852 ( .A1(n7570), .A2(n7569), .A3(n7568), .A4(n7567), .ZN(n7571)
         );
  OAI22_X1 U9853 ( .A1(n7572), .A2(n7571), .B1(keyinput_f63), .B2(
        P3_REG3_REG_15__SCAN_IN), .ZN(n7573) );
  AOI21_X1 U9854 ( .B1(keyinput_f63), .B2(P3_REG3_REG_15__SCAN_IN), .A(n7573), 
        .ZN(n7661) );
  AOI22_X1 U9855 ( .A1(n10837), .A2(keyinput_g35), .B1(keyinput_g59), .B2(
        n7575), .ZN(n7574) );
  OAI221_X1 U9856 ( .B1(n10837), .B2(keyinput_g35), .C1(n7575), .C2(
        keyinput_g59), .A(n7574), .ZN(n7584) );
  INV_X1 U9857 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n7577) );
  AOI22_X1 U9858 ( .A1(n11645), .A2(keyinput_g6), .B1(n7577), .B2(keyinput_g44), .ZN(n7576) );
  OAI221_X1 U9859 ( .B1(n11645), .B2(keyinput_g6), .C1(n7577), .C2(
        keyinput_g44), .A(n7576), .ZN(n7583) );
  AOI22_X1 U9860 ( .A1(n9460), .A2(keyinput_g55), .B1(keyinput_g17), .B2(n9898), .ZN(n7578) );
  OAI221_X1 U9861 ( .B1(n9460), .B2(keyinput_g55), .C1(n9898), .C2(
        keyinput_g17), .A(n7578), .ZN(n7582) );
  XNOR2_X1 U9862 ( .A(SI_7_), .B(keyinput_g25), .ZN(n7580) );
  XNOR2_X1 U9863 ( .A(keyinput_g54), .B(P3_REG3_REG_0__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9864 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  NOR4_X1 U9865 ( .A1(n7584), .A2(n7583), .A3(n7582), .A4(n7581), .ZN(n7618)
         );
  INV_X1 U9866 ( .A(SI_23_), .ZN(n10917) );
  AOI22_X1 U9867 ( .A1(n10917), .A2(keyinput_g9), .B1(n9491), .B2(keyinput_g10), .ZN(n7585) );
  OAI221_X1 U9868 ( .B1(n10917), .B2(keyinput_g9), .C1(n9491), .C2(
        keyinput_g10), .A(n7585), .ZN(n7593) );
  AOI22_X1 U9869 ( .A1(n9745), .A2(keyinput_g21), .B1(n9991), .B2(keyinput_g16), .ZN(n7586) );
  OAI221_X1 U9870 ( .B1(n9745), .B2(keyinput_g21), .C1(n9991), .C2(
        keyinput_g16), .A(n7586), .ZN(n7592) );
  INV_X1 U9871 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U9872 ( .A1(n11760), .A2(keyinput_g48), .B1(n12378), .B2(
        keyinput_g62), .ZN(n7587) );
  OAI221_X1 U9873 ( .B1(n11760), .B2(keyinput_g48), .C1(n12378), .C2(
        keyinput_g62), .A(n7587), .ZN(n7591) );
  INV_X1 U9874 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9564) );
  INV_X1 U9875 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n7589) );
  AOI22_X1 U9876 ( .A1(n9564), .A2(keyinput_g36), .B1(keyinput_g57), .B2(n7589), .ZN(n7588) );
  OAI221_X1 U9877 ( .B1(n9564), .B2(keyinput_g36), .C1(n7589), .C2(
        keyinput_g57), .A(n7588), .ZN(n7590) );
  NOR4_X1 U9878 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n7617)
         );
  INV_X1 U9879 ( .A(SI_30_), .ZN(n12528) );
  AOI22_X1 U9880 ( .A1(n12528), .A2(keyinput_g2), .B1(keyinput_g0), .B2(n7595), 
        .ZN(n7594) );
  OAI221_X1 U9881 ( .B1(n12528), .B2(keyinput_g2), .C1(n7595), .C2(keyinput_g0), .A(n7594), .ZN(n7604) );
  AOI22_X1 U9882 ( .A1(n7597), .A2(keyinput_g60), .B1(keyinput_g50), .B2(n9403), .ZN(n7596) );
  OAI221_X1 U9883 ( .B1(n7597), .B2(keyinput_g60), .C1(n9403), .C2(
        keyinput_g50), .A(n7596), .ZN(n7603) );
  AOI22_X1 U9884 ( .A1(n10465), .A2(keyinput_g13), .B1(n10401), .B2(
        keyinput_g52), .ZN(n7598) );
  OAI221_X1 U9885 ( .B1(n10465), .B2(keyinput_g13), .C1(n10401), .C2(
        keyinput_g52), .A(n7598), .ZN(n7602) );
  XNOR2_X1 U9886 ( .A(SI_2_), .B(keyinput_g30), .ZN(n7600) );
  XNOR2_X1 U9887 ( .A(SI_31_), .B(keyinput_g1), .ZN(n7599) );
  NAND2_X1 U9888 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  NOR4_X1 U9889 ( .A1(n7604), .A2(n7603), .A3(n7602), .A4(n7601), .ZN(n7616)
         );
  XNOR2_X1 U9890 ( .A(SI_9_), .B(keyinput_g23), .ZN(n7608) );
  XNOR2_X1 U9891 ( .A(SI_28_), .B(keyinput_g4), .ZN(n7607) );
  XNOR2_X1 U9892 ( .A(SI_3_), .B(keyinput_g29), .ZN(n7606) );
  XNOR2_X1 U9893 ( .A(SI_24_), .B(keyinput_g8), .ZN(n7605) );
  NAND4_X1 U9894 ( .A1(n7608), .A2(n7607), .A3(n7606), .A4(n7605), .ZN(n7614)
         );
  XNOR2_X1 U9895 ( .A(SI_6_), .B(keyinput_g26), .ZN(n7612) );
  XNOR2_X1 U9896 ( .A(SI_25_), .B(keyinput_g7), .ZN(n7611) );
  XNOR2_X1 U9897 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n7610)
         );
  XNOR2_X1 U9898 ( .A(SI_4_), .B(keyinput_g28), .ZN(n7609) );
  NAND4_X1 U9899 ( .A1(n7612), .A2(n7611), .A3(n7610), .A4(n7609), .ZN(n7613)
         );
  NOR2_X1 U9900 ( .A1(n7614), .A2(n7613), .ZN(n7615) );
  NAND4_X1 U9901 ( .A1(n7618), .A2(n7617), .A3(n7616), .A4(n7615), .ZN(n7659)
         );
  AOI22_X1 U9902 ( .A1(SI_18_), .A2(keyinput_g14), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n7619) );
  OAI221_X1 U9903 ( .B1(SI_18_), .B2(keyinput_g14), .C1(SI_21_), .C2(
        keyinput_g11), .A(n7619), .ZN(n7626) );
  AOI22_X1 U9904 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n7620) );
  OAI221_X1 U9905 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n7620), .ZN(n7625) );
  AOI22_X1 U9906 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .ZN(n7621) );
  OAI221_X1 U9907 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P3_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n7621), .ZN(n7624) );
  AOI22_X1 U9908 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n7622) );
  OAI221_X1 U9909 ( .B1(SI_10_), .B2(keyinput_g22), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n7622), .ZN(n7623) );
  NOR4_X1 U9910 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n7657)
         );
  AOI22_X1 U9911 ( .A1(SI_29_), .A2(keyinput_g3), .B1(n7628), .B2(keyinput_g32), .ZN(n7627) );
  OAI221_X1 U9912 ( .B1(SI_29_), .B2(keyinput_g3), .C1(n7628), .C2(
        keyinput_g32), .A(n7627), .ZN(n7634) );
  AOI22_X1 U9913 ( .A1(SI_12_), .A2(keyinput_g20), .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n7629) );
  OAI221_X1 U9914 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n7629), .ZN(n7633) );
  AOI22_X1 U9915 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n7630) );
  OAI221_X1 U9916 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n7630), .ZN(n7632) );
  XNOR2_X1 U9917 ( .A(SI_5_), .B(keyinput_g27), .ZN(n7631) );
  NOR4_X1 U9918 ( .A1(n7634), .A2(n7633), .A3(n7632), .A4(n7631), .ZN(n7656)
         );
  INV_X1 U9919 ( .A(SI_27_), .ZN(n11736) );
  AOI22_X1 U9920 ( .A1(n11736), .A2(keyinput_g5), .B1(P3_U3151), .B2(
        keyinput_g34), .ZN(n7635) );
  OAI221_X1 U9921 ( .B1(n11736), .B2(keyinput_g5), .C1(P3_U3151), .C2(
        keyinput_g34), .A(n7635), .ZN(n7645) );
  INV_X1 U9922 ( .A(SI_17_), .ZN(n7638) );
  INV_X1 U9923 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n7637) );
  AOI22_X1 U9924 ( .A1(n7638), .A2(keyinput_g15), .B1(n7637), .B2(keyinput_g42), .ZN(n7636) );
  OAI221_X1 U9925 ( .B1(n7638), .B2(keyinput_g15), .C1(n7637), .C2(
        keyinput_g42), .A(n7636), .ZN(n7644) );
  AOI22_X1 U9926 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n7639) );
  OAI221_X1 U9927 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7639), .ZN(n7643) );
  XNOR2_X1 U9928 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n7641) );
  XNOR2_X1 U9929 ( .A(SI_1_), .B(keyinput_g31), .ZN(n7640) );
  NAND2_X1 U9930 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NOR4_X1 U9931 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n7655)
         );
  AOI22_X1 U9932 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(SI_20_), 
        .B2(keyinput_g12), .ZN(n7646) );
  OAI221_X1 U9933 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(SI_20_), 
        .C2(keyinput_g12), .A(n7646), .ZN(n7653) );
  AOI22_X1 U9934 ( .A1(SI_14_), .A2(keyinput_g18), .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n7647) );
  OAI221_X1 U9935 ( .B1(SI_14_), .B2(keyinput_g18), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n7647), .ZN(n7652) );
  AOI22_X1 U9936 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n7648) );
  OAI221_X1 U9937 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n7648), .ZN(n7651) );
  AOI22_X1 U9938 ( .A1(SI_8_), .A2(keyinput_g24), .B1(SI_13_), .B2(
        keyinput_g19), .ZN(n7649) );
  OAI221_X1 U9939 ( .B1(SI_8_), .B2(keyinput_g24), .C1(SI_13_), .C2(
        keyinput_g19), .A(n7649), .ZN(n7650) );
  NOR4_X1 U9940 ( .A1(n7653), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n7654)
         );
  NAND4_X1 U9941 ( .A1(n7657), .A2(n7656), .A3(n7655), .A4(n7654), .ZN(n7658)
         );
  OAI22_X1 U9942 ( .A1(keyinput_g63), .A2(n11677), .B1(n7659), .B2(n7658), 
        .ZN(n7660) );
  AOI211_X1 U9943 ( .C1(keyinput_g63), .C2(n11677), .A(n7661), .B(n7660), .ZN(
        n7662) );
  NOR2_X1 U9944 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n7668) );
  NOR2_X2 U9945 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8034) );
  NOR2_X1 U9946 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7673) );
  NOR2_X1 U9947 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7672) );
  NOR2_X1 U9948 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7671) );
  NOR2_X1 U9949 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7676) );
  NAND2_X1 U9950 ( .A1(n7679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7680) );
  INV_X1 U9951 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7684) );
  AND2_X4 U9952 ( .A1(n7813), .A2(n14120), .ZN(n8332) );
  NAND2_X1 U9953 ( .A1(n8332), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7683) );
  INV_X1 U9954 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7681) );
  OR2_X1 U9955 ( .A1(n8184), .A2(n7681), .ZN(n7682) );
  OAI211_X1 U9956 ( .C1(n8205), .C2(n7684), .A(n7683), .B(n7682), .ZN(n13821)
         );
  NAND2_X1 U9957 ( .A1(n7799), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7686) );
  NAND2_X1 U9958 ( .A1(n8429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7689) );
  INV_X1 U9959 ( .A(n11297), .ZN(n10571) );
  NAND2_X1 U9960 ( .A1(n10284), .A2(n10571), .ZN(n10471) );
  INV_X1 U9961 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9962 ( .A1(n8332), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9963 ( .A1(n6485), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7690) );
  OAI211_X1 U9964 ( .C1(n6482), .C2(n7692), .A(n7691), .B(n7690), .ZN(n13842)
         );
  OAI21_X1 U9965 ( .B1(n13821), .B2(n10471), .A(n13842), .ZN(n7805) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9733), .Z(n8862) );
  MUX2_X1 U9967 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7697), .Z(n7698) );
  NAND2_X1 U9968 ( .A1(n7698), .A2(SI_0_), .ZN(n7834) );
  INV_X1 U9969 ( .A(n7699), .ZN(n7700) );
  INV_X1 U9970 ( .A(SI_1_), .ZN(n9754) );
  INV_X1 U9971 ( .A(SI_2_), .ZN(n9716) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8501), .Z(n7867) );
  AND2_X1 U9973 ( .A1(n7867), .A2(n6805), .ZN(n7701) );
  NAND2_X1 U9974 ( .A1(n7705), .A2(SI_3_), .ZN(n7895) );
  MUX2_X1 U9975 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8501), .Z(n7708) );
  NAND2_X1 U9976 ( .A1(n7708), .A2(SI_4_), .ZN(n7707) );
  AND2_X1 U9977 ( .A1(n7895), .A2(n7707), .ZN(n7712) );
  INV_X1 U9978 ( .A(n7707), .ZN(n7710) );
  INV_X1 U9979 ( .A(n7896), .ZN(n7709) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8501), .Z(n7713) );
  XNOR2_X1 U9981 ( .A(n7713), .B(SI_5_), .ZN(n7911) );
  NAND2_X1 U9982 ( .A1(n7713), .A2(SI_5_), .ZN(n7935) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8501), .Z(n7715) );
  NAND2_X1 U9984 ( .A1(n7715), .A2(SI_6_), .ZN(n7714) );
  AND2_X1 U9985 ( .A1(n7935), .A2(n7714), .ZN(n7718) );
  INV_X1 U9986 ( .A(n7714), .ZN(n7717) );
  XNOR2_X1 U9987 ( .A(n7715), .B(SI_6_), .ZN(n7937) );
  INV_X1 U9988 ( .A(n7937), .ZN(n7716) );
  MUX2_X1 U9989 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n6627), .Z(n7720) );
  XNOR2_X1 U9990 ( .A(n7720), .B(SI_7_), .ZN(n7951) );
  INV_X1 U9991 ( .A(n7951), .ZN(n7719) );
  NAND2_X1 U9992 ( .A1(n7720), .A2(SI_7_), .ZN(n7968) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6627), .Z(n7722) );
  NAND2_X1 U9994 ( .A1(n7722), .A2(SI_8_), .ZN(n7721) );
  AND2_X1 U9995 ( .A1(n7968), .A2(n7721), .ZN(n7725) );
  INV_X1 U9996 ( .A(n7721), .ZN(n7724) );
  XNOR2_X1 U9997 ( .A(n7722), .B(SI_8_), .ZN(n7970) );
  INV_X1 U9998 ( .A(n7970), .ZN(n7723) );
  AOI21_X2 U9999 ( .B1(n7969), .B2(n7725), .A(n7378), .ZN(n7995) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6627), .Z(n7727) );
  XNOR2_X1 U10001 ( .A(n7727), .B(SI_9_), .ZN(n7994) );
  INV_X1 U10002 ( .A(n7994), .ZN(n7726) );
  NAND2_X1 U10003 ( .A1(n7995), .A2(n7726), .ZN(n7729) );
  NAND2_X1 U10004 ( .A1(n7727), .A2(SI_9_), .ZN(n7728) );
  NAND2_X1 U10005 ( .A1(n7729), .A2(n7728), .ZN(n8013) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6627), .Z(n8011) );
  INV_X1 U10007 ( .A(n8011), .ZN(n7730) );
  NAND2_X1 U10008 ( .A1(n7730), .A2(n9740), .ZN(n7731) );
  NAND2_X1 U10009 ( .A1(n8013), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U10010 ( .A1(n8011), .A2(SI_10_), .ZN(n7732) );
  MUX2_X1 U10011 ( .A(n9903), .B(n9901), .S(n6627), .Z(n7734) );
  INV_X1 U10012 ( .A(n7734), .ZN(n7735) );
  NAND2_X1 U10013 ( .A1(n7735), .A2(SI_11_), .ZN(n7736) );
  NAND2_X1 U10014 ( .A1(n7737), .A2(n7736), .ZN(n8032) );
  MUX2_X1 U10015 ( .A(n9324), .B(n10221), .S(n6627), .Z(n7738) );
  INV_X1 U10016 ( .A(n7738), .ZN(n7739) );
  NAND2_X1 U10017 ( .A1(n7739), .A2(SI_12_), .ZN(n7740) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n6627), .Z(n8071) );
  INV_X1 U10019 ( .A(n8071), .ZN(n7742) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6627), .Z(n8090) );
  INV_X1 U10021 ( .A(n8090), .ZN(n8103) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6627), .Z(n7745) );
  NAND2_X1 U10023 ( .A1(n7745), .A2(SI_15_), .ZN(n7746) );
  OAI21_X1 U10024 ( .B1(n8103), .B2(n9822), .A(n7746), .ZN(n7743) );
  INV_X1 U10025 ( .A(n7743), .ZN(n7744) );
  NOR2_X1 U10026 ( .A1(n8090), .A2(SI_14_), .ZN(n7747) );
  INV_X1 U10027 ( .A(n7745), .ZN(n8108) );
  AOI22_X1 U10028 ( .A1(n7747), .A2(n7746), .B1(n9898), .B2(n8108), .ZN(n7748)
         );
  MUX2_X1 U10029 ( .A(n10534), .B(n10532), .S(n6627), .Z(n7749) );
  XNOR2_X1 U10030 ( .A(n7749), .B(SI_16_), .ZN(n8133) );
  NAND2_X1 U10031 ( .A1(n7749), .A2(n9991), .ZN(n7750) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n6627), .Z(n8148) );
  NOR2_X1 U10033 ( .A1(n8148), .A2(SI_17_), .ZN(n7751) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9733), .Z(n8173) );
  NAND2_X1 U10035 ( .A1(n7752), .A2(SI_18_), .ZN(n7753) );
  MUX2_X1 U10036 ( .A(n10884), .B(n10886), .S(n9733), .Z(n7755) );
  INV_X1 U10037 ( .A(n7755), .ZN(n7756) );
  NAND2_X1 U10038 ( .A1(n7756), .A2(SI_19_), .ZN(n7757) );
  NAND2_X1 U10039 ( .A1(n7758), .A2(n7757), .ZN(n8164) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9733), .Z(n8228) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9733), .Z(n8223) );
  NOR2_X1 U10042 ( .A1(n8223), .A2(SI_20_), .ZN(n7759) );
  INV_X1 U10043 ( .A(n8223), .ZN(n7760) );
  NOR2_X1 U10044 ( .A1(n7760), .A2(n10724), .ZN(n7763) );
  INV_X1 U10045 ( .A(n7761), .ZN(n7762) );
  AOI22_X1 U10046 ( .A1(n7763), .A2(n7762), .B1(n8228), .B2(SI_21_), .ZN(n8242) );
  NAND2_X1 U10047 ( .A1(n7764), .A2(n9491), .ZN(n7765) );
  INV_X1 U10048 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7767) );
  INV_X1 U10049 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11628) );
  MUX2_X1 U10050 ( .A(n7767), .B(n11628), .S(n9733), .Z(n7769) );
  INV_X1 U10051 ( .A(n7768), .ZN(n7771) );
  INV_X1 U10052 ( .A(n7769), .ZN(n7770) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9733), .Z(n8273) );
  NAND2_X1 U10054 ( .A1(n7773), .A2(n8273), .ZN(n7776) );
  NAND2_X1 U10055 ( .A1(n7774), .A2(SI_24_), .ZN(n7775) );
  INV_X1 U10056 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11987) );
  MUX2_X1 U10057 ( .A(n11987), .B(n11882), .S(n9733), .Z(n7777) );
  NAND2_X1 U10058 ( .A1(n7777), .A2(n11631), .ZN(n7780) );
  INV_X1 U10059 ( .A(n7777), .ZN(n7778) );
  NAND2_X1 U10060 ( .A1(n7778), .A2(SI_25_), .ZN(n7779) );
  NAND2_X1 U10061 ( .A1(n7780), .A2(n7779), .ZN(n8290) );
  MUX2_X1 U10062 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9733), .Z(n8304) );
  INV_X1 U10063 ( .A(n8304), .ZN(n7781) );
  INV_X1 U10064 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14124) );
  INV_X1 U10065 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13577) );
  MUX2_X1 U10066 ( .A(n14124), .B(n13577), .S(n9733), .Z(n8324) );
  INV_X1 U10067 ( .A(n8324), .ZN(n7782) );
  NOR2_X1 U10068 ( .A1(n7782), .A2(SI_27_), .ZN(n7784) );
  NAND2_X1 U10069 ( .A1(n7782), .A2(SI_27_), .ZN(n7783) );
  MUX2_X1 U10070 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9733), .Z(n7785) );
  XNOR2_X1 U10071 ( .A(n7785), .B(SI_28_), .ZN(n8338) );
  INV_X1 U10072 ( .A(n7785), .ZN(n7786) );
  INV_X1 U10073 ( .A(SI_28_), .ZN(n11924) );
  NAND2_X1 U10074 ( .A1(n7786), .A2(n11924), .ZN(n7787) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9733), .Z(n7788) );
  XNOR2_X1 U10076 ( .A(n7788), .B(n13057), .ZN(n7823) );
  INV_X1 U10077 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U10078 ( .A1(n7789), .A2(n13057), .ZN(n7790) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9733), .Z(n8365) );
  XNOR2_X1 U10080 ( .A(n8365), .B(SI_30_), .ZN(n8367) );
  INV_X1 U10081 ( .A(n8367), .ZN(n7792) );
  XNOR2_X2 U10082 ( .A(n7794), .B(n7793), .ZN(n11928) );
  NAND2_X1 U10083 ( .A1(n7795), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7796) );
  INV_X1 U10084 ( .A(n10284), .ZN(n11511) );
  NAND2_X1 U10085 ( .A1(n7801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7802) );
  MUX2_X1 U10086 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7802), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n7803) );
  NAND2_X1 U10087 ( .A1(n8362), .A2(n13897), .ZN(n10282) );
  OR2_X1 U10088 ( .A1(n8362), .A2(n13897), .ZN(n7804) );
  NAND2_X1 U10089 ( .A1(n10282), .A2(n7804), .ZN(n7806) );
  MUX2_X1 U10090 ( .A(n10571), .B(n11511), .S(n7806), .Z(n7882) );
  MUX2_X1 U10091 ( .A(n7805), .B(n14019), .S(n8377), .Z(n8353) );
  INV_X4 U10092 ( .A(n7882), .ZN(n8375) );
  NAND2_X1 U10093 ( .A1(n13824), .A2(n8375), .ZN(n7810) );
  INV_X1 U10094 ( .A(n13821), .ZN(n8392) );
  INV_X1 U10095 ( .A(n7806), .ZN(n7807) );
  OAI22_X1 U10096 ( .A1(n8375), .A2(n8392), .B1(n10284), .B2(n7807), .ZN(n7808) );
  NAND2_X1 U10097 ( .A1(n7808), .A2(n13842), .ZN(n7809) );
  NAND2_X1 U10098 ( .A1(n7810), .A2(n7809), .ZN(n8358) );
  NAND2_X1 U10099 ( .A1(n8331), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7822) );
  INV_X1 U10100 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7811) );
  OR2_X1 U10101 ( .A1(n7876), .A2(n7811), .ZN(n7821) );
  INV_X2 U10102 ( .A(n7842), .ZN(n7889) );
  NAND2_X1 U10103 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7905) );
  INV_X1 U10104 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7904) );
  NOR2_X1 U10105 ( .A1(n7905), .A2(n7904), .ZN(n7929) );
  NAND2_X1 U10106 ( .A1(n7929), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10107 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n7814) );
  NAND2_X1 U10108 ( .A1(n8025), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10109 ( .A1(n8096), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8116) );
  INV_X1 U10110 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10111 ( .A1(n8217), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10112 ( .A1(n8268), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U10113 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n8285), .ZN(n8298) );
  INV_X1 U10114 ( .A(n8298), .ZN(n7815) );
  NAND2_X1 U10115 ( .A1(n7815), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8318) );
  INV_X1 U10116 ( .A(n8318), .ZN(n7816) );
  NAND2_X1 U10117 ( .A1(n7816), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8333) );
  INV_X1 U10118 ( .A(n8333), .ZN(n7817) );
  NAND2_X1 U10119 ( .A1(n7817), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13844) );
  OR2_X1 U10120 ( .A1(n7889), .A2(n13844), .ZN(n7820) );
  INV_X1 U10121 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7818) );
  OR2_X1 U10122 ( .A1(n8184), .A2(n7818), .ZN(n7819) );
  AND4_X1 U10123 ( .A1(n7822), .A2(n7821), .A3(n7820), .A4(n7819), .ZN(n7827)
         );
  NAND2_X1 U10124 ( .A1(n13569), .A2(n8372), .ZN(n7826) );
  NAND2_X1 U10125 ( .A1(n8178), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7825) );
  MUX2_X1 U10126 ( .A(n7827), .B(n14022), .S(n8377), .Z(n8352) );
  MUX2_X1 U10127 ( .A(n13665), .B(n13841), .S(n8375), .Z(n8351) );
  OAI22_X1 U10128 ( .A1(n8353), .A2(n8358), .B1(n8352), .B2(n8351), .ZN(n7828)
         );
  INV_X1 U10129 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13691) );
  OR2_X1 U10130 ( .A1(n6487), .A2(n13691), .ZN(n7833) );
  INV_X1 U10131 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10132 ( .A1(n8332), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7830) );
  XNOR2_X1 U10133 ( .A(n7835), .B(n7834), .ZN(n9736) );
  INV_X1 U10134 ( .A(n9736), .ZN(n7836) );
  NAND2_X1 U10135 ( .A1(n7837), .A2(n7836), .ZN(n7841) );
  NAND2_X1 U10136 ( .A1(n7862), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10137 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7838) );
  XNOR2_X1 U10138 ( .A(n7838), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13693) );
  NAND2_X1 U10139 ( .A1(n6488), .A2(n13693), .ZN(n7839) );
  INV_X1 U10140 ( .A(n10578), .ZN(n8402) );
  MUX2_X1 U10141 ( .A(n8402), .B(n6511), .S(n7882), .Z(n7866) );
  NAND2_X1 U10142 ( .A1(n7842), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7847) );
  INV_X1 U10143 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7843) );
  NAND4_X2 U10144 ( .A1(n7847), .A2(n7846), .A3(n7845), .A4(n7844), .ZN(n13690) );
  INV_X1 U10145 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10360) );
  NOR2_X1 U10146 ( .A1(n9733), .A2(n7628), .ZN(n7848) );
  XNOR2_X1 U10147 ( .A(n7848), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14132) );
  MUX2_X1 U10148 ( .A(n10360), .B(n14132), .S(n9896), .Z(n10622) );
  NOR2_X1 U10149 ( .A1(n10576), .A2(n8375), .ZN(n7850) );
  NAND2_X1 U10150 ( .A1(n6511), .A2(n8402), .ZN(n7849) );
  NOR2_X1 U10151 ( .A1(n7850), .A2(n7849), .ZN(n7854) );
  NAND2_X1 U10152 ( .A1(n13690), .A2(n10622), .ZN(n8403) );
  NAND2_X1 U10153 ( .A1(n8403), .A2(n10468), .ZN(n7851) );
  NAND2_X1 U10154 ( .A1(n7851), .A2(n10576), .ZN(n7852) );
  INV_X1 U10155 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10347) );
  OR2_X1 U10156 ( .A1(n6487), .A2(n10347), .ZN(n7860) );
  NAND2_X1 U10157 ( .A1(n8332), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10158 ( .A1(n7855), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7858) );
  INV_X1 U10159 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10160 ( .A1(n9728), .A2(n7837), .ZN(n7865) );
  OR2_X1 U10161 ( .A1(n7863), .A2(n8135), .ZN(n7864) );
  XNOR2_X1 U10162 ( .A(n7864), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U10163 ( .A1(n7868), .A2(n7867), .ZN(n7870) );
  NAND2_X1 U10164 ( .A1(n7870), .A2(n7869), .ZN(n7872) );
  NAND2_X1 U10165 ( .A1(n9737), .A2(n7837), .ZN(n7875) );
  OR2_X1 U10166 ( .A1(n7898), .A2(n8135), .ZN(n7873) );
  XNOR2_X1 U10167 ( .A(n7873), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U10168 ( .A1(n7862), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n8177), .B2(
        n13711), .ZN(n7874) );
  NAND2_X1 U10169 ( .A1(n6485), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7881) );
  OR2_X1 U10170 ( .A1(n7889), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7880) );
  INV_X1 U10171 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n13703) );
  INV_X1 U10172 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7877) );
  OR2_X1 U10173 ( .A1(n8205), .A2(n7877), .ZN(n7878) );
  OR2_X1 U10174 ( .A1(n14447), .A2(n10732), .ZN(n7886) );
  NAND2_X1 U10175 ( .A1(n10637), .A2(n10374), .ZN(n14436) );
  MUX2_X1 U10176 ( .A(n14436), .B(n7883), .S(n8375), .Z(n7884) );
  MUX2_X1 U10177 ( .A(n7886), .B(n10585), .S(n8375), .Z(n7887) );
  INV_X2 U10178 ( .A(n6482), .ZN(n8331) );
  NAND2_X1 U10179 ( .A1(n8331), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7894) );
  INV_X1 U10180 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7888) );
  OR2_X1 U10181 ( .A1(n7876), .A2(n7888), .ZN(n7893) );
  OAI21_X1 U10182 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7905), .ZN(n10754) );
  OR2_X1 U10183 ( .A1(n7889), .A2(n10754), .ZN(n7892) );
  INV_X1 U10184 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7890) );
  OR2_X1 U10185 ( .A1(n8184), .A2(n7890), .ZN(n7891) );
  NAND2_X1 U10186 ( .A1(n8545), .A2(n8372), .ZN(n7901) );
  NAND2_X1 U10187 ( .A1(n7898), .A2(n7897), .ZN(n7913) );
  NAND2_X1 U10188 ( .A1(n7913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7899) );
  XNOR2_X1 U10189 ( .A(n7899), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U10190 ( .A1(n8178), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8177), .B2(
        n13719), .ZN(n7900) );
  MUX2_X1 U10191 ( .A(n14357), .B(n14516), .S(n7882), .Z(n7903) );
  INV_X1 U10192 ( .A(n14357), .ZN(n13686) );
  MUX2_X1 U10193 ( .A(n13686), .B(n10751), .S(n8375), .Z(n7902) );
  INV_X1 U10194 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9929) );
  OR2_X1 U10195 ( .A1(n7876), .A2(n9929), .ZN(n7910) );
  AND2_X1 U10196 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  OR2_X1 U10197 ( .A1(n7906), .A2(n7929), .ZN(n14423) );
  OR2_X1 U10198 ( .A1(n7889), .A2(n14423), .ZN(n7909) );
  INV_X1 U10199 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9908) );
  OR2_X1 U10200 ( .A1(n8184), .A2(n9908), .ZN(n7908) );
  NAND2_X1 U10201 ( .A1(n8331), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7907) );
  NAND4_X1 U10202 ( .A1(n7910), .A2(n7909), .A3(n7908), .A4(n7907), .ZN(n13685) );
  NAND2_X1 U10203 ( .A1(n9755), .A2(n8372), .ZN(n7920) );
  NAND2_X1 U10204 ( .A1(n7915), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7914) );
  MUX2_X1 U10205 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7914), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7918) );
  INV_X1 U10206 ( .A(n7915), .ZN(n7917) );
  INV_X1 U10207 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10208 ( .A1(n7917), .A2(n7916), .ZN(n7953) );
  NAND2_X1 U10209 ( .A1(n7918), .A2(n7953), .ZN(n9946) );
  INV_X1 U10210 ( .A(n9946), .ZN(n9930) );
  AOI22_X1 U10211 ( .A1(n8178), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8177), .B2(
        n9930), .ZN(n7919) );
  MUX2_X1 U10212 ( .A(n13685), .B(n14431), .S(n8375), .Z(n7924) );
  NAND2_X1 U10213 ( .A1(n7923), .A2(n7924), .ZN(n7922) );
  MUX2_X1 U10214 ( .A(n13685), .B(n14431), .S(n8377), .Z(n7921) );
  NAND2_X1 U10215 ( .A1(n7922), .A2(n7921), .ZN(n7928) );
  INV_X1 U10216 ( .A(n7923), .ZN(n7926) );
  INV_X1 U10217 ( .A(n7924), .ZN(n7925) );
  NAND2_X1 U10218 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  NAND2_X1 U10219 ( .A1(n8332), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10220 ( .A1(n8331), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7933) );
  OR2_X1 U10221 ( .A1(n7929), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10222 ( .A1(n7945), .A2(n7930), .ZN(n10859) );
  OR2_X1 U10223 ( .A1(n7889), .A2(n10859), .ZN(n7932) );
  NAND2_X1 U10224 ( .A1(n6485), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7931) );
  NAND4_X1 U10225 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n13684) );
  NAND2_X1 U10226 ( .A1(n7936), .A2(n7935), .ZN(n7938) );
  XNOR2_X1 U10227 ( .A(n7938), .B(n7937), .ZN(n9762) );
  NAND2_X1 U10228 ( .A1(n9762), .A2(n8372), .ZN(n7941) );
  NAND2_X1 U10229 ( .A1(n7953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7939) );
  XNOR2_X1 U10230 ( .A(n7939), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U10231 ( .A1(n8178), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8177), .B2(
        n9931), .ZN(n7940) );
  NAND2_X1 U10232 ( .A1(n7941), .A2(n7940), .ZN(n14533) );
  MUX2_X1 U10233 ( .A(n13684), .B(n14533), .S(n8377), .Z(n7943) );
  MUX2_X1 U10234 ( .A(n13684), .B(n14533), .S(n8375), .Z(n7942) );
  INV_X1 U10235 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9933) );
  OR2_X1 U10236 ( .A1(n7876), .A2(n9933), .ZN(n7950) );
  NAND2_X1 U10237 ( .A1(n8331), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10238 ( .A1(n7945), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U10239 ( .A1(n7988), .A2(n7946), .ZN(n14409) );
  OR2_X1 U10240 ( .A1(n7889), .A2(n14409), .ZN(n7948) );
  NAND2_X1 U10241 ( .A1(n6485), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7947) );
  NAND4_X1 U10242 ( .A1(n7950), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n13683) );
  XNOR2_X1 U10243 ( .A(n7952), .B(n7951), .ZN(n9794) );
  NAND2_X1 U10244 ( .A1(n9794), .A2(n8372), .ZN(n7956) );
  NAND2_X1 U10245 ( .A1(n7972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7954) );
  XNOR2_X1 U10246 ( .A(n7954), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U10247 ( .A1(n8178), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8177), .B2(
        n9934), .ZN(n7955) );
  NAND2_X1 U10248 ( .A1(n7956), .A2(n7955), .ZN(n11027) );
  MUX2_X1 U10249 ( .A(n13683), .B(n11027), .S(n8375), .Z(n7960) );
  NAND2_X1 U10250 ( .A1(n7959), .A2(n7960), .ZN(n7958) );
  MUX2_X1 U10251 ( .A(n13683), .B(n11027), .S(n8377), .Z(n7957) );
  NAND2_X1 U10252 ( .A1(n7958), .A2(n7957), .ZN(n7979) );
  INV_X1 U10253 ( .A(n7959), .ZN(n7962) );
  INV_X1 U10254 ( .A(n7960), .ZN(n7961) );
  NAND2_X1 U10255 ( .A1(n7962), .A2(n7961), .ZN(n7982) );
  NAND2_X1 U10256 ( .A1(n7979), .A2(n7982), .ZN(n7976) );
  NAND2_X1 U10257 ( .A1(n8331), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7967) );
  INV_X1 U10258 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7987) );
  XNOR2_X1 U10259 ( .A(n7988), .B(n7987), .ZN(n11555) );
  OR2_X1 U10260 ( .A1(n7889), .A2(n11555), .ZN(n7966) );
  INV_X1 U10261 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7963) );
  OR2_X1 U10262 ( .A1(n8184), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U10263 ( .A1(n8332), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7964) );
  NAND4_X1 U10264 ( .A1(n7967), .A2(n7966), .A3(n7965), .A4(n7964), .ZN(n13682) );
  NAND2_X1 U10265 ( .A1(n7969), .A2(n7968), .ZN(n7971) );
  XNOR2_X1 U10266 ( .A(n7971), .B(n7970), .ZN(n9800) );
  NAND2_X1 U10267 ( .A1(n9800), .A2(n8372), .ZN(n7975) );
  NAND2_X1 U10268 ( .A1(n7996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7973) );
  XNOR2_X1 U10269 ( .A(n7973), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U10270 ( .A1(n8178), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9954), .B2(
        n8177), .ZN(n7974) );
  NAND2_X1 U10271 ( .A1(n7975), .A2(n7974), .ZN(n14550) );
  MUX2_X1 U10272 ( .A(n13682), .B(n14550), .S(n8377), .Z(n7980) );
  NAND2_X1 U10273 ( .A1(n7976), .A2(n7980), .ZN(n7978) );
  MUX2_X1 U10274 ( .A(n13682), .B(n14550), .S(n8375), .Z(n7977) );
  NAND2_X1 U10275 ( .A1(n7978), .A2(n7977), .ZN(n7985) );
  INV_X1 U10276 ( .A(n7980), .ZN(n7981) );
  AND2_X1 U10277 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  NAND2_X1 U10278 ( .A1(n7979), .A2(n7983), .ZN(n7984) );
  NAND2_X1 U10279 ( .A1(n7985), .A2(n7984), .ZN(n8002) );
  INV_X1 U10280 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9967) );
  OR2_X1 U10281 ( .A1(n7876), .A2(n9967), .ZN(n7993) );
  INV_X1 U10282 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9957) );
  OR2_X1 U10283 ( .A1(n8184), .A2(n9957), .ZN(n7992) );
  INV_X1 U10284 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7986) );
  OAI21_X1 U10285 ( .B1(n7988), .B2(n7987), .A(n7986), .ZN(n7989) );
  NAND2_X1 U10286 ( .A1(n7989), .A2(n8004), .ZN(n11400) );
  OR2_X1 U10287 ( .A1(n7889), .A2(n11400), .ZN(n7991) );
  NAND2_X1 U10288 ( .A1(n8331), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7990) );
  NAND4_X1 U10289 ( .A1(n7993), .A2(n7992), .A3(n7991), .A4(n7990), .ZN(n13681) );
  XNOR2_X1 U10290 ( .A(n7995), .B(n7994), .ZN(n9818) );
  NAND2_X1 U10291 ( .A1(n9818), .A2(n8372), .ZN(n8000) );
  OAI21_X1 U10292 ( .B1(n7996), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8036) );
  INV_X1 U10293 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U10294 ( .A1(n8036), .A2(n7997), .ZN(n8014) );
  OR2_X1 U10295 ( .A1(n8036), .A2(n7997), .ZN(n7998) );
  AOI22_X1 U10296 ( .A1(n9968), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n7999) );
  MUX2_X1 U10297 ( .A(n13681), .B(n14557), .S(n8375), .Z(n8003) );
  MUX2_X1 U10298 ( .A(n13681), .B(n14557), .S(n8377), .Z(n8001) );
  NAND2_X1 U10299 ( .A1(n8332), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U10300 ( .A1(n6485), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8009) );
  INV_X1 U10301 ( .A(n8025), .ZN(n8006) );
  NAND2_X1 U10302 ( .A1(n8004), .A2(n9980), .ZN(n8005) );
  NAND2_X1 U10303 ( .A1(n8006), .A2(n8005), .ZN(n11598) );
  OR2_X1 U10304 ( .A1(n7889), .A2(n11598), .ZN(n8008) );
  NAND2_X1 U10305 ( .A1(n8331), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8007) );
  NAND4_X1 U10306 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n13680) );
  XNOR2_X1 U10307 ( .A(n8011), .B(SI_10_), .ZN(n8012) );
  XNOR2_X1 U10308 ( .A(n8013), .B(n8012), .ZN(n9890) );
  NAND2_X1 U10309 ( .A1(n9890), .A2(n8372), .ZN(n8017) );
  NAND2_X1 U10310 ( .A1(n8014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U10311 ( .A(n8015), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U10312 ( .A1(n9969), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8016) );
  MUX2_X1 U10313 ( .A(n13680), .B(n11591), .S(n8377), .Z(n8021) );
  MUX2_X1 U10314 ( .A(n13680), .B(n11591), .S(n8375), .Z(n8018) );
  NAND2_X1 U10315 ( .A1(n8019), .A2(n8018), .ZN(n8024) );
  INV_X1 U10316 ( .A(n8020), .ZN(n8022) );
  NAND2_X1 U10317 ( .A1(n8022), .A2(n7028), .ZN(n8023) );
  NAND2_X1 U10318 ( .A1(n8024), .A2(n8023), .ZN(n8042) );
  OR2_X1 U10319 ( .A1(n8025), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10320 ( .A1(n8049), .A2(n8026), .ZN(n14281) );
  OR2_X1 U10321 ( .A1(n7889), .A2(n14281), .ZN(n8031) );
  NAND2_X1 U10322 ( .A1(n8332), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8030) );
  INV_X1 U10323 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8027) );
  OR2_X1 U10324 ( .A1(n8184), .A2(n8027), .ZN(n8029) );
  NAND2_X1 U10325 ( .A1(n8331), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8028) );
  NAND4_X1 U10326 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n13679) );
  XNOR2_X1 U10327 ( .A(n8033), .B(n8032), .ZN(n9900) );
  NAND2_X1 U10328 ( .A1(n9900), .A2(n8372), .ZN(n8039) );
  OR2_X1 U10329 ( .A1(n8034), .A2(n8135), .ZN(n8035) );
  NAND2_X1 U10330 ( .A1(n8036), .A2(n8035), .ZN(n8056) );
  INV_X1 U10331 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8037) );
  XNOR2_X1 U10332 ( .A(n8056), .B(n8037), .ZN(n10150) );
  AOI22_X1 U10333 ( .A1(n10150), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n8038) );
  MUX2_X1 U10334 ( .A(n13679), .B(n14276), .S(n8375), .Z(n8043) );
  NAND2_X1 U10335 ( .A1(n8042), .A2(n8043), .ZN(n8041) );
  MUX2_X1 U10336 ( .A(n13679), .B(n14276), .S(n8377), .Z(n8040) );
  NAND2_X1 U10337 ( .A1(n8041), .A2(n8040), .ZN(n8047) );
  INV_X1 U10338 ( .A(n8042), .ZN(n8045) );
  INV_X1 U10339 ( .A(n8043), .ZN(n8044) );
  NAND2_X1 U10340 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  OR2_X1 U10341 ( .A1(n7876), .A2(n10143), .ZN(n8054) );
  INV_X1 U10342 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10149) );
  OR2_X1 U10343 ( .A1(n8184), .A2(n10149), .ZN(n8053) );
  NAND2_X1 U10344 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U10345 ( .A1(n8064), .A2(n8050), .ZN(n11707) );
  OR2_X1 U10346 ( .A1(n7889), .A2(n11707), .ZN(n8052) );
  NAND2_X1 U10347 ( .A1(n8331), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8051) );
  NAND4_X1 U10348 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n13678) );
  XNOR2_X1 U10349 ( .A(n8055), .B(n7386), .ZN(n10067) );
  NAND2_X1 U10350 ( .A1(n10067), .A2(n8372), .ZN(n8059) );
  NAND2_X1 U10351 ( .A1(n8057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8075) );
  XNOR2_X1 U10352 ( .A(n8075), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U10353 ( .A1(n10387), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8058) );
  MUX2_X1 U10354 ( .A(n13678), .B(n11701), .S(n8377), .Z(n8061) );
  MUX2_X1 U10355 ( .A(n13678), .B(n11701), .S(n8375), .Z(n8060) );
  INV_X1 U10356 ( .A(n8061), .ZN(n8062) );
  NAND2_X1 U10357 ( .A1(n8332), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10358 ( .A1(n6485), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8069) );
  INV_X1 U10359 ( .A(n8096), .ZN(n8066) );
  NAND2_X1 U10360 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  NAND2_X1 U10361 ( .A1(n8066), .A2(n8065), .ZN(n11822) );
  OR2_X1 U10362 ( .A1(n7889), .A2(n11822), .ZN(n8068) );
  NAND2_X1 U10363 ( .A1(n8331), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8067) );
  NAND4_X1 U10364 ( .A1(n8070), .A2(n8069), .A3(n8068), .A4(n8067), .ZN(n13677) );
  XNOR2_X1 U10365 ( .A(n8071), .B(n9798), .ZN(n8072) );
  XNOR2_X1 U10366 ( .A(n8073), .B(n8072), .ZN(n10304) );
  NAND2_X1 U10367 ( .A1(n10304), .A2(n8372), .ZN(n8081) );
  INV_X1 U10368 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10369 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  NAND2_X1 U10370 ( .A1(n8076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8078) );
  INV_X1 U10371 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10372 ( .A1(n8078), .A2(n8077), .ZN(n8091) );
  OR2_X1 U10373 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  AOI22_X1 U10374 ( .A1(n10497), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8080) );
  MUX2_X1 U10375 ( .A(n13677), .B(n11824), .S(n8375), .Z(n8085) );
  MUX2_X1 U10376 ( .A(n13677), .B(n11824), .S(n8377), .Z(n8082) );
  NAND2_X1 U10377 ( .A1(n8083), .A2(n8082), .ZN(n8089) );
  INV_X1 U10378 ( .A(n8084), .ZN(n8087) );
  INV_X1 U10379 ( .A(n8085), .ZN(n8086) );
  NAND2_X1 U10380 ( .A1(n8087), .A2(n8086), .ZN(n8088) );
  NAND2_X1 U10381 ( .A1(n8089), .A2(n8088), .ZN(n8101) );
  XNOR2_X1 U10382 ( .A(n8102), .B(n8090), .ZN(n10613) );
  NAND2_X1 U10383 ( .A1(n10613), .A2(n8372), .ZN(n8094) );
  NAND2_X1 U10384 ( .A1(n8091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8092) );
  XNOR2_X1 U10385 ( .A(n8092), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U10386 ( .A1(n10967), .A2(n8177), .B1(n8178), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8093) );
  INV_X1 U10387 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10959) );
  INV_X1 U10388 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8095) );
  OAI22_X1 U10389 ( .A1(n7876), .A2(n10959), .B1(n8184), .B2(n8095), .ZN(n8100) );
  OR2_X1 U10390 ( .A1(n8096), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10391 ( .A1(n8116), .A2(n8097), .ZN(n14252) );
  NAND2_X1 U10392 ( .A1(n8331), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8098) );
  OAI21_X1 U10393 ( .B1(n14252), .B2(n7889), .A(n8098), .ZN(n8099) );
  INV_X1 U10394 ( .A(n13676), .ZN(n12041) );
  NAND2_X1 U10395 ( .A1(n14247), .A2(n12041), .ZN(n8123) );
  NAND2_X1 U10396 ( .A1(n8101), .A2(n11615), .ZN(n8127) );
  INV_X1 U10397 ( .A(n8102), .ZN(n8104) );
  NAND2_X1 U10398 ( .A1(n8104), .A2(n8103), .ZN(n8107) );
  NAND2_X1 U10399 ( .A1(n8105), .A2(n9822), .ZN(n8106) );
  NAND2_X1 U10400 ( .A1(n8107), .A2(n8106), .ZN(n8110) );
  XNOR2_X1 U10401 ( .A(n8108), .B(SI_15_), .ZN(n8109) );
  XNOR2_X1 U10402 ( .A(n8110), .B(n8109), .ZN(n10679) );
  NAND2_X1 U10403 ( .A1(n10679), .A2(n8372), .ZN(n8114) );
  NAND2_X1 U10404 ( .A1(n8111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8112) );
  XNOR2_X1 U10405 ( .A(n8112), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U10406 ( .A1(n8178), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8177), 
        .B2(n10970), .ZN(n8113) );
  NAND2_X1 U10407 ( .A1(n8116), .A2(n8115), .ZN(n8117) );
  NAND2_X1 U10408 ( .A1(n8129), .A2(n8117), .ZN(n14302) );
  OR2_X1 U10409 ( .A1(n14302), .A2(n7889), .ZN(n8122) );
  NAND2_X1 U10410 ( .A1(n6485), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10411 ( .A1(n8331), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8118) );
  AND2_X1 U10412 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  INV_X1 U10413 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11668) );
  OR2_X1 U10414 ( .A1(n7876), .A2(n11668), .ZN(n8120) );
  NAND2_X1 U10415 ( .A1(n14298), .A2(n12055), .ZN(n8397) );
  AND2_X1 U10416 ( .A1(n8397), .A2(n8123), .ZN(n8125) );
  AND2_X1 U10417 ( .A1(n11795), .A2(n11662), .ZN(n8124) );
  MUX2_X1 U10418 ( .A(n8125), .B(n8124), .S(n8375), .Z(n8126) );
  NAND2_X1 U10419 ( .A1(n8127), .A2(n8126), .ZN(n8145) );
  MUX2_X1 U10420 ( .A(n8397), .B(n11795), .S(n8377), .Z(n8144) );
  AND2_X1 U10421 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  OR2_X1 U10422 ( .A1(n8130), .A2(n8160), .ZN(n14261) );
  AOI22_X1 U10423 ( .A1(n8331), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6485), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n8132) );
  INV_X1 U10424 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10963) );
  OR2_X1 U10425 ( .A1(n7876), .A2(n10963), .ZN(n8131) );
  OAI211_X1 U10426 ( .C1(n14261), .C2(n7889), .A(n8132), .B(n8131), .ZN(n13674) );
  XNOR2_X1 U10427 ( .A(n8134), .B(n8133), .ZN(n10531) );
  NAND2_X1 U10428 ( .A1(n10531), .A2(n8372), .ZN(n8138) );
  NOR2_X1 U10429 ( .A1(n8111), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8152) );
  OR2_X1 U10430 ( .A1(n8152), .A2(n8135), .ZN(n8136) );
  XNOR2_X1 U10431 ( .A(n8136), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U10432 ( .A1(n8178), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8177), 
        .B2(n13763), .ZN(n8137) );
  MUX2_X1 U10433 ( .A(n13674), .B(n14256), .S(n8377), .Z(n8140) );
  AND2_X1 U10434 ( .A1(n8144), .A2(n8140), .ZN(n8139) );
  NAND2_X1 U10435 ( .A1(n8145), .A2(n8139), .ZN(n8143) );
  INV_X1 U10436 ( .A(n8140), .ZN(n8141) );
  MUX2_X1 U10437 ( .A(n13674), .B(n14256), .S(n8375), .Z(n8146) );
  OR2_X1 U10438 ( .A1(n8141), .A2(n8146), .ZN(n8142) );
  INV_X1 U10439 ( .A(n8146), .ZN(n8147) );
  XNOR2_X1 U10440 ( .A(n8148), .B(n7638), .ZN(n8149) );
  XNOR2_X1 U10441 ( .A(n8150), .B(n8149), .ZN(n10675) );
  NAND2_X1 U10442 ( .A1(n10675), .A2(n8372), .ZN(n8159) );
  INV_X1 U10443 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10444 ( .A1(n8152), .A2(n8151), .ZN(n8154) );
  NAND2_X1 U10445 ( .A1(n8154), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8153) );
  MUX2_X1 U10446 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8153), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8157) );
  INV_X1 U10447 ( .A(n8154), .ZN(n8156) );
  INV_X1 U10448 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10449 ( .A1(n8156), .A2(n8155), .ZN(n8175) );
  AOI22_X1 U10450 ( .A1(n8178), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8177), 
        .B2(n13789), .ZN(n8158) );
  NOR2_X1 U10451 ( .A1(n8160), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8161) );
  OR2_X1 U10452 ( .A1(n8181), .A2(n8161), .ZN(n14272) );
  AOI22_X1 U10453 ( .A1(n8332), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n6485), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10454 ( .A1(n8331), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8162) );
  OAI211_X1 U10455 ( .C1(n14272), .C2(n7889), .A(n8163), .B(n8162), .ZN(n14002) );
  NAND2_X1 U10456 ( .A1(n12068), .A2(n14002), .ZN(n12008) );
  AOI22_X1 U10457 ( .A1(n8178), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13964), 
        .B2(n8177), .ZN(n8165) );
  NAND2_X1 U10458 ( .A1(n8183), .A2(n8166), .ZN(n8167) );
  NAND2_X1 U10459 ( .A1(n8199), .A2(n8167), .ZN(n13986) );
  OR2_X1 U10460 ( .A1(n13986), .A2(n7889), .ZN(n8172) );
  INV_X1 U10461 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13801) );
  NAND2_X1 U10462 ( .A1(n8331), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10463 ( .A1(n8332), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U10464 ( .C1(n13801), .C2(n8184), .A(n8169), .B(n8168), .ZN(n8170)
         );
  INV_X1 U10465 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U10466 ( .A1(n8172), .A2(n8171), .ZN(n14004) );
  XNOR2_X1 U10467 ( .A(n14085), .B(n14004), .ZN(n13982) );
  XNOR2_X1 U10468 ( .A(n8174), .B(n8173), .ZN(n10843) );
  NAND2_X1 U10469 ( .A1(n10843), .A2(n8372), .ZN(n8180) );
  NAND2_X1 U10470 ( .A1(n8175), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8176) );
  XNOR2_X1 U10471 ( .A(n8176), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U10472 ( .A1(n8178), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8177), 
        .B2(n13804), .ZN(n8179) );
  OR2_X1 U10473 ( .A1(n8181), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10474 ( .A1(n8183), .A2(n8182), .ZN(n14292) );
  OR2_X1 U10475 ( .A1(n14292), .A2(n7889), .ZN(n8189) );
  INV_X1 U10476 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14009) );
  NAND2_X1 U10477 ( .A1(n8331), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8186) );
  INV_X1 U10478 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13791) );
  OR2_X1 U10479 ( .A1(n8184), .A2(n13791), .ZN(n8185) );
  OAI211_X1 U10480 ( .C1(n7876), .C2(n14009), .A(n8186), .B(n8185), .ZN(n8187)
         );
  INV_X1 U10481 ( .A(n8187), .ZN(n8188) );
  NAND2_X1 U10482 ( .A1(n8189), .A2(n8188), .ZN(n13673) );
  XNOR2_X1 U10483 ( .A(n14092), .B(n13673), .ZN(n14000) );
  MUX2_X1 U10484 ( .A(n14002), .B(n12068), .S(n8377), .Z(n8190) );
  INV_X1 U10485 ( .A(n13673), .ZN(n13600) );
  NAND3_X1 U10486 ( .A1(n14092), .A2(n13600), .A3(n8377), .ZN(n8192) );
  OR3_X1 U10487 ( .A1(n14092), .A2(n13600), .A3(n8377), .ZN(n8191) );
  NAND2_X1 U10488 ( .A1(n8192), .A2(n8191), .ZN(n8193) );
  NAND2_X1 U10489 ( .A1(n13982), .A2(n8193), .ZN(n8197) );
  NAND2_X1 U10490 ( .A1(n14004), .A2(n8375), .ZN(n8195) );
  INV_X1 U10491 ( .A(n14004), .ZN(n11992) );
  NAND2_X1 U10492 ( .A1(n11992), .A2(n8377), .ZN(n8194) );
  MUX2_X1 U10493 ( .A(n8195), .B(n8194), .S(n14085), .Z(n8196) );
  AND2_X1 U10494 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  NAND2_X1 U10495 ( .A1(n8199), .A2(n13639), .ZN(n8201) );
  INV_X1 U10496 ( .A(n8217), .ZN(n8200) );
  NAND2_X1 U10497 ( .A1(n8201), .A2(n8200), .ZN(n13974) );
  OR2_X1 U10498 ( .A1(n13974), .A2(n7889), .ZN(n8208) );
  INV_X1 U10499 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U10500 ( .A1(n6485), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U10501 ( .A1(n8332), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8202) );
  OAI211_X1 U10502 ( .C1(n6482), .C2(n8204), .A(n8203), .B(n8202), .ZN(n8206)
         );
  INV_X1 U10503 ( .A(n8206), .ZN(n8207) );
  XNOR2_X1 U10504 ( .A(n8225), .B(n10724), .ZN(n8222) );
  XNOR2_X1 U10505 ( .A(n8222), .B(n8223), .ZN(n11296) );
  NAND2_X1 U10506 ( .A1(n11296), .A2(n8372), .ZN(n8210) );
  NAND2_X1 U10507 ( .A1(n8178), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8209) );
  MUX2_X1 U10508 ( .A(n13614), .B(n14077), .S(n8375), .Z(n8212) );
  INV_X1 U10509 ( .A(n13614), .ZN(n13672) );
  MUX2_X1 U10510 ( .A(n13672), .B(n8395), .S(n8377), .Z(n8211) );
  OAI21_X1 U10511 ( .B1(n8213), .B2(n8212), .A(n8211), .ZN(n8215) );
  NAND2_X1 U10512 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U10513 ( .A1(n8331), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U10514 ( .A1(n8332), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8220) );
  OAI21_X1 U10515 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n8217), .A(n8216), .ZN(
        n13958) );
  OR2_X1 U10516 ( .A1(n7889), .A2(n13958), .ZN(n8219) );
  NAND2_X1 U10517 ( .A1(n6485), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8218) );
  NAND4_X1 U10518 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n13671) );
  INV_X1 U10519 ( .A(n8222), .ZN(n8224) );
  NAND2_X1 U10520 ( .A1(n8224), .A2(n8223), .ZN(n8227) );
  OR2_X1 U10521 ( .A1(n8225), .A2(n10724), .ZN(n8226) );
  NAND2_X1 U10522 ( .A1(n8227), .A2(n8226), .ZN(n8230) );
  XNOR2_X1 U10523 ( .A(n8228), .B(SI_21_), .ZN(n8229) );
  NAND2_X1 U10524 ( .A1(n11509), .A2(n8372), .ZN(n8232) );
  NAND2_X1 U10525 ( .A1(n8178), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8231) );
  NAND2_X2 U10526 ( .A1(n8232), .A2(n8231), .ZN(n14071) );
  MUX2_X1 U10527 ( .A(n13671), .B(n14071), .S(n8377), .Z(n8234) );
  MUX2_X1 U10528 ( .A(n13671), .B(n14071), .S(n8375), .Z(n8233) );
  INV_X1 U10529 ( .A(n8234), .ZN(n8235) );
  NAND2_X1 U10530 ( .A1(n8332), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10531 ( .A1(n6485), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8240) );
  OAI21_X1 U10532 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8237), .A(n8236), .ZN(
        n13948) );
  OR2_X1 U10533 ( .A1(n7889), .A2(n13948), .ZN(n8239) );
  NAND2_X1 U10534 ( .A1(n8331), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8238) );
  NAND4_X1 U10535 ( .A1(n8241), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n13670) );
  NAND2_X1 U10536 ( .A1(n8243), .A2(n8242), .ZN(n8244) );
  XNOR2_X1 U10537 ( .A(n8245), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14130) );
  MUX2_X1 U10538 ( .A(n13670), .B(n13947), .S(n8375), .Z(n8249) );
  MUX2_X1 U10539 ( .A(n13670), .B(n13947), .S(n8377), .Z(n8246) );
  NAND2_X1 U10540 ( .A1(n8247), .A2(n8246), .ZN(n8253) );
  INV_X1 U10541 ( .A(n8248), .ZN(n8251) );
  INV_X1 U10542 ( .A(n8249), .ZN(n8250) );
  NAND2_X1 U10543 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  NAND2_X1 U10544 ( .A1(n8253), .A2(n8252), .ZN(n8264) );
  NAND2_X1 U10545 ( .A1(n8331), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10546 ( .A1(n8332), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8258) );
  OAI21_X1 U10547 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8255), .A(n8254), .ZN(
        n13935) );
  OR2_X1 U10548 ( .A1(n7889), .A2(n13935), .ZN(n8257) );
  NAND2_X1 U10549 ( .A1(n6485), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8256) );
  NAND4_X1 U10550 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n13669) );
  XNOR2_X1 U10551 ( .A(n8260), .B(SI_23_), .ZN(n11625) );
  NAND2_X1 U10552 ( .A1(n11625), .A2(n8372), .ZN(n8262) );
  NAND2_X1 U10553 ( .A1(n8178), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8261) );
  MUX2_X1 U10554 ( .A(n13669), .B(n14058), .S(n8377), .Z(n8265) );
  MUX2_X1 U10555 ( .A(n13669), .B(n14058), .S(n8375), .Z(n8263) );
  INV_X1 U10556 ( .A(n8265), .ZN(n8266) );
  NAND2_X1 U10557 ( .A1(n8331), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8272) );
  NAND2_X1 U10558 ( .A1(n8332), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8271) );
  OAI21_X1 U10559 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n8268), .A(n8267), .ZN(
        n13913) );
  OR2_X1 U10560 ( .A1(n7889), .A2(n13913), .ZN(n8270) );
  NAND2_X1 U10561 ( .A1(n6485), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8269) );
  NAND4_X1 U10562 ( .A1(n8272), .A2(n8271), .A3(n8270), .A4(n8269), .ZN(n13668) );
  XNOR2_X1 U10563 ( .A(n8274), .B(n8273), .ZN(n11777) );
  NAND2_X1 U10564 ( .A1(n11777), .A2(n8372), .ZN(n8276) );
  NAND2_X1 U10565 ( .A1(n8178), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8275) );
  MUX2_X1 U10566 ( .A(n13668), .B(n13920), .S(n8375), .Z(n8280) );
  MUX2_X1 U10567 ( .A(n13668), .B(n13920), .S(n8377), .Z(n8277) );
  NAND2_X1 U10568 ( .A1(n8278), .A2(n8277), .ZN(n8284) );
  INV_X1 U10569 ( .A(n8279), .ZN(n8282) );
  INV_X1 U10570 ( .A(n8280), .ZN(n8281) );
  NAND2_X1 U10571 ( .A1(n8282), .A2(n8281), .ZN(n8283) );
  NAND2_X1 U10572 ( .A1(n8331), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10573 ( .A1(n8332), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8288) );
  OAI21_X1 U10574 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n8285), .A(n8298), .ZN(
        n13895) );
  OR2_X1 U10575 ( .A1(n7889), .A2(n13895), .ZN(n8287) );
  NAND2_X1 U10576 ( .A1(n6485), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8286) );
  NAND4_X1 U10577 ( .A1(n8289), .A2(n8288), .A3(n8287), .A4(n8286), .ZN(n13667) );
  XNOR2_X1 U10578 ( .A(n8291), .B(n8290), .ZN(n11880) );
  NAND2_X1 U10579 ( .A1(n11880), .A2(n8372), .ZN(n8293) );
  NAND2_X1 U10580 ( .A1(n8178), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8292) );
  MUX2_X1 U10581 ( .A(n13667), .B(n14045), .S(n8377), .Z(n8295) );
  MUX2_X1 U10582 ( .A(n13667), .B(n14045), .S(n8375), .Z(n8294) );
  INV_X1 U10583 ( .A(n8295), .ZN(n8296) );
  NAND2_X1 U10584 ( .A1(n8331), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U10585 ( .A1(n8332), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8302) );
  INV_X1 U10586 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10587 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  NAND2_X1 U10588 ( .A1(n8318), .A2(n8299), .ZN(n13875) );
  OR2_X1 U10589 ( .A1(n7889), .A2(n13875), .ZN(n8301) );
  NAND2_X1 U10590 ( .A1(n6485), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8300) );
  NAND4_X1 U10591 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n13666) );
  XNOR2_X1 U10592 ( .A(n8304), .B(n11645), .ZN(n8305) );
  NAND2_X1 U10593 ( .A1(n13579), .A2(n8372), .ZN(n8308) );
  NAND2_X1 U10594 ( .A1(n8178), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8307) );
  NAND2_X2 U10595 ( .A1(n8308), .A2(n8307), .ZN(n14039) );
  MUX2_X1 U10596 ( .A(n13666), .B(n14039), .S(n8375), .Z(n8312) );
  NAND2_X1 U10597 ( .A1(n8311), .A2(n8312), .ZN(n8310) );
  MUX2_X1 U10598 ( .A(n13666), .B(n14039), .S(n8377), .Z(n8309) );
  NAND2_X1 U10599 ( .A1(n8310), .A2(n8309), .ZN(n8316) );
  INV_X1 U10600 ( .A(n8312), .ZN(n8313) );
  NAND2_X1 U10601 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U10602 ( .A1(n8332), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10603 ( .A1(n6485), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8322) );
  INV_X1 U10604 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10605 ( .A1(n8318), .A2(n8317), .ZN(n8319) );
  NAND2_X1 U10606 ( .A1(n8333), .A2(n8319), .ZN(n13588) );
  OR2_X1 U10607 ( .A1(n7889), .A2(n13588), .ZN(n8321) );
  NAND2_X1 U10608 ( .A1(n8331), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8320) );
  NAND4_X1 U10609 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n13834) );
  XNOR2_X1 U10610 ( .A(n8324), .B(SI_27_), .ZN(n8325) );
  XNOR2_X1 U10611 ( .A(n8326), .B(n8325), .ZN(n13575) );
  NAND2_X1 U10612 ( .A1(n13575), .A2(n8372), .ZN(n8328) );
  NAND2_X1 U10613 ( .A1(n8178), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8327) );
  MUX2_X1 U10614 ( .A(n13834), .B(n14033), .S(n8377), .Z(n8330) );
  MUX2_X1 U10615 ( .A(n13834), .B(n14033), .S(n8375), .Z(n8329) );
  NAND2_X1 U10616 ( .A1(n8331), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10617 ( .A1(n8332), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8336) );
  INV_X1 U10618 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12146) );
  XNOR2_X1 U10619 ( .A(n8333), .B(n12146), .ZN(n13864) );
  OR2_X1 U10620 ( .A1(n7889), .A2(n13864), .ZN(n8335) );
  NAND2_X1 U10621 ( .A1(n6485), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8334) );
  NAND4_X1 U10622 ( .A1(n8337), .A2(n8336), .A3(n8335), .A4(n8334), .ZN(n13846) );
  NAND2_X1 U10623 ( .A1(n11927), .A2(n8372), .ZN(n8341) );
  NAND2_X1 U10624 ( .A1(n8178), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8340) );
  MUX2_X1 U10625 ( .A(n13846), .B(n14028), .S(n8375), .Z(n8345) );
  INV_X1 U10626 ( .A(n14028), .ZN(n13832) );
  MUX2_X1 U10627 ( .A(n13831), .B(n13832), .S(n8377), .Z(n8342) );
  AOI21_X1 U10628 ( .B1(n8344), .B2(n8345), .A(n8342), .ZN(n8343) );
  INV_X1 U10629 ( .A(n8344), .ZN(n8347) );
  INV_X1 U10630 ( .A(n8345), .ZN(n8346) );
  INV_X1 U10631 ( .A(n8358), .ZN(n8355) );
  NAND2_X1 U10632 ( .A1(n8352), .A2(n8351), .ZN(n8357) );
  INV_X1 U10633 ( .A(n8353), .ZN(n8354) );
  AOI21_X1 U10634 ( .B1(n8355), .B2(n8357), .A(n8354), .ZN(n8356) );
  INV_X1 U10635 ( .A(n8357), .ZN(n8359) );
  NAND2_X1 U10636 ( .A1(n14131), .A2(n10284), .ZN(n10295) );
  NAND2_X1 U10637 ( .A1(n8363), .A2(n11297), .ZN(n10470) );
  NAND2_X1 U10638 ( .A1(n10295), .A2(n10470), .ZN(n8364) );
  OR2_X1 U10639 ( .A1(n10281), .A2(n13897), .ZN(n10559) );
  AND2_X1 U10640 ( .A1(n8364), .A2(n10559), .ZN(n8379) );
  INV_X1 U10641 ( .A(n8365), .ZN(n8366) );
  OAI22_X1 U10642 ( .A1(n8368), .A2(n8367), .B1(n8366), .B2(n12528), .ZN(n8371) );
  MUX2_X1 U10643 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9733), .Z(n8369) );
  XNOR2_X1 U10644 ( .A(n8369), .B(SI_31_), .ZN(n8370) );
  XNOR2_X1 U10645 ( .A(n8371), .B(n8370), .ZN(n13565) );
  NAND2_X1 U10646 ( .A1(n13565), .A2(n8372), .ZN(n8374) );
  NAND2_X1 U10647 ( .A1(n8178), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8373) );
  XOR2_X1 U10648 ( .A(n13821), .B(n8378), .Z(n8414) );
  NOR2_X1 U10649 ( .A1(n14016), .A2(n8375), .ZN(n8388) );
  INV_X1 U10650 ( .A(n8379), .ZN(n8387) );
  NOR4_X1 U10651 ( .A1(n8388), .A2(n14016), .A3(n13821), .A4(n8387), .ZN(n8384) );
  INV_X1 U10652 ( .A(n8388), .ZN(n8376) );
  NOR3_X1 U10653 ( .A1(n8376), .A2(n8379), .A3(n13821), .ZN(n8383) );
  NOR2_X1 U10654 ( .A1(n8378), .A2(n8377), .ZN(n8386) );
  NAND3_X1 U10655 ( .A1(n14016), .A2(n8379), .A3(n13821), .ZN(n8381) );
  NAND3_X1 U10656 ( .A1(n8386), .A2(n13821), .A3(n8387), .ZN(n8380) );
  NAND2_X1 U10657 ( .A1(n11511), .A2(n10571), .ZN(n8416) );
  OAI211_X1 U10658 ( .C1(n8386), .C2(n8381), .A(n8380), .B(n8416), .ZN(n8382)
         );
  NOR4_X1 U10659 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), .ZN(n8419)
         );
  INV_X1 U10660 ( .A(n8386), .ZN(n8391) );
  AOI21_X1 U10661 ( .B1(n8388), .B2(n8392), .A(n8387), .ZN(n8389) );
  OAI211_X1 U10662 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8389), .ZN(n8418)
         );
  INV_X1 U10663 ( .A(n13834), .ZN(n13830) );
  XNOR2_X1 U10664 ( .A(n14033), .B(n13830), .ZN(n12006) );
  NAND2_X1 U10665 ( .A1(n14028), .A2(n13831), .ZN(n13837) );
  OR2_X1 U10666 ( .A1(n14028), .A2(n13831), .ZN(n8393) );
  NAND2_X1 U10667 ( .A1(n13837), .A2(n8393), .ZN(n13861) );
  NAND2_X1 U10668 ( .A1(n14039), .A2(n13621), .ZN(n12002) );
  OR2_X1 U10669 ( .A1(n14039), .A2(n13621), .ZN(n8394) );
  NAND2_X1 U10670 ( .A1(n12002), .A2(n8394), .ZN(n13878) );
  INV_X1 U10671 ( .A(n13668), .ZN(n13622) );
  XNOR2_X1 U10672 ( .A(n13920), .B(n13622), .ZN(n13905) );
  INV_X1 U10673 ( .A(n13667), .ZN(n13659) );
  XNOR2_X1 U10674 ( .A(n14045), .B(n13659), .ZN(n13888) );
  INV_X1 U10675 ( .A(n13669), .ZN(n11999) );
  XNOR2_X1 U10676 ( .A(n14058), .B(n11999), .ZN(n13926) );
  XNOR2_X1 U10677 ( .A(n14063), .B(n13670), .ZN(n13944) );
  NAND2_X1 U10678 ( .A1(n8395), .A2(n13614), .ZN(n8396) );
  NAND2_X1 U10679 ( .A1(n11994), .A2(n8396), .ZN(n13972) );
  NAND2_X1 U10680 ( .A1(n11795), .A2(n8397), .ZN(n11667) );
  NAND2_X1 U10681 ( .A1(n6513), .A2(n12008), .ZN(n11865) );
  XNOR2_X1 U10682 ( .A(n11824), .B(n13677), .ZN(n11609) );
  XNOR2_X1 U10683 ( .A(n11701), .B(n11699), .ZN(n11374) );
  INV_X1 U10684 ( .A(n13682), .ZN(n11390) );
  XNOR2_X1 U10685 ( .A(n14550), .B(n11390), .ZN(n10902) );
  XNOR2_X1 U10686 ( .A(n11027), .B(n13683), .ZN(n14405) );
  INV_X1 U10687 ( .A(n13684), .ZN(n10856) );
  NAND2_X1 U10688 ( .A1(n14533), .A2(n10856), .ZN(n10755) );
  OR2_X1 U10689 ( .A1(n14533), .A2(n10856), .ZN(n8399) );
  INV_X1 U10690 ( .A(n13685), .ZN(n8400) );
  NAND2_X1 U10691 ( .A1(n14431), .A2(n8400), .ZN(n10599) );
  OR2_X1 U10692 ( .A1(n14431), .A2(n8400), .ZN(n8401) );
  AND2_X1 U10693 ( .A1(n10576), .A2(n8403), .ZN(n10649) );
  NAND4_X1 U10694 ( .A1(n10581), .A2(n10618), .A3(n10649), .A4(n10579), .ZN(
        n8404) );
  NOR2_X1 U10695 ( .A1(n8404), .A2(n6937), .ZN(n8405) );
  NAND4_X1 U10696 ( .A1(n14405), .A2(n10596), .A3(n10595), .A4(n8405), .ZN(
        n8406) );
  NOR2_X1 U10697 ( .A1(n10902), .A2(n8406), .ZN(n8407) );
  XNOR2_X1 U10698 ( .A(n11591), .B(n13680), .ZN(n10901) );
  XNOR2_X1 U10699 ( .A(n14557), .B(n13681), .ZN(n14388) );
  NAND4_X1 U10700 ( .A1(n11227), .A2(n8407), .A3(n10901), .A4(n14388), .ZN(
        n8408) );
  NOR2_X1 U10701 ( .A1(n11374), .A2(n8408), .ZN(n8409) );
  AND2_X1 U10702 ( .A1(n11609), .A2(n8409), .ZN(n8410) );
  XNOR2_X1 U10703 ( .A(n14256), .B(n13674), .ZN(n11797) );
  NAND4_X1 U10704 ( .A1(n11865), .A2(n11615), .A3(n8410), .A4(n11797), .ZN(
        n8411) );
  INV_X1 U10705 ( .A(n13671), .ZN(n11995) );
  XNOR2_X1 U10706 ( .A(n14071), .B(n11995), .ZN(n13961) );
  OR4_X1 U10707 ( .A1(n13878), .A2(n13905), .A3(n13888), .A4(n8412), .ZN(n8413) );
  XNOR2_X1 U10708 ( .A(n13824), .B(n13842), .ZN(n8415) );
  INV_X1 U10709 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U10710 ( .A1(n8424), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8422) );
  INV_X1 U10711 ( .A(n9894), .ZN(n8423) );
  NAND2_X1 U10712 ( .A1(n8423), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11622) );
  NAND2_X1 U10713 ( .A1(n8425), .A2(n8421), .ZN(n8432) );
  INV_X1 U10714 ( .A(n8427), .ZN(n8428) );
  OAI21_X1 U10715 ( .B1(n8429), .B2(n8428), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8430) );
  MUX2_X1 U10716 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8430), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8431) );
  NAND2_X1 U10717 ( .A1(n10257), .A2(n10262), .ZN(n8435) );
  XNOR2_X1 U10718 ( .A(n8434), .B(n8433), .ZN(n10256) );
  OR2_X1 U10719 ( .A1(n10295), .A2(n10275), .ZN(n10727) );
  NAND2_X1 U10720 ( .A1(n10558), .A2(n10727), .ZN(n10293) );
  OR2_X1 U10721 ( .A1(n10295), .A2(n11928), .ZN(n13658) );
  NOR3_X1 U10722 ( .A1(n10293), .A2(n14122), .A3(n13658), .ZN(n8437) );
  OAI21_X1 U10723 ( .B1(n11622), .B2(n14131), .A(P1_B_REG_SCAN_IN), .ZN(n8436)
         );
  OR2_X1 U10724 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  OAI21_X1 U10725 ( .B1(n8439), .B2(n11622), .A(n8438), .ZN(P1_U3242) );
  NOR2_X1 U10726 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8442) );
  NOR2_X1 U10727 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8441) );
  NOR2_X1 U10728 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8446) );
  NOR2_X1 U10729 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8445) );
  NOR2_X1 U10730 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8444) );
  NAND2_X1 U10731 ( .A1(n6478), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8462) );
  INV_X1 U10732 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8454) );
  OR2_X1 U10733 ( .A1(n8966), .A2(n8454), .ZN(n8461) );
  INV_X1 U10734 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8456) );
  INV_X1 U10735 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10829) );
  INV_X1 U10736 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8464) );
  INV_X1 U10737 ( .A(n8467), .ZN(n8470) );
  INV_X1 U10738 ( .A(n8468), .ZN(n8469) );
  INV_X1 U10739 ( .A(n9040), .ZN(n8478) );
  AND3_X1 U10740 ( .A1(n11346), .A2(n10181), .A3(n8487), .ZN(n8481) );
  NAND2_X1 U10741 ( .A1(n9020), .A2(n8490), .ZN(n8493) );
  NAND2_X1 U10742 ( .A1(n9733), .A2(SI_0_), .ZN(n8482) );
  XNOR2_X1 U10743 ( .A(n8482), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13583) );
  NAND2_X1 U10744 ( .A1(n9053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8484) );
  MUX2_X1 U10745 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13583), .S(n9770), .Z(n10241)
         );
  NAND2_X2 U10746 ( .A1(n11346), .A2(n10181), .ZN(n10244) );
  AOI21_X1 U10747 ( .B1(n10202), .B2(n8487), .A(n10244), .ZN(n8488) );
  OAI21_X1 U10748 ( .B1(n8493), .B2(n10241), .A(n8488), .ZN(n8496) );
  NAND2_X1 U10749 ( .A1(n8492), .A2(n8491), .ZN(n8494) );
  NAND2_X1 U10750 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  NAND2_X1 U10751 ( .A1(n8496), .A2(n8495), .ZN(n8510) );
  INV_X1 U10752 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13415) );
  INV_X1 U10753 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13412) );
  INV_X1 U10754 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9777) );
  INV_X1 U10755 ( .A(n8501), .ZN(n9727) );
  INV_X1 U10756 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9734) );
  OR2_X1 U10757 ( .A1(n8990), .A2(n9734), .ZN(n8506) );
  NAND2_X1 U10758 ( .A1(n9770), .A2(n9733), .ZN(n8518) );
  OR2_X1 U10759 ( .A1(n8518), .A2(n9736), .ZN(n8504) );
  INV_X1 U10760 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10761 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8502) );
  XNOR2_X1 U10762 ( .A(n8503), .B(n8502), .ZN(n14600) );
  MUX2_X1 U10763 ( .A(n13200), .B(n10654), .S(n6512), .Z(n8507) );
  INV_X1 U10764 ( .A(n8507), .ZN(n8509) );
  MUX2_X1 U10765 ( .A(n13200), .B(n10654), .S(n8490), .Z(n8508) );
  OAI21_X1 U10766 ( .B1(n8510), .B2(n8509), .A(n8508), .ZN(n8512) );
  NAND2_X1 U10767 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10768 ( .A1(n6478), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8517) );
  INV_X1 U10769 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11350) );
  OR2_X1 U10770 ( .A1(n6476), .A2(n11350), .ZN(n8516) );
  INV_X1 U10771 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8513) );
  OR2_X1 U10772 ( .A1(n8966), .A2(n8513), .ZN(n8515) );
  INV_X1 U10773 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9778) );
  OR2_X1 U10774 ( .A1(n8526), .A2(n9778), .ZN(n8514) );
  OR2_X1 U10775 ( .A1(n8519), .A2(n8728), .ZN(n8520) );
  XNOR2_X1 U10776 ( .A(n8520), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9779) );
  MUX2_X1 U10777 ( .A(n13198), .B(n11356), .S(n8490), .Z(n8523) );
  NAND2_X1 U10778 ( .A1(n8524), .A2(n8523), .ZN(n8522) );
  MUX2_X1 U10779 ( .A(n13198), .B(n11356), .S(n8996), .Z(n8521) );
  NAND2_X1 U10780 ( .A1(n8522), .A2(n8521), .ZN(n8525) );
  OR2_X1 U10781 ( .A1(n6476), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8531) );
  INV_X1 U10782 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8527) );
  OR2_X1 U10783 ( .A1(n8526), .A2(n8527), .ZN(n8530) );
  INV_X1 U10784 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10785 ( .A1(n9737), .A2(n6489), .ZN(n8535) );
  OR2_X1 U10786 ( .A1(n8547), .A2(n8728), .ZN(n8533) );
  XNOR2_X1 U10787 ( .A(n8533), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U10788 ( .A1(n8814), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8815), .B2(
        n9780), .ZN(n8534) );
  MUX2_X1 U10789 ( .A(n13197), .B(n10694), .S(n6512), .Z(n8537) );
  MUX2_X1 U10790 ( .A(n13197), .B(n10694), .S(n8490), .Z(n8536) );
  INV_X1 U10791 ( .A(n8537), .ZN(n8538) );
  NAND2_X1 U10792 ( .A1(n6479), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8544) );
  INV_X1 U10793 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8539) );
  OR2_X1 U10794 ( .A1(n8966), .A2(n8539), .ZN(n8543) );
  AND2_X1 U10795 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8559) );
  INV_X1 U10796 ( .A(n8559), .ZN(n8561) );
  OAI21_X1 U10797 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8561), .ZN(n10998) );
  OR2_X1 U10798 ( .A1(n6476), .A2(n10998), .ZN(n8542) );
  INV_X1 U10799 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8540) );
  OR2_X1 U10800 ( .A1(n8526), .A2(n8540), .ZN(n8541) );
  NAND4_X1 U10801 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n13196) );
  NAND2_X1 U10802 ( .A1(n8545), .A2(n6490), .ZN(n8550) );
  INV_X1 U10803 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U10804 ( .A1(n8547), .A2(n8546), .ZN(n8569) );
  NAND2_X1 U10805 ( .A1(n8569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U10806 ( .A(n8548), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10807 ( .A1(n8814), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8815), .B2(
        n9781), .ZN(n8549) );
  MUX2_X1 U10808 ( .A(n13196), .B(n10994), .S(n8490), .Z(n8554) );
  NAND2_X1 U10809 ( .A1(n8553), .A2(n8554), .ZN(n8552) );
  MUX2_X1 U10810 ( .A(n13196), .B(n10994), .S(n8996), .Z(n8551) );
  NAND2_X1 U10811 ( .A1(n8552), .A2(n8551), .ZN(n8558) );
  INV_X1 U10812 ( .A(n8553), .ZN(n8556) );
  INV_X1 U10813 ( .A(n8554), .ZN(n8555) );
  NAND2_X1 U10814 ( .A1(n8556), .A2(n8555), .ZN(n8557) );
  NAND2_X1 U10815 ( .A1(n6478), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8567) );
  INV_X1 U10816 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11034) );
  OR2_X1 U10817 ( .A1(n8966), .A2(n11034), .ZN(n8566) );
  AND2_X1 U10818 ( .A1(n8559), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8576) );
  INV_X1 U10819 ( .A(n8576), .ZN(n8578) );
  INV_X1 U10820 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10821 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U10822 ( .A1(n8578), .A2(n8562), .ZN(n11035) );
  OR2_X1 U10823 ( .A1(n6476), .A2(n11035), .ZN(n8565) );
  INV_X1 U10824 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8563) );
  OR2_X1 U10825 ( .A1(n8526), .A2(n8563), .ZN(n8564) );
  NAND4_X1 U10826 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n13195) );
  NAND2_X1 U10827 ( .A1(n9755), .A2(n6489), .ZN(n8572) );
  NAND2_X1 U10828 ( .A1(n8586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8570) );
  XNOR2_X1 U10829 ( .A(n8570), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9782) );
  AOI22_X1 U10830 ( .A1(n8814), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8815), .B2(
        n9782), .ZN(n8571) );
  NAND2_X1 U10831 ( .A1(n8572), .A2(n8571), .ZN(n11052) );
  MUX2_X1 U10832 ( .A(n13195), .B(n11052), .S(n8996), .Z(n8574) );
  MUX2_X1 U10833 ( .A(n13195), .B(n11052), .S(n8490), .Z(n8573) );
  INV_X1 U10834 ( .A(n8574), .ZN(n8575) );
  NAND2_X1 U10835 ( .A1(n8986), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8585) );
  INV_X1 U10836 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11063) );
  OR2_X1 U10837 ( .A1(n8966), .A2(n11063), .ZN(n8584) );
  INV_X1 U10838 ( .A(n8601), .ZN(n8603) );
  INV_X1 U10839 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U10840 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  NAND2_X1 U10841 ( .A1(n8603), .A2(n8579), .ZN(n11067) );
  OR2_X1 U10842 ( .A1(n6476), .A2(n11067), .ZN(n8583) );
  INV_X1 U10843 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8581) );
  OR2_X1 U10844 ( .A1(n8580), .A2(n8581), .ZN(n8582) );
  NAND4_X1 U10845 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n13194) );
  NAND2_X1 U10846 ( .A1(n9762), .A2(n6490), .ZN(n8591) );
  INV_X1 U10847 ( .A(n8586), .ZN(n8588) );
  INV_X1 U10848 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U10849 ( .A1(n8588), .A2(n8587), .ZN(n8609) );
  NAND2_X1 U10850 ( .A1(n8609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10851 ( .A(n8589), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10852 ( .A1(n8814), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8815), .B2(
        n9848), .ZN(n8590) );
  NAND2_X1 U10853 ( .A1(n8591), .A2(n8590), .ZN(n14706) );
  MUX2_X1 U10854 ( .A(n13194), .B(n14706), .S(n8490), .Z(n8595) );
  NAND2_X1 U10855 ( .A1(n8594), .A2(n8595), .ZN(n8593) );
  MUX2_X1 U10856 ( .A(n13194), .B(n14706), .S(n8996), .Z(n8592) );
  NAND2_X1 U10857 ( .A1(n8593), .A2(n8592), .ZN(n8599) );
  INV_X1 U10858 ( .A(n8594), .ZN(n8597) );
  INV_X1 U10859 ( .A(n8595), .ZN(n8596) );
  NAND2_X1 U10860 ( .A1(n8597), .A2(n8596), .ZN(n8598) );
  INV_X1 U10861 ( .A(n8966), .ZN(n8985) );
  NAND2_X1 U10862 ( .A1(n8985), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8608) );
  INV_X1 U10863 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8600) );
  OR2_X1 U10864 ( .A1(n8580), .A2(n8600), .ZN(n8607) );
  NAND2_X1 U10865 ( .A1(n8601), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8618) );
  INV_X1 U10866 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U10867 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  NAND2_X1 U10868 ( .A1(n8618), .A2(n8604), .ZN(n11461) );
  OR2_X1 U10869 ( .A1(n6476), .A2(n11461), .ZN(n8606) );
  INV_X1 U10870 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9842) );
  OR2_X1 U10871 ( .A1(n8526), .A2(n9842), .ZN(n8605) );
  NAND4_X1 U10872 ( .A1(n8608), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(n13193) );
  NAND2_X1 U10873 ( .A1(n9794), .A2(n6490), .ZN(n8614) );
  INV_X1 U10874 ( .A(n8609), .ZN(n8611) );
  INV_X1 U10875 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10876 ( .A1(n8611), .A2(n8610), .ZN(n8625) );
  NAND2_X1 U10877 ( .A1(n8625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8612) );
  XNOR2_X1 U10878 ( .A(n8612), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10879 ( .A1(n8814), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8815), .B2(
        n9850), .ZN(n8613) );
  NAND2_X1 U10880 ( .A1(n8614), .A2(n8613), .ZN(n14714) );
  MUX2_X1 U10881 ( .A(n13193), .B(n14714), .S(n8996), .Z(n8616) );
  MUX2_X1 U10882 ( .A(n13193), .B(n14714), .S(n8490), .Z(n8615) );
  NAND2_X1 U10883 ( .A1(n6479), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8624) );
  INV_X1 U10884 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11482) );
  OR2_X1 U10885 ( .A1(n8966), .A2(n11482), .ZN(n8623) );
  INV_X1 U10886 ( .A(n8635), .ZN(n8637) );
  NAND2_X1 U10887 ( .A1(n8618), .A2(n8617), .ZN(n8619) );
  NAND2_X1 U10888 ( .A1(n8637), .A2(n8619), .ZN(n11481) );
  OR2_X1 U10889 ( .A1(n6476), .A2(n11481), .ZN(n8622) );
  INV_X1 U10890 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8620) );
  OR2_X1 U10891 ( .A1(n8526), .A2(n8620), .ZN(n8621) );
  NAND4_X1 U10892 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n13192) );
  NAND2_X1 U10893 ( .A1(n9800), .A2(n6490), .ZN(n8628) );
  NAND2_X1 U10894 ( .A1(n8644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8626) );
  XNOR2_X1 U10895 ( .A(n8626), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9876) );
  AOI22_X1 U10896 ( .A1(n8814), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8815), .B2(
        n9876), .ZN(n8627) );
  MUX2_X1 U10897 ( .A(n13192), .B(n11484), .S(n8490), .Z(n8632) );
  NAND2_X1 U10898 ( .A1(n8631), .A2(n8632), .ZN(n8630) );
  MUX2_X1 U10899 ( .A(n13192), .B(n11484), .S(n8996), .Z(n8629) );
  NAND2_X1 U10900 ( .A1(n8630), .A2(n8629), .ZN(n8651) );
  NAND2_X1 U10901 ( .A1(n8634), .A2(n8633), .ZN(n8650) );
  NAND2_X1 U10902 ( .A1(n6478), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8643) );
  INV_X1 U10903 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11338) );
  OR2_X1 U10904 ( .A1(n8966), .A2(n11338), .ZN(n8642) );
  NAND2_X1 U10905 ( .A1(n8635), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8655) );
  INV_X1 U10906 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10907 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  NAND2_X1 U10908 ( .A1(n8655), .A2(n8638), .ZN(n11337) );
  OR2_X1 U10909 ( .A1(n6476), .A2(n11337), .ZN(n8641) );
  INV_X1 U10910 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8639) );
  OR2_X1 U10911 ( .A1(n8526), .A2(n8639), .ZN(n8640) );
  NAND4_X1 U10912 ( .A1(n8643), .A2(n8642), .A3(n8641), .A4(n8640), .ZN(n13191) );
  NAND2_X1 U10913 ( .A1(n9818), .A2(n6489), .ZN(n8648) );
  INV_X1 U10914 ( .A(n8644), .ZN(n8645) );
  NAND2_X1 U10915 ( .A1(n8645), .A2(n7341), .ZN(n8661) );
  NAND2_X1 U10916 ( .A1(n8661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8646) );
  XNOR2_X1 U10917 ( .A(n8646), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U10918 ( .A1(n8814), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8815), .B2(
        n10127), .ZN(n8647) );
  MUX2_X1 U10919 ( .A(n13191), .B(n14727), .S(n8996), .Z(n8652) );
  MUX2_X1 U10920 ( .A(n13191), .B(n14727), .S(n8490), .Z(n8649) );
  INV_X1 U10921 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U10922 ( .A1(n6479), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8660) );
  INV_X1 U10923 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11502) );
  OR2_X1 U10924 ( .A1(n8966), .A2(n11502), .ZN(n8659) );
  INV_X1 U10925 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10926 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  NAND2_X1 U10927 ( .A1(n8674), .A2(n8656), .ZN(n11501) );
  OR2_X1 U10928 ( .A1(n6476), .A2(n11501), .ZN(n8658) );
  INV_X1 U10929 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10133) );
  OR2_X1 U10930 ( .A1(n8526), .A2(n10133), .ZN(n8657) );
  NAND4_X1 U10931 ( .A1(n8660), .A2(n8659), .A3(n8658), .A4(n8657), .ZN(n13190) );
  NAND2_X1 U10932 ( .A1(n9890), .A2(n6489), .ZN(n8664) );
  NAND2_X1 U10933 ( .A1(n8681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8662) );
  XNOR2_X1 U10934 ( .A(n8662), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U10935 ( .A1(n8814), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10171), 
        .B2(n8815), .ZN(n8663) );
  MUX2_X1 U10936 ( .A(n13190), .B(n14736), .S(n8490), .Z(n8668) );
  NAND2_X1 U10937 ( .A1(n8667), .A2(n8668), .ZN(n8666) );
  MUX2_X1 U10938 ( .A(n13190), .B(n14736), .S(n8996), .Z(n8665) );
  NAND2_X1 U10939 ( .A1(n8666), .A2(n8665), .ZN(n8672) );
  INV_X1 U10940 ( .A(n8667), .ZN(n8670) );
  INV_X1 U10941 ( .A(n8668), .ZN(n8669) );
  NAND2_X1 U10942 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  NAND2_X1 U10943 ( .A1(n8985), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8680) );
  INV_X1 U10944 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8673) );
  OR2_X1 U10945 ( .A1(n8526), .A2(n8673), .ZN(n8679) );
  INV_X1 U10946 ( .A(n8688), .ZN(n8690) );
  NAND2_X1 U10947 ( .A1(n8674), .A2(n11107), .ZN(n8675) );
  NAND2_X1 U10948 ( .A1(n8690), .A2(n8675), .ZN(n11288) );
  OR2_X1 U10949 ( .A1(n6476), .A2(n11288), .ZN(n8678) );
  INV_X1 U10950 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8676) );
  OR2_X1 U10951 ( .A1(n8580), .A2(n8676), .ZN(n8677) );
  NAND4_X1 U10952 ( .A1(n8680), .A2(n8679), .A3(n8678), .A4(n8677), .ZN(n13189) );
  NAND2_X1 U10953 ( .A1(n9900), .A2(n6490), .ZN(n8684) );
  OAI21_X1 U10954 ( .B1(n8681), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8682) );
  XNOR2_X1 U10955 ( .A(n8682), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U10956 ( .A1(n10172), .A2(n8815), .B1(n8814), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8683) );
  MUX2_X1 U10957 ( .A(n13189), .B(n11302), .S(n8996), .Z(n8686) );
  MUX2_X1 U10958 ( .A(n13189), .B(n11302), .S(n8490), .Z(n8685) );
  INV_X1 U10959 ( .A(n8686), .ZN(n8687) );
  NAND2_X1 U10960 ( .A1(n6478), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8696) );
  INV_X1 U10961 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11309) );
  OR2_X1 U10962 ( .A1(n8966), .A2(n11309), .ZN(n8695) );
  INV_X1 U10963 ( .A(n8704), .ZN(n8706) );
  INV_X1 U10964 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U10965 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  NAND2_X1 U10966 ( .A1(n8706), .A2(n8691), .ZN(n11423) );
  OR2_X1 U10967 ( .A1(n6476), .A2(n11423), .ZN(n8694) );
  INV_X1 U10968 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8692) );
  OR2_X1 U10969 ( .A1(n8526), .A2(n8692), .ZN(n8693) );
  NAND4_X1 U10970 ( .A1(n8696), .A2(n8695), .A3(n8694), .A4(n8693), .ZN(n13188) );
  NAND2_X1 U10971 ( .A1(n10067), .A2(n6489), .ZN(n8700) );
  NAND2_X1 U10972 ( .A1(n8697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8698) );
  XNOR2_X1 U10973 ( .A(n8698), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U10974 ( .A1(n8814), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8815), 
        .B2(n10516), .ZN(n8699) );
  MUX2_X1 U10975 ( .A(n13188), .B(n11520), .S(n8490), .Z(n8702) );
  INV_X1 U10976 ( .A(n13188), .ZN(n11519) );
  MUX2_X1 U10977 ( .A(n11519), .B(n6823), .S(n8996), .Z(n8701) );
  AOI21_X1 U10978 ( .B1(n8703), .B2(n8702), .A(n8701), .ZN(n8720) );
  NOR2_X1 U10979 ( .A1(n8703), .A2(n8702), .ZN(n8719) );
  NAND2_X1 U10980 ( .A1(n8986), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8712) );
  INV_X1 U10981 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U10982 ( .A1(n8706), .A2(n8705), .ZN(n8707) );
  NAND2_X1 U10983 ( .A1(n8722), .A2(n8707), .ZN(n11547) );
  OR2_X1 U10984 ( .A1(n6476), .A2(n11547), .ZN(n8711) );
  INV_X1 U10985 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11114) );
  OR2_X1 U10986 ( .A1(n8966), .A2(n11114), .ZN(n8710) );
  INV_X1 U10987 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8708) );
  OR2_X1 U10988 ( .A1(n8580), .A2(n8708), .ZN(n8709) );
  NAND2_X1 U10989 ( .A1(n10304), .A2(n6489), .ZN(n8718) );
  NAND2_X1 U10990 ( .A1(n8713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8714) );
  MUX2_X1 U10991 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8714), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8715) );
  INV_X1 U10992 ( .A(n8715), .ZN(n8716) );
  NOR2_X1 U10993 ( .A1(n8716), .A2(n8467), .ZN(n11123) );
  AOI22_X1 U10994 ( .A1(n8814), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8815), 
        .B2(n11123), .ZN(n8717) );
  MUX2_X1 U10995 ( .A(n11648), .B(n13539), .S(n8490), .Z(n8733) );
  INV_X1 U10996 ( .A(n11648), .ZN(n13187) );
  MUX2_X1 U10997 ( .A(n13187), .B(n11649), .S(n8996), .Z(n8732) );
  OAI22_X1 U10998 ( .A1(n8720), .A2(n8719), .B1(n8733), .B2(n8732), .ZN(n8735)
         );
  NAND2_X1 U10999 ( .A1(n6478), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8727) );
  INV_X1 U11000 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11652) );
  OR2_X1 U11001 ( .A1(n8966), .A2(n11652), .ZN(n8726) );
  INV_X1 U11002 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11126) );
  OR2_X1 U11003 ( .A1(n8526), .A2(n11126), .ZN(n8725) );
  NAND2_X1 U11004 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  NAND2_X1 U11005 ( .A1(n8766), .A2(n8723), .ZN(n14242) );
  OR2_X1 U11006 ( .A1(n6476), .A2(n14242), .ZN(n8724) );
  AND4_X1 U11007 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n11846)
         );
  NAND2_X1 U11008 ( .A1(n10613), .A2(n6490), .ZN(n8731) );
  OR2_X1 U11009 ( .A1(n8467), .A2(n8728), .ZN(n8729) );
  XNOR2_X1 U11010 ( .A(n8729), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U11011 ( .A1(n8814), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8815), 
        .B2(n11124), .ZN(n8730) );
  MUX2_X1 U11012 ( .A(n11846), .B(n13532), .S(n8490), .Z(n8737) );
  MUX2_X1 U11013 ( .A(n13186), .B(n14239), .S(n8996), .Z(n8736) );
  AOI22_X1 U11014 ( .A1(n8737), .A2(n8736), .B1(n8733), .B2(n8732), .ZN(n8734)
         );
  NAND2_X1 U11015 ( .A1(n8735), .A2(n8734), .ZN(n8782) );
  INV_X1 U11016 ( .A(n8736), .ZN(n8739) );
  INV_X1 U11017 ( .A(n8737), .ZN(n8738) );
  NAND2_X1 U11018 ( .A1(n8739), .A2(n8738), .ZN(n8781) );
  INV_X1 U11019 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11020 ( .A1(n8740), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8795) );
  INV_X1 U11021 ( .A(n8740), .ZN(n8753) );
  INV_X1 U11022 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11023 ( .A1(n8753), .A2(n8741), .ZN(n8742) );
  NAND2_X1 U11024 ( .A1(n8795), .A2(n8742), .ZN(n13401) );
  OR2_X1 U11025 ( .A1(n13401), .A2(n6476), .ZN(n8744) );
  AOI22_X1 U11026 ( .A1(n8985), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8986), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n8743) );
  OAI211_X1 U11027 ( .C1(n8580), .C2(n8745), .A(n8744), .B(n8743), .ZN(n13183)
         );
  NAND2_X1 U11028 ( .A1(n10675), .A2(n6490), .ZN(n8750) );
  NAND2_X1 U11029 ( .A1(n8746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8747) );
  MUX2_X1 U11030 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8747), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8748) );
  AOI22_X1 U11031 ( .A1(n8814), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n13201), 
        .B2(n8815), .ZN(n8749) );
  MUX2_X1 U11032 ( .A(n13183), .B(n13400), .S(n8996), .Z(n8788) );
  NAND2_X1 U11033 ( .A1(n13400), .A2(n13183), .ZN(n11931) );
  INV_X1 U11034 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U11035 ( .A1(n8768), .A2(n8751), .ZN(n8752) );
  NAND2_X1 U11036 ( .A1(n8753), .A2(n8752), .ZN(n13103) );
  OR2_X1 U11037 ( .A1(n13103), .A2(n6476), .ZN(n8757) );
  NAND2_X1 U11038 ( .A1(n6479), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11039 ( .A1(n8985), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8754) );
  AND2_X1 U11040 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  OAI211_X1 U11041 ( .C1(n8526), .C2(n11317), .A(n8757), .B(n8756), .ZN(n13184) );
  AND2_X1 U11042 ( .A1(n13184), .A2(n8490), .ZN(n8764) );
  NOR2_X1 U11043 ( .A1(n13184), .A2(n8490), .ZN(n8763) );
  NAND2_X1 U11044 ( .A1(n10531), .A2(n6489), .ZN(n8762) );
  INV_X1 U11045 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8758) );
  AND2_X1 U11046 ( .A1(n8775), .A2(n8758), .ZN(n8759) );
  OR2_X1 U11047 ( .A1(n8759), .A2(n8728), .ZN(n8760) );
  XNOR2_X1 U11048 ( .A(n8760), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U11049 ( .A1(n8814), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8815), 
        .B2(n11119), .ZN(n8761) );
  MUX2_X1 U11050 ( .A(n8764), .B(n8763), .S(n12157), .Z(n8765) );
  AOI21_X1 U11051 ( .B1(n8788), .B2(n11931), .A(n8765), .ZN(n8787) );
  NAND2_X1 U11052 ( .A1(n8766), .A2(n11855), .ZN(n8767) );
  AND2_X1 U11053 ( .A1(n8768), .A2(n8767), .ZN(n11858) );
  NAND2_X1 U11054 ( .A1(n11858), .A2(n6475), .ZN(n8774) );
  INV_X1 U11055 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8769) );
  OR2_X1 U11056 ( .A1(n8580), .A2(n8769), .ZN(n8773) );
  INV_X1 U11057 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11746) );
  OR2_X1 U11058 ( .A1(n8966), .A2(n11746), .ZN(n8772) );
  INV_X1 U11059 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8770) );
  OR2_X1 U11060 ( .A1(n8526), .A2(n8770), .ZN(n8771) );
  NAND2_X1 U11061 ( .A1(n10679), .A2(n6489), .ZN(n8778) );
  OR2_X1 U11062 ( .A1(n8775), .A2(n8728), .ZN(n8776) );
  XNOR2_X1 U11063 ( .A(n8776), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U11064 ( .A1(n8814), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8815), 
        .B2(n14653), .ZN(n8777) );
  AND2_X2 U11065 ( .A1(n8778), .A2(n8777), .ZN(n13523) );
  MUX2_X1 U11066 ( .A(n11854), .B(n13523), .S(n8490), .Z(n8784) );
  MUX2_X1 U11067 ( .A(n13185), .B(n11748), .S(n8996), .Z(n8783) );
  NAND2_X1 U11068 ( .A1(n8784), .A2(n8783), .ZN(n8779) );
  NAND2_X1 U11069 ( .A1(n8787), .A2(n8779), .ZN(n8780) );
  AOI21_X1 U11070 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8793) );
  INV_X1 U11071 ( .A(n8783), .ZN(n8786) );
  INV_X1 U11072 ( .A(n8784), .ZN(n8785) );
  INV_X1 U11073 ( .A(n13184), .ZN(n11947) );
  XNOR2_X1 U11074 ( .A(n12157), .B(n11947), .ZN(n11949) );
  AOI21_X1 U11075 ( .B1(n8786), .B2(n8785), .A(n11949), .ZN(n8791) );
  INV_X1 U11076 ( .A(n8787), .ZN(n8790) );
  NOR2_X1 U11077 ( .A1(n13400), .A2(n13183), .ZN(n8789) );
  OAI22_X1 U11078 ( .A1(n8791), .A2(n8790), .B1(n8789), .B2(n8788), .ZN(n8792)
         );
  INV_X1 U11079 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11080 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  NAND2_X1 U11081 ( .A1(n8805), .A2(n8796), .ZN(n13380) );
  AOI22_X1 U11082 ( .A1(n8985), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8986), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11083 ( .A1(n6479), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U11084 ( .C1(n13380), .C2(n6476), .A(n8798), .B(n8797), .ZN(n13182) );
  NAND2_X1 U11085 ( .A1(n10843), .A2(n6490), .ZN(n8802) );
  NAND2_X1 U11086 ( .A1(n8799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8800) );
  XNOR2_X1 U11087 ( .A(n8800), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14674) );
  AOI22_X1 U11088 ( .A1(n14674), .A2(n8815), .B1(n8814), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8801) );
  MUX2_X1 U11089 ( .A(n13182), .B(n13503), .S(n8490), .Z(n8804) );
  MUX2_X1 U11090 ( .A(n13182), .B(n13503), .S(n8996), .Z(n8803) );
  INV_X1 U11091 ( .A(n8826), .ZN(n8807) );
  NAND2_X1 U11092 ( .A1(n8805), .A2(n13078), .ZN(n8806) );
  NAND2_X1 U11093 ( .A1(n8807), .A2(n8806), .ZN(n13367) );
  OR2_X1 U11094 ( .A1(n13367), .A2(n6476), .ZN(n8813) );
  INV_X1 U11095 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11096 ( .A1(n6478), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11097 ( .A1(n8986), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8808) );
  OAI211_X1 U11098 ( .C1(n8966), .C2(n8810), .A(n8809), .B(n8808), .ZN(n8811)
         );
  INV_X1 U11099 ( .A(n8811), .ZN(n8812) );
  NAND2_X1 U11100 ( .A1(n8813), .A2(n8812), .ZN(n13181) );
  NAND2_X1 U11101 ( .A1(n10883), .A2(n6489), .ZN(n8817) );
  AOI22_X1 U11102 ( .A1(n10202), .A2(n8815), .B1(n8814), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8816) );
  MUX2_X1 U11103 ( .A(n13181), .B(n13498), .S(n8996), .Z(n8821) );
  NAND2_X1 U11104 ( .A1(n8820), .A2(n8821), .ZN(n8819) );
  MUX2_X1 U11105 ( .A(n13181), .B(n13498), .S(n8490), .Z(n8818) );
  NAND2_X1 U11106 ( .A1(n8819), .A2(n8818), .ZN(n8825) );
  INV_X1 U11107 ( .A(n8820), .ZN(n8823) );
  INV_X1 U11108 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U11109 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U11110 ( .A1(n8825), .A2(n8824), .ZN(n8837) );
  NOR2_X1 U11111 ( .A1(n8826), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8827) );
  OR2_X1 U11112 ( .A1(n8843), .A2(n8827), .ZN(n13353) );
  INV_X1 U11113 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U11114 ( .A1(n8985), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11115 ( .A1(n8986), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8828) );
  OAI211_X1 U11116 ( .C1(n8580), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8831)
         );
  INV_X1 U11117 ( .A(n8831), .ZN(n8832) );
  OAI21_X1 U11118 ( .B1(n13353), .B2(n6476), .A(n8832), .ZN(n13180) );
  NAND2_X1 U11119 ( .A1(n11296), .A2(n6490), .ZN(n8834) );
  OR2_X1 U11120 ( .A1(n8990), .A2(n7164), .ZN(n8833) );
  MUX2_X1 U11121 ( .A(n13180), .B(n12181), .S(n8490), .Z(n8838) );
  NAND2_X1 U11122 ( .A1(n8837), .A2(n8838), .ZN(n8836) );
  MUX2_X1 U11123 ( .A(n13180), .B(n12181), .S(n6512), .Z(n8835) );
  NAND2_X1 U11124 ( .A1(n8836), .A2(n8835), .ZN(n8842) );
  INV_X1 U11125 ( .A(n8837), .ZN(n8840) );
  INV_X1 U11126 ( .A(n8838), .ZN(n8839) );
  NAND2_X1 U11127 ( .A1(n8840), .A2(n8839), .ZN(n8841) );
  OR2_X1 U11128 ( .A1(n8843), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8844) );
  AND2_X1 U11129 ( .A1(n8844), .A2(n8855), .ZN(n13342) );
  NAND2_X1 U11130 ( .A1(n13342), .A2(n6475), .ZN(n8850) );
  INV_X1 U11131 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U11132 ( .A1(n8986), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U11133 ( .A1(n8985), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8845) );
  OAI211_X1 U11134 ( .C1(n8580), .C2(n8847), .A(n8846), .B(n8845), .ZN(n8848)
         );
  INV_X1 U11135 ( .A(n8848), .ZN(n8849) );
  NAND2_X1 U11136 ( .A1(n8850), .A2(n8849), .ZN(n13179) );
  NAND2_X1 U11137 ( .A1(n11509), .A2(n6490), .ZN(n8852) );
  INV_X1 U11138 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11510) );
  OR2_X1 U11139 ( .A1(n8990), .A2(n11510), .ZN(n8851) );
  MUX2_X1 U11140 ( .A(n13179), .B(n13346), .S(n8996), .Z(n8854) );
  MUX2_X1 U11141 ( .A(n13179), .B(n13346), .S(n8490), .Z(n8853) );
  NAND2_X1 U11142 ( .A1(n6479), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8861) );
  INV_X1 U11143 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13330) );
  OR2_X1 U11144 ( .A1(n8966), .A2(n13330), .ZN(n8860) );
  INV_X1 U11145 ( .A(n8874), .ZN(n8876) );
  OAI21_X1 U11146 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n8856), .A(n8876), .ZN(
        n13326) );
  OR2_X1 U11147 ( .A1(n6476), .A2(n13326), .ZN(n8859) );
  INV_X1 U11148 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8857) );
  OR2_X1 U11149 ( .A1(n8526), .A2(n8857), .ZN(n8858) );
  NAND4_X1 U11150 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(n13178) );
  XNOR2_X1 U11151 ( .A(n8863), .B(n8862), .ZN(n11563) );
  NAND2_X1 U11152 ( .A1(n11563), .A2(n6489), .ZN(n8865) );
  INV_X1 U11153 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11565) );
  OR2_X1 U11154 ( .A1(n8990), .A2(n11565), .ZN(n8864) );
  MUX2_X1 U11155 ( .A(n13178), .B(n13474), .S(n8490), .Z(n8869) );
  NAND2_X1 U11156 ( .A1(n8868), .A2(n8869), .ZN(n8867) );
  MUX2_X1 U11157 ( .A(n13178), .B(n13474), .S(n6512), .Z(n8866) );
  NAND2_X1 U11158 ( .A1(n8867), .A2(n8866), .ZN(n8873) );
  INV_X1 U11159 ( .A(n8868), .ZN(n8871) );
  INV_X1 U11160 ( .A(n8869), .ZN(n8870) );
  NAND2_X1 U11161 ( .A1(n8871), .A2(n8870), .ZN(n8872) );
  NAND2_X1 U11162 ( .A1(n6479), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8883) );
  INV_X1 U11163 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13309) );
  OR2_X1 U11164 ( .A1(n8966), .A2(n13309), .ZN(n8882) );
  INV_X1 U11165 ( .A(n8889), .ZN(n8878) );
  INV_X1 U11166 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11167 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  NAND2_X1 U11168 ( .A1(n8878), .A2(n8877), .ZN(n13308) );
  OR2_X1 U11169 ( .A1(n6476), .A2(n13308), .ZN(n8881) );
  INV_X1 U11170 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8879) );
  OR2_X1 U11171 ( .A1(n8526), .A2(n8879), .ZN(n8880) );
  NAND4_X1 U11172 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n13177) );
  NAND2_X1 U11173 ( .A1(n11625), .A2(n6489), .ZN(n8885) );
  OR2_X1 U11174 ( .A1(n8990), .A2(n11628), .ZN(n8884) );
  MUX2_X1 U11175 ( .A(n13177), .B(n13468), .S(n8996), .Z(n8887) );
  MUX2_X1 U11176 ( .A(n13177), .B(n13468), .S(n8490), .Z(n8886) );
  INV_X1 U11177 ( .A(n8887), .ZN(n8888) );
  NAND2_X1 U11178 ( .A1(n6478), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8894) );
  INV_X1 U11179 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13299) );
  OR2_X1 U11180 ( .A1(n8966), .A2(n13299), .ZN(n8893) );
  OAI21_X1 U11181 ( .B1(n8889), .B2(P2_REG3_REG_24__SCAN_IN), .A(n8907), .ZN(
        n13298) );
  OR2_X1 U11182 ( .A1(n6476), .A2(n13298), .ZN(n8892) );
  INV_X1 U11183 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8890) );
  OR2_X1 U11184 ( .A1(n8526), .A2(n8890), .ZN(n8891) );
  NAND4_X1 U11185 ( .A1(n8894), .A2(n8893), .A3(n8892), .A4(n8891), .ZN(n13176) );
  NAND2_X1 U11186 ( .A1(n11777), .A2(n6490), .ZN(n8896) );
  INV_X1 U11187 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11839) );
  OR2_X1 U11188 ( .A1(n8990), .A2(n11839), .ZN(n8895) );
  MUX2_X1 U11189 ( .A(n13176), .B(n13462), .S(n8490), .Z(n8900) );
  NAND2_X1 U11190 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  MUX2_X1 U11191 ( .A(n13176), .B(n13462), .S(n6512), .Z(n8897) );
  NAND2_X1 U11192 ( .A1(n8898), .A2(n8897), .ZN(n8904) );
  INV_X1 U11193 ( .A(n8899), .ZN(n8902) );
  INV_X1 U11194 ( .A(n8900), .ZN(n8901) );
  NAND2_X1 U11195 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  NAND2_X1 U11196 ( .A1(n6478), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8914) );
  INV_X1 U11197 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8905) );
  OR2_X1 U11198 ( .A1(n8966), .A2(n8905), .ZN(n8913) );
  INV_X1 U11199 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U11200 ( .A1(n8907), .A2(n8906), .ZN(n8909) );
  INV_X1 U11201 ( .A(n8919), .ZN(n8908) );
  NAND2_X1 U11202 ( .A1(n8909), .A2(n8908), .ZN(n13284) );
  OR2_X1 U11203 ( .A1(n6476), .A2(n13284), .ZN(n8912) );
  INV_X1 U11204 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8910) );
  OR2_X1 U11205 ( .A1(n8526), .A2(n8910), .ZN(n8911) );
  NAND4_X1 U11206 ( .A1(n8914), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n13175) );
  OR2_X1 U11207 ( .A1(n8990), .A2(n11882), .ZN(n8915) );
  MUX2_X1 U11208 ( .A(n13175), .B(n13457), .S(n6512), .Z(n8917) );
  MUX2_X1 U11209 ( .A(n13175), .B(n13457), .S(n8490), .Z(n8916) );
  INV_X1 U11210 ( .A(n8917), .ZN(n8918) );
  NAND2_X1 U11211 ( .A1(n6478), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8924) );
  INV_X1 U11212 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13269) );
  OR2_X1 U11213 ( .A1(n8966), .A2(n13269), .ZN(n8923) );
  NAND2_X1 U11214 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8919), .ZN(n8938) );
  OAI21_X1 U11215 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n8919), .A(n8938), .ZN(
        n13271) );
  OR2_X1 U11216 ( .A1(n6476), .A2(n13271), .ZN(n8922) );
  INV_X1 U11217 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8920) );
  OR2_X1 U11218 ( .A1(n8526), .A2(n8920), .ZN(n8921) );
  NAND4_X1 U11219 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n13174) );
  NAND2_X1 U11220 ( .A1(n13579), .A2(n6489), .ZN(n8926) );
  OR2_X1 U11221 ( .A1(n8990), .A2(n13580), .ZN(n8925) );
  MUX2_X1 U11222 ( .A(n13174), .B(n13274), .S(n8490), .Z(n8930) );
  NAND2_X1 U11223 ( .A1(n8929), .A2(n8930), .ZN(n8928) );
  MUX2_X1 U11224 ( .A(n13174), .B(n13274), .S(n6512), .Z(n8927) );
  NAND2_X1 U11225 ( .A1(n8928), .A2(n8927), .ZN(n8934) );
  INV_X1 U11226 ( .A(n8929), .ZN(n8932) );
  INV_X1 U11227 ( .A(n8930), .ZN(n8931) );
  NAND2_X1 U11228 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NAND2_X1 U11229 ( .A1(n8934), .A2(n8933), .ZN(n8949) );
  NAND2_X1 U11230 ( .A1(n6479), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8944) );
  INV_X1 U11231 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13259) );
  OR2_X1 U11232 ( .A1(n8966), .A2(n13259), .ZN(n8943) );
  INV_X1 U11233 ( .A(n8938), .ZN(n8936) );
  NAND2_X1 U11234 ( .A1(n8936), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8953) );
  INV_X1 U11235 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11236 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U11237 ( .A1(n8953), .A2(n8939), .ZN(n13258) );
  OR2_X1 U11238 ( .A1(n6476), .A2(n13258), .ZN(n8942) );
  INV_X1 U11239 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8940) );
  OR2_X1 U11240 ( .A1(n8526), .A2(n8940), .ZN(n8941) );
  NAND4_X1 U11241 ( .A1(n8944), .A2(n8943), .A3(n8942), .A4(n8941), .ZN(n13173) );
  NAND2_X1 U11242 ( .A1(n13575), .A2(n6490), .ZN(n8946) );
  OR2_X1 U11243 ( .A1(n8990), .A2(n13577), .ZN(n8945) );
  MUX2_X1 U11244 ( .A(n13173), .B(n13442), .S(n6512), .Z(n8948) );
  INV_X1 U11245 ( .A(n13173), .ZN(n13162) );
  INV_X1 U11246 ( .A(n13442), .ZN(n11970) );
  MUX2_X1 U11247 ( .A(n13162), .B(n11970), .S(n8490), .Z(n8947) );
  NAND2_X1 U11248 ( .A1(n8985), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8959) );
  INV_X1 U11249 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8950) );
  OR2_X1 U11250 ( .A1(n8580), .A2(n8950), .ZN(n8958) );
  INV_X1 U11251 ( .A(n8953), .ZN(n8951) );
  NAND2_X1 U11252 ( .A1(n8951), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11942) );
  INV_X1 U11253 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U11254 ( .A1(n8953), .A2(n8952), .ZN(n8954) );
  NAND2_X1 U11255 ( .A1(n11942), .A2(n8954), .ZN(n13247) );
  OR2_X1 U11256 ( .A1(n6476), .A2(n13247), .ZN(n8957) );
  INV_X1 U11257 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8955) );
  OR2_X1 U11258 ( .A1(n8526), .A2(n8955), .ZN(n8956) );
  INV_X1 U11259 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9589) );
  OR2_X1 U11260 ( .A1(n8990), .A2(n9589), .ZN(n8960) );
  MUX2_X1 U11261 ( .A(n13061), .B(n13240), .S(n6512), .Z(n8980) );
  MUX2_X1 U11262 ( .A(n13172), .B(n13436), .S(n8490), .Z(n8979) );
  NAND2_X1 U11263 ( .A1(n13565), .A2(n6490), .ZN(n8963) );
  INV_X1 U11264 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8961) );
  OR2_X1 U11265 ( .A1(n8990), .A2(n8961), .ZN(n8962) );
  INV_X1 U11266 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U11267 ( .A1(n8526), .A2(n8964), .ZN(n8970) );
  INV_X1 U11268 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8965) );
  NOR2_X1 U11269 ( .A1(n8966), .A2(n8965), .ZN(n8969) );
  INV_X1 U11270 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8967) );
  NOR2_X1 U11271 ( .A1(n8580), .A2(n8967), .ZN(n8968) );
  OR3_X1 U11272 ( .A1(n8970), .A2(n8969), .A3(n8968), .ZN(n13226) );
  XNOR2_X1 U11273 ( .A(n13227), .B(n13226), .ZN(n9035) );
  NAND2_X1 U11274 ( .A1(n8985), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8977) );
  INV_X1 U11275 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8971) );
  OR2_X1 U11276 ( .A1(n8526), .A2(n8971), .ZN(n8976) );
  OR2_X1 U11277 ( .A1(n6476), .A2(n11942), .ZN(n8975) );
  INV_X1 U11278 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8973) );
  OR2_X1 U11279 ( .A1(n8580), .A2(n8973), .ZN(n8974) );
  INV_X1 U11280 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13570) );
  NOR2_X1 U11281 ( .A1(n8990), .A2(n13570), .ZN(n8978) );
  MUX2_X1 U11282 ( .A(n12218), .B(n11945), .S(n6512), .Z(n8998) );
  INV_X1 U11283 ( .A(n12218), .ZN(n13171) );
  MUX2_X1 U11284 ( .A(n13171), .B(n13432), .S(n8490), .Z(n8997) );
  AOI22_X1 U11285 ( .A1(n8998), .A2(n8997), .B1(n8980), .B2(n8979), .ZN(n8981)
         );
  INV_X1 U11286 ( .A(n13226), .ZN(n9004) );
  NAND2_X1 U11287 ( .A1(n13227), .A2(n9004), .ZN(n8984) );
  OR2_X1 U11288 ( .A1(n13227), .A2(n9004), .ZN(n8983) );
  MUX2_X1 U11289 ( .A(n8984), .B(n8983), .S(n8490), .Z(n9000) );
  INV_X1 U11290 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11291 ( .A1(n8985), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11292 ( .A1(n8986), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8987) );
  OAI211_X1 U11293 ( .C1(n8580), .C2(n8989), .A(n8988), .B(n8987), .ZN(n13170)
         );
  NAND2_X1 U11294 ( .A1(n12273), .A2(n6489), .ZN(n8992) );
  INV_X1 U11295 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12533) );
  OR2_X1 U11296 ( .A1(n8990), .A2(n12533), .ZN(n8991) );
  MUX2_X1 U11297 ( .A(n13170), .B(n9033), .S(n8490), .Z(n9003) );
  NAND2_X1 U11298 ( .A1(n13226), .A2(n8490), .ZN(n8993) );
  OR2_X1 U11299 ( .A1(n10828), .A2(n8487), .ZN(n9012) );
  NAND4_X1 U11300 ( .A1(n8993), .A2(n10181), .A3(n9012), .A4(n10232), .ZN(
        n8994) );
  AND2_X1 U11301 ( .A1(n8994), .A2(n13170), .ZN(n8995) );
  AOI21_X1 U11302 ( .B1(n9033), .B2(n8996), .A(n8995), .ZN(n9002) );
  OAI22_X1 U11303 ( .A1(n9003), .A2(n9002), .B1(n8998), .B2(n8997), .ZN(n8999)
         );
  NAND2_X1 U11304 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  NAND2_X1 U11305 ( .A1(n9003), .A2(n9002), .ZN(n9008) );
  NAND3_X1 U11306 ( .A1(n13227), .A2(n9004), .A3(n8490), .ZN(n9006) );
  OR3_X1 U11307 ( .A1(n13227), .A2(n9004), .A3(n8490), .ZN(n9005) );
  NAND2_X1 U11308 ( .A1(n9006), .A2(n9005), .ZN(n9007) );
  INV_X1 U11309 ( .A(n9038), .ZN(n9016) );
  NAND2_X1 U11310 ( .A1(n13217), .A2(n10181), .ZN(n9010) );
  OAI211_X1 U11311 ( .C1(n10205), .C2(n10244), .A(n10232), .B(n9010), .ZN(
        n9011) );
  INV_X1 U11312 ( .A(n9011), .ZN(n9015) );
  INV_X1 U11313 ( .A(n6472), .ZN(n9022) );
  NAND2_X1 U11314 ( .A1(n9022), .A2(n10181), .ZN(n10206) );
  OAI21_X1 U11315 ( .B1(n10206), .B2(n13217), .A(n9012), .ZN(n9013) );
  NAND2_X1 U11316 ( .A1(n9016), .A2(n9013), .ZN(n9014) );
  OAI21_X1 U11317 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9045) );
  INV_X1 U11318 ( .A(n10828), .ZN(n9037) );
  NAND2_X1 U11319 ( .A1(n13436), .A2(n13172), .ZN(n11940) );
  OR2_X1 U11320 ( .A1(n13436), .A2(n13172), .ZN(n9017) );
  INV_X1 U11321 ( .A(n13175), .ZN(n13164) );
  OR2_X1 U11322 ( .A1(n13274), .A2(n13093), .ZN(n11969) );
  NAND2_X1 U11323 ( .A1(n13274), .A2(n13093), .ZN(n11967) );
  XOR2_X1 U11324 ( .A(n13179), .B(n13346), .Z(n13338) );
  INV_X1 U11325 ( .A(n13178), .ZN(n11963) );
  XNOR2_X1 U11326 ( .A(n13474), .B(n11963), .ZN(n13332) );
  INV_X1 U11327 ( .A(n13180), .ZN(n13077) );
  XNOR2_X1 U11328 ( .A(n12181), .B(n13077), .ZN(n11957) );
  XNOR2_X1 U11329 ( .A(n13498), .B(n13181), .ZN(n13363) );
  XOR2_X1 U11330 ( .A(n13186), .B(n14239), .Z(n11659) );
  INV_X1 U11331 ( .A(n13183), .ZN(n13153) );
  XNOR2_X1 U11332 ( .A(n13400), .B(n13153), .ZN(n13393) );
  XNOR2_X1 U11333 ( .A(n11649), .B(n13187), .ZN(n11521) );
  INV_X1 U11334 ( .A(n13190), .ZN(n11282) );
  XNOR2_X1 U11335 ( .A(n14736), .B(n11282), .ZN(n11494) );
  INV_X1 U11336 ( .A(n13191), .ZN(n11281) );
  XNOR2_X1 U11337 ( .A(n14727), .B(n11281), .ZN(n11333) );
  INV_X1 U11338 ( .A(n13192), .ZN(n11278) );
  XNOR2_X1 U11339 ( .A(n11484), .B(n11278), .ZN(n11477) );
  XNOR2_X1 U11340 ( .A(n14714), .B(n13193), .ZN(n11455) );
  XNOR2_X1 U11341 ( .A(n11044), .B(n13197), .ZN(n10663) );
  INV_X1 U11342 ( .A(n13195), .ZN(n9018) );
  NAND2_X1 U11343 ( .A1(n11052), .A2(n9018), .ZN(n11057) );
  OR2_X1 U11344 ( .A1(n11052), .A2(n9018), .ZN(n9019) );
  NAND2_X1 U11345 ( .A1(n11057), .A2(n9019), .ZN(n10704) );
  NAND2_X1 U11346 ( .A1(n9020), .A2(n10241), .ZN(n10199) );
  OR2_X1 U11347 ( .A1(n9020), .A2(n10241), .ZN(n9021) );
  NAND2_X1 U11348 ( .A1(n10199), .A2(n9021), .ZN(n14687) );
  NAND2_X1 U11349 ( .A1(n13198), .A2(n14693), .ZN(n9023) );
  NOR4_X1 U11350 ( .A1(n10663), .A2(n10704), .A3(n9024), .A4(n11348), .ZN(
        n9025) );
  XNOR2_X1 U11351 ( .A(n14706), .B(n13194), .ZN(n11059) );
  XNOR2_X1 U11352 ( .A(n10994), .B(n13196), .ZN(n10986) );
  NAND4_X1 U11353 ( .A1(n11455), .A2(n9025), .A3(n11059), .A4(n10986), .ZN(
        n9026) );
  NOR4_X1 U11354 ( .A1(n11494), .A2(n11333), .A3(n11477), .A4(n9026), .ZN(
        n9027) );
  XNOR2_X1 U11355 ( .A(n11520), .B(n13188), .ZN(n11304) );
  XNOR2_X1 U11356 ( .A(n11302), .B(n13189), .ZN(n11300) );
  NAND4_X1 U11357 ( .A1(n11521), .A2(n9027), .A3(n11304), .A4(n11300), .ZN(
        n9028) );
  NOR4_X1 U11358 ( .A1(n11659), .A2(n13393), .A3(n11949), .A4(n9028), .ZN(
        n9029) );
  XNOR2_X1 U11359 ( .A(n13503), .B(n13182), .ZN(n13387) );
  NAND4_X1 U11360 ( .A1(n13363), .A2(n9029), .A3(n13387), .A4(n11742), .ZN(
        n9030) );
  NOR4_X1 U11361 ( .A1(n13338), .A2(n13332), .A3(n11957), .A4(n9030), .ZN(
        n9031) );
  XNOR2_X1 U11362 ( .A(n13468), .B(n13177), .ZN(n13314) );
  XNOR2_X1 U11363 ( .A(n13462), .B(n13176), .ZN(n13292) );
  NAND4_X1 U11364 ( .A1(n13266), .A2(n9031), .A3(n13314), .A4(n13292), .ZN(
        n9032) );
  XOR2_X1 U11365 ( .A(n13170), .B(n13430), .Z(n9034) );
  XNOR2_X1 U11366 ( .A(n13432), .B(n13171), .ZN(n11971) );
  AOI211_X1 U11367 ( .C1(n9038), .C2(n9037), .A(n10181), .B(n9036), .ZN(n9044)
         );
  NAND2_X1 U11368 ( .A1(n9040), .A2(n9039), .ZN(n9042) );
  NAND2_X1 U11369 ( .A1(n9042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U11370 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9041), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n9043) );
  NOR2_X1 U11371 ( .A1(n9768), .A2(P2_U3088), .ZN(n9062) );
  OAI21_X1 U11372 ( .B1(n9045), .B2(n9044), .A(n9062), .ZN(n9066) );
  NAND2_X1 U11373 ( .A1(n9046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9047) );
  MUX2_X1 U11374 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9047), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9049) );
  INV_X1 U11375 ( .A(n11837), .ZN(n9060) );
  NAND2_X1 U11376 ( .A1(n9051), .A2(n9050), .ZN(n9057) );
  NAND2_X1 U11377 ( .A1(n9057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9052) );
  MUX2_X1 U11378 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9052), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9054) );
  NAND2_X1 U11379 ( .A1(n9054), .A2(n9053), .ZN(n13582) );
  NAND2_X1 U11380 ( .A1(n9055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9056) );
  MUX2_X1 U11381 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9056), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9058) );
  NOR2_X1 U11382 ( .A1(n13582), .A2(n11881), .ZN(n9059) );
  NAND2_X1 U11383 ( .A1(n9060), .A2(n9059), .ZN(n9706) );
  INV_X1 U11384 ( .A(n10209), .ZN(n9061) );
  NAND2_X1 U11385 ( .A1(n9061), .A2(n10228), .ZN(n13163) );
  NOR4_X1 U11386 ( .A1(n14683), .A2(n10232), .A3(n13576), .A4(n13163), .ZN(
        n9064) );
  INV_X1 U11387 ( .A(n9062), .ZN(n11626) );
  OAI21_X1 U11388 ( .B1(n11626), .B2(n10205), .A(P2_B_REG_SCAN_IN), .ZN(n9063)
         );
  OR2_X1 U11389 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U11390 ( .A1(n9066), .A2(n9065), .ZN(P2_U3328) );
  NAND3_X1 U11391 ( .A1(n9070), .A2(n9256), .A3(n9069), .ZN(n9071) );
  INV_X1 U11392 ( .A(n9084), .ZN(n9081) );
  NAND2_X1 U11393 ( .A1(n9081), .A2(n9080), .ZN(n13050) );
  XNOR2_X2 U11394 ( .A(n9083), .B(n9082), .ZN(n9090) );
  AND2_X4 U11395 ( .A1(n9090), .A2(n9088), .ZN(n12538) );
  NAND2_X1 U11396 ( .A1(n12538), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U11397 ( .A1(n9086), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9093) );
  INV_X1 U11398 ( .A(n9090), .ZN(n9087) );
  INV_X1 U11399 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10020) );
  OR2_X1 U11400 ( .A1(n9139), .A2(n10020), .ZN(n9092) );
  OR2_X2 U11401 ( .A1(n9157), .A2(n7577), .ZN(n9091) );
  XNOR2_X2 U11402 ( .A(n9097), .B(n9096), .ZN(n11925) );
  OR2_X1 U11403 ( .A1(n9099), .A2(n9098), .ZN(n9101) );
  XNOR2_X2 U11404 ( .A(n9101), .B(n9100), .ZN(n9616) );
  INV_X1 U11405 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9102) );
  OR2_X1 U11406 ( .A1(n9561), .A2(n9754), .ZN(n9106) );
  INV_X1 U11407 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U11408 ( .A1(n9104), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9125) );
  XNOR2_X1 U11409 ( .A(n9127), .B(n9125), .ZN(n9753) );
  OR2_X1 U11410 ( .A1(n9113), .A2(n9753), .ZN(n9105) );
  OAI211_X1 U11411 ( .C1(n9103), .C2(n10028), .A(n9106), .B(n9105), .ZN(n9107)
         );
  INV_X1 U11412 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U11413 ( .A1(n9086), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11414 ( .A1(n9312), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9109) );
  INV_X1 U11415 ( .A(n14772), .ZN(n14776) );
  OR2_X1 U11416 ( .A1(n6480), .A2(n7628), .ZN(n9117) );
  INV_X1 U11417 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11418 ( .A1(n9114), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9115) );
  AND2_X1 U11419 ( .A1(n9125), .A2(n9115), .ZN(n9711) );
  OR2_X1 U11420 ( .A1(n9475), .A2(n9711), .ZN(n9116) );
  OAI211_X1 U11421 ( .C1(n14776), .C2(n9103), .A(n9117), .B(n9116), .ZN(n15014) );
  NAND2_X1 U11422 ( .A1(n10119), .A2(n14995), .ZN(n9120) );
  NAND2_X1 U11423 ( .A1(n9118), .A2(n14992), .ZN(n9119) );
  NAND2_X1 U11424 ( .A1(n9120), .A2(n9119), .ZN(n14981) );
  NAND2_X1 U11425 ( .A1(n12538), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9124) );
  INV_X1 U11426 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10046) );
  OR2_X1 U11427 ( .A1(n9139), .A2(n10046), .ZN(n9121) );
  OR2_X1 U11428 ( .A1(n6480), .A2(SI_2_), .ZN(n9135) );
  INV_X1 U11429 ( .A(n9125), .ZN(n9126) );
  NAND2_X1 U11430 ( .A1(n9127), .A2(n9126), .ZN(n9129) );
  NAND2_X1 U11431 ( .A1(n9734), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9128) );
  NAND2_X1 U11432 ( .A1(n9752), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9146) );
  INV_X1 U11433 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U11434 ( .A1(n9730), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U11435 ( .A(n9145), .B(n9144), .ZN(n9715) );
  OR2_X1 U11436 ( .A1(n9475), .A2(n9715), .ZN(n9134) );
  OR2_X1 U11437 ( .A1(n9103), .A2(n10056), .ZN(n9133) );
  NAND2_X1 U11438 ( .A1(n14997), .A2(n10093), .ZN(n12399) );
  INV_X1 U11439 ( .A(n14997), .ZN(n14964) );
  INV_X1 U11440 ( .A(n10093), .ZN(n14977) );
  NAND2_X1 U11441 ( .A1(n14964), .A2(n14977), .ZN(n12391) );
  NAND2_X1 U11442 ( .A1(n14981), .A2(n12392), .ZN(n9137) );
  NAND2_X1 U11443 ( .A1(n14997), .A2(n14977), .ZN(n9136) );
  NAND2_X1 U11444 ( .A1(n12538), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9143) );
  OR2_X1 U11445 ( .A1(n9157), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9142) );
  INV_X1 U11446 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9138) );
  OR2_X1 U11447 ( .A1(n9387), .A2(n9138), .ZN(n9141) );
  INV_X1 U11448 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11167) );
  OR2_X1 U11449 ( .A1(n9139), .A2(n11167), .ZN(n9140) );
  OR2_X1 U11450 ( .A1(n6481), .A2(SI_3_), .ZN(n9152) );
  NAND2_X1 U11451 ( .A1(n9748), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9165) );
  INV_X1 U11452 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9739) );
  NAND2_X1 U11453 ( .A1(n9739), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9147) );
  XNOR2_X1 U11454 ( .A(n9164), .B(n9163), .ZN(n9721) );
  OR2_X1 U11455 ( .A1(n9475), .A2(n9721), .ZN(n9151) );
  OR2_X1 U11456 ( .A1(n9148), .A2(n9098), .ZN(n9149) );
  XNOR2_X1 U11457 ( .A(n9149), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11168) );
  OR2_X1 U11458 ( .A1(n9103), .A2(n11168), .ZN(n9150) );
  INV_X1 U11459 ( .A(n14970), .ZN(n9153) );
  NAND2_X1 U11460 ( .A1(n12611), .A2(n9153), .ZN(n12404) );
  NAND2_X1 U11461 ( .A1(n14983), .A2(n14970), .ZN(n12400) );
  AND2_X1 U11462 ( .A1(n12404), .A2(n12400), .ZN(n14960) );
  INV_X1 U11463 ( .A(n14960), .ZN(n9154) );
  NAND2_X1 U11464 ( .A1(n12611), .A2(n14970), .ZN(n9155) );
  NAND2_X1 U11465 ( .A1(n9156), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9162) );
  INV_X1 U11466 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11174) );
  OR2_X1 U11467 ( .A1(n12540), .A2(n11174), .ZN(n9161) );
  INV_X1 U11468 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11173) );
  AND2_X1 U11469 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9158) );
  NOR2_X1 U11470 ( .A1(n9175), .A2(n9158), .ZN(n10920) );
  OR2_X1 U11471 ( .A1(n9157), .A2(n10920), .ZN(n9159) );
  OR2_X1 U11472 ( .A1(n6481), .A2(SI_4_), .ZN(n9172) );
  NAND2_X1 U11473 ( .A1(n9750), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9184) );
  INV_X1 U11474 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U11475 ( .A1(n9742), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9166) );
  XNOR2_X1 U11476 ( .A(n9183), .B(n9182), .ZN(n9712) );
  OR2_X1 U11477 ( .A1(n9475), .A2(n9712), .ZN(n9171) );
  NAND2_X1 U11478 ( .A1(n9148), .A2(n9167), .ZN(n9187) );
  NAND2_X1 U11479 ( .A1(n9187), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9169) );
  INV_X1 U11480 ( .A(n14807), .ZN(n11175) );
  OR2_X1 U11481 ( .A1(n9103), .A2(n11175), .ZN(n9170) );
  NAND2_X1 U11482 ( .A1(n10794), .A2(n10919), .ZN(n12409) );
  INV_X1 U11483 ( .A(n10919), .ZN(n9173) );
  NAND2_X1 U11484 ( .A1(n14963), .A2(n9173), .ZN(n12412) );
  NAND2_X1 U11485 ( .A1(n12409), .A2(n12412), .ZN(n12406) );
  NAND2_X1 U11486 ( .A1(n14963), .A2(n10919), .ZN(n9174) );
  NAND2_X1 U11487 ( .A1(n9156), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9181) );
  INV_X1 U11488 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11180) );
  OR2_X1 U11489 ( .A1(n12540), .A2(n11180), .ZN(n9180) );
  INV_X1 U11490 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11179) );
  OR2_X1 U11491 ( .A1(n9369), .A2(n11179), .ZN(n9179) );
  INV_X1 U11492 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11493 ( .A1(n9175), .A2(n9176), .ZN(n9194) );
  OR2_X1 U11494 ( .A1(n9176), .A2(n9175), .ZN(n9177) );
  AND2_X1 U11495 ( .A1(n9194), .A2(n9177), .ZN(n10799) );
  OR2_X1 U11496 ( .A1(n9157), .A2(n10799), .ZN(n9178) );
  AND4_X2 U11497 ( .A1(n9181), .A2(n9180), .A3(n9179), .A4(n9178), .ZN(n10690)
         );
  NAND2_X1 U11498 ( .A1(n9185), .A2(n9184), .ZN(n9204) );
  NAND2_X1 U11499 ( .A1(n9758), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11500 ( .A1(n9756), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9186) );
  XNOR2_X1 U11501 ( .A(n9204), .B(n9203), .ZN(n9718) );
  OR2_X1 U11502 ( .A1(n9475), .A2(n9718), .ZN(n9191) );
  OR2_X1 U11503 ( .A1(n6481), .A2(SI_5_), .ZN(n9190) );
  NOR2_X1 U11504 ( .A1(n9187), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9201) );
  OR2_X1 U11505 ( .A1(n9201), .A2(n9098), .ZN(n9188) );
  XNOR2_X1 U11506 ( .A(n9188), .B(n9200), .ZN(n14824) );
  INV_X1 U11507 ( .A(n14824), .ZN(n11181) );
  OR2_X1 U11508 ( .A1(n9103), .A2(n11181), .ZN(n9189) );
  NAND2_X1 U11509 ( .A1(n10690), .A2(n10511), .ZN(n12414) );
  INV_X1 U11510 ( .A(n10511), .ZN(n10798) );
  NAND2_X1 U11511 ( .A1(n12610), .A2(n10798), .ZN(n12410) );
  INV_X1 U11512 ( .A(n12565), .ZN(n9192) );
  NAND2_X1 U11513 ( .A1(n10690), .A2(n10798), .ZN(n9193) );
  NAND2_X1 U11514 ( .A1(n9156), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9199) );
  INV_X1 U11515 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11187) );
  OR2_X1 U11516 ( .A1(n12540), .A2(n11187), .ZN(n9198) );
  INV_X1 U11517 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11186) );
  OR2_X1 U11518 ( .A1(n9369), .A2(n11186), .ZN(n9197) );
  NAND2_X1 U11519 ( .A1(n9194), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9195) );
  AND2_X1 U11520 ( .A1(n9211), .A2(n9195), .ZN(n10931) );
  OR2_X1 U11521 ( .A1(n9157), .A2(n10931), .ZN(n9196) );
  NAND2_X1 U11522 ( .A1(n9201), .A2(n9200), .ZN(n9217) );
  NAND2_X1 U11523 ( .A1(n9217), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U11524 ( .A(n9202), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U11525 ( .A1(n9204), .A2(n9203), .ZN(n9206) );
  NAND2_X1 U11526 ( .A1(n9206), .A2(n9205), .ZN(n9221) );
  XNOR2_X1 U11527 ( .A(n9765), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9207) );
  XNOR2_X1 U11528 ( .A(n9221), .B(n9207), .ZN(n9710) );
  OR2_X1 U11529 ( .A1(n9475), .A2(n9710), .ZN(n9209) );
  INV_X1 U11530 ( .A(SI_6_), .ZN(n9709) );
  OR2_X1 U11531 ( .A1(n6480), .A2(n9709), .ZN(n9208) );
  OAI211_X1 U11532 ( .C1(n9103), .C2(n14842), .A(n9209), .B(n9208), .ZN(n10930) );
  NAND2_X1 U11533 ( .A1(n10838), .A2(n10930), .ZN(n12422) );
  INV_X1 U11534 ( .A(n10838), .ZN(n14949) );
  INV_X1 U11535 ( .A(n10930), .ZN(n10685) );
  NAND2_X1 U11536 ( .A1(n14949), .A2(n10685), .ZN(n12415) );
  NAND2_X1 U11537 ( .A1(n12422), .A2(n12415), .ZN(n10933) );
  NAND2_X1 U11538 ( .A1(n14949), .A2(n10930), .ZN(n9210) );
  NAND2_X1 U11539 ( .A1(n10932), .A2(n9210), .ZN(n14948) );
  INV_X1 U11540 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11192) );
  OR2_X1 U11541 ( .A1(n9369), .A2(n11192), .ZN(n9216) );
  AND2_X1 U11542 ( .A1(n9211), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9212) );
  NOR2_X1 U11543 ( .A1(n9231), .A2(n9212), .ZN(n14955) );
  OR2_X1 U11544 ( .A1(n9157), .A2(n14955), .ZN(n9215) );
  NAND2_X1 U11545 ( .A1(n9610), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9214) );
  NAND2_X1 U11546 ( .A1(n9156), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9213) );
  NAND4_X1 U11547 ( .A1(n9216), .A2(n9215), .A3(n9214), .A4(n9213), .ZN(n12609) );
  OAI21_X1 U11548 ( .B1(n9217), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9219) );
  INV_X1 U11549 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9218) );
  XNOR2_X1 U11550 ( .A(n9219), .B(n9218), .ZN(n14859) );
  OR2_X1 U11551 ( .A1(n6480), .A2(SI_7_), .ZN(n9229) );
  NAND2_X1 U11552 ( .A1(n9763), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11553 ( .A1(n9221), .A2(n9220), .ZN(n9223) );
  NAND2_X1 U11554 ( .A1(n9765), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11555 ( .A1(n9797), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U11556 ( .A1(n9795), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11557 ( .A1(n9237), .A2(n9224), .ZN(n9225) );
  NAND2_X1 U11558 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  AND2_X1 U11559 ( .A1(n9238), .A2(n9227), .ZN(n9724) );
  OR2_X1 U11560 ( .A1(n9475), .A2(n9724), .ZN(n9228) );
  OAI211_X1 U11561 ( .C1(n11193), .C2(n9103), .A(n9229), .B(n9228), .ZN(n14954) );
  XNOR2_X1 U11562 ( .A(n12609), .B(n14954), .ZN(n14947) );
  INV_X1 U11563 ( .A(n14954), .ZN(n10840) );
  NAND2_X1 U11564 ( .A1(n12609), .A2(n10840), .ZN(n9230) );
  NAND2_X1 U11565 ( .A1(n9156), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9236) );
  INV_X1 U11566 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11199) );
  OR2_X1 U11567 ( .A1(n12540), .A2(n11199), .ZN(n9235) );
  INV_X1 U11568 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11198) );
  OR2_X1 U11569 ( .A1(n9369), .A2(n11198), .ZN(n9234) );
  NOR2_X1 U11570 ( .A1(n9231), .A2(n12299), .ZN(n9232) );
  OR2_X1 U11571 ( .A1(n9262), .A2(n9232), .ZN(n12301) );
  INV_X1 U11572 ( .A(n12301), .ZN(n11094) );
  OR2_X1 U11573 ( .A1(n9157), .A2(n11094), .ZN(n9233) );
  INV_X1 U11574 ( .A(SI_8_), .ZN(n9743) );
  NAND2_X1 U11575 ( .A1(n9804), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U11576 ( .A1(n9802), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9239) );
  OR2_X1 U11577 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  NAND2_X1 U11578 ( .A1(n9251), .A2(n9242), .ZN(n9744) );
  OR2_X1 U11579 ( .A1(n9744), .A2(n9475), .ZN(n9247) );
  OR2_X1 U11580 ( .A1(n9244), .A2(n9098), .ZN(n9245) );
  XNOR2_X1 U11581 ( .A(n9245), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11200) );
  OR2_X1 U11582 ( .A1(n9103), .A2(n14876), .ZN(n9246) );
  OAI211_X1 U11583 ( .C1(n6481), .C2(n9743), .A(n9247), .B(n9246), .ZN(n12300)
         );
  NAND2_X1 U11584 ( .A1(n10946), .A2(n12300), .ZN(n12429) );
  INV_X1 U11585 ( .A(n12300), .ZN(n15048) );
  NAND2_X1 U11586 ( .A1(n14950), .A2(n15048), .ZN(n12428) );
  NAND2_X1 U11587 ( .A1(n10946), .A2(n15048), .ZN(n9249) );
  NAND2_X1 U11588 ( .A1(n9821), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11589 ( .A1(n9819), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9252) );
  OR2_X1 U11590 ( .A1(n9254), .A2(n9253), .ZN(n9255) );
  NAND2_X1 U11591 ( .A1(n9270), .A2(n9255), .ZN(n9732) );
  NAND2_X1 U11592 ( .A1(n9732), .A2(n12537), .ZN(n9261) );
  INV_X1 U11593 ( .A(SI_9_), .ZN(n9731) );
  NAND2_X1 U11594 ( .A1(n9244), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U11595 ( .A1(n9258), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9257) );
  MUX2_X1 U11596 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9257), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9259) );
  NAND2_X1 U11597 ( .A1(n9259), .A2(n9383), .ZN(n14895) );
  AOI22_X1 U11598 ( .A1(n9439), .A2(n9731), .B1(n10013), .B2(n14895), .ZN(
        n9260) );
  INV_X1 U11599 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11204) );
  OR2_X1 U11600 ( .A1(n9369), .A2(n11204), .ZN(n9267) );
  OR2_X1 U11601 ( .A1(n9262), .A2(n10952), .ZN(n9263) );
  AND2_X1 U11602 ( .A1(n9279), .A2(n9263), .ZN(n11250) );
  OR2_X1 U11603 ( .A1(n9157), .A2(n11250), .ZN(n9266) );
  NAND2_X1 U11604 ( .A1(n9610), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11605 ( .A1(n9086), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9264) );
  NAND4_X1 U11606 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(n14935) );
  NAND2_X1 U11607 ( .A1(n12432), .A2(n14935), .ZN(n12433) );
  INV_X1 U11608 ( .A(n14935), .ZN(n11072) );
  NAND2_X1 U11609 ( .A1(n11072), .A2(n11249), .ZN(n9268) );
  NAND2_X1 U11610 ( .A1(n9891), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11611 ( .A1(n9893), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9271) );
  OR2_X1 U11612 ( .A1(n9273), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U11613 ( .A1(n9294), .A2(n9274), .ZN(n9741) );
  NAND2_X1 U11614 ( .A1(n9741), .A2(n12537), .ZN(n9278) );
  NAND2_X1 U11615 ( .A1(n9383), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9276) );
  XNOR2_X1 U11616 ( .A(n9276), .B(n9275), .ZN(n11213) );
  AOI22_X1 U11617 ( .A1(n9439), .A2(n9740), .B1(n10013), .B2(n11213), .ZN(
        n9277) );
  NAND2_X1 U11618 ( .A1(n9278), .A2(n9277), .ZN(n14940) );
  INV_X1 U11619 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11211) );
  OR2_X1 U11620 ( .A1(n12540), .A2(n11211), .ZN(n9284) );
  INV_X1 U11621 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11210) );
  OR2_X1 U11622 ( .A1(n9369), .A2(n11210), .ZN(n9283) );
  NAND2_X1 U11623 ( .A1(n9279), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9280) );
  AND2_X1 U11624 ( .A1(n9286), .A2(n9280), .ZN(n11079) );
  OR2_X1 U11625 ( .A1(n9157), .A2(n11079), .ZN(n9282) );
  NAND2_X1 U11626 ( .A1(n9156), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9281) );
  NAND4_X1 U11627 ( .A1(n9284), .A2(n9283), .A3(n9282), .A4(n9281), .ZN(n12608) );
  OR2_X1 U11628 ( .A1(n14940), .A2(n12608), .ZN(n12437) );
  NAND2_X1 U11629 ( .A1(n14940), .A2(n12608), .ZN(n12438) );
  NAND2_X1 U11630 ( .A1(n12437), .A2(n12438), .ZN(n14933) );
  INV_X1 U11631 ( .A(n12608), .ZN(n14201) );
  OR2_X1 U11632 ( .A1(n14940), .A2(n14201), .ZN(n9285) );
  NAND2_X1 U11633 ( .A1(n9286), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9287) );
  AND2_X1 U11634 ( .A1(n9306), .A2(n9287), .ZN(n14203) );
  OR2_X1 U11635 ( .A1(n9157), .A2(n14203), .ZN(n9292) );
  INV_X1 U11636 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9288) );
  OR2_X1 U11637 ( .A1(n9369), .A2(n9288), .ZN(n9291) );
  NAND2_X1 U11638 ( .A1(n9156), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11639 ( .A1(n9610), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9289) );
  NAND4_X1 U11640 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n14936) );
  XNOR2_X1 U11641 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9295) );
  XNOR2_X1 U11642 ( .A(n9299), .B(n9295), .ZN(n9746) );
  NOR2_X1 U11643 ( .A1(n9383), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11644 ( .A1(n9301), .A2(n9098), .ZN(n9296) );
  XNOR2_X1 U11645 ( .A(n9296), .B(n9300), .ZN(n11435) );
  INV_X1 U11646 ( .A(n11435), .ZN(n11441) );
  OAI22_X1 U11647 ( .A1(n6481), .A2(SI_11_), .B1(n11441), .B2(n9103), .ZN(
        n9297) );
  AOI21_X1 U11648 ( .B1(n9746), .B2(n12537), .A(n9297), .ZN(n11261) );
  NAND2_X1 U11649 ( .A1(n9901), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9298) );
  XNOR2_X1 U11650 ( .A(n10221), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n9321) );
  XNOR2_X1 U11651 ( .A(n9323), .B(n9321), .ZN(n9759) );
  NAND2_X1 U11652 ( .A1(n9759), .A2(n12537), .ZN(n9304) );
  OR2_X1 U11653 ( .A1(n9328), .A2(n9098), .ZN(n9302) );
  XNOR2_X1 U11654 ( .A(n9302), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U11655 ( .A1(n9439), .A2(SI_12_), .B1(n10013), .B2(n11721), .ZN(
        n9303) );
  NAND2_X1 U11656 ( .A1(n9304), .A2(n9303), .ZN(n14221) );
  NAND2_X1 U11657 ( .A1(n9086), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9311) );
  INV_X1 U11658 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11773) );
  OR2_X1 U11659 ( .A1(n12540), .A2(n11773), .ZN(n9310) );
  INV_X1 U11660 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n9305) );
  OR2_X1 U11661 ( .A1(n9369), .A2(n9305), .ZN(n9309) );
  AND2_X1 U11662 ( .A1(n9306), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9307) );
  NOR2_X1 U11663 ( .A1(n9314), .A2(n9307), .ZN(n11772) );
  OR2_X1 U11664 ( .A1(n9157), .A2(n11772), .ZN(n9308) );
  OR2_X1 U11665 ( .A1(n14221), .A2(n14202), .ZN(n12447) );
  NAND2_X1 U11666 ( .A1(n14221), .A2(n14202), .ZN(n12448) );
  NAND2_X1 U11667 ( .A1(n12447), .A2(n12448), .ZN(n11769) );
  NAND2_X1 U11668 ( .A1(n14221), .A2(n12607), .ZN(n9332) );
  OR2_X1 U11669 ( .A1(n9314), .A2(n9313), .ZN(n9315) );
  NAND2_X1 U11670 ( .A1(n9314), .A2(n9313), .ZN(n9347) );
  AND2_X1 U11671 ( .A1(n9315), .A2(n9347), .ZN(n14189) );
  INV_X1 U11672 ( .A(n14189), .ZN(n11582) );
  NAND2_X1 U11673 ( .A1(n9594), .A2(n11582), .ZN(n9320) );
  INV_X1 U11674 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9316) );
  OR2_X1 U11675 ( .A1(n9369), .A2(n9316), .ZN(n9319) );
  NAND2_X1 U11676 ( .A1(n9156), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11677 ( .A1(n9610), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9317) );
  NAND4_X1 U11678 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(n12606) );
  INV_X1 U11679 ( .A(n9321), .ZN(n9322) );
  NAND2_X1 U11680 ( .A1(n9323), .A2(n9322), .ZN(n9326) );
  NAND2_X1 U11681 ( .A1(n9324), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9325) );
  XNOR2_X1 U11682 ( .A(n9335), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U11683 ( .A1(n9799), .A2(n12537), .ZN(n9331) );
  INV_X1 U11684 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9327) );
  AND2_X1 U11685 ( .A1(n9328), .A2(n9327), .ZN(n9342) );
  OR2_X1 U11686 ( .A1(n9342), .A2(n9098), .ZN(n9329) );
  INV_X1 U11687 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9341) );
  XNOR2_X1 U11688 ( .A(n9329), .B(n9341), .ZN(n12617) );
  AOI22_X1 U11689 ( .A1(n9439), .A2(n9798), .B1(n12617), .B2(n10013), .ZN(
        n9330) );
  AND2_X1 U11690 ( .A1(n9332), .A2(n7359), .ZN(n9333) );
  INV_X1 U11691 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11692 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  XNOR2_X1 U11693 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9340) );
  XNOR2_X1 U11694 ( .A(n9356), .B(n9340), .ZN(n9823) );
  NAND2_X1 U11695 ( .A1(n9823), .A2(n12537), .ZN(n9346) );
  NAND2_X1 U11696 ( .A1(n9342), .A2(n9341), .ZN(n9362) );
  NAND2_X1 U11697 ( .A1(n9362), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9344) );
  XNOR2_X1 U11698 ( .A(n9344), .B(n9343), .ZN(n12644) );
  AOI22_X1 U11699 ( .A1(n12644), .A2(n10013), .B1(n9439), .B2(n9822), .ZN(
        n9345) );
  NAND2_X1 U11700 ( .A1(n9610), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U11701 ( .A1(n12538), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11702 ( .A1(n9347), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U11703 ( .A1(n9367), .A2(n9348), .ZN(n11832) );
  NAND2_X1 U11704 ( .A1(n9594), .A2(n11832), .ZN(n9350) );
  NAND2_X1 U11705 ( .A1(n9156), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9349) );
  NAND4_X1 U11706 ( .A1(n9352), .A2(n9351), .A3(n9350), .A4(n9349), .ZN(n12605) );
  OR2_X1 U11707 ( .A1(n11912), .A2(n12605), .ZN(n12459) );
  NAND2_X1 U11708 ( .A1(n11912), .A2(n12605), .ZN(n12463) );
  INV_X1 U11709 ( .A(n12605), .ZN(n14188) );
  OR2_X1 U11710 ( .A1(n11912), .A2(n14188), .ZN(n9354) );
  NAND2_X1 U11711 ( .A1(n10616), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11712 ( .A1(n10682), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11713 ( .A1(n10680), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11714 ( .A1(n9376), .A2(n9358), .ZN(n9359) );
  NAND2_X1 U11715 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  NAND2_X1 U11716 ( .A1(n9377), .A2(n9361), .ZN(n9899) );
  OR2_X1 U11717 ( .A1(n9899), .A2(n9475), .ZN(n9366) );
  OAI21_X1 U11718 ( .B1(n9362), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9363) );
  XNOR2_X1 U11719 ( .A(n9363), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12674) );
  NOR2_X1 U11720 ( .A1(n6481), .A2(n9898), .ZN(n9364) );
  AOI21_X1 U11721 ( .B1(n12674), .B2(n10013), .A(n9364), .ZN(n9365) );
  NAND2_X1 U11722 ( .A1(n9366), .A2(n9365), .ZN(n11889) );
  AND2_X1 U11723 ( .A1(n9367), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9368) );
  OR2_X1 U11724 ( .A1(n9368), .A2(n9388), .ZN(n11890) );
  NAND2_X1 U11725 ( .A1(n11890), .A2(n9594), .ZN(n9374) );
  INV_X1 U11726 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12641) );
  INV_X1 U11727 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n11918) );
  OR2_X1 U11728 ( .A1(n9369), .A2(n11918), .ZN(n9370) );
  OAI21_X1 U11729 ( .B1(n12540), .B2(n12641), .A(n9370), .ZN(n9371) );
  INV_X1 U11730 ( .A(n9371), .ZN(n9373) );
  NAND2_X1 U11731 ( .A1(n9156), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9372) );
  OR2_X1 U11732 ( .A1(n11889), .A2(n12921), .ZN(n12462) );
  NAND2_X1 U11733 ( .A1(n11889), .A2(n12921), .ZN(n12467) );
  NAND2_X1 U11734 ( .A1(n12462), .A2(n12467), .ZN(n12575) );
  NAND2_X1 U11735 ( .A1(n11889), .A2(n12604), .ZN(n9375) );
  NAND2_X1 U11736 ( .A1(n10534), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U11737 ( .A1(n10532), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9378) );
  OR2_X1 U11738 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  NAND2_X1 U11739 ( .A1(n9396), .A2(n9381), .ZN(n9992) );
  OR2_X1 U11740 ( .A1(n9992), .A2(n9475), .ZN(n9386) );
  OAI21_X1 U11741 ( .B1(n9383), .B2(n9382), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9384) );
  XNOR2_X1 U11742 ( .A(n9384), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U11743 ( .A1(n9439), .A2(SI_16_), .B1(n10013), .B2(n12682), .ZN(
        n9385) );
  INV_X1 U11744 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13041) );
  NOR2_X1 U11745 ( .A1(n9388), .A2(n11760), .ZN(n9389) );
  OR2_X1 U11746 ( .A1(n9404), .A2(n9389), .ZN(n12926) );
  NAND2_X1 U11747 ( .A1(n12926), .A2(n9594), .ZN(n9391) );
  AOI22_X1 U11748 ( .A1(n9610), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12538), 
        .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n9390) );
  OAI211_X1 U11749 ( .C1(n12543), .C2(n13041), .A(n9391), .B(n9390), .ZN(
        n12909) );
  OR2_X1 U11750 ( .A1(n12925), .A2(n12909), .ZN(n9392) );
  NAND2_X1 U11751 ( .A1(n12919), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11752 ( .A1(n12925), .A2(n12909), .ZN(n9393) );
  NAND2_X1 U11753 ( .A1(n9394), .A2(n9393), .ZN(n12908) );
  NAND2_X1 U11754 ( .A1(n10678), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9414) );
  INV_X1 U11755 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U11756 ( .A1(n10676), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11757 ( .A1(n9414), .A2(n9397), .ZN(n9411) );
  XNOR2_X1 U11758 ( .A(n9413), .B(n9411), .ZN(n10316) );
  NAND2_X1 U11759 ( .A1(n10316), .A2(n12537), .ZN(n9402) );
  MUX2_X1 U11760 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9399), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9400) );
  NAND2_X1 U11761 ( .A1(n9400), .A2(n9646), .ZN(n12709) );
  INV_X1 U11762 ( .A(n12709), .ZN(n14173) );
  AOI22_X1 U11763 ( .A1(n9439), .A2(SI_17_), .B1(n10013), .B2(n14173), .ZN(
        n9401) );
  OR2_X1 U11764 ( .A1(n9404), .A2(n9403), .ZN(n9405) );
  NAND2_X1 U11765 ( .A1(n9422), .A2(n9405), .ZN(n12914) );
  NAND2_X1 U11766 ( .A1(n12914), .A2(n9594), .ZN(n9408) );
  AOI22_X1 U11767 ( .A1(n9610), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12538), 
        .B2(P3_REG1_REG_17__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U11768 ( .A1(n9156), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9406) );
  OR2_X1 U11769 ( .A1(n12988), .A2(n12922), .ZN(n12473) );
  NAND2_X1 U11770 ( .A1(n12988), .A2(n12922), .ZN(n12472) );
  NAND2_X1 U11771 ( .A1(n12473), .A2(n12472), .ZN(n9631) );
  INV_X1 U11772 ( .A(n12922), .ZN(n12602) );
  NAND2_X1 U11773 ( .A1(n12988), .A2(n12602), .ZN(n9409) );
  INV_X1 U11774 ( .A(n9411), .ZN(n9412) );
  NAND2_X1 U11775 ( .A1(n10847), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9431) );
  INV_X1 U11776 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U11777 ( .A1(n10845), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9415) );
  OR2_X1 U11778 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U11779 ( .A1(n9432), .A2(n9418), .ZN(n10326) );
  OR2_X1 U11780 ( .A1(n10326), .A2(n9475), .ZN(n9421) );
  NAND2_X1 U11781 ( .A1(n9646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9419) );
  XNOR2_X1 U11782 ( .A(n9419), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U11783 ( .A1(n9439), .A2(SI_18_), .B1(n10013), .B2(n12726), .ZN(
        n9420) );
  NAND2_X1 U11784 ( .A1(n9421), .A2(n9420), .ZN(n12367) );
  NAND2_X1 U11785 ( .A1(n9422), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11786 ( .A1(n9442), .A2(n9423), .ZN(n12903) );
  NAND2_X1 U11787 ( .A1(n12903), .A2(n9594), .ZN(n9428) );
  INV_X1 U11788 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U11789 ( .A1(n9610), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11790 ( .A1(n12538), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9424) );
  OAI211_X1 U11791 ( .C1(n13036), .C2(n12543), .A(n9425), .B(n9424), .ZN(n9426) );
  INV_X1 U11792 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U11793 ( .A1(n12367), .A2(n12886), .ZN(n12479) );
  OR2_X1 U11794 ( .A1(n12367), .A2(n12910), .ZN(n9430) );
  NAND2_X1 U11795 ( .A1(n10884), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U11796 ( .A1(n10886), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9433) );
  OR2_X1 U11797 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  NAND2_X1 U11798 ( .A1(n9454), .A2(n9436), .ZN(n10464) );
  OR2_X1 U11799 ( .A1(n10464), .A2(n9475), .ZN(n9441) );
  INV_X1 U11800 ( .A(n9603), .ZN(n9437) );
  NAND2_X1 U11801 ( .A1(n9437), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9438) );
  AOI22_X1 U11802 ( .A1(n9439), .A2(SI_19_), .B1(n12723), .B2(n10013), .ZN(
        n9440) );
  AND2_X1 U11803 ( .A1(n9442), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9443) );
  OR2_X1 U11804 ( .A1(n9443), .A2(n9461), .ZN(n12889) );
  NAND2_X1 U11805 ( .A1(n12889), .A2(n9594), .ZN(n9449) );
  INV_X1 U11806 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11807 ( .A1(n12538), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11808 ( .A1(n9156), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9444) );
  OAI211_X1 U11809 ( .C1(n9446), .C2(n12540), .A(n9445), .B(n9444), .ZN(n9447)
         );
  INV_X1 U11810 ( .A(n9447), .ZN(n9448) );
  NAND2_X1 U11811 ( .A1(n9449), .A2(n9448), .ZN(n12866) );
  NAND2_X1 U11812 ( .A1(n12561), .A2(n12866), .ZN(n9450) );
  OR2_X1 U11813 ( .A1(n12561), .A2(n12866), .ZN(n9451) );
  NAND2_X1 U11814 ( .A1(n9456), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U11815 ( .A1(n9470), .A2(n9457), .ZN(n10723) );
  OR2_X1 U11816 ( .A1(n10723), .A2(n9475), .ZN(n9459) );
  OR2_X1 U11817 ( .A1(n6481), .A2(n10724), .ZN(n9458) );
  NOR2_X1 U11818 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  OR2_X1 U11819 ( .A1(n9479), .A2(n9462), .ZN(n12877) );
  NAND2_X1 U11820 ( .A1(n12877), .A2(n9594), .ZN(n9468) );
  INV_X1 U11821 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U11822 ( .A1(n9610), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11823 ( .A1(n12538), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9463) );
  OAI211_X1 U11824 ( .C1(n9465), .C2(n12543), .A(n9464), .B(n9463), .ZN(n9466)
         );
  INV_X1 U11825 ( .A(n9466), .ZN(n9467) );
  NAND2_X1 U11826 ( .A1(n12976), .A2(n12885), .ZN(n12489) );
  NAND2_X1 U11827 ( .A1(n12976), .A2(n12601), .ZN(n9469) );
  INV_X1 U11828 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11513) );
  NAND2_X1 U11829 ( .A1(n11513), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U11830 ( .A1(n11510), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9471) );
  OR2_X1 U11831 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  NAND2_X1 U11832 ( .A1(n9490), .A2(n9474), .ZN(n11921) );
  OR2_X1 U11833 ( .A1(n11921), .A2(n9475), .ZN(n9477) );
  OR2_X1 U11834 ( .A1(n6481), .A2(n11922), .ZN(n9476) );
  OR2_X1 U11835 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  NAND2_X1 U11836 ( .A1(n9494), .A2(n9480), .ZN(n12861) );
  NAND2_X1 U11837 ( .A1(n12861), .A2(n9594), .ZN(n9485) );
  INV_X1 U11838 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U11839 ( .A1(n9610), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U11840 ( .A1(n12538), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9481) );
  OAI211_X1 U11841 ( .C1(n13027), .C2(n12543), .A(n9482), .B(n9481), .ZN(n9483) );
  INV_X1 U11842 ( .A(n9483), .ZN(n9484) );
  OR2_X1 U11843 ( .A1(n12860), .A2(n12872), .ZN(n9486) );
  NAND2_X1 U11844 ( .A1(n12855), .A2(n9486), .ZN(n9488) );
  NAND2_X1 U11845 ( .A1(n12860), .A2(n12872), .ZN(n9487) );
  XNOR2_X1 U11846 ( .A(n11565), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9503) );
  XNOR2_X1 U11847 ( .A(n9504), .B(n9503), .ZN(n10848) );
  NAND2_X1 U11848 ( .A1(n10848), .A2(n12537), .ZN(n9493) );
  OR2_X1 U11849 ( .A1(n6481), .A2(n9491), .ZN(n9492) );
  NAND2_X1 U11850 ( .A1(n9494), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U11851 ( .A1(n9508), .A2(n9495), .ZN(n12850) );
  NAND2_X1 U11852 ( .A1(n12850), .A2(n9594), .ZN(n9500) );
  INV_X1 U11853 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13023) );
  NAND2_X1 U11854 ( .A1(n9610), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11855 ( .A1(n12538), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9496) );
  OAI211_X1 U11856 ( .C1(n13023), .C2(n12543), .A(n9497), .B(n9496), .ZN(n9498) );
  INV_X1 U11857 ( .A(n9498), .ZN(n9499) );
  AND2_X1 U11858 ( .A1(n12849), .A2(n12831), .ZN(n9502) );
  OR2_X1 U11859 ( .A1(n12849), .A2(n12831), .ZN(n9501) );
  NAND2_X1 U11860 ( .A1(n11565), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9505) );
  XNOR2_X1 U11861 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9517) );
  XNOR2_X1 U11862 ( .A(n9518), .B(n9517), .ZN(n10915) );
  NAND2_X1 U11863 ( .A1(n10915), .A2(n12537), .ZN(n9507) );
  OR2_X1 U11864 ( .A1(n6481), .A2(n10917), .ZN(n9506) );
  AND2_X1 U11865 ( .A1(n9508), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9509) );
  OR2_X1 U11866 ( .A1(n9509), .A2(n9523), .ZN(n12835) );
  NAND2_X1 U11867 ( .A1(n12835), .A2(n9594), .ZN(n9515) );
  INV_X1 U11868 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11869 ( .A1(n9610), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11870 ( .A1(n12538), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9510) );
  OAI211_X1 U11871 ( .C1(n9512), .C2(n12543), .A(n9511), .B(n9510), .ZN(n9513)
         );
  INV_X1 U11872 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U11873 ( .A1(n12963), .A2(n12845), .ZN(n12501) );
  OR2_X2 U11874 ( .A1(n12829), .A2(n12839), .ZN(n12828) );
  NAND2_X1 U11875 ( .A1(n12963), .A2(n12818), .ZN(n9516) );
  NAND2_X1 U11876 ( .A1(n9519), .A2(n11839), .ZN(n9520) );
  NAND2_X1 U11877 ( .A1(n9521), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11878 ( .A1(n9533), .A2(n9522), .ZN(n11294) );
  OR2_X1 U11879 ( .A1(n9523), .A2(n12341), .ZN(n9524) );
  NAND2_X1 U11880 ( .A1(n9537), .A2(n9524), .ZN(n12822) );
  NAND2_X1 U11881 ( .A1(n12822), .A2(n9594), .ZN(n9530) );
  INV_X1 U11882 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11883 ( .A1(n12538), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U11884 ( .A1(n9610), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9525) );
  OAI211_X1 U11885 ( .C1(n9527), .C2(n12543), .A(n9526), .B(n9525), .ZN(n9528)
         );
  INV_X1 U11886 ( .A(n9528), .ZN(n9529) );
  NAND2_X1 U11887 ( .A1(n12958), .A2(n12832), .ZN(n9531) );
  XNOR2_X1 U11888 ( .A(n11882), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U11889 ( .A(n9545), .B(n9534), .ZN(n11629) );
  NAND2_X1 U11890 ( .A1(n11629), .A2(n12537), .ZN(n9536) );
  OR2_X1 U11891 ( .A1(n6481), .A2(n11631), .ZN(n9535) );
  NAND2_X1 U11892 ( .A1(n9537), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U11893 ( .A1(n9566), .A2(n9538), .ZN(n12805) );
  NAND2_X1 U11894 ( .A1(n12805), .A2(n9594), .ZN(n9543) );
  INV_X1 U11895 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U11896 ( .A1(n9610), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11897 ( .A1(n12538), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9539) );
  OAI211_X1 U11898 ( .C1(n13017), .C2(n12543), .A(n9540), .B(n9539), .ZN(n9541) );
  INV_X1 U11899 ( .A(n9541), .ZN(n9542) );
  OR2_X1 U11900 ( .A1(n12315), .A2(n12821), .ZN(n12509) );
  NAND2_X1 U11901 ( .A1(n12315), .A2(n12821), .ZN(n12510) );
  NAND2_X1 U11902 ( .A1(n12509), .A2(n12510), .ZN(n12800) );
  INV_X1 U11903 ( .A(n12821), .ZN(n12600) );
  NAND2_X1 U11904 ( .A1(n11882), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U11905 ( .A1(n11987), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9546) );
  XNOR2_X1 U11906 ( .A(n13580), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9548) );
  XNOR2_X1 U11907 ( .A(n9558), .B(n9548), .ZN(n11643) );
  NAND2_X1 U11908 ( .A1(n11643), .A2(n12537), .ZN(n9550) );
  OR2_X1 U11909 ( .A1(n6481), .A2(n11645), .ZN(n9549) );
  XNOR2_X1 U11910 ( .A(n9566), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U11911 ( .A1(n12790), .A2(n9594), .ZN(n9555) );
  INV_X1 U11912 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U11913 ( .A1(n9610), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U11914 ( .A1(n12538), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9551) );
  OAI211_X1 U11915 ( .C1(n13013), .C2(n12543), .A(n9552), .B(n9551), .ZN(n9553) );
  INV_X1 U11916 ( .A(n9553), .ZN(n9554) );
  OR2_X1 U11917 ( .A1(n12791), .A2(n12802), .ZN(n9556) );
  NOR2_X1 U11918 ( .A1(n13580), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U11919 ( .A1(n13580), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9559) );
  XNOR2_X1 U11920 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9560) );
  XNOR2_X1 U11921 ( .A(n9576), .B(n9560), .ZN(n11735) );
  NAND2_X1 U11922 ( .A1(n11735), .A2(n12537), .ZN(n9563) );
  OR2_X1 U11923 ( .A1(n6481), .A2(n11736), .ZN(n9562) );
  OAI21_X1 U11924 ( .B1(n9566), .B2(P3_REG3_REG_26__SCAN_IN), .A(
        P3_REG3_REG_27__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U11925 ( .A1(n12378), .A2(n9564), .ZN(n9565) );
  NAND2_X1 U11926 ( .A1(n9567), .A2(n9581), .ZN(n12777) );
  NAND2_X1 U11927 ( .A1(n12777), .A2(n9594), .ZN(n9572) );
  INV_X1 U11928 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U11929 ( .A1(n9610), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U11930 ( .A1(n12538), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9568) );
  OAI211_X1 U11931 ( .C1(n13009), .C2(n12543), .A(n9569), .B(n9568), .ZN(n9570) );
  INV_X1 U11932 ( .A(n9570), .ZN(n9571) );
  OR2_X1 U11933 ( .A1(n12778), .A2(n12786), .ZN(n12518) );
  NAND2_X1 U11934 ( .A1(n12778), .A2(n12786), .ZN(n12752) );
  OR2_X1 U11935 ( .A1(n12778), .A2(n12758), .ZN(n9574) );
  AND2_X1 U11936 ( .A1(n13577), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U11937 ( .A1(n14124), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9577) );
  XNOR2_X1 U11938 ( .A(n9589), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U11939 ( .A(n9588), .B(n9578), .ZN(n11923) );
  NAND2_X1 U11940 ( .A1(n11923), .A2(n12537), .ZN(n9580) );
  OR2_X1 U11941 ( .A1(n6481), .A2(n11924), .ZN(n9579) );
  AND2_X1 U11942 ( .A1(n9581), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9582) );
  INV_X1 U11943 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U11944 ( .A1(n9610), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U11945 ( .A1(n12538), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9583) );
  OAI211_X1 U11946 ( .C1(n13005), .C2(n12543), .A(n9584), .B(n9583), .ZN(n9585) );
  NAND2_X1 U11947 ( .A1(n12268), .A2(n12773), .ZN(n12387) );
  INV_X1 U11948 ( .A(n12773), .ZN(n12599) );
  NOR2_X1 U11949 ( .A1(n9589), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U11950 ( .A1(n9589), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9590) );
  XNOR2_X1 U11951 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12223) );
  XNOR2_X1 U11952 ( .A(n12225), .B(n12223), .ZN(n13054) );
  NAND2_X1 U11953 ( .A1(n13054), .A2(n12537), .ZN(n9593) );
  OR2_X1 U11954 ( .A1(n6481), .A2(n13057), .ZN(n9592) );
  INV_X1 U11955 ( .A(n11982), .ZN(n9600) );
  NAND2_X1 U11956 ( .A1(n12744), .A2(n9594), .ZN(n12547) );
  INV_X1 U11957 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U11958 ( .A1(n9610), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11959 ( .A1(n12538), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9595) );
  OAI211_X1 U11960 ( .C1(n9597), .C2(n12543), .A(n9596), .B(n9595), .ZN(n9598)
         );
  INV_X1 U11961 ( .A(n9598), .ZN(n9599) );
  NAND2_X1 U11962 ( .A1(n12547), .A2(n9599), .ZN(n12757) );
  INV_X1 U11963 ( .A(n12757), .ZN(n12267) );
  NAND2_X1 U11964 ( .A1(n9600), .A2(n12267), .ZN(n12531) );
  NAND2_X1 U11965 ( .A1(n11982), .A2(n12757), .ZN(n12550) );
  XNOR2_X1 U11966 ( .A(n9601), .B(n12584), .ZN(n9620) );
  NAND2_X1 U11967 ( .A1(n9661), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9604) );
  NAND2_X1 U11968 ( .A1(n12595), .A2(n12723), .ZN(n9693) );
  NAND2_X1 U11969 ( .A1(n9605), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9606) );
  MUX2_X1 U11970 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9606), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9607) );
  NAND2_X1 U11971 ( .A1(n9608), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U11972 ( .A1(n10791), .A2(n9692), .ZN(n12560) );
  INV_X1 U11973 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U11974 ( .A1(n9610), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9612) );
  NAND2_X1 U11975 ( .A1(n12538), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9611) );
  OAI211_X1 U11976 ( .C1(n9613), .C2(n12543), .A(n9612), .B(n9611), .ZN(n9614)
         );
  INV_X1 U11977 ( .A(n9614), .ZN(n9615) );
  AND2_X1 U11978 ( .A1(n12547), .A2(n9615), .ZN(n12548) );
  INV_X1 U11979 ( .A(n11925), .ZN(n12592) );
  NAND2_X1 U11980 ( .A1(n12592), .A2(n12627), .ZN(n10014) );
  AND2_X1 U11981 ( .A1(n9103), .A2(n10014), .ZN(n10111) );
  INV_X1 U11982 ( .A(n10111), .ZN(n10114) );
  NAND2_X1 U11983 ( .A1(n12592), .A2(P3_B_REG_SCAN_IN), .ZN(n9617) );
  NAND2_X1 U11984 ( .A1(n14962), .A2(n9617), .ZN(n12745) );
  NAND2_X1 U11985 ( .A1(n12599), .A2(n14965), .ZN(n9618) );
  OAI21_X1 U11986 ( .B1(n12548), .B2(n12745), .A(n9618), .ZN(n9619) );
  NAND2_X1 U11987 ( .A1(n14993), .A2(n12394), .ZN(n9622) );
  NAND2_X1 U11988 ( .A1(n9622), .A2(n10094), .ZN(n14975) );
  INV_X1 U11989 ( .A(n12406), .ZN(n12562) );
  NAND2_X1 U11990 ( .A1(n10918), .A2(n12562), .ZN(n9623) );
  INV_X1 U11991 ( .A(n10933), .ZN(n12563) );
  NAND2_X1 U11992 ( .A1(n14945), .A2(n14944), .ZN(n9624) );
  INV_X1 U11993 ( .A(n12609), .ZN(n10689) );
  NAND2_X1 U11994 ( .A1(n10689), .A2(n10840), .ZN(n12424) );
  NAND2_X1 U11995 ( .A1(n9624), .A2(n12424), .ZN(n11086) );
  NAND2_X1 U11996 ( .A1(n11086), .A2(n12569), .ZN(n9625) );
  NOR2_X1 U11997 ( .A1(n11249), .A2(n14935), .ZN(n9626) );
  NAND2_X1 U11998 ( .A1(n11249), .A2(n14935), .ZN(n9627) );
  INV_X1 U11999 ( .A(n12438), .ZN(n9628) );
  INV_X1 U12000 ( .A(n11261), .ZN(n14207) );
  OR2_X1 U12001 ( .A1(n14207), .A2(n14936), .ZN(n12442) );
  NAND2_X1 U12002 ( .A1(n14207), .A2(n14936), .ZN(n12443) );
  INV_X1 U12003 ( .A(n11769), .ZN(n12573) );
  NAND2_X1 U12004 ( .A1(n11767), .A2(n12573), .ZN(n9629) );
  NOR2_X1 U12005 ( .A1(n14193), .A2(n12606), .ZN(n12453) );
  NAND2_X1 U12006 ( .A1(n14193), .A2(n12606), .ZN(n12446) );
  INV_X1 U12007 ( .A(n12575), .ZN(n12460) );
  INV_X1 U12008 ( .A(n12909), .ZN(n12229) );
  OR2_X1 U12009 ( .A1(n12925), .A2(n12229), .ZN(n12469) );
  NAND2_X1 U12010 ( .A1(n12925), .A2(n12229), .ZN(n12468) );
  NAND2_X1 U12011 ( .A1(n12913), .A2(n12912), .ZN(n9632) );
  OR2_X1 U12012 ( .A1(n12561), .A2(n12899), .ZN(n12485) );
  AND2_X1 U12013 ( .A1(n12561), .A2(n12899), .ZN(n12484) );
  NAND2_X1 U12014 ( .A1(n12876), .A2(n12488), .ZN(n12858) );
  NAND2_X1 U12015 ( .A1(n12860), .A2(n12846), .ZN(n12492) );
  OR2_X1 U12016 ( .A1(n12860), .A2(n12846), .ZN(n12493) );
  NAND2_X1 U12017 ( .A1(n12849), .A2(n12857), .ZN(n12498) );
  NAND2_X1 U12018 ( .A1(n12958), .A2(n7179), .ZN(n12388) );
  NAND2_X1 U12019 ( .A1(n12798), .A2(n12797), .ZN(n9633) );
  INV_X1 U12020 ( .A(n12802), .ZN(n12772) );
  OR2_X1 U12021 ( .A1(n12791), .A2(n12772), .ZN(n12515) );
  NAND2_X1 U12022 ( .A1(n12783), .A2(n12515), .ZN(n9634) );
  NAND2_X1 U12023 ( .A1(n12791), .A2(n12772), .ZN(n12516) );
  NAND2_X1 U12024 ( .A1(n9634), .A2(n12516), .ZN(n12766) );
  AND2_X1 U12025 ( .A1(n12387), .A2(n12752), .ZN(n12523) );
  NAND2_X1 U12026 ( .A1(n12768), .A2(n12523), .ZN(n9635) );
  NAND2_X1 U12027 ( .A1(n9635), .A2(n12521), .ZN(n12552) );
  INV_X1 U12028 ( .A(n12584), .ZN(n9636) );
  XNOR2_X1 U12029 ( .A(n12552), .B(n9636), .ZN(n11984) );
  OAI21_X1 U12030 ( .B1(n9644), .B2(n9692), .A(n12723), .ZN(n9637) );
  NAND2_X1 U12031 ( .A1(n9637), .A2(n12393), .ZN(n9640) );
  NAND2_X1 U12032 ( .A1(n12393), .A2(n10725), .ZN(n9638) );
  NAND2_X1 U12033 ( .A1(n9644), .A2(n9638), .ZN(n9639) );
  NAND2_X1 U12034 ( .A1(n9640), .A2(n9639), .ZN(n10106) );
  AND2_X1 U12035 ( .A1(n15047), .A2(n9694), .ZN(n9641) );
  NAND2_X1 U12036 ( .A1(n10106), .A2(n9641), .ZN(n9643) );
  AND2_X1 U12037 ( .A1(n9692), .A2(n12740), .ZN(n9642) );
  NAND2_X1 U12038 ( .A1(n12595), .A2(n9642), .ZN(n9683) );
  NAND2_X1 U12039 ( .A1(n9644), .A2(n14979), .ZN(n15049) );
  NAND2_X1 U12040 ( .A1(n11984), .A2(n15063), .ZN(n9645) );
  INV_X1 U12041 ( .A(n9646), .ZN(n9648) );
  XNOR2_X1 U12042 ( .A(n9655), .B(P3_B_REG_SCAN_IN), .ZN(n9653) );
  OAI21_X1 U12043 ( .B1(n9649), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9650) );
  MUX2_X1 U12044 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9650), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9652) );
  NAND2_X1 U12045 ( .A1(n9651), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9654) );
  INV_X1 U12046 ( .A(n9664), .ZN(n11646) );
  NAND2_X1 U12047 ( .A1(n9655), .A2(n11646), .ZN(n9656) );
  NAND2_X1 U12048 ( .A1(n11632), .A2(n11646), .ZN(n9659) );
  AND2_X1 U12049 ( .A1(n9657), .A2(n10332), .ZN(n9699) );
  INV_X1 U12050 ( .A(n9699), .ZN(n9679) );
  AND2_X1 U12051 ( .A1(n9665), .A2(n9664), .ZN(n9666) );
  NAND2_X1 U12052 ( .A1(n9667), .A2(n9666), .ZN(n10080) );
  NOR2_X1 U12053 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9671) );
  NOR4_X1 U12054 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9670) );
  NOR4_X1 U12055 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9669) );
  NOR4_X1 U12056 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9668) );
  NAND4_X1 U12057 ( .A1(n9671), .A2(n9670), .A3(n9669), .A4(n9668), .ZN(n9677)
         );
  NOR4_X1 U12058 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9675) );
  NOR4_X1 U12059 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9674) );
  NOR4_X1 U12060 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9673) );
  NOR4_X1 U12061 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9672) );
  NAND4_X1 U12062 ( .A1(n9675), .A2(n9674), .A3(n9673), .A4(n9672), .ZN(n9676)
         );
  NOR2_X1 U12063 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  NAND3_X1 U12064 ( .A1(n9679), .A2(n10337), .A3(n9698), .ZN(n9680) );
  NAND2_X1 U12065 ( .A1(n12595), .A2(n12740), .ZN(n9681) );
  OAI21_X1 U12066 ( .B1(n15047), .B2(n9692), .A(n9681), .ZN(n9682) );
  INV_X1 U12067 ( .A(n9694), .ZN(n12587) );
  AOI21_X1 U12068 ( .B1(n9682), .B2(n12587), .A(n12525), .ZN(n9686) );
  NAND2_X1 U12069 ( .A1(n12514), .A2(n9683), .ZN(n10331) );
  NAND2_X1 U12070 ( .A1(n12525), .A2(n12587), .ZN(n10334) );
  NAND2_X1 U12071 ( .A1(n10331), .A2(n10334), .ZN(n9684) );
  NAND2_X1 U12072 ( .A1(n9684), .A2(n13045), .ZN(n9685) );
  OAI21_X1 U12073 ( .B1(n9686), .B2(n13045), .A(n9685), .ZN(n9687) );
  INV_X1 U12074 ( .A(n9687), .ZN(n9688) );
  NAND2_X1 U12075 ( .A1(n9600), .A2(n9689), .ZN(n9690) );
  NAND2_X1 U12076 ( .A1(n9691), .A2(n9690), .ZN(P3_U3488) );
  NAND2_X1 U12077 ( .A1(n12393), .A2(n9692), .ZN(n12588) );
  NOR2_X1 U12078 ( .A1(n9693), .A2(n12588), .ZN(n10078) );
  NAND2_X1 U12079 ( .A1(n10337), .A2(n10078), .ZN(n10104) );
  INV_X1 U12080 ( .A(n10337), .ZN(n9695) );
  NAND2_X1 U12081 ( .A1(n12525), .A2(n9694), .ZN(n10338) );
  OR2_X1 U12082 ( .A1(n9695), .A2(n10338), .ZN(n10085) );
  NAND2_X1 U12083 ( .A1(n10104), .A2(n10085), .ZN(n9697) );
  AND2_X1 U12084 ( .A1(n9696), .A2(n9698), .ZN(n10113) );
  NAND2_X1 U12085 ( .A1(n9697), .A2(n10113), .ZN(n9701) );
  AND2_X1 U12086 ( .A1(n9699), .A2(n9698), .ZN(n10110) );
  NAND3_X1 U12087 ( .A1(n10110), .A2(n10337), .A3(n10106), .ZN(n9700) );
  NAND2_X1 U12088 ( .A1(n15066), .A2(n15015), .ZN(n13043) );
  NAND2_X1 U12089 ( .A1(n9704), .A2(n9703), .ZN(P3_U3456) );
  INV_X1 U12090 ( .A(n10328), .ZN(n9705) );
  INV_X1 U12091 ( .A(n9706), .ZN(n9707) );
  NAND2_X1 U12092 ( .A1(n9707), .A2(n9768), .ZN(n9772) );
  INV_X1 U12093 ( .A(n10080), .ZN(n9708) );
  NOR2_X1 U12094 ( .A1(n9733), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13048) );
  INV_X2 U12095 ( .A(n13048), .ZN(n13056) );
  OAI222_X1 U12096 ( .A1(n14842), .A2(P3_U3151), .B1(n13056), .B2(n9710), .C1(
        n9709), .C2(n13058), .ZN(P3_U3289) );
  OAI222_X1 U12097 ( .A1(n14776), .A2(P3_U3151), .B1(n13056), .B2(n9711), .C1(
        n7628), .C2(n13058), .ZN(P3_U3295) );
  INV_X1 U12098 ( .A(n9712), .ZN(n9714) );
  INV_X1 U12099 ( .A(SI_4_), .ZN(n9713) );
  OAI222_X1 U12100 ( .A1(n13056), .A2(n9714), .B1(n13058), .B2(n9713), .C1(
        n14807), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12101 ( .A(n9715), .ZN(n9717) );
  INV_X1 U12102 ( .A(n10056), .ZN(n11152) );
  OAI222_X1 U12103 ( .A1(n13056), .A2(n9717), .B1(n13058), .B2(n9716), .C1(
        n11152), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12104 ( .A(n9718), .ZN(n9720) );
  INV_X1 U12105 ( .A(SI_5_), .ZN(n9719) );
  OAI222_X1 U12106 ( .A1(n13056), .A2(n9720), .B1(n13058), .B2(n9719), .C1(
        n14824), .C2(P3_U3151), .ZN(P3_U3290) );
  INV_X1 U12107 ( .A(n9721), .ZN(n9723) );
  INV_X1 U12108 ( .A(SI_3_), .ZN(n9722) );
  INV_X1 U12109 ( .A(n11168), .ZN(n14792) );
  OAI222_X1 U12110 ( .A1(n13056), .A2(n9723), .B1(n13058), .B2(n9722), .C1(
        n14792), .C2(P3_U3151), .ZN(P3_U3292) );
  INV_X1 U12111 ( .A(n9724), .ZN(n9726) );
  INV_X1 U12112 ( .A(SI_7_), .ZN(n9725) );
  OAI222_X1 U12113 ( .A1(n13056), .A2(n9726), .B1(n13058), .B2(n9725), .C1(
        n14859), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12114 ( .A(n9728), .ZN(n9751) );
  INV_X1 U12115 ( .A(n10357), .ZN(n9729) );
  OAI222_X1 U12116 ( .A1(n14125), .A2(n9730), .B1(n14128), .B2(n9751), .C1(
        P1_U3086), .C2(n9729), .ZN(P1_U3353) );
  OAI222_X1 U12117 ( .A1(n13056), .A2(n9732), .B1(n13058), .B2(n9731), .C1(
        n14895), .C2(P3_U3151), .ZN(P3_U3286) );
  NOR2_X1 U12118 ( .A1(n9733), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13572) );
  INV_X2 U12119 ( .A(n13572), .ZN(n13578) );
  AND2_X1 U12120 ( .A1(n9733), .A2(P2_U3088), .ZN(n11624) );
  INV_X2 U12121 ( .A(n11624), .ZN(n13581) );
  OAI222_X1 U12122 ( .A1(n13578), .A2(n9734), .B1(n13581), .B2(n9736), .C1(
        n14600), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U12123 ( .A(n13693), .ZN(n9735) );
  OAI222_X1 U12124 ( .A1(n14125), .A2(n6648), .B1(n14128), .B2(n9736), .C1(
        n9735), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U12125 ( .A(n9737), .ZN(n9747) );
  INV_X1 U12126 ( .A(n13711), .ZN(n9738) );
  OAI222_X1 U12127 ( .A1(n14125), .A2(n9739), .B1(n14128), .B2(n9747), .C1(
        P1_U3086), .C2(n9738), .ZN(P1_U3352) );
  OAI222_X1 U12128 ( .A1(n13056), .A2(n9741), .B1(n13058), .B2(n9740), .C1(
        n11213), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12129 ( .A(n8545), .ZN(n9749) );
  INV_X1 U12130 ( .A(n13719), .ZN(n9928) );
  OAI222_X1 U12131 ( .A1(n14125), .A2(n9742), .B1(n14128), .B2(n9749), .C1(
        P1_U3086), .C2(n9928), .ZN(P1_U3351) );
  OAI222_X1 U12132 ( .A1(n13056), .A2(n9744), .B1(n13058), .B2(n9743), .C1(
        n14876), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12133 ( .A1(n13056), .A2(n9746), .B1(n13058), .B2(n9745), .C1(
        n11435), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12134 ( .A(n9780), .ZN(n9873) );
  OAI222_X1 U12135 ( .A1(n13578), .A2(n9748), .B1(n13581), .B2(n9747), .C1(
        P2_U3088), .C2(n9873), .ZN(P2_U3324) );
  INV_X1 U12136 ( .A(n9781), .ZN(n9817) );
  OAI222_X1 U12137 ( .A1(n13578), .A2(n9750), .B1(n13581), .B2(n9749), .C1(
        P2_U3088), .C2(n9817), .ZN(P2_U3323) );
  INV_X1 U12138 ( .A(n9779), .ZN(n14613) );
  OAI222_X1 U12139 ( .A1(n13578), .A2(n9752), .B1(n13581), .B2(n9751), .C1(
        P2_U3088), .C2(n14613), .ZN(P2_U3325) );
  OAI222_X1 U12140 ( .A1(P3_U3151), .A2(n10028), .B1(n13058), .B2(n9754), .C1(
        n13056), .C2(n9753), .ZN(P3_U3294) );
  INV_X1 U12141 ( .A(n9755), .ZN(n9757) );
  OAI222_X1 U12142 ( .A1(n14125), .A2(n9756), .B1(n14128), .B2(n9757), .C1(
        P1_U3086), .C2(n9946), .ZN(P1_U3350) );
  INV_X1 U12143 ( .A(n9782), .ZN(n9839) );
  OAI222_X1 U12144 ( .A1(n13578), .A2(n9758), .B1(n13581), .B2(n9757), .C1(
        P2_U3088), .C2(n9839), .ZN(P2_U3322) );
  AND2_X1 U12145 ( .A1(n9824), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12146 ( .A1(n9824), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12147 ( .A1(n9824), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12148 ( .A1(n9824), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12149 ( .A1(n9824), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12150 ( .A1(n9824), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12151 ( .A1(n9824), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12152 ( .A1(n9824), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12153 ( .A1(n9824), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12154 ( .A1(n9824), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12155 ( .A1(n9824), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12156 ( .A1(n9824), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12157 ( .A1(n9824), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12158 ( .A1(n9824), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12159 ( .A1(n9824), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12160 ( .A1(n9824), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  INV_X1 U12161 ( .A(n9759), .ZN(n9761) );
  OAI222_X1 U12162 ( .A1(n13056), .A2(n9761), .B1(n13058), .B2(n9760), .C1(
        n11714), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12163 ( .A(n9762), .ZN(n9764) );
  INV_X1 U12164 ( .A(n9931), .ZN(n13734) );
  OAI222_X1 U12165 ( .A1(n14125), .A2(n9763), .B1(n14128), .B2(n9764), .C1(
        P1_U3086), .C2(n13734), .ZN(P1_U3349) );
  INV_X1 U12166 ( .A(n9848), .ZN(n9841) );
  OAI222_X1 U12167 ( .A1(n13578), .A2(n9765), .B1(n13581), .B2(n9764), .C1(
        P2_U3088), .C2(n9841), .ZN(P2_U3321) );
  NAND2_X1 U12168 ( .A1(n9020), .A2(P2_U3947), .ZN(n9766) );
  OAI21_X1 U12169 ( .B1(P2_U3947), .B2(n9114), .A(n9766), .ZN(P2_U3531) );
  INV_X1 U12170 ( .A(n14600), .ZN(n9767) );
  MUX2_X1 U12171 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n13412), .S(n14600), .Z(
        n14604) );
  NAND2_X1 U12172 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n14603) );
  AOI21_X1 U12173 ( .B1(n9767), .B2(P2_REG2_REG_1__SCAN_IN), .A(n14602), .ZN(
        n14621) );
  MUX2_X1 U12174 ( .A(n8513), .B(P2_REG2_REG_2__SCAN_IN), .S(n9779), .Z(n14620) );
  NOR2_X1 U12175 ( .A1(n14613), .A2(n8513), .ZN(n9861) );
  INV_X1 U12176 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U12177 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11043), .S(n9780), .Z(n9860) );
  OAI21_X1 U12178 ( .B1(n14619), .B2(n9861), .A(n9860), .ZN(n9859) );
  NAND2_X1 U12179 ( .A1(n9780), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9812) );
  MUX2_X1 U12180 ( .A(n8539), .B(P2_REG2_REG_4__SCAN_IN), .S(n9781), .Z(n9811)
         );
  NOR2_X1 U12181 ( .A1(n9817), .A2(n8539), .ZN(n9832) );
  MUX2_X1 U12182 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11034), .S(n9782), .Z(n9831) );
  OAI21_X1 U12183 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9830) );
  NAND2_X1 U12184 ( .A1(n9782), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9775) );
  MUX2_X1 U12185 ( .A(n11063), .B(P2_REG2_REG_6__SCAN_IN), .S(n9848), .Z(n9774) );
  AOI21_X1 U12186 ( .B1(n9830), .B2(n9775), .A(n9774), .ZN(n9847) );
  NAND2_X1 U12187 ( .A1(n10228), .A2(n9768), .ZN(n9769) );
  NAND2_X1 U12188 ( .A1(n9770), .A2(n9769), .ZN(n9771) );
  NAND2_X1 U12189 ( .A1(n9772), .A2(n9771), .ZN(n9789) );
  NOR2_X1 U12190 ( .A1(n10209), .A2(P2_U3088), .ZN(n13571) );
  NAND2_X1 U12191 ( .A1(n9789), .A2(n13571), .ZN(n9787) );
  INV_X1 U12192 ( .A(n9787), .ZN(n9773) );
  INV_X1 U12193 ( .A(n13576), .ZN(n11973) );
  NAND3_X1 U12194 ( .A1(n9830), .A2(n9775), .A3(n9774), .ZN(n9776) );
  NAND2_X1 U12195 ( .A1(n14655), .A2(n9776), .ZN(n9793) );
  MUX2_X1 U12196 ( .A(n9777), .B(P2_REG1_REG_1__SCAN_IN), .S(n14600), .Z(
        n14607) );
  NAND3_X1 U12197 ( .A1(n14607), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .ZN(n14606) );
  OAI21_X1 U12198 ( .B1(n9777), .B2(n14600), .A(n14606), .ZN(n14618) );
  MUX2_X1 U12199 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9778), .S(n9779), .Z(n14617) );
  NAND2_X1 U12200 ( .A1(n14618), .A2(n14617), .ZN(n14616) );
  NAND2_X1 U12201 ( .A1(n9779), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9868) );
  MUX2_X1 U12202 ( .A(n8527), .B(P2_REG1_REG_3__SCAN_IN), .S(n9780), .Z(n9867)
         );
  AOI21_X1 U12203 ( .B1(n14616), .B2(n9868), .A(n9867), .ZN(n9866) );
  AOI21_X1 U12204 ( .B1(n9780), .B2(P2_REG1_REG_3__SCAN_IN), .A(n9866), .ZN(
        n9807) );
  MUX2_X1 U12205 ( .A(n8540), .B(P2_REG1_REG_4__SCAN_IN), .S(n9781), .Z(n9806)
         );
  NOR2_X1 U12206 ( .A1(n9807), .A2(n9806), .ZN(n9805) );
  AOI21_X1 U12207 ( .B1(n9781), .B2(P2_REG1_REG_4__SCAN_IN), .A(n9805), .ZN(
        n9827) );
  MUX2_X1 U12208 ( .A(n8563), .B(P2_REG1_REG_5__SCAN_IN), .S(n9782), .Z(n9826)
         );
  NOR2_X1 U12209 ( .A1(n9827), .A2(n9826), .ZN(n9825) );
  INV_X1 U12210 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14760) );
  MUX2_X1 U12211 ( .A(n14760), .B(P2_REG1_REG_6__SCAN_IN), .S(n9848), .Z(n9784) );
  NOR2_X1 U12212 ( .A1(n9839), .A2(n8563), .ZN(n9786) );
  INV_X1 U12213 ( .A(n9786), .ZN(n9783) );
  NAND2_X1 U12214 ( .A1(n9784), .A2(n9783), .ZN(n9788) );
  MUX2_X1 U12215 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14760), .S(n9848), .Z(n9785) );
  OAI21_X1 U12216 ( .B1(n9825), .B2(n9786), .A(n9785), .ZN(n9840) );
  OAI211_X1 U12217 ( .C1(n9825), .C2(n9788), .A(n9840), .B(n14658), .ZN(n9792)
         );
  AND2_X1 U12218 ( .A1(n9789), .A2(n10209), .ZN(n14599) );
  AND2_X1 U12219 ( .A1(n14599), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14673) );
  OR2_X1 U12220 ( .A1(n9789), .A2(P2_U3088), .ZN(n14677) );
  NAND2_X1 U12221 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10550) );
  OAI21_X1 U12222 ( .B1(n14677), .B2(n6949), .A(n10550), .ZN(n9790) );
  AOI21_X1 U12223 ( .B1(n9848), .B2(n14673), .A(n9790), .ZN(n9791) );
  OAI211_X1 U12224 ( .C1(n9847), .C2(n9793), .A(n9792), .B(n9791), .ZN(
        P2_U3220) );
  INV_X1 U12225 ( .A(n9794), .ZN(n9796) );
  INV_X1 U12226 ( .A(n9850), .ZN(n14627) );
  OAI222_X1 U12227 ( .A1(n13578), .A2(n9795), .B1(n13581), .B2(n9796), .C1(
        P2_U3088), .C2(n14627), .ZN(P2_U3320) );
  INV_X1 U12228 ( .A(n9934), .ZN(n13748) );
  OAI222_X1 U12229 ( .A1(n14125), .A2(n9797), .B1(n14128), .B2(n9796), .C1(
        P1_U3086), .C2(n13748), .ZN(P1_U3348) );
  OAI222_X1 U12230 ( .A1(n13056), .A2(n9799), .B1(n13058), .B2(n9798), .C1(
        n12617), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12231 ( .A(n9800), .ZN(n9803) );
  INV_X1 U12232 ( .A(n9876), .ZN(n9801) );
  OAI222_X1 U12233 ( .A1(n13578), .A2(n9802), .B1(n13581), .B2(n9803), .C1(
        P2_U3088), .C2(n9801), .ZN(P2_U3319) );
  INV_X1 U12234 ( .A(n9954), .ZN(n9966) );
  OAI222_X1 U12235 ( .A1(n14125), .A2(n9804), .B1(n14128), .B2(n9803), .C1(
        P1_U3086), .C2(n9966), .ZN(P1_U3347) );
  INV_X1 U12236 ( .A(n14677), .ZN(n14652) );
  NAND2_X1 U12237 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10438) );
  AOI211_X1 U12238 ( .C1(n9807), .C2(n9806), .A(n9805), .B(n14668), .ZN(n9808)
         );
  INV_X1 U12239 ( .A(n9808), .ZN(n9809) );
  NAND2_X1 U12240 ( .A1(n10438), .A2(n9809), .ZN(n9810) );
  AOI21_X1 U12241 ( .B1(n14652), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9810), .ZN(
        n9816) );
  INV_X1 U12242 ( .A(n9833), .ZN(n9814) );
  NAND3_X1 U12243 ( .A1(n9859), .A2(n9812), .A3(n9811), .ZN(n9813) );
  NAND3_X1 U12244 ( .A1(n14655), .A2(n9814), .A3(n9813), .ZN(n9815) );
  OAI211_X1 U12245 ( .C1(n14644), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P2_U3218) );
  INV_X1 U12246 ( .A(n9818), .ZN(n9820) );
  INV_X1 U12247 ( .A(n10127), .ZN(n10132) );
  OAI222_X1 U12248 ( .A1(n13578), .A2(n9819), .B1(n13581), .B2(n9820), .C1(
        P2_U3088), .C2(n10132), .ZN(P2_U3318) );
  INV_X1 U12249 ( .A(n9968), .ZN(n9998) );
  OAI222_X1 U12250 ( .A1(n14125), .A2(n9821), .B1(n14128), .B2(n9820), .C1(
        P1_U3086), .C2(n9998), .ZN(P1_U3346) );
  OAI222_X1 U12251 ( .A1(n13056), .A2(n9823), .B1(n13058), .B2(n9822), .C1(
        n12644), .C2(P3_U3151), .ZN(P3_U3281) );
  AND2_X1 U12252 ( .A1(n9824), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12253 ( .A1(n9824), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12254 ( .A1(n9824), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12255 ( .A1(n9824), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12256 ( .A1(n9824), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12257 ( .A1(n9824), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12258 ( .A1(n9824), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12259 ( .A1(n9824), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12260 ( .A1(n9824), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12261 ( .A1(n9824), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12262 ( .A1(n9824), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12263 ( .A1(n9824), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12264 ( .A1(n9824), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12265 ( .A1(n9824), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  NAND2_X1 U12266 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10486) );
  AOI211_X1 U12267 ( .C1(n9827), .C2(n9826), .A(n9825), .B(n14668), .ZN(n9828)
         );
  INV_X1 U12268 ( .A(n9828), .ZN(n9829) );
  NAND2_X1 U12269 ( .A1(n10486), .A2(n9829), .ZN(n9837) );
  INV_X1 U12270 ( .A(n9830), .ZN(n9835) );
  NOR3_X1 U12271 ( .A1(n9833), .A2(n9832), .A3(n9831), .ZN(n9834) );
  NOR3_X1 U12272 ( .A1(n14670), .A2(n9835), .A3(n9834), .ZN(n9836) );
  AOI211_X1 U12273 ( .C1(n14652), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9837), .B(
        n9836), .ZN(n9838) );
  OAI21_X1 U12274 ( .B1(n9839), .B2(n14644), .A(n9838), .ZN(P2_U3219) );
  OAI21_X1 U12275 ( .B1(n14760), .B2(n9841), .A(n9840), .ZN(n14636) );
  MUX2_X1 U12276 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9842), .S(n9850), .Z(n14635) );
  NAND2_X1 U12277 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  NAND2_X1 U12278 ( .A1(n9850), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U12279 ( .A(n8620), .B(P2_REG1_REG_8__SCAN_IN), .S(n9876), .Z(n9843)
         );
  AOI21_X1 U12280 ( .B1(n14634), .B2(n9844), .A(n9843), .ZN(n9874) );
  NAND3_X1 U12281 ( .A1(n14634), .A2(n9844), .A3(n9843), .ZN(n9845) );
  NAND2_X1 U12282 ( .A1(n9845), .A2(n14658), .ZN(n9857) );
  INV_X1 U12283 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U12284 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10786) );
  OAI21_X1 U12285 ( .B1(n14677), .B2(n9846), .A(n10786), .ZN(n9855) );
  AOI21_X1 U12286 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9848), .A(n9847), .ZN(
        n14631) );
  INV_X1 U12287 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9849) );
  MUX2_X1 U12288 ( .A(n9849), .B(P2_REG2_REG_7__SCAN_IN), .S(n9850), .Z(n14630) );
  OR2_X1 U12289 ( .A1(n14631), .A2(n14630), .ZN(n14632) );
  NAND2_X1 U12290 ( .A1(n9850), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9852) );
  MUX2_X1 U12291 ( .A(n11482), .B(P2_REG2_REG_8__SCAN_IN), .S(n9876), .Z(n9851) );
  AND3_X1 U12292 ( .A1(n14632), .A2(n9852), .A3(n9851), .ZN(n9853) );
  NOR3_X1 U12293 ( .A1(n9875), .A2(n9853), .A3(n14670), .ZN(n9854) );
  AOI211_X1 U12294 ( .C1(n14673), .C2(n9876), .A(n9855), .B(n9854), .ZN(n9856)
         );
  OAI21_X1 U12295 ( .B1(n9874), .B2(n9857), .A(n9856), .ZN(P2_U3222) );
  INV_X1 U12296 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U12297 ( .A1(n14677), .A2(n9858), .ZN(n9865) );
  INV_X1 U12298 ( .A(n9859), .ZN(n9863) );
  NOR3_X1 U12299 ( .A1(n14619), .A2(n9861), .A3(n9860), .ZN(n9862) );
  NOR3_X1 U12300 ( .A1(n14670), .A2(n9863), .A3(n9862), .ZN(n9864) );
  AOI211_X1 U12301 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n9865), 
        .B(n9864), .ZN(n9872) );
  INV_X1 U12302 ( .A(n9866), .ZN(n9870) );
  NAND3_X1 U12303 ( .A1(n14616), .A2(n9868), .A3(n9867), .ZN(n9869) );
  NAND3_X1 U12304 ( .A1(n14658), .A2(n9870), .A3(n9869), .ZN(n9871) );
  OAI211_X1 U12305 ( .C1(n14644), .C2(n9873), .A(n9872), .B(n9871), .ZN(
        P2_U3217) );
  AOI21_X1 U12306 ( .B1(n9876), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9874), .ZN(
        n9885) );
  NOR3_X1 U12307 ( .A1(n9885), .A2(n8639), .A3(n14668), .ZN(n9878) );
  AOI21_X1 U12308 ( .B1(n9876), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9875), .ZN(
        n9881) );
  NOR3_X1 U12309 ( .A1(n9881), .A2(n11338), .A3(n14670), .ZN(n9877) );
  NOR3_X1 U12310 ( .A1(n9878), .A2(n9877), .A3(n14673), .ZN(n9889) );
  NAND2_X1 U12311 ( .A1(n10132), .A2(n11338), .ZN(n9880) );
  MUX2_X1 U12312 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11338), .S(n10127), .Z(
        n9879) );
  NAND2_X1 U12313 ( .A1(n9881), .A2(n9879), .ZN(n10126) );
  OAI21_X1 U12314 ( .B1(n9881), .B2(n9880), .A(n10126), .ZN(n9883) );
  NAND2_X1 U12315 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10878) );
  OAI21_X1 U12316 ( .B1(n14677), .B2(n14150), .A(n10878), .ZN(n9882) );
  AOI21_X1 U12317 ( .B1(n9883), .B2(n14655), .A(n9882), .ZN(n9888) );
  NOR3_X1 U12318 ( .A1(n9885), .A2(n10127), .A3(P2_REG1_REG_9__SCAN_IN), .ZN(
        n9886) );
  MUX2_X1 U12319 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8639), .S(n10127), .Z(n9884) );
  AND2_X1 U12320 ( .A1(n9885), .A2(n9884), .ZN(n10131) );
  OAI21_X1 U12321 ( .B1(n9886), .B2(n10131), .A(n14658), .ZN(n9887) );
  OAI211_X1 U12322 ( .C1(n9889), .C2(n10132), .A(n9888), .B(n9887), .ZN(
        P2_U3223) );
  INV_X1 U12323 ( .A(n9890), .ZN(n9892) );
  INV_X1 U12324 ( .A(n9969), .ZN(n9981) );
  OAI222_X1 U12325 ( .A1(n14125), .A2(n9891), .B1(n14128), .B2(n9892), .C1(
        P1_U3086), .C2(n9981), .ZN(P1_U3345) );
  INV_X1 U12326 ( .A(n10171), .ZN(n10140) );
  OAI222_X1 U12327 ( .A1(n13578), .A2(n9893), .B1(n13581), .B2(n9892), .C1(
        P2_U3088), .C2(n10140), .ZN(P2_U3317) );
  NAND2_X1 U12328 ( .A1(n7082), .A2(n11622), .ZN(n9919) );
  INV_X1 U12329 ( .A(n10295), .ZN(n9895) );
  NAND2_X1 U12330 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  NAND2_X1 U12331 ( .A1(n9897), .A2(n9896), .ZN(n9917) );
  NAND2_X1 U12332 ( .A1(n9919), .A2(n9917), .ZN(n14384) );
  INV_X1 U12333 ( .A(n14384), .ZN(n13787) );
  CLKBUF_X2 U12334 ( .A(P1_U4016), .Z(n13689) );
  NOR2_X1 U12335 ( .A1(n13787), .A2(n13689), .ZN(P1_U3085) );
  INV_X1 U12336 ( .A(n12674), .ZN(n12667) );
  OAI222_X1 U12337 ( .A1(n13056), .A2(n9899), .B1(n13058), .B2(n9898), .C1(
        n12667), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12338 ( .A(n9900), .ZN(n9902) );
  INV_X1 U12339 ( .A(n10172), .ZN(n10449) );
  OAI222_X1 U12340 ( .A1(n13578), .A2(n9901), .B1(n13581), .B2(n9902), .C1(
        P2_U3088), .C2(n10449), .ZN(P2_U3316) );
  INV_X1 U12341 ( .A(n10150), .ZN(n10142) );
  OAI222_X1 U12342 ( .A1(n9903), .A2(n14125), .B1(P1_U3086), .B2(n10142), .C1(
        n14128), .C2(n9902), .ZN(P1_U3344) );
  MUX2_X1 U12343 ( .A(n7963), .B(P1_REG1_REG_8__SCAN_IN), .S(n9954), .Z(n9916)
         );
  INV_X1 U12344 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14581) );
  MUX2_X1 U12345 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14581), .S(n10357), .Z(
        n10352) );
  INV_X1 U12346 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14579) );
  MUX2_X1 U12347 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14579), .S(n13693), .Z(
        n13699) );
  AND2_X1 U12348 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13698) );
  NAND2_X1 U12349 ( .A1(n13699), .A2(n13698), .ZN(n13697) );
  NAND2_X1 U12350 ( .A1(n13693), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12351 ( .A1(n13697), .A2(n9904), .ZN(n10351) );
  NAND2_X1 U12352 ( .A1(n10352), .A2(n10351), .ZN(n10350) );
  NAND2_X1 U12353 ( .A1(n10357), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U12354 ( .A1(n10350), .A2(n9905), .ZN(n13708) );
  INV_X1 U12355 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14583) );
  MUX2_X1 U12356 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n14583), .S(n13711), .Z(
        n13709) );
  NAND2_X1 U12357 ( .A1(n13708), .A2(n13709), .ZN(n13707) );
  NAND2_X1 U12358 ( .A1(n13711), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U12359 ( .A1(n13707), .A2(n9906), .ZN(n13721) );
  MUX2_X1 U12360 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7890), .S(n13719), .Z(
        n13722) );
  NAND2_X1 U12361 ( .A1(n13721), .A2(n13722), .ZN(n13720) );
  NAND2_X1 U12362 ( .A1(n13719), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U12363 ( .A1(n13720), .A2(n9907), .ZN(n9944) );
  XNOR2_X1 U12364 ( .A(n9946), .B(n9908), .ZN(n9945) );
  OR2_X1 U12365 ( .A1(n9944), .A2(n9945), .ZN(n9942) );
  NAND2_X1 U12366 ( .A1(n9946), .A2(n9908), .ZN(n9909) );
  AND2_X1 U12367 ( .A1(n9942), .A2(n9909), .ZN(n13743) );
  INV_X1 U12368 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9910) );
  XNOR2_X1 U12369 ( .A(n9931), .B(n9910), .ZN(n13744) );
  NAND2_X1 U12370 ( .A1(n13743), .A2(n13744), .ZN(n13742) );
  NAND2_X1 U12371 ( .A1(n9931), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9911) );
  NAND2_X1 U12372 ( .A1(n13742), .A2(n9911), .ZN(n13752) );
  INV_X1 U12373 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9912) );
  XNOR2_X1 U12374 ( .A(n9934), .B(n9912), .ZN(n13753) );
  NAND2_X1 U12375 ( .A1(n13752), .A2(n13753), .ZN(n13751) );
  NAND2_X1 U12376 ( .A1(n9934), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U12377 ( .A1(n13751), .A2(n9913), .ZN(n9915) );
  OR2_X1 U12378 ( .A1(n9915), .A2(n9916), .ZN(n9956) );
  INV_X1 U12379 ( .A(n9956), .ZN(n9914) );
  AOI21_X1 U12380 ( .B1(n9916), .B2(n9915), .A(n9914), .ZN(n9941) );
  INV_X1 U12381 ( .A(n9917), .ZN(n9918) );
  NAND2_X1 U12382 ( .A1(n9919), .A2(n9918), .ZN(n10074) );
  INV_X1 U12383 ( .A(n10074), .ZN(n9920) );
  AND2_X1 U12384 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11553) );
  INV_X1 U12385 ( .A(n11928), .ZN(n10294) );
  NOR2_X1 U12386 ( .A1(n14380), .A2(n9966), .ZN(n9921) );
  AOI211_X1 U12387 ( .C1(n13787), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11553), .B(
        n9921), .ZN(n9940) );
  INV_X1 U12388 ( .A(n14122), .ZN(n10358) );
  NAND2_X1 U12389 ( .A1(n10294), .A2(n10358), .ZN(n9922) );
  OR2_X1 U12390 ( .A1(n10074), .A2(n9922), .ZN(n14370) );
  INV_X1 U12391 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9923) );
  MUX2_X1 U12392 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9923), .S(n10357), .Z(
        n10349) );
  INV_X1 U12393 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9924) );
  MUX2_X1 U12394 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9924), .S(n13693), .Z(
        n13696) );
  AND2_X1 U12395 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9925) );
  NAND2_X1 U12396 ( .A1(n13696), .A2(n9925), .ZN(n13695) );
  NAND2_X1 U12397 ( .A1(n13693), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12398 ( .A1(n13695), .A2(n9926), .ZN(n10348) );
  AOI22_X1 U12399 ( .A1(n10349), .A2(n10348), .B1(n10357), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n13704) );
  MUX2_X1 U12400 ( .A(n13703), .B(P1_REG2_REG_3__SCAN_IN), .S(n13711), .Z(
        n9927) );
  OR2_X1 U12401 ( .A1(n13704), .A2(n9927), .ZN(n13726) );
  NAND2_X1 U12402 ( .A1(n13711), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13725) );
  MUX2_X1 U12403 ( .A(n7888), .B(P1_REG2_REG_4__SCAN_IN), .S(n13719), .Z(
        n13724) );
  AOI21_X1 U12404 ( .B1(n13726), .B2(n13725), .A(n13724), .ZN(n13723) );
  NOR2_X1 U12405 ( .A1(n9928), .A2(n7888), .ZN(n9948) );
  MUX2_X1 U12406 ( .A(n9929), .B(P1_REG2_REG_5__SCAN_IN), .S(n9946), .Z(n9949)
         );
  OAI21_X1 U12407 ( .B1(n13723), .B2(n9948), .A(n9949), .ZN(n13739) );
  NAND2_X1 U12408 ( .A1(n9930), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13738) );
  INV_X1 U12409 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9932) );
  MUX2_X1 U12410 ( .A(n9932), .B(P1_REG2_REG_6__SCAN_IN), .S(n9931), .Z(n13737) );
  AOI21_X1 U12411 ( .B1(n13739), .B2(n13738), .A(n13737), .ZN(n13756) );
  NOR2_X1 U12412 ( .A1(n13734), .A2(n9932), .ZN(n13755) );
  MUX2_X1 U12413 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9933), .S(n9934), .Z(n13754) );
  OAI21_X1 U12414 ( .B1(n13756), .B2(n13755), .A(n13754), .ZN(n13758) );
  NAND2_X1 U12415 ( .A1(n9934), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9936) );
  INV_X1 U12416 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9965) );
  MUX2_X1 U12417 ( .A(n9965), .B(P1_REG2_REG_8__SCAN_IN), .S(n9954), .Z(n9935)
         );
  AOI21_X1 U12418 ( .B1(n13758), .B2(n9936), .A(n9935), .ZN(n10002) );
  INV_X1 U12419 ( .A(n10002), .ZN(n9938) );
  NAND3_X1 U12420 ( .A1(n13758), .A2(n9936), .A3(n9935), .ZN(n9937) );
  NAND3_X1 U12421 ( .A1(n13811), .A2(n9938), .A3(n9937), .ZN(n9939) );
  OAI211_X1 U12422 ( .C1(n9941), .C2(n13767), .A(n9940), .B(n9939), .ZN(
        P1_U3251) );
  INV_X1 U12423 ( .A(n9942), .ZN(n9943) );
  AOI21_X1 U12424 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9953) );
  AND2_X1 U12425 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10815) );
  NOR2_X1 U12426 ( .A1(n14380), .A2(n9946), .ZN(n9947) );
  AOI211_X1 U12427 ( .C1(n13787), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10815), .B(
        n9947), .ZN(n9952) );
  OR3_X1 U12428 ( .A1(n13723), .A2(n9949), .A3(n9948), .ZN(n9950) );
  NAND3_X1 U12429 ( .A1(n13811), .A2(n13739), .A3(n9950), .ZN(n9951) );
  OAI211_X1 U12430 ( .C1(n9953), .C2(n13767), .A(n9952), .B(n9951), .ZN(
        P1_U3248) );
  MUX2_X1 U12431 ( .A(n8027), .B(P1_REG1_REG_11__SCAN_IN), .S(n10150), .Z(
        n9962) );
  OR2_X1 U12432 ( .A1(n9954), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U12433 ( .A1(n9956), .A2(n9955), .ZN(n9994) );
  MUX2_X1 U12434 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9957), .S(n9968), .Z(n9995)
         );
  NAND2_X1 U12435 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  NAND2_X1 U12436 ( .A1(n9998), .A2(n9957), .ZN(n9958) );
  AND2_X1 U12437 ( .A1(n9993), .A2(n9958), .ZN(n9986) );
  INV_X1 U12438 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14592) );
  MUX2_X1 U12439 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14592), .S(n9969), .Z(
        n9985) );
  NAND2_X1 U12440 ( .A1(n9986), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U12441 ( .A1(n9969), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U12442 ( .A1(n9984), .A2(n9959), .ZN(n9961) );
  OR2_X1 U12443 ( .A1(n9961), .A2(n9962), .ZN(n10152) );
  INV_X1 U12444 ( .A(n10152), .ZN(n9960) );
  AOI21_X1 U12445 ( .B1(n9962), .B2(n9961), .A(n9960), .ZN(n9976) );
  NAND2_X1 U12446 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14279)
         );
  INV_X1 U12447 ( .A(n14279), .ZN(n9964) );
  NOR2_X1 U12448 ( .A1(n14380), .A2(n10142), .ZN(n9963) );
  AOI211_X1 U12449 ( .C1(n13787), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9964), .B(
        n9963), .ZN(n9975) );
  NOR2_X1 U12450 ( .A1(n9966), .A2(n9965), .ZN(n10001) );
  MUX2_X1 U12451 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9967), .S(n9968), .Z(n10000) );
  OAI21_X1 U12452 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n9999) );
  NAND2_X1 U12453 ( .A1(n9968), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9978) );
  INV_X1 U12454 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U12455 ( .A(n9970), .B(P1_REG2_REG_10__SCAN_IN), .S(n9969), .Z(n9977) );
  AOI21_X1 U12456 ( .B1(n9999), .B2(n9978), .A(n9977), .ZN(n9990) );
  NOR2_X1 U12457 ( .A1(n9981), .A2(n9970), .ZN(n9972) );
  INV_X1 U12458 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11010) );
  MUX2_X1 U12459 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11010), .S(n10150), .Z(
        n9971) );
  OAI21_X1 U12460 ( .B1(n9990), .B2(n9972), .A(n9971), .ZN(n10141) );
  OR3_X1 U12461 ( .A1(n9990), .A2(n9972), .A3(n9971), .ZN(n9973) );
  NAND3_X1 U12462 ( .A1(n10141), .A2(n13811), .A3(n9973), .ZN(n9974) );
  OAI211_X1 U12463 ( .C1(n9976), .C2(n13767), .A(n9975), .B(n9974), .ZN(
        P1_U3254) );
  NAND3_X1 U12464 ( .A1(n9999), .A2(n9978), .A3(n9977), .ZN(n9979) );
  NAND2_X1 U12465 ( .A1(n9979), .A2(n13811), .ZN(n9989) );
  NOR2_X1 U12466 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9980), .ZN(n9983) );
  NOR2_X1 U12467 ( .A1(n14380), .A2(n9981), .ZN(n9982) );
  AOI211_X1 U12468 ( .C1(n13787), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n9983), .B(
        n9982), .ZN(n9988) );
  OAI211_X1 U12469 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n14375), .ZN(n9987)
         );
  OAI211_X1 U12470 ( .C1(n9990), .C2(n9989), .A(n9988), .B(n9987), .ZN(
        P1_U3253) );
  INV_X1 U12471 ( .A(n12682), .ZN(n12706) );
  OAI222_X1 U12472 ( .A1(n13056), .A2(n9992), .B1(n12706), .B2(P3_U3151), .C1(
        n9991), .C2(n13058), .ZN(P3_U3279) );
  OAI21_X1 U12473 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n10007) );
  NAND2_X1 U12474 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11403) );
  INV_X1 U12475 ( .A(n11403), .ZN(n9996) );
  AOI21_X1 U12476 ( .B1(n13787), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9996), .ZN(
        n9997) );
  OAI21_X1 U12477 ( .B1(n9998), .B2(n14380), .A(n9997), .ZN(n10006) );
  INV_X1 U12478 ( .A(n9999), .ZN(n10004) );
  NOR3_X1 U12479 ( .A1(n10002), .A2(n10001), .A3(n10000), .ZN(n10003) );
  NOR3_X1 U12480 ( .A1(n10004), .A2(n10003), .A3(n14370), .ZN(n10005) );
  AOI211_X1 U12481 ( .C1(n14375), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10008) );
  INV_X1 U12482 ( .A(n10008), .ZN(P1_U3252) );
  NOR2_X1 U12483 ( .A1(n10342), .A2(n14772), .ZN(n10009) );
  NAND2_X1 U12484 ( .A1(n9131), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10010) );
  AOI21_X1 U12485 ( .B1(n10020), .B2(n10011), .A(n10042), .ZN(n10040) );
  OR2_X1 U12486 ( .A1(n10079), .A2(P3_U3151), .ZN(n12597) );
  INV_X1 U12487 ( .A(n12597), .ZN(n10012) );
  AOI21_X1 U12488 ( .B1(n12525), .B2(n10079), .A(n10013), .ZN(n10016) );
  INV_X1 U12489 ( .A(n10014), .ZN(n10015) );
  INV_X1 U12490 ( .A(n10016), .ZN(n10017) );
  AND2_X1 U12491 ( .A1(P3_U3897), .A2(n11925), .ZN(n14892) );
  INV_X1 U12492 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10019) );
  MUX2_X1 U12493 ( .A(n10342), .B(n10019), .S(n12729), .Z(n14771) );
  NAND2_X1 U12494 ( .A1(n14771), .A2(n14772), .ZN(n14770) );
  INV_X1 U12495 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U12496 ( .A(n10020), .B(n10031), .S(n12729), .Z(n10021) );
  INV_X1 U12497 ( .A(n10028), .ZN(n10037) );
  NAND2_X1 U12498 ( .A1(n10021), .A2(n10037), .ZN(n10053) );
  INV_X1 U12499 ( .A(n10021), .ZN(n10022) );
  NAND2_X1 U12500 ( .A1(n10022), .A2(n10028), .ZN(n10023) );
  NAND2_X1 U12501 ( .A1(n10053), .A2(n10023), .ZN(n10025) );
  OR2_X1 U12502 ( .A1(n10025), .A2(n14770), .ZN(n10052) );
  INV_X1 U12503 ( .A(n10052), .ZN(n10024) );
  AOI21_X1 U12504 ( .B1(n14770), .B2(n10025), .A(n10024), .ZN(n10026) );
  OAI22_X1 U12505 ( .A1(n14915), .A2(n10026), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n7577), .ZN(n10034) );
  NAND2_X1 U12506 ( .A1(n10035), .A2(n12729), .ZN(n14769) );
  NOR3_X1 U12507 ( .A1(n10019), .A2(P3_IR_REG_1__SCAN_IN), .A3(n14772), .ZN(
        n10058) );
  AND2_X1 U12508 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n14776), .ZN(n10027) );
  NOR2_X1 U12509 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  OR2_X1 U12510 ( .A1(n10058), .A2(n10029), .ZN(n10030) );
  AOI21_X1 U12511 ( .B1(n10031), .B2(n10030), .A(n10057), .ZN(n10032) );
  NOR2_X1 U12512 ( .A1(n14769), .A2(n10032), .ZN(n10033) );
  AOI211_X1 U12513 ( .C1(n14899), .C2(P3_ADDR_REG_1__SCAN_IN), .A(n10034), .B(
        n10033), .ZN(n10039) );
  INV_X1 U12514 ( .A(n10035), .ZN(n10036) );
  INV_X1 U12515 ( .A(P3_U3897), .ZN(n12603) );
  MUX2_X1 U12516 ( .A(n10036), .B(n12603), .S(n12592), .Z(n14896) );
  NAND2_X1 U12517 ( .A1(n14926), .A2(n10037), .ZN(n10038) );
  OAI211_X1 U12518 ( .C1(n10040), .C2(n14921), .A(n10039), .B(n10038), .ZN(
        P3_U3183) );
  INV_X1 U12519 ( .A(n14921), .ZN(n12702) );
  XNOR2_X1 U12520 ( .A(n10056), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10044) );
  AND2_X1 U12521 ( .A1(n9131), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U12522 ( .A1(n10043), .A2(n10044), .ZN(n11137) );
  OAI21_X1 U12523 ( .B1(n10044), .B2(n10043), .A(n11137), .ZN(n10065) );
  NAND2_X1 U12524 ( .A1(n10052), .A2(n10053), .ZN(n10050) );
  INV_X1 U12525 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10045) );
  MUX2_X1 U12526 ( .A(n10046), .B(n10045), .S(n12729), .Z(n10047) );
  NAND2_X1 U12527 ( .A1(n10047), .A2(n10056), .ZN(n14787) );
  INV_X1 U12528 ( .A(n10047), .ZN(n10048) );
  NAND2_X1 U12529 ( .A1(n10048), .A2(n11152), .ZN(n10049) );
  AND2_X1 U12530 ( .A1(n14787), .A2(n10049), .ZN(n10051) );
  NAND2_X1 U12531 ( .A1(n10050), .A2(n10051), .ZN(n14788) );
  INV_X1 U12532 ( .A(n10051), .ZN(n10054) );
  NAND3_X1 U12533 ( .A1(n10054), .A2(n10053), .A3(n10052), .ZN(n10055) );
  AOI21_X1 U12534 ( .B1(n14788), .B2(n10055), .A(n14915), .ZN(n10064) );
  MUX2_X1 U12535 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10045), .S(n10056), .Z(
        n10060) );
  AOI21_X1 U12536 ( .B1(n10060), .B2(n10059), .A(n11151), .ZN(n10062) );
  AOI22_X1 U12537 ( .A1(n14899), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10061) );
  OAI21_X1 U12538 ( .B1(n10062), .B2(n14769), .A(n10061), .ZN(n10063) );
  AOI211_X1 U12539 ( .C1(n12702), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10066) );
  OAI21_X1 U12540 ( .B1(n11152), .B2(n14896), .A(n10066), .ZN(P3_U3184) );
  INV_X1 U12541 ( .A(n10067), .ZN(n10220) );
  INV_X1 U12542 ( .A(n14125), .ZN(n14114) );
  AOI22_X1 U12543 ( .A1(n10387), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14114), .ZN(n10068) );
  OAI21_X1 U12544 ( .B1(n10220), .B2(n14128), .A(n10068), .ZN(P1_U3343) );
  INV_X1 U12545 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12546 ( .A1(n10358), .A2(n10069), .ZN(n10070) );
  NAND2_X1 U12547 ( .A1(n10294), .A2(n10070), .ZN(n10361) );
  INV_X1 U12548 ( .A(n10361), .ZN(n10071) );
  OAI21_X1 U12549 ( .B1(n10358), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10071), .ZN(
        n10072) );
  MUX2_X1 U12550 ( .A(n10072), .B(n10071), .S(P1_IR_REG_0__SCAN_IN), .Z(n10073) );
  INV_X1 U12551 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10643) );
  OAI22_X1 U12552 ( .A1(n10074), .A2(n10073), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10643), .ZN(n10076) );
  NOR3_X1 U12553 ( .A1(n13767), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10360), .ZN(
        n10075) );
  AOI211_X1 U12554 ( .C1(n13787), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10076), .B(
        n10075), .ZN(n10077) );
  INV_X1 U12555 ( .A(n10077), .ZN(P1_U3243) );
  INV_X1 U12556 ( .A(n10106), .ZN(n10083) );
  INV_X1 U12557 ( .A(n10110), .ZN(n10086) );
  NAND2_X1 U12558 ( .A1(n10086), .A2(n10078), .ZN(n10082) );
  AND3_X1 U12559 ( .A1(n10334), .A2(n10080), .A3(n10079), .ZN(n10081) );
  OAI211_X1 U12560 ( .C1(n10113), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10084) );
  NAND2_X1 U12561 ( .A1(n10084), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10088) );
  INV_X1 U12562 ( .A(n10085), .ZN(n12593) );
  NAND2_X1 U12563 ( .A1(n10086), .A2(n12593), .ZN(n10087) );
  NOR2_X1 U12564 ( .A1(n12383), .A2(P3_U3151), .ZN(n10161) );
  INV_X1 U12565 ( .A(n12588), .ZN(n10089) );
  NAND2_X1 U12566 ( .A1(n12393), .A2(n12723), .ZN(n10090) );
  NAND2_X1 U12567 ( .A1(n10090), .A2(n10725), .ZN(n10091) );
  NAND2_X2 U12568 ( .A1(n10092), .A2(n10091), .ZN(n10097) );
  XNOR2_X1 U12569 ( .A(n10097), .B(n10093), .ZN(n10306) );
  XNOR2_X1 U12570 ( .A(n14964), .B(n10306), .ZN(n10103) );
  INV_X1 U12571 ( .A(n10094), .ZN(n10095) );
  OAI21_X1 U12572 ( .B1(n10095), .B2(n14993), .A(n10097), .ZN(n10099) );
  NOR3_X1 U12573 ( .A1(n9118), .A2(n10097), .A3(n14992), .ZN(n10098) );
  INV_X1 U12574 ( .A(n10100), .ZN(n10101) );
  NAND2_X1 U12575 ( .A1(n10121), .A2(n10101), .ZN(n10102) );
  NAND2_X1 U12576 ( .A1(n10102), .A2(n10103), .ZN(n10309) );
  OAI21_X1 U12577 ( .B1(n10103), .B2(n10102), .A(n10309), .ZN(n10109) );
  INV_X1 U12578 ( .A(n10104), .ZN(n10105) );
  NAND2_X1 U12579 ( .A1(n10105), .A2(n10110), .ZN(n10108) );
  NAND4_X1 U12580 ( .A1(n10113), .A2(n10337), .A3(n15047), .A4(n10106), .ZN(
        n10107) );
  NAND2_X1 U12581 ( .A1(n10109), .A2(n12376), .ZN(n10118) );
  AND2_X1 U12582 ( .A1(n10337), .A2(n15015), .ZN(n10112) );
  OAI21_X2 U12583 ( .B1(n10113), .B2(n14979), .A(n10112), .ZN(n12386) );
  OAI22_X1 U12584 ( .A1(n12386), .A2(n14977), .B1(n12380), .B2(n14983), .ZN(
        n10116) );
  AOI21_X1 U12585 ( .B1(n12355), .B2(n12612), .A(n10116), .ZN(n10117) );
  OAI211_X1 U12586 ( .C1(n10161), .C2(n7575), .A(n10118), .B(n10117), .ZN(
        P3_U3177) );
  NAND3_X1 U12587 ( .A1(n10119), .A2(n10097), .A3(n14993), .ZN(n10120) );
  OAI211_X1 U12588 ( .C1(n10122), .C2(n14995), .A(n10121), .B(n10120), .ZN(
        n10123) );
  NAND2_X1 U12589 ( .A1(n10123), .A2(n12376), .ZN(n10125) );
  OAI22_X1 U12590 ( .A1(n14992), .A2(n12386), .B1(n12380), .B2(n14997), .ZN(
        n10124) );
  OAI211_X1 U12591 ( .C1(n10161), .C2(n7577), .A(n10125), .B(n6603), .ZN(
        P3_U3162) );
  OAI21_X1 U12592 ( .B1(n10127), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10126), .ZN(
        n10129) );
  MUX2_X1 U12593 ( .A(n11502), .B(P2_REG2_REG_10__SCAN_IN), .S(n10171), .Z(
        n10128) );
  AOI211_X1 U12594 ( .C1(n10129), .C2(n10128), .A(n14670), .B(n10162), .ZN(
        n10130) );
  INV_X1 U12595 ( .A(n10130), .ZN(n10139) );
  NAND2_X1 U12596 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10891)
         );
  AOI21_X1 U12597 ( .B1(n8639), .B2(n10132), .A(n10131), .ZN(n10135) );
  MUX2_X1 U12598 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10133), .S(n10171), .Z(
        n10134) );
  NAND2_X1 U12599 ( .A1(n10135), .A2(n10134), .ZN(n10175) );
  OAI211_X1 U12600 ( .C1(n10135), .C2(n10134), .A(n14658), .B(n10175), .ZN(
        n10136) );
  NAND2_X1 U12601 ( .A1(n10891), .A2(n10136), .ZN(n10137) );
  AOI21_X1 U12602 ( .B1(n14652), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10137), 
        .ZN(n10138) );
  OAI211_X1 U12603 ( .C1(n14644), .C2(n10140), .A(n10139), .B(n10138), .ZN(
        P2_U3224) );
  OAI21_X1 U12604 ( .B1(n10142), .B2(n11010), .A(n10141), .ZN(n10146) );
  INV_X1 U12605 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10143) );
  MUX2_X1 U12606 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10143), .S(n10387), .Z(
        n10144) );
  INV_X1 U12607 ( .A(n10144), .ZN(n10145) );
  NOR2_X1 U12608 ( .A1(n10145), .A2(n10146), .ZN(n10385) );
  AOI21_X1 U12609 ( .B1(n10146), .B2(n10145), .A(n10385), .ZN(n10158) );
  AND2_X1 U12610 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11709) );
  INV_X1 U12611 ( .A(n10387), .ZN(n10147) );
  NOR2_X1 U12612 ( .A1(n14380), .A2(n10147), .ZN(n10148) );
  AOI211_X1 U12613 ( .C1(n13787), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n11709), 
        .B(n10148), .ZN(n10157) );
  MUX2_X1 U12614 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10149), .S(n10387), .Z(
        n10154) );
  OR2_X1 U12615 ( .A1(n10150), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U12616 ( .A1(n10152), .A2(n10151), .ZN(n10153) );
  NAND2_X1 U12617 ( .A1(n10153), .A2(n10154), .ZN(n10380) );
  OAI21_X1 U12618 ( .B1(n10154), .B2(n10153), .A(n10380), .ZN(n10155) );
  NAND2_X1 U12619 ( .A1(n10155), .A2(n14375), .ZN(n10156) );
  OAI211_X1 U12620 ( .C1(n10158), .C2(n14370), .A(n10157), .B(n10156), .ZN(
        P1_U3255) );
  INV_X1 U12621 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14775) );
  INV_X1 U12622 ( .A(n12380), .ZN(n12365) );
  INV_X1 U12623 ( .A(n15014), .ZN(n10344) );
  AND2_X1 U12624 ( .A1(n14993), .A2(n12389), .ZN(n12564) );
  OAI22_X1 U12625 ( .A1(n12371), .A2(n12564), .B1(n12386), .B2(n10344), .ZN(
        n10159) );
  AOI21_X1 U12626 ( .B1(n12365), .B2(n12612), .A(n10159), .ZN(n10160) );
  OAI21_X1 U12627 ( .B1(n10161), .B2(n14775), .A(n10160), .ZN(P3_U3172) );
  AOI21_X1 U12628 ( .B1(n10171), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10162), 
        .ZN(n10165) );
  INV_X1 U12629 ( .A(n10165), .ZN(n10168) );
  INV_X1 U12630 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10163) );
  MUX2_X1 U12631 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10163), .S(n10172), .Z(
        n10164) );
  INV_X1 U12632 ( .A(n10164), .ZN(n10167) );
  NAND2_X1 U12633 ( .A1(n10165), .A2(n10164), .ZN(n10452) );
  INV_X1 U12634 ( .A(n10452), .ZN(n10166) );
  AOI21_X1 U12635 ( .B1(n10168), .B2(n10167), .A(n10166), .ZN(n10180) );
  NOR2_X1 U12636 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11107), .ZN(n10170) );
  NOR2_X1 U12637 ( .A1(n14644), .A2(n10449), .ZN(n10169) );
  AOI211_X1 U12638 ( .C1(n14652), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10170), 
        .B(n10169), .ZN(n10179) );
  NAND2_X1 U12639 ( .A1(n10171), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10174) );
  MUX2_X1 U12640 ( .A(n8673), .B(P2_REG1_REG_11__SCAN_IN), .S(n10172), .Z(
        n10173) );
  AOI21_X1 U12641 ( .B1(n10175), .B2(n10174), .A(n10173), .ZN(n10444) );
  INV_X1 U12642 ( .A(n10444), .ZN(n10177) );
  NAND3_X1 U12643 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10176) );
  NAND3_X1 U12644 ( .A1(n10177), .A2(n14658), .A3(n10176), .ZN(n10178) );
  OAI211_X1 U12645 ( .C1(n10180), .C2(n14670), .A(n10179), .B(n10178), .ZN(
        P2_U3225) );
  XNOR2_X1 U12646 ( .A(n11837), .B(P2_B_REG_SCAN_IN), .ZN(n10182) );
  INV_X1 U12647 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U12648 ( .A1(n14679), .A2(n14684), .ZN(n10184) );
  NAND2_X1 U12649 ( .A1(n13582), .A2(n11881), .ZN(n10183) );
  NAND2_X1 U12650 ( .A1(n10184), .A2(n10183), .ZN(n14685) );
  NOR2_X1 U12651 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10188) );
  NOR4_X1 U12652 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10187) );
  NOR4_X1 U12653 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n10186) );
  NOR4_X1 U12654 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n10185) );
  AND4_X1 U12655 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10194) );
  NOR4_X1 U12656 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n10192) );
  NOR4_X1 U12657 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n10191) );
  NOR4_X1 U12658 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10190) );
  NOR4_X1 U12659 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n10189) );
  AND4_X1 U12660 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  NAND2_X1 U12661 ( .A1(n10194), .A2(n10193), .ZN(n10195) );
  AND2_X1 U12662 ( .A1(n14679), .A2(n10195), .ZN(n10222) );
  INV_X1 U12663 ( .A(n10222), .ZN(n10196) );
  NAND3_X1 U12664 ( .A1(n10238), .A2(n14685), .A3(n10196), .ZN(n10653) );
  INV_X1 U12665 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14682) );
  AND2_X1 U12666 ( .A1(n11837), .A2(n13582), .ZN(n10197) );
  AOI21_X1 U12667 ( .B1(n14679), .B2(n14682), .A(n10197), .ZN(n10227) );
  INV_X1 U12668 ( .A(n10227), .ZN(n10223) );
  NAND2_X1 U12669 ( .A1(n10232), .A2(n10228), .ZN(n10651) );
  NAND3_X1 U12670 ( .A1(n10223), .A2(n14686), .A3(n10651), .ZN(n10821) );
  INV_X1 U12671 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U12672 ( .A1(n10656), .A2(n10200), .ZN(n13419) );
  INV_X1 U12673 ( .A(n13419), .ZN(n10217) );
  XNOR2_X1 U12674 ( .A(n10244), .B(n8487), .ZN(n10201) );
  INV_X1 U12675 ( .A(n10245), .ZN(n14745) );
  NAND2_X1 U12676 ( .A1(n13419), .A2(n14745), .ZN(n10213) );
  NOR2_X1 U12677 ( .A1(n9020), .A2(n8489), .ZN(n10204) );
  NAND2_X1 U12678 ( .A1(n10202), .A2(n10205), .ZN(n10207) );
  NAND2_X1 U12679 ( .A1(n10208), .A2(n13541), .ZN(n10212) );
  NAND2_X1 U12680 ( .A1(n9020), .A2(n13141), .ZN(n10211) );
  NAND2_X1 U12681 ( .A1(n10209), .A2(n10228), .ZN(n13161) );
  INV_X1 U12682 ( .A(n13161), .ZN(n13139) );
  NAND2_X1 U12683 ( .A1(n13198), .A2(n13139), .ZN(n10210) );
  AND2_X1 U12684 ( .A1(n10211), .A2(n10210), .ZN(n10459) );
  AND3_X1 U12685 ( .A1(n10213), .A2(n10212), .A3(n10459), .ZN(n13413) );
  NOR2_X1 U12686 ( .A1(n10654), .A2(n10241), .ZN(n11351) );
  NAND2_X1 U12687 ( .A1(n10654), .A2(n10241), .ZN(n10214) );
  NAND2_X1 U12688 ( .A1(n10214), .A2(n6486), .ZN(n10215) );
  NOR2_X1 U12689 ( .A1(n11351), .A2(n10215), .ZN(n13421) );
  AOI21_X1 U12690 ( .B1(n14735), .B2(n10654), .A(n13421), .ZN(n10216) );
  OAI211_X1 U12691 ( .C1(n10217), .C2(n14739), .A(n13413), .B(n10216), .ZN(
        n13545) );
  NAND2_X1 U12692 ( .A1(n13545), .A2(n14756), .ZN(n10218) );
  OAI21_X1 U12693 ( .B1(n14756), .B2(n10219), .A(n10218), .ZN(P2_U3433) );
  INV_X1 U12694 ( .A(n10516), .ZN(n10524) );
  OAI222_X1 U12695 ( .A1(n13578), .A2(n10221), .B1(n13581), .B2(n10220), .C1(
        n10524), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI21_X1 U12696 ( .B1(n10223), .B2(n10822), .A(n10238), .ZN(n10226) );
  AND2_X1 U12697 ( .A1(n10651), .A2(n10224), .ZN(n10225) );
  NAND2_X1 U12698 ( .A1(n10226), .A2(n10225), .ZN(n10421) );
  NOR2_X1 U12699 ( .A1(n10421), .A2(P2_U3088), .ZN(n10458) );
  NAND2_X1 U12700 ( .A1(n10227), .A2(n14686), .ZN(n14681) );
  NOR2_X1 U12701 ( .A1(n14681), .A2(n10822), .ZN(n10237) );
  INV_X1 U12702 ( .A(n10237), .ZN(n10229) );
  NAND2_X1 U12703 ( .A1(n9020), .A2(n10230), .ZN(n10231) );
  NAND2_X1 U12704 ( .A1(n10231), .A2(n10241), .ZN(n10247) );
  OAI21_X1 U12705 ( .B1(n10241), .B2(n10231), .A(n10247), .ZN(n10235) );
  INV_X1 U12706 ( .A(n10232), .ZN(n10233) );
  NAND2_X1 U12707 ( .A1(n13200), .A2(n13139), .ZN(n10826) );
  INV_X1 U12708 ( .A(n10826), .ZN(n10234) );
  AOI22_X1 U12709 ( .A1(n14235), .A2(n10235), .B1(n14237), .B2(n10234), .ZN(
        n10243) );
  INV_X1 U12710 ( .A(n10236), .ZN(n10825) );
  NOR2_X1 U12711 ( .A1(n10825), .A2(n6472), .ZN(n10993) );
  NAND2_X1 U12712 ( .A1(n10237), .A2(n10993), .ZN(n10240) );
  NAND2_X1 U12713 ( .A1(n14240), .A2(n10241), .ZN(n10242) );
  OAI211_X1 U12714 ( .C1(n10458), .C2(n10829), .A(n10243), .B(n10242), .ZN(
        P2_U3204) );
  NAND2_X1 U12715 ( .A1(n12213), .A2(n8489), .ZN(n10246) );
  NAND2_X1 U12716 ( .A1(n10247), .A2(n10246), .ZN(n10457) );
  NAND2_X1 U12717 ( .A1(n13200), .A2(n10230), .ZN(n10249) );
  XNOR2_X1 U12718 ( .A(n10248), .B(n10249), .ZN(n10456) );
  NAND2_X1 U12719 ( .A1(n10457), .A2(n10456), .ZN(n10252) );
  INV_X1 U12720 ( .A(n10248), .ZN(n10250) );
  NAND2_X1 U12721 ( .A1(n10250), .A2(n10249), .ZN(n10251) );
  NAND2_X1 U12722 ( .A1(n10252), .A2(n10251), .ZN(n10408) );
  XNOR2_X1 U12723 ( .A(n10426), .B(n11356), .ZN(n10409) );
  NAND2_X1 U12724 ( .A1(n13198), .A2(n10230), .ZN(n10410) );
  XNOR2_X1 U12725 ( .A(n10409), .B(n10410), .ZN(n10407) );
  XOR2_X1 U12726 ( .A(n10408), .B(n10407), .Z(n10255) );
  INV_X1 U12727 ( .A(n14237), .ZN(n13143) );
  AOI22_X1 U12728 ( .A1(n13141), .A2(n13200), .B1(n13197), .B2(n13139), .ZN(
        n11361) );
  OAI22_X1 U12729 ( .A1(n10458), .A2(n11350), .B1(n13143), .B2(n11361), .ZN(
        n10253) );
  AOI21_X1 U12730 ( .B1(n11356), .B2(n14240), .A(n10253), .ZN(n10254) );
  OAI21_X1 U12731 ( .B1(n10255), .B2(n13168), .A(n10254), .ZN(P2_U3209) );
  NAND2_X1 U12732 ( .A1(n10256), .A2(P1_B_REG_SCAN_IN), .ZN(n10258) );
  MUX2_X1 U12733 ( .A(n10258), .B(P1_B_REG_SCAN_IN), .S(n10257), .Z(n10259) );
  AND2_X1 U12734 ( .A1(n10259), .A2(n10262), .ZN(n10327) );
  INV_X1 U12735 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U12736 ( .A1(n10257), .A2(n10262), .ZN(n10260) );
  INV_X1 U12737 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10264) );
  INV_X1 U12738 ( .A(n10262), .ZN(n14129) );
  AND2_X1 U12739 ( .A1(n10256), .A2(n14129), .ZN(n10263) );
  AND2_X1 U12740 ( .A1(n10554), .A2(n10555), .ZN(n10298) );
  NOR4_X1 U12741 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10268) );
  NOR4_X1 U12742 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10267) );
  NOR4_X1 U12743 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10266) );
  NOR4_X1 U12744 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10265) );
  NAND4_X1 U12745 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10274) );
  NOR2_X1 U12746 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10272) );
  NOR4_X1 U12747 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10271) );
  NOR4_X1 U12748 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10270) );
  NOR4_X1 U12749 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10269) );
  NAND4_X1 U12750 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  OAI21_X1 U12751 ( .B1(n10274), .B2(n10273), .A(n10327), .ZN(n10297) );
  NAND2_X1 U12752 ( .A1(n10298), .A2(n10297), .ZN(n10292) );
  NAND3_X1 U12753 ( .A1(n10558), .A2(n14570), .A3(n10295), .ZN(n10276) );
  INV_X1 U12754 ( .A(n10285), .ZN(n10277) );
  AND2_X2 U12755 ( .A1(n10278), .A2(n10468), .ZN(n10811) );
  INV_X1 U12756 ( .A(n13688), .ZN(n10623) );
  INV_X2 U12757 ( .A(n10811), .ZN(n12139) );
  XNOR2_X1 U12758 ( .A(n10367), .B(n10368), .ZN(n10369) );
  NAND2_X1 U12759 ( .A1(n10811), .A2(n13690), .ZN(n10288) );
  INV_X1 U12760 ( .A(n10622), .ZN(n10646) );
  NAND2_X1 U12761 ( .A1(n10807), .A2(n10646), .ZN(n10287) );
  NAND2_X1 U12762 ( .A1(n10289), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10286) );
  INV_X1 U12763 ( .A(n13690), .ZN(n10291) );
  AOI22_X1 U12764 ( .A1(n10811), .A2(n10646), .B1(n10289), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10290) );
  AOI21_X1 U12765 ( .B1(n10318), .B2(n10733), .A(n10320), .ZN(n10370) );
  XOR2_X1 U12766 ( .A(n10369), .B(n10370), .Z(n10303) );
  NAND2_X1 U12767 ( .A1(n10292), .A2(n10466), .ZN(n10728) );
  AND2_X1 U12768 ( .A1(n10728), .A2(n10558), .ZN(n14352) );
  INV_X1 U12769 ( .A(n10293), .ZN(n10296) );
  NAND2_X1 U12770 ( .A1(n10728), .A2(n10296), .ZN(n10376) );
  INV_X1 U12771 ( .A(n10376), .ZN(n10300) );
  AND2_X1 U12772 ( .A1(n14354), .A2(n14003), .ZN(n10620) );
  AOI21_X1 U12773 ( .B1(n14353), .B2(n13690), .A(n10620), .ZN(n10299) );
  NAND2_X1 U12774 ( .A1(n10298), .A2(n10556), .ZN(n14284) );
  OAI22_X1 U12775 ( .A1(n10300), .A2(n13691), .B1(n10299), .B2(n14284), .ZN(
        n10301) );
  AOI21_X1 U12776 ( .B1(n14297), .B2(n10277), .A(n10301), .ZN(n10302) );
  OAI21_X1 U12777 ( .B1(n13663), .B2(n10303), .A(n10302), .ZN(P1_U3222) );
  INV_X1 U12778 ( .A(n10304), .ZN(n10366) );
  AOI22_X1 U12779 ( .A1(n10497), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n14114), .ZN(n10305) );
  OAI21_X1 U12780 ( .B1(n10366), .B2(n14128), .A(n10305), .ZN(P1_U3342) );
  NAND2_X1 U12781 ( .A1(n10306), .A2(n14997), .ZN(n10307) );
  AND2_X1 U12782 ( .A1(n10309), .A2(n10307), .ZN(n10311) );
  OAI211_X1 U12783 ( .C1(n10311), .C2(n10310), .A(n12376), .B(n10397), .ZN(
        n10315) );
  INV_X1 U12784 ( .A(n12386), .ZN(n12359) );
  INV_X1 U12785 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10312) );
  NOR2_X1 U12786 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10312), .ZN(n14785) );
  INV_X1 U12787 ( .A(n12355), .ZN(n12379) );
  OAI22_X1 U12788 ( .A1(n12379), .A2(n14997), .B1(n10794), .B2(n12380), .ZN(
        n10313) );
  AOI211_X1 U12789 ( .C1(n12359), .C2(n14970), .A(n14785), .B(n10313), .ZN(
        n10314) );
  OAI211_X1 U12790 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n10956), .A(n10315), .B(
        n10314), .ZN(P3_U3158) );
  INV_X1 U12791 ( .A(n10316), .ZN(n10317) );
  OAI222_X1 U12792 ( .A1(n12709), .A2(P3_U3151), .B1(n13056), .B2(n10317), 
        .C1(n7638), .C2(n13058), .ZN(P3_U3278) );
  AND2_X1 U12793 ( .A1(n10319), .A2(n10318), .ZN(n10321) );
  OR2_X1 U12794 ( .A1(n10321), .A2(n10320), .ZN(n10359) );
  NAND2_X1 U12795 ( .A1(n13688), .A2(n14003), .ZN(n10644) );
  NAND2_X1 U12796 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10376), .ZN(n10322) );
  OAI21_X1 U12797 ( .B1(n14284), .B2(n10644), .A(n10322), .ZN(n10323) );
  AOI21_X1 U12798 ( .B1(n14359), .B2(n10359), .A(n10323), .ZN(n10324) );
  OAI21_X1 U12799 ( .B1(n14286), .B2(n10622), .A(n10324), .ZN(P1_U3232) );
  INV_X1 U12800 ( .A(n12726), .ZN(n12734) );
  OAI222_X1 U12801 ( .A1(n13056), .A2(n10326), .B1(n13058), .B2(n10325), .C1(
        n12734), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U12802 ( .A(n10256), .ZN(n10329) );
  NAND2_X1 U12803 ( .A1(n10328), .A2(n14129), .ZN(n10345) );
  OAI22_X1 U12804 ( .A1(n14488), .A2(P1_D_REG_1__SCAN_IN), .B1(n10329), .B2(
        n10345), .ZN(n10330) );
  INV_X1 U12805 ( .A(n10330), .ZN(P1_U3446) );
  XNOR2_X1 U12806 ( .A(n10332), .B(n10331), .ZN(n10333) );
  NAND3_X1 U12807 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10340) );
  INV_X1 U12808 ( .A(n14979), .ZN(n15005) );
  NOR2_X1 U12809 ( .A1(n15047), .A2(n15005), .ZN(n10336) );
  NAND2_X1 U12810 ( .A1(n10338), .A2(n15047), .ZN(n10339) );
  OAI22_X1 U12811 ( .A1(n12564), .A2(n10339), .B1(n9118), .B2(n14996), .ZN(
        n15013) );
  AOI21_X1 U12812 ( .B1(n15007), .B2(P3_REG3_REG_0__SCAN_IN), .A(n15013), .ZN(
        n10341) );
  MUX2_X1 U12813 ( .A(n10342), .B(n10341), .S(n15010), .Z(n10343) );
  OAI21_X1 U12814 ( .B1(n10344), .B2(n12928), .A(n10343), .ZN(P3_U3233) );
  OAI22_X1 U12815 ( .A1(n14488), .A2(P1_D_REG_0__SCAN_IN), .B1(n10257), .B2(
        n10345), .ZN(n10346) );
  INV_X1 U12816 ( .A(n10346), .ZN(P1_U3445) );
  INV_X1 U12817 ( .A(n14380), .ZN(n13718) );
  OAI22_X1 U12818 ( .A1(n14384), .A2(n7392), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10347), .ZN(n10356) );
  XNOR2_X1 U12819 ( .A(n10349), .B(n10348), .ZN(n10354) );
  OAI211_X1 U12820 ( .C1(n10352), .C2(n10351), .A(n14375), .B(n10350), .ZN(
        n10353) );
  OAI21_X1 U12821 ( .B1(n10354), .B2(n14370), .A(n10353), .ZN(n10355) );
  AOI211_X1 U12822 ( .C1(n10357), .C2(n13718), .A(n10356), .B(n10355), .ZN(
        n10364) );
  NAND2_X1 U12823 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13694) );
  MUX2_X1 U12824 ( .A(n10359), .B(n13694), .S(n10358), .Z(n10363) );
  NAND2_X1 U12825 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  OAI211_X1 U12826 ( .C1(n10363), .C2(n11928), .A(n13689), .B(n10362), .ZN(
        n13732) );
  NAND2_X1 U12827 ( .A1(n10364), .A2(n13732), .ZN(P1_U3245) );
  INV_X1 U12828 ( .A(n11123), .ZN(n11113) );
  INV_X1 U12829 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10365) );
  OAI222_X1 U12830 ( .A1(P2_U3088), .A2(n11113), .B1(n13581), .B2(n10366), 
        .C1(n10365), .C2(n13578), .ZN(P2_U3314) );
  OAI22_X1 U12831 ( .A1(n10370), .A2(n10369), .B1(n10368), .B2(n10367), .ZN(
        n10739) );
  INV_X1 U12832 ( .A(n10371), .ZN(n10372) );
  INV_X1 U12833 ( .A(n10733), .ZN(n12039) );
  XNOR2_X1 U12834 ( .A(n10372), .B(n12039), .ZN(n10737) );
  OAI22_X1 U12835 ( .A1(n10373), .A2(n10374), .B1(n14503), .B2(n12139), .ZN(
        n10735) );
  XNOR2_X1 U12836 ( .A(n10737), .B(n10735), .ZN(n10738) );
  XNOR2_X1 U12837 ( .A(n10739), .B(n10738), .ZN(n10375) );
  NAND2_X1 U12838 ( .A1(n10375), .A2(n14359), .ZN(n10378) );
  OAI22_X1 U12839 ( .A1(n10623), .A2(n13658), .B1(n10732), .B2(n14356), .ZN(
        n10635) );
  AOI22_X1 U12840 ( .A1(n10376), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14364), 
        .B2(n10635), .ZN(n10377) );
  OAI211_X1 U12841 ( .C1(n14503), .C2(n14286), .A(n10378), .B(n10377), .ZN(
        P1_U3237) );
  OR2_X1 U12842 ( .A1(n10387), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10379) );
  AND2_X1 U12843 ( .A1(n10380), .A2(n10379), .ZN(n10382) );
  INV_X1 U12844 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14318) );
  MUX2_X1 U12845 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14318), .S(n10497), .Z(
        n10381) );
  NAND2_X1 U12846 ( .A1(n10382), .A2(n10381), .ZN(n10492) );
  OAI211_X1 U12847 ( .C1(n10382), .C2(n10381), .A(n10492), .B(n14375), .ZN(
        n10394) );
  NAND2_X1 U12848 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11821)
         );
  INV_X1 U12849 ( .A(n11821), .ZN(n10383) );
  AOI21_X1 U12850 ( .B1(n13787), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10383), 
        .ZN(n10384) );
  INV_X1 U12851 ( .A(n10384), .ZN(n10392) );
  INV_X1 U12852 ( .A(n10385), .ZN(n10386) );
  OAI21_X1 U12853 ( .B1(n10387), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10386), 
        .ZN(n10390) );
  INV_X1 U12854 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10388) );
  MUX2_X1 U12855 ( .A(n10388), .B(P1_REG2_REG_13__SCAN_IN), .S(n10497), .Z(
        n10389) );
  NOR2_X1 U12856 ( .A1(n10389), .A2(n10390), .ZN(n10496) );
  AOI211_X1 U12857 ( .C1(n10390), .C2(n10389), .A(n10496), .B(n14370), .ZN(
        n10391) );
  AOI211_X1 U12858 ( .C1(n13718), .C2(n10497), .A(n10392), .B(n10391), .ZN(
        n10393) );
  NAND2_X1 U12859 ( .A1(n10394), .A2(n10393), .ZN(P1_U3256) );
  XNOR2_X1 U12860 ( .A(n10097), .B(n10919), .ZN(n10398) );
  NAND2_X1 U12861 ( .A1(n10398), .A2(n10794), .ZN(n10505) );
  OAI21_X1 U12862 ( .B1(n10398), .B2(n10794), .A(n10505), .ZN(n10399) );
  AOI21_X1 U12863 ( .B1(n10400), .B2(n10399), .A(n10507), .ZN(n10406) );
  NOR2_X1 U12864 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10401), .ZN(n14809) );
  OAI22_X1 U12865 ( .A1(n12379), .A2(n14983), .B1(n10690), .B2(n12380), .ZN(
        n10402) );
  AOI211_X1 U12866 ( .C1(n12359), .C2(n10919), .A(n14809), .B(n10402), .ZN(
        n10405) );
  INV_X1 U12867 ( .A(n10920), .ZN(n10403) );
  NAND2_X1 U12868 ( .A1(n12383), .A2(n10403), .ZN(n10404) );
  OAI211_X1 U12869 ( .C1(n10406), .C2(n12371), .A(n10405), .B(n10404), .ZN(
        P3_U3170) );
  INV_X1 U12870 ( .A(n14240), .ZN(n13149) );
  NAND2_X1 U12871 ( .A1(n10408), .A2(n10407), .ZN(n10413) );
  INV_X1 U12872 ( .A(n10409), .ZN(n10411) );
  NAND2_X1 U12873 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  INV_X1 U12874 ( .A(n10416), .ZN(n10414) );
  NAND2_X1 U12875 ( .A1(n10416), .A2(n10415), .ZN(n10427) );
  AOI21_X1 U12876 ( .B1(n10417), .B2(n10418), .A(n13168), .ZN(n10420) );
  NAND2_X1 U12877 ( .A1(n10420), .A2(n10428), .ZN(n10425) );
  INV_X1 U12878 ( .A(n13196), .ZN(n10700) );
  OAI22_X1 U12879 ( .A1(n7235), .A2(n13163), .B1(n10700), .B2(n13161), .ZN(
        n10667) );
  INV_X1 U12880 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U12881 ( .A1(n14243), .A2(n10422), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10423) );
  AOI21_X1 U12882 ( .B1(n14237), .B2(n10667), .A(n10423), .ZN(n10424) );
  OAI211_X1 U12883 ( .C1(n11044), .C2(n13149), .A(n10425), .B(n10424), .ZN(
        P2_U3190) );
  INV_X2 U12884 ( .A(n10426), .ZN(n12205) );
  XNOR2_X1 U12885 ( .A(n10994), .B(n12205), .ZN(n10478) );
  NAND2_X1 U12886 ( .A1(n13196), .A2(n10230), .ZN(n10477) );
  XNOR2_X1 U12887 ( .A(n10478), .B(n10477), .ZN(n10433) );
  INV_X1 U12888 ( .A(n10432), .ZN(n10430) );
  INV_X1 U12889 ( .A(n10433), .ZN(n10429) );
  NAND2_X1 U12890 ( .A1(n10430), .A2(n10429), .ZN(n10480) );
  INV_X1 U12891 ( .A(n10480), .ZN(n10431) );
  AOI21_X1 U12892 ( .B1(n10433), .B2(n10432), .A(n10431), .ZN(n10441) );
  NAND2_X1 U12893 ( .A1(n13197), .A2(n13141), .ZN(n10435) );
  NAND2_X1 U12894 ( .A1(n13195), .A2(n13139), .ZN(n10434) );
  AND2_X1 U12895 ( .A1(n10435), .A2(n10434), .ZN(n10989) );
  INV_X1 U12896 ( .A(n10989), .ZN(n10436) );
  NAND2_X1 U12897 ( .A1(n14237), .A2(n10436), .ZN(n10437) );
  OAI211_X1 U12898 ( .C1(n14243), .C2(n10998), .A(n10438), .B(n10437), .ZN(
        n10439) );
  AOI21_X1 U12899 ( .B1(n10994), .B2(n14240), .A(n10439), .ZN(n10440) );
  OAI21_X1 U12900 ( .B1(n10441), .B2(n13168), .A(n10440), .ZN(P2_U3202) );
  INV_X1 U12901 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14334) );
  NAND2_X1 U12902 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11422)
         );
  OAI21_X1 U12903 ( .B1(n14677), .B2(n14334), .A(n11422), .ZN(n10448) );
  NOR2_X1 U12904 ( .A1(n10449), .A2(n8673), .ZN(n10443) );
  XNOR2_X1 U12905 ( .A(n10516), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n10442) );
  NOR3_X1 U12906 ( .A1(n10444), .A2(n10443), .A3(n10442), .ZN(n10518) );
  INV_X1 U12907 ( .A(n10518), .ZN(n10446) );
  OAI21_X1 U12908 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(n10445) );
  AOI21_X1 U12909 ( .B1(n10446), .B2(n10445), .A(n14668), .ZN(n10447) );
  AOI211_X1 U12910 ( .C1(n14673), .C2(n10516), .A(n10448), .B(n10447), .ZN(
        n10455) );
  NAND2_X1 U12911 ( .A1(n10449), .A2(n10163), .ZN(n10450) );
  MUX2_X1 U12912 ( .A(n11309), .B(P2_REG2_REG_12__SCAN_IN), .S(n10516), .Z(
        n10451) );
  AOI21_X1 U12913 ( .B1(n10452), .B2(n10450), .A(n10451), .ZN(n10523) );
  AND3_X1 U12914 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n10453) );
  OAI21_X1 U12915 ( .B1(n10523), .B2(n10453), .A(n14655), .ZN(n10454) );
  NAND2_X1 U12916 ( .A1(n10455), .A2(n10454), .ZN(P2_U3226) );
  XOR2_X1 U12917 ( .A(n10456), .B(n10457), .Z(n10463) );
  INV_X1 U12918 ( .A(n10458), .ZN(n10461) );
  INV_X1 U12919 ( .A(n10654), .ZN(n13416) );
  OAI22_X1 U12920 ( .A1(n13416), .A2(n13149), .B1(n13143), .B2(n10459), .ZN(
        n10460) );
  AOI21_X1 U12921 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10461), .A(n10460), .ZN(
        n10462) );
  OAI21_X1 U12922 ( .B1(n10463), .B2(n13168), .A(n10462), .ZN(P2_U3194) );
  OAI222_X1 U12923 ( .A1(n12740), .A2(P3_U3151), .B1(n13058), .B2(n10465), 
        .C1(n13056), .C2(n10464), .ZN(P3_U3276) );
  NOR2_X1 U12924 ( .A1(n10555), .A2(n10557), .ZN(n10467) );
  INV_X1 U12925 ( .A(n10649), .ZN(n10475) );
  AOI21_X1 U12926 ( .B1(n10468), .B2(n14131), .A(n13964), .ZN(n10469) );
  NAND2_X1 U12927 ( .A1(n12140), .A2(n10469), .ZN(n14497) );
  OR2_X1 U12928 ( .A1(n10470), .A2(n13897), .ZN(n14095) );
  NAND2_X1 U12929 ( .A1(n14131), .A2(n13964), .ZN(n10472) );
  NAND2_X1 U12930 ( .A1(n14517), .A2(n14566), .ZN(n10474) );
  OAI21_X1 U12931 ( .B1(n10570), .B2(n10622), .A(n10644), .ZN(n10473) );
  AOI21_X1 U12932 ( .B1(n10475), .B2(n10474), .A(n10473), .ZN(n14489) );
  NAND2_X1 U12933 ( .A1(n14591), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10476) );
  OAI21_X1 U12934 ( .B1(n14591), .B2(n14489), .A(n10476), .ZN(P1_U3528) );
  XNOR2_X1 U12935 ( .A(n11052), .B(n12213), .ZN(n10535) );
  NAND2_X1 U12936 ( .A1(n13195), .A2(n10230), .ZN(n10536) );
  XNOR2_X1 U12937 ( .A(n10535), .B(n10536), .ZN(n10482) );
  NAND2_X1 U12938 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  NAND2_X1 U12939 ( .A1(n10480), .A2(n10479), .ZN(n10481) );
  OAI21_X1 U12940 ( .B1(n10482), .B2(n10481), .A(n10539), .ZN(n10489) );
  INV_X1 U12941 ( .A(n11052), .ZN(n11036) );
  NOR2_X1 U12942 ( .A1(n13149), .A2(n11036), .ZN(n10488) );
  NAND2_X1 U12943 ( .A1(n13196), .A2(n13141), .ZN(n10484) );
  NAND2_X1 U12944 ( .A1(n13194), .A2(n13139), .ZN(n10483) );
  NAND2_X1 U12945 ( .A1(n10484), .A2(n10483), .ZN(n10707) );
  NAND2_X1 U12946 ( .A1(n14237), .A2(n10707), .ZN(n10485) );
  OAI211_X1 U12947 ( .C1(n14243), .C2(n11035), .A(n10486), .B(n10485), .ZN(
        n10487) );
  AOI211_X1 U12948 ( .C1(n10489), .C2(n14235), .A(n10488), .B(n10487), .ZN(
        n10490) );
  INV_X1 U12949 ( .A(n10490), .ZN(P2_U3199) );
  NAND2_X1 U12950 ( .A1(n10497), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U12951 ( .A1(n10492), .A2(n10491), .ZN(n10494) );
  MUX2_X1 U12952 ( .A(n8095), .B(P1_REG1_REG_14__SCAN_IN), .S(n10967), .Z(
        n10493) );
  NAND2_X1 U12953 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  AOI21_X1 U12954 ( .B1(n10969), .B2(n10495), .A(n13767), .ZN(n10504) );
  AOI21_X1 U12955 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10497), .A(n10496), 
        .ZN(n10499) );
  MUX2_X1 U12956 ( .A(n10959), .B(P1_REG2_REG_14__SCAN_IN), .S(n10967), .Z(
        n10498) );
  NOR2_X1 U12957 ( .A1(n10499), .A2(n10498), .ZN(n10957) );
  AOI211_X1 U12958 ( .C1(n10499), .C2(n10498), .A(n14370), .B(n10957), .ZN(
        n10503) );
  INV_X1 U12959 ( .A(n10967), .ZN(n10960) );
  NAND2_X1 U12960 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14250)
         );
  INV_X1 U12961 ( .A(n14250), .ZN(n10500) );
  AOI21_X1 U12962 ( .B1(n13787), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10500), 
        .ZN(n10501) );
  OAI21_X1 U12963 ( .B1(n10960), .B2(n14380), .A(n10501), .ZN(n10502) );
  OR3_X1 U12964 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(P1_U3257) );
  INV_X1 U12965 ( .A(n10505), .ZN(n10506) );
  XNOR2_X1 U12966 ( .A(n10097), .B(n10511), .ZN(n10683) );
  XNOR2_X1 U12967 ( .A(n10683), .B(n10690), .ZN(n10508) );
  AOI21_X1 U12968 ( .B1(n10509), .B2(n10508), .A(n10684), .ZN(n10515) );
  AND2_X1 U12969 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14826) );
  OAI22_X1 U12970 ( .A1(n12379), .A2(n10794), .B1(n10838), .B2(n12380), .ZN(
        n10510) );
  AOI211_X1 U12971 ( .C1(n12359), .C2(n10511), .A(n14826), .B(n10510), .ZN(
        n10514) );
  INV_X1 U12972 ( .A(n10799), .ZN(n10512) );
  NAND2_X1 U12973 ( .A1(n12383), .A2(n10512), .ZN(n10513) );
  OAI211_X1 U12974 ( .C1(n10515), .C2(n12371), .A(n10514), .B(n10513), .ZN(
        P3_U3167) );
  NAND2_X1 U12975 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11548)
         );
  OAI21_X1 U12976 ( .B1(n14677), .B2(n7482), .A(n11548), .ZN(n10522) );
  XNOR2_X1 U12977 ( .A(n11123), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n10520) );
  NOR2_X1 U12978 ( .A1(n10516), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10517) );
  OR2_X1 U12979 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  NOR3_X1 U12980 ( .A1(n10518), .A2(n10517), .A3(n10520), .ZN(n11122) );
  AOI211_X1 U12981 ( .C1(n10520), .C2(n10519), .A(n14668), .B(n11122), .ZN(
        n10521) );
  AOI211_X1 U12982 ( .C1(n14673), .C2(n11123), .A(n10522), .B(n10521), .ZN(
        n10530) );
  NAND2_X1 U12983 ( .A1(n11123), .A2(n11114), .ZN(n10525) );
  OAI21_X1 U12984 ( .B1(n11123), .B2(n11114), .A(n10525), .ZN(n10527) );
  NAND2_X1 U12985 ( .A1(n11113), .A2(n11114), .ZN(n10526) );
  OAI211_X1 U12986 ( .C1(n11114), .C2(n11113), .A(n10528), .B(n10526), .ZN(
        n11112) );
  OAI211_X1 U12987 ( .C1(n10528), .C2(n10527), .A(n11112), .B(n14655), .ZN(
        n10529) );
  NAND2_X1 U12988 ( .A1(n10530), .A2(n10529), .ZN(P2_U3227) );
  INV_X1 U12989 ( .A(n11119), .ZN(n11326) );
  INV_X1 U12990 ( .A(n10531), .ZN(n10533) );
  OAI222_X1 U12991 ( .A1(P2_U3088), .A2(n11326), .B1(n13581), .B2(n10533), 
        .C1(n10532), .C2(n13578), .ZN(P2_U3311) );
  INV_X1 U12992 ( .A(n13763), .ZN(n13776) );
  OAI222_X1 U12993 ( .A1(n14125), .A2(n10534), .B1(n14128), .B2(n10533), .C1(
        n13776), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12994 ( .A(n10535), .ZN(n10537) );
  NAND2_X1 U12995 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  XNOR2_X1 U12996 ( .A(n14706), .B(n12213), .ZN(n10540) );
  AND2_X1 U12997 ( .A1(n13194), .A2(n10230), .ZN(n10541) );
  NAND2_X1 U12998 ( .A1(n10540), .A2(n10541), .ZN(n10716) );
  INV_X1 U12999 ( .A(n10540), .ZN(n10543) );
  INV_X1 U13000 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U13001 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  AND2_X1 U13002 ( .A1(n10716), .A2(n10544), .ZN(n10545) );
  OAI211_X1 U13003 ( .C1(n10546), .C2(n10545), .A(n10717), .B(n14235), .ZN(
        n10553) );
  NAND2_X1 U13004 ( .A1(n13195), .A2(n13141), .ZN(n10548) );
  NAND2_X1 U13005 ( .A1(n13193), .A2(n13139), .ZN(n10547) );
  NAND2_X1 U13006 ( .A1(n10548), .A2(n10547), .ZN(n11061) );
  NAND2_X1 U13007 ( .A1(n14237), .A2(n11061), .ZN(n10549) );
  OAI211_X1 U13008 ( .C1(n14243), .C2(n11067), .A(n10550), .B(n10549), .ZN(
        n10551) );
  AOI21_X1 U13009 ( .B1(n14706), .B2(n14240), .A(n10551), .ZN(n10552) );
  NAND2_X1 U13010 ( .A1(n10553), .A2(n10552), .ZN(P2_U3211) );
  INV_X1 U13011 ( .A(n10554), .ZN(n11683) );
  NAND3_X1 U13012 ( .A1(n11683), .A2(n10556), .A3(n10555), .ZN(n13845) );
  NAND2_X2 U13013 ( .A1(n10558), .A2(n10557), .ZN(n14439) );
  OR2_X1 U13014 ( .A1(n14395), .A2(n14497), .ZN(n10560) );
  AND2_X1 U13015 ( .A1(n13690), .A2(n10646), .ZN(n10617) );
  NAND2_X1 U13016 ( .A1(n10623), .A2(n10285), .ZN(n10561) );
  OAI21_X2 U13017 ( .B1(n10618), .B2(n10617), .A(n10561), .ZN(n10629) );
  OR2_X1 U13018 ( .A1(n14354), .A2(n10637), .ZN(n10562) );
  NAND2_X1 U13019 ( .A1(n14435), .A2(n14437), .ZN(n10565) );
  INV_X1 U13020 ( .A(n10732), .ZN(n13687) );
  OR2_X1 U13021 ( .A1(n14447), .A2(n13687), .ZN(n10564) );
  XNOR2_X1 U13022 ( .A(n10589), .B(n10583), .ZN(n14518) );
  NAND2_X1 U13023 ( .A1(n10285), .A2(n10622), .ZN(n10636) );
  OAI211_X1 U13024 ( .C1(n14516), .C2(n14451), .A(n14448), .B(n14430), .ZN(
        n14515) );
  NAND2_X1 U13025 ( .A1(n13687), .A2(n14353), .ZN(n10567) );
  NAND2_X1 U13026 ( .A1(n13685), .A2(n14003), .ZN(n10566) );
  AND2_X1 U13027 ( .A1(n10567), .A2(n10566), .ZN(n14514) );
  INV_X1 U13028 ( .A(n14439), .ZN(n14394) );
  INV_X1 U13029 ( .A(n10754), .ZN(n10568) );
  NAND2_X1 U13030 ( .A1(n14394), .A2(n10568), .ZN(n10569) );
  OAI211_X1 U13031 ( .C1(n14515), .C2(n13964), .A(n14514), .B(n10569), .ZN(
        n10575) );
  INV_X1 U13032 ( .A(n10570), .ZN(n10572) );
  NAND2_X1 U13033 ( .A1(n10572), .A2(n10571), .ZN(n10573) );
  OAI22_X1 U13034 ( .A1(n14516), .A2(n14444), .B1(n14010), .B2(n7888), .ZN(
        n10574) );
  AOI21_X1 U13035 ( .B1(n14010), .B2(n10575), .A(n10574), .ZN(n10588) );
  INV_X1 U13036 ( .A(n13955), .ZN(n13995) );
  INV_X1 U13037 ( .A(n10576), .ZN(n10577) );
  OAI21_X1 U13038 ( .B1(n10578), .B2(n10577), .A(n6511), .ZN(n10632) );
  INV_X1 U13039 ( .A(n10632), .ZN(n10580) );
  NAND2_X1 U13040 ( .A1(n10630), .A2(n14436), .ZN(n10582) );
  NAND2_X1 U13041 ( .A1(n10582), .A2(n10581), .ZN(n10584) );
  NAND3_X1 U13042 ( .A1(n10584), .A2(n6937), .A3(n10585), .ZN(n10586) );
  NAND2_X1 U13043 ( .A1(n10594), .A2(n10586), .ZN(n14521) );
  NAND2_X1 U13044 ( .A1(n13995), .A2(n14521), .ZN(n10587) );
  OAI211_X1 U13045 ( .C1(n13998), .C2(n14518), .A(n10588), .B(n10587), .ZN(
        P1_U3289) );
  NAND2_X1 U13046 ( .A1(n10589), .A2(n6937), .ZN(n10591) );
  NAND2_X1 U13047 ( .A1(n14516), .A2(n14357), .ZN(n10590) );
  NAND2_X1 U13048 ( .A1(n10591), .A2(n10590), .ZN(n14419) );
  INV_X1 U13049 ( .A(n10595), .ZN(n14421) );
  NAND2_X1 U13050 ( .A1(n14419), .A2(n14421), .ZN(n10593) );
  OR2_X1 U13051 ( .A1(n14431), .A2(n13685), .ZN(n10592) );
  XNOR2_X1 U13052 ( .A(n10767), .B(n10766), .ZN(n14532) );
  INV_X1 U13053 ( .A(n14532), .ZN(n10612) );
  NAND2_X1 U13054 ( .A1(n10598), .A2(n10599), .ZN(n10597) );
  NAND2_X1 U13055 ( .A1(n10597), .A2(n10596), .ZN(n10756) );
  NAND3_X1 U13056 ( .A1(n10766), .A2(n10599), .A3(n10598), .ZN(n10600) );
  NAND2_X1 U13057 ( .A1(n10756), .A2(n10600), .ZN(n10604) );
  NAND2_X1 U13058 ( .A1(n13685), .A2(n14353), .ZN(n10602) );
  NAND2_X1 U13059 ( .A1(n13683), .A2(n14003), .ZN(n10601) );
  AND2_X1 U13060 ( .A1(n10602), .A2(n10601), .ZN(n10860) );
  INV_X1 U13061 ( .A(n10860), .ZN(n10603) );
  AOI21_X1 U13062 ( .B1(n10604), .B2(n14522), .A(n10603), .ZN(n14539) );
  MUX2_X1 U13063 ( .A(n9932), .B(n14539), .S(n14010), .Z(n10611) );
  NAND2_X1 U13064 ( .A1(n14533), .A2(n14428), .ZN(n10605) );
  NAND2_X1 U13065 ( .A1(n10605), .A2(n14448), .ZN(n10606) );
  OR2_X1 U13066 ( .A1(n14415), .A2(n10606), .ZN(n14535) );
  INV_X1 U13067 ( .A(n14535), .ZN(n10609) );
  INV_X1 U13068 ( .A(n14533), .ZN(n10607) );
  OAI22_X1 U13069 ( .A1(n14444), .A2(n10607), .B1(n10859), .B2(n14439), .ZN(
        n10608) );
  AOI21_X1 U13070 ( .B1(n14452), .B2(n10609), .A(n10608), .ZN(n10610) );
  OAI211_X1 U13071 ( .C1(n13998), .C2(n10612), .A(n10611), .B(n10610), .ZN(
        P1_U3287) );
  INV_X1 U13072 ( .A(n10613), .ZN(n10615) );
  OAI222_X1 U13073 ( .A1(n14125), .A2(n10614), .B1(n14128), .B2(n10615), .C1(
        n10960), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13074 ( .A(n11124), .ZN(n14643) );
  OAI222_X1 U13075 ( .A1(n13578), .A2(n10616), .B1(n13581), .B2(n10615), .C1(
        n14643), .C2(P2_U3088), .ZN(P2_U3313) );
  XOR2_X1 U13076 ( .A(n10618), .B(n10617), .Z(n14498) );
  INV_X1 U13077 ( .A(n14010), .ZN(n14441) );
  NAND2_X1 U13078 ( .A1(n10618), .A2(n13690), .ZN(n10619) );
  AOI21_X1 U13079 ( .B1(n10619), .B2(n14522), .A(n14353), .ZN(n14491) );
  INV_X1 U13080 ( .A(n14491), .ZN(n10621) );
  AOI21_X1 U13081 ( .B1(n10621), .B2(n13690), .A(n10620), .ZN(n14496) );
  OAI22_X1 U13082 ( .A1(n14441), .A2(n14496), .B1(n13691), .B2(n14439), .ZN(
        n10625) );
  OAI21_X1 U13083 ( .B1(n6620), .B2(n10622), .A(n10636), .ZN(n14493) );
  XNOR2_X1 U13084 ( .A(n14493), .B(n10623), .ZN(n14490) );
  NOR3_X1 U13085 ( .A1(n13955), .A2(n14491), .A3(n14490), .ZN(n10624) );
  AOI211_X1 U13086 ( .C1(n14441), .C2(P1_REG2_REG_1__SCAN_IN), .A(n10625), .B(
        n10624), .ZN(n10628) );
  NOR2_X1 U13087 ( .A1(n13917), .A2(n14492), .ZN(n13979) );
  INV_X1 U13088 ( .A(n14493), .ZN(n10626) );
  AOI22_X1 U13089 ( .A1(n14396), .A2(n10277), .B1(n13979), .B2(n10626), .ZN(
        n10627) );
  OAI211_X1 U13090 ( .C1(n13998), .C2(n14498), .A(n10628), .B(n10627), .ZN(
        P1_U3292) );
  INV_X1 U13091 ( .A(n14497), .ZN(n14531) );
  XNOR2_X1 U13092 ( .A(n10629), .B(n10631), .ZN(n14507) );
  NAND2_X1 U13093 ( .A1(n10632), .A2(n10631), .ZN(n10633) );
  AOI21_X1 U13094 ( .B1(n10630), .B2(n10633), .A(n14566), .ZN(n10634) );
  AOI211_X1 U13095 ( .C1(n14531), .C2(n14507), .A(n10635), .B(n10634), .ZN(
        n14504) );
  AOI21_X1 U13096 ( .B1(n10637), .B2(n10636), .A(n14492), .ZN(n10638) );
  NAND2_X1 U13097 ( .A1(n10638), .A2(n14446), .ZN(n14502) );
  NOR2_X1 U13098 ( .A1(n13917), .A2(n14502), .ZN(n10641) );
  AOI22_X1 U13099 ( .A1(n14441), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14394), .ZN(n10639) );
  OAI21_X1 U13100 ( .B1(n14444), .B2(n14503), .A(n10639), .ZN(n10640) );
  AOI211_X1 U13101 ( .C1(n14507), .C2(n14453), .A(n10641), .B(n10640), .ZN(
        n10642) );
  OAI21_X1 U13102 ( .B1(n14395), .B2(n14504), .A(n10642), .ZN(P1_U3291) );
  INV_X1 U13103 ( .A(n13998), .ZN(n13953) );
  NOR2_X1 U13104 ( .A1(n13953), .A2(n13995), .ZN(n10650) );
  OAI22_X1 U13105 ( .A1(n14395), .A2(n10644), .B1(n10643), .B2(n14439), .ZN(
        n10645) );
  AOI21_X1 U13106 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14395), .A(n10645), .ZN(
        n10648) );
  OAI21_X1 U13107 ( .B1(n14396), .B2(n13979), .A(n10646), .ZN(n10647) );
  OAI211_X1 U13108 ( .C1(n10650), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        P1_U3293) );
  INV_X1 U13109 ( .A(n10651), .ZN(n10652) );
  OR2_X1 U13110 ( .A1(n13198), .A2(n11356), .ZN(n10657) );
  NAND2_X1 U13111 ( .A1(n11347), .A2(n10657), .ZN(n10658) );
  NAND2_X1 U13112 ( .A1(n10658), .A2(n10663), .ZN(n10696) );
  OAI21_X1 U13113 ( .B1(n10658), .B2(n10663), .A(n10696), .ZN(n10659) );
  INV_X1 U13114 ( .A(n10659), .ZN(n11049) );
  OR2_X1 U13115 ( .A1(n13200), .A2(n13416), .ZN(n10660) );
  NAND2_X1 U13116 ( .A1(n10661), .A2(n10660), .ZN(n11357) );
  INV_X1 U13117 ( .A(n11348), .ZN(n11358) );
  INV_X1 U13118 ( .A(n10663), .ZN(n10664) );
  NAND2_X1 U13119 ( .A1(n10665), .A2(n10664), .ZN(n10699) );
  OAI21_X1 U13120 ( .B1(n10665), .B2(n10664), .A(n10699), .ZN(n10668) );
  NOR2_X1 U13121 ( .A1(n11049), .A2(n10245), .ZN(n10666) );
  AOI211_X1 U13122 ( .C1(n13541), .C2(n10668), .A(n10667), .B(n10666), .ZN(
        n11042) );
  AND2_X1 U13123 ( .A1(n11351), .A2(n14693), .ZN(n11352) );
  INV_X1 U13124 ( .A(n11352), .ZN(n10670) );
  NAND2_X1 U13125 ( .A1(n11352), .A2(n11044), .ZN(n10995) );
  INV_X1 U13126 ( .A(n10995), .ZN(n10669) );
  AOI211_X1 U13127 ( .C1(n10694), .C2(n10670), .A(n10230), .B(n10669), .ZN(
        n11046) );
  AOI21_X1 U13128 ( .B1(n14735), .B2(n10694), .A(n11046), .ZN(n10671) );
  OAI211_X1 U13129 ( .C1(n11049), .C2(n14739), .A(n11042), .B(n10671), .ZN(
        n10673) );
  NAND2_X1 U13130 ( .A1(n10673), .A2(n14768), .ZN(n10672) );
  OAI21_X1 U13131 ( .B1(n14768), .B2(n8527), .A(n10672), .ZN(P2_U3502) );
  NAND2_X1 U13132 ( .A1(n10673), .A2(n14756), .ZN(n10674) );
  OAI21_X1 U13133 ( .B1(n14756), .B2(n8528), .A(n10674), .ZN(P2_U3439) );
  INV_X1 U13134 ( .A(n10675), .ZN(n10677) );
  INV_X1 U13135 ( .A(n13201), .ZN(n13208) );
  OAI222_X1 U13136 ( .A1(n13578), .A2(n10676), .B1(n13581), .B2(n10677), .C1(
        n13208), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13137 ( .A(n13789), .ZN(n13771) );
  OAI222_X1 U13138 ( .A1(n14125), .A2(n10678), .B1(n14128), .B2(n10677), .C1(
        n13771), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13139 ( .A(n10679), .ZN(n10681) );
  INV_X1 U13140 ( .A(n14653), .ZN(n11128) );
  OAI222_X1 U13141 ( .A1(n13578), .A2(n10680), .B1(n13581), .B2(n10681), .C1(
        n11128), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U13142 ( .A(n10970), .ZN(n14379) );
  OAI222_X1 U13143 ( .A1(n14125), .A2(n10682), .B1(n14128), .B2(n10681), .C1(
        n14379), .C2(P1_U3086), .ZN(P1_U3340) );
  XNOR2_X1 U13144 ( .A(n10097), .B(n10685), .ZN(n10833) );
  XNOR2_X1 U13145 ( .A(n10833), .B(n10838), .ZN(n10686) );
  OAI211_X1 U13146 ( .C1(n10687), .C2(n10686), .A(n10835), .B(n12376), .ZN(
        n10693) );
  NOR2_X1 U13147 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10688), .ZN(n14844) );
  OAI22_X1 U13148 ( .A1(n12379), .A2(n10690), .B1(n10689), .B2(n12380), .ZN(
        n10691) );
  AOI211_X1 U13149 ( .C1(n12359), .C2(n10930), .A(n14844), .B(n10691), .ZN(
        n10692) );
  OAI211_X1 U13150 ( .C1(n10931), .C2(n10956), .A(n10693), .B(n10692), .ZN(
        P3_U3179) );
  OR2_X1 U13151 ( .A1(n13197), .A2(n10694), .ZN(n10695) );
  INV_X1 U13152 ( .A(n10986), .ZN(n10981) );
  OR2_X1 U13153 ( .A1(n10994), .A2(n13196), .ZN(n10697) );
  XNOR2_X1 U13154 ( .A(n11054), .B(n10704), .ZN(n10708) );
  INV_X1 U13155 ( .A(n10708), .ZN(n11041) );
  OR2_X1 U13156 ( .A1(n11044), .A2(n13197), .ZN(n10698) );
  NAND2_X1 U13157 ( .A1(n10699), .A2(n10698), .ZN(n10987) );
  NAND2_X1 U13158 ( .A1(n10994), .A2(n10700), .ZN(n10703) );
  NAND2_X1 U13159 ( .A1(n10985), .A2(n10703), .ZN(n10702) );
  INV_X1 U13160 ( .A(n10704), .ZN(n10701) );
  NAND3_X1 U13161 ( .A1(n10985), .A2(n10704), .A3(n10703), .ZN(n10705) );
  AOI21_X1 U13162 ( .B1(n11058), .B2(n10705), .A(n13529), .ZN(n10706) );
  AOI211_X1 U13163 ( .C1(n14745), .C2(n10708), .A(n10707), .B(n10706), .ZN(
        n11033) );
  OR2_X1 U13164 ( .A1(n10995), .A2(n10994), .ZN(n10996) );
  NAND2_X1 U13165 ( .A1(n10996), .A2(n11052), .ZN(n10709) );
  NAND2_X1 U13166 ( .A1(n10709), .A2(n6486), .ZN(n10710) );
  NOR2_X1 U13167 ( .A1(n11064), .A2(n10710), .ZN(n11038) );
  AOI21_X1 U13168 ( .B1(n14735), .B2(n11052), .A(n11038), .ZN(n10711) );
  OAI211_X1 U13169 ( .C1(n11041), .C2(n14739), .A(n11033), .B(n10711), .ZN(
        n10713) );
  NAND2_X1 U13170 ( .A1(n10713), .A2(n14768), .ZN(n10712) );
  OAI21_X1 U13171 ( .B1(n14768), .B2(n8563), .A(n10712), .ZN(P2_U3504) );
  INV_X1 U13172 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U13173 ( .A1(n10713), .A2(n14756), .ZN(n10714) );
  OAI21_X1 U13174 ( .B1(n14756), .B2(n10715), .A(n10714), .ZN(P2_U3445) );
  INV_X1 U13175 ( .A(n14714), .ZN(n11464) );
  XNOR2_X1 U13176 ( .A(n14714), .B(n12213), .ZN(n10781) );
  NAND2_X1 U13177 ( .A1(n13193), .A2(n10230), .ZN(n10779) );
  XNOR2_X1 U13178 ( .A(n10781), .B(n10779), .ZN(n10718) );
  NAND2_X1 U13179 ( .A1(n10719), .A2(n10718), .ZN(n10783) );
  OAI211_X1 U13180 ( .C1(n10719), .C2(n10718), .A(n10783), .B(n14235), .ZN(
        n10722) );
  INV_X1 U13181 ( .A(n13194), .ZN(n11274) );
  OAI22_X1 U13182 ( .A1(n11278), .A2(n13161), .B1(n11274), .B2(n13163), .ZN(
        n11457) );
  AND2_X1 U13183 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14629) );
  NOR2_X1 U13184 ( .A1(n14243), .A2(n11461), .ZN(n10720) );
  AOI211_X1 U13185 ( .C1(n14237), .C2(n11457), .A(n14629), .B(n10720), .ZN(
        n10721) );
  OAI211_X1 U13186 ( .C1(n11464), .C2(n13149), .A(n10722), .B(n10721), .ZN(
        P2_U3185) );
  OAI222_X1 U13187 ( .A1(n10725), .A2(P3_U3151), .B1(n13058), .B2(n10724), 
        .C1(n13056), .C2(n10723), .ZN(P3_U3275) );
  NAND2_X1 U13188 ( .A1(n12603), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10726) );
  OAI21_X1 U13189 ( .B1(n12548), .B2(n12603), .A(n10726), .ZN(P3_U3521) );
  NAND2_X1 U13190 ( .A1(n10729), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10730) );
  INV_X1 U13191 ( .A(n14447), .ZN(n14443) );
  OAI22_X1 U13192 ( .A1(n10732), .A2(n10373), .B1(n14443), .B2(n12139), .ZN(
        n10741) );
  INV_X1 U13193 ( .A(n10741), .ZN(n10743) );
  XNOR2_X1 U13194 ( .A(n10734), .B(n10733), .ZN(n10740) );
  INV_X1 U13195 ( .A(n10740), .ZN(n10742) );
  INV_X1 U13196 ( .A(n10735), .ZN(n10736) );
  AOI22_X1 U13197 ( .A1(n10739), .A2(n10738), .B1(n10737), .B2(n10736), .ZN(
        n14361) );
  XOR2_X1 U13198 ( .A(n10741), .B(n10740), .Z(n14360) );
  NAND2_X1 U13199 ( .A1(n14361), .A2(n14360), .ZN(n14358) );
  OAI22_X1 U13200 ( .A1(n14516), .A2(n12139), .B1(n14357), .B2(n10373), .ZN(
        n10744) );
  NOR2_X2 U13201 ( .A1(n10745), .A2(n10744), .ZN(n10804) );
  NAND2_X1 U13202 ( .A1(n10745), .A2(n10744), .ZN(n10805) );
  INV_X1 U13203 ( .A(n10805), .ZN(n10746) );
  NOR2_X1 U13204 ( .A1(n10804), .A2(n10746), .ZN(n10748) );
  OAI22_X1 U13205 ( .A1(n14516), .A2(n10731), .B1(n14357), .B2(n12139), .ZN(
        n10747) );
  XOR2_X1 U13206 ( .A(n12140), .B(n10747), .Z(n10806) );
  XNOR2_X1 U13207 ( .A(n10748), .B(n10806), .ZN(n10749) );
  NAND2_X1 U13208 ( .A1(n10749), .A2(n14359), .ZN(n10753) );
  NAND2_X1 U13209 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U13210 ( .B1(n14284), .B2(n14514), .A(n13716), .ZN(n10750) );
  AOI21_X1 U13211 ( .B1(n14297), .B2(n10751), .A(n10750), .ZN(n10752) );
  OAI211_X1 U13212 ( .C1(n14367), .C2(n10754), .A(n10753), .B(n10752), .ZN(
        P1_U3230) );
  NAND2_X1 U13213 ( .A1(n10756), .A2(n10755), .ZN(n14403) );
  NAND2_X1 U13214 ( .A1(n14403), .A2(n14405), .ZN(n14402) );
  INV_X1 U13215 ( .A(n13683), .ZN(n11017) );
  NAND2_X1 U13216 ( .A1(n11027), .A2(n11017), .ZN(n10757) );
  INV_X1 U13217 ( .A(n10902), .ZN(n10758) );
  OAI21_X1 U13218 ( .B1(n6600), .B2(n10758), .A(n10897), .ZN(n14553) );
  NAND2_X1 U13219 ( .A1(n13683), .A2(n14353), .ZN(n10760) );
  NAND2_X1 U13220 ( .A1(n13681), .A2(n14003), .ZN(n10759) );
  NAND2_X1 U13221 ( .A1(n10760), .A2(n10759), .ZN(n14548) );
  INV_X1 U13222 ( .A(n14548), .ZN(n10761) );
  MUX2_X1 U13223 ( .A(n10761), .B(n9965), .S(n14395), .Z(n10762) );
  OAI21_X1 U13224 ( .B1(n14439), .B2(n11555), .A(n10762), .ZN(n10765) );
  INV_X1 U13225 ( .A(n11027), .ZN(n14542) );
  NAND2_X1 U13226 ( .A1(n14542), .A2(n14415), .ZN(n14414) );
  AOI21_X1 U13227 ( .B1(n14414), .B2(n14550), .A(n14492), .ZN(n10763) );
  OR2_X1 U13228 ( .A1(n14414), .A2(n14550), .ZN(n14397) );
  NAND2_X1 U13229 ( .A1(n10763), .A2(n14397), .ZN(n14551) );
  NOR2_X1 U13230 ( .A1(n14551), .A2(n13917), .ZN(n10764) );
  AOI211_X1 U13231 ( .C1(n14396), .C2(n14550), .A(n10765), .B(n10764), .ZN(
        n10774) );
  NAND2_X1 U13232 ( .A1(n10767), .A2(n10766), .ZN(n10769) );
  OR2_X1 U13233 ( .A1(n14533), .A2(n13684), .ZN(n10768) );
  NAND2_X1 U13234 ( .A1(n10769), .A2(n10768), .ZN(n14404) );
  INV_X1 U13235 ( .A(n14405), .ZN(n10770) );
  NAND2_X1 U13236 ( .A1(n14404), .A2(n10770), .ZN(n10772) );
  OR2_X1 U13237 ( .A1(n11027), .A2(n13683), .ZN(n10771) );
  NAND2_X1 U13238 ( .A1(n10772), .A2(n10771), .ZN(n10903) );
  XNOR2_X1 U13239 ( .A(n10903), .B(n10902), .ZN(n14555) );
  NAND2_X1 U13240 ( .A1(n14555), .A2(n13953), .ZN(n10773) );
  OAI211_X1 U13241 ( .C1(n14553), .C2(n13955), .A(n10774), .B(n10773), .ZN(
        P1_U3285) );
  XNOR2_X1 U13242 ( .A(n11484), .B(n12205), .ZN(n10775) );
  NAND2_X1 U13243 ( .A1(n13192), .A2(n10230), .ZN(n10776) );
  NAND2_X1 U13244 ( .A1(n10775), .A2(n10776), .ZN(n10871) );
  INV_X1 U13245 ( .A(n10775), .ZN(n10778) );
  INV_X1 U13246 ( .A(n10776), .ZN(n10777) );
  NAND2_X1 U13247 ( .A1(n10778), .A2(n10777), .ZN(n10873) );
  NAND2_X1 U13248 ( .A1(n10871), .A2(n10873), .ZN(n10784) );
  INV_X1 U13249 ( .A(n10779), .ZN(n10780) );
  NAND2_X1 U13250 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  XOR2_X1 U13251 ( .A(n10784), .B(n10872), .Z(n10789) );
  INV_X1 U13252 ( .A(n13193), .ZN(n11276) );
  OAI22_X1 U13253 ( .A1(n11276), .A2(n13163), .B1(n11281), .B2(n13161), .ZN(
        n11474) );
  NAND2_X1 U13254 ( .A1(n14237), .A2(n11474), .ZN(n10785) );
  OAI211_X1 U13255 ( .C1(n14243), .C2(n11481), .A(n10786), .B(n10785), .ZN(
        n10787) );
  AOI21_X1 U13256 ( .B1(n11484), .B2(n14240), .A(n10787), .ZN(n10788) );
  OAI21_X1 U13257 ( .B1(n10789), .B2(n13168), .A(n10788), .ZN(P2_U3193) );
  XNOR2_X1 U13258 ( .A(n10790), .B(n9192), .ZN(n15033) );
  NAND2_X1 U13259 ( .A1(n10791), .A2(n14979), .ZN(n11766) );
  INV_X1 U13260 ( .A(n11766), .ZN(n14990) );
  NAND2_X1 U13261 ( .A1(n15010), .A2(n14990), .ZN(n12794) );
  OAI21_X1 U13262 ( .B1(n6604), .B2(n9192), .A(n10793), .ZN(n10796) );
  OAI22_X1 U13263 ( .A1(n10794), .A2(n14998), .B1(n10838), .B2(n14996), .ZN(
        n10795) );
  AOI21_X1 U13264 ( .B1(n10796), .B2(n15001), .A(n10795), .ZN(n10797) );
  OAI21_X1 U13265 ( .B1(n15004), .B2(n15033), .A(n10797), .ZN(n15034) );
  NAND2_X1 U13266 ( .A1(n15034), .A2(n15010), .ZN(n10803) );
  NOR2_X1 U13267 ( .A1(n10798), .A2(n15047), .ZN(n15035) );
  INV_X1 U13268 ( .A(n15035), .ZN(n10800) );
  OAI22_X1 U13269 ( .A1(n14939), .A2(n10800), .B1(n10799), .B2(n14978), .ZN(
        n10801) );
  AOI21_X1 U13270 ( .B1(n15012), .B2(P3_REG2_REG_5__SCAN_IN), .A(n10801), .ZN(
        n10802) );
  OAI211_X1 U13271 ( .C1(n15033), .C2(n12794), .A(n10803), .B(n10802), .ZN(
        P3_U3228) );
  NAND2_X1 U13272 ( .A1(n14431), .A2(n12130), .ZN(n10809) );
  INV_X2 U13273 ( .A(n12139), .ZN(n12131) );
  NAND2_X1 U13274 ( .A1(n12131), .A2(n13685), .ZN(n10808) );
  NAND2_X1 U13275 ( .A1(n10809), .A2(n10808), .ZN(n10810) );
  XNOR2_X1 U13276 ( .A(n10810), .B(n12140), .ZN(n10852) );
  NAND2_X1 U13277 ( .A1(n14431), .A2(n12131), .ZN(n10813) );
  NAND2_X1 U13278 ( .A1(n12135), .A2(n13685), .ZN(n10812) );
  NAND2_X1 U13279 ( .A1(n10813), .A2(n10812), .ZN(n10851) );
  NAND2_X1 U13280 ( .A1(n13684), .A2(n14003), .ZN(n10814) );
  OAI21_X1 U13281 ( .B1(n14357), .B2(n13658), .A(n10814), .ZN(n14524) );
  AOI21_X1 U13282 ( .B1(n14364), .B2(n14524), .A(n10815), .ZN(n10817) );
  AND2_X1 U13283 ( .A1(n14431), .A2(n14549), .ZN(n14525) );
  NAND2_X1 U13284 ( .A1(n14352), .A2(n14525), .ZN(n10816) );
  OAI211_X1 U13285 ( .C1(n14367), .C2(n14423), .A(n10817), .B(n10816), .ZN(
        n10818) );
  AOI21_X1 U13286 ( .B1(n10819), .B2(n14359), .A(n10818), .ZN(n10820) );
  INV_X1 U13287 ( .A(n10820), .ZN(P1_U3227) );
  OR2_X1 U13288 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  OR2_X1 U13289 ( .A1(n10828), .A2(n8479), .ZN(n11050) );
  INV_X1 U13290 ( .A(n11050), .ZN(n10824) );
  NAND2_X1 U13291 ( .A1(n13406), .A2(n10824), .ZN(n11364) );
  NOR2_X1 U13292 ( .A1(n8489), .A2(n10825), .ZN(n14689) );
  NOR2_X1 U13293 ( .A1(n14745), .A2(n13541), .ZN(n10827) );
  OAI21_X1 U13294 ( .B1(n14687), .B2(n10827), .A(n10826), .ZN(n14688) );
  AOI21_X1 U13295 ( .B1(n14689), .B2(n10828), .A(n14688), .ZN(n10830) );
  OAI22_X1 U13296 ( .A1(n10830), .A2(n13402), .B1(n10829), .B2(n13414), .ZN(
        n10831) );
  AOI21_X1 U13297 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13402), .A(n10831), .ZN(
        n10832) );
  OAI21_X1 U13298 ( .B1(n14687), .B2(n11364), .A(n10832), .ZN(P2_U3265) );
  INV_X1 U13299 ( .A(n10833), .ZN(n10834) );
  XNOR2_X1 U13300 ( .A(n14944), .B(n10097), .ZN(n10942) );
  XOR2_X1 U13301 ( .A(n10941), .B(n10942), .Z(n10836) );
  NAND2_X1 U13302 ( .A1(n10836), .A2(n12376), .ZN(n10842) );
  NOR2_X1 U13303 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10837), .ZN(n14861) );
  OAI22_X1 U13304 ( .A1(n12379), .A2(n10838), .B1(n10946), .B2(n12380), .ZN(
        n10839) );
  AOI211_X1 U13305 ( .C1(n12359), .C2(n10840), .A(n14861), .B(n10839), .ZN(
        n10841) );
  OAI211_X1 U13306 ( .C1(n14955), .C2(n10956), .A(n10842), .B(n10841), .ZN(
        P3_U3153) );
  INV_X1 U13307 ( .A(n10843), .ZN(n10846) );
  INV_X1 U13308 ( .A(n14674), .ZN(n10844) );
  OAI222_X1 U13309 ( .A1(n13578), .A2(n10845), .B1(n13581), .B2(n10846), .C1(
        P2_U3088), .C2(n10844), .ZN(P2_U3309) );
  INV_X1 U13310 ( .A(n13804), .ZN(n13797) );
  OAI222_X1 U13311 ( .A1(n14125), .A2(n10847), .B1(n14128), .B2(n10846), .C1(
        P1_U3086), .C2(n13797), .ZN(P1_U3337) );
  INV_X1 U13312 ( .A(n10848), .ZN(n10850) );
  OAI22_X1 U13313 ( .A1(n12595), .A2(P3_U3151), .B1(SI_22_), .B2(n13058), .ZN(
        n10849) );
  AOI21_X1 U13314 ( .B1(n10850), .B2(n13048), .A(n10849), .ZN(P3_U3273) );
  INV_X1 U13315 ( .A(n10852), .ZN(n10855) );
  INV_X1 U13316 ( .A(n10851), .ZN(n10854) );
  NOR2_X1 U13317 ( .A1(n10373), .A2(n10856), .ZN(n10857) );
  AOI21_X1 U13318 ( .B1(n14533), .B2(n12131), .A(n10857), .ZN(n11019) );
  AOI22_X1 U13319 ( .A1(n14533), .A2(n12130), .B1(n12131), .B2(n13684), .ZN(
        n10858) );
  INV_X2 U13320 ( .A(n12039), .ZN(n12140) );
  XNOR2_X1 U13321 ( .A(n10858), .B(n12140), .ZN(n11020) );
  XOR2_X1 U13322 ( .A(n11019), .B(n11020), .Z(n11023) );
  XNOR2_X1 U13323 ( .A(n11024), .B(n11023), .ZN(n10865) );
  INV_X1 U13324 ( .A(n14367), .ZN(n13653) );
  INV_X1 U13325 ( .A(n10859), .ZN(n10862) );
  INV_X1 U13326 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n13733) );
  OAI22_X1 U13327 ( .A1(n14284), .A2(n10860), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13733), .ZN(n10861) );
  AOI21_X1 U13328 ( .B1(n13653), .B2(n10862), .A(n10861), .ZN(n10864) );
  NAND2_X1 U13329 ( .A1(n14297), .A2(n14533), .ZN(n10863) );
  OAI211_X1 U13330 ( .C1(n10865), .C2(n13663), .A(n10864), .B(n10863), .ZN(
        P1_U3239) );
  XNOR2_X1 U13331 ( .A(n14727), .B(n12205), .ZN(n10866) );
  NAND2_X1 U13332 ( .A1(n13191), .A2(n10230), .ZN(n10867) );
  NAND2_X1 U13333 ( .A1(n10866), .A2(n10867), .ZN(n10887) );
  INV_X1 U13334 ( .A(n10866), .ZN(n10869) );
  INV_X1 U13335 ( .A(n10867), .ZN(n10868) );
  NAND2_X1 U13336 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  NAND2_X1 U13337 ( .A1(n10887), .A2(n10870), .ZN(n10877) );
  INV_X1 U13338 ( .A(n10888), .ZN(n10875) );
  AOI21_X1 U13339 ( .B1(n10877), .B2(n10876), .A(n10875), .ZN(n10882) );
  NOR2_X1 U13340 ( .A1(n14243), .A2(n11337), .ZN(n10880) );
  AOI22_X1 U13341 ( .A1(n13141), .A2(n13192), .B1(n13190), .B2(n13139), .ZN(
        n11335) );
  OAI21_X1 U13342 ( .B1(n13143), .B2(n11335), .A(n10878), .ZN(n10879) );
  AOI211_X1 U13343 ( .C1(n14727), .C2(n14240), .A(n10880), .B(n10879), .ZN(
        n10881) );
  OAI21_X1 U13344 ( .B1(n10882), .B2(n13168), .A(n10881), .ZN(P2_U3203) );
  INV_X1 U13345 ( .A(n10883), .ZN(n10885) );
  OAI222_X1 U13346 ( .A1(n14125), .A2(n10884), .B1(n14128), .B2(n10885), .C1(
        P1_U3086), .C2(n13897), .ZN(P1_U3336) );
  OAI222_X1 U13347 ( .A1(n13578), .A2(n10886), .B1(n13581), .B2(n10885), .C1(
        n13217), .C2(P2_U3088), .ZN(P2_U3308) );
  XNOR2_X1 U13348 ( .A(n14736), .B(n12205), .ZN(n11098) );
  NAND2_X1 U13349 ( .A1(n13190), .A2(n10230), .ZN(n11099) );
  XNOR2_X1 U13350 ( .A(n11098), .B(n11099), .ZN(n11103) );
  XNOR2_X1 U13351 ( .A(n11104), .B(n11103), .ZN(n10895) );
  NOR2_X1 U13352 ( .A1(n14243), .A2(n11501), .ZN(n10893) );
  NAND2_X1 U13353 ( .A1(n13191), .A2(n13141), .ZN(n10890) );
  NAND2_X1 U13354 ( .A1(n13189), .A2(n13139), .ZN(n10889) );
  AND2_X1 U13355 ( .A1(n10890), .A2(n10889), .ZN(n11492) );
  OAI21_X1 U13356 ( .B1(n13143), .B2(n11492), .A(n10891), .ZN(n10892) );
  AOI211_X1 U13357 ( .C1(n14736), .C2(n14240), .A(n10893), .B(n10892), .ZN(
        n10894) );
  OAI21_X1 U13358 ( .B1(n10895), .B2(n13168), .A(n10894), .ZN(P2_U3189) );
  OR2_X1 U13359 ( .A1(n14550), .A2(n11390), .ZN(n10896) );
  INV_X1 U13360 ( .A(n13681), .ZN(n10898) );
  NAND2_X1 U13361 ( .A1(n14557), .A2(n10898), .ZN(n10899) );
  NAND2_X1 U13362 ( .A1(n10900), .A2(n10899), .ZN(n11004) );
  XNOR2_X1 U13363 ( .A(n11004), .B(n11007), .ZN(n14567) );
  NAND2_X1 U13364 ( .A1(n10903), .A2(n10902), .ZN(n10905) );
  OR2_X1 U13365 ( .A1(n14550), .A2(n13682), .ZN(n10904) );
  OR2_X1 U13366 ( .A1(n14557), .A2(n13681), .ZN(n10906) );
  XNOR2_X1 U13367 ( .A(n11008), .B(n11007), .ZN(n14575) );
  AOI211_X1 U13368 ( .C1(n11591), .C2(n6519), .A(n14492), .B(n11009), .ZN(
        n10908) );
  NAND2_X1 U13369 ( .A1(n13679), .A2(n14003), .ZN(n11597) );
  INV_X1 U13370 ( .A(n11597), .ZN(n10907) );
  NOR2_X1 U13371 ( .A1(n10908), .A2(n10907), .ZN(n14569) );
  NOR2_X1 U13372 ( .A1(n14441), .A2(n13964), .ZN(n13992) );
  INV_X1 U13373 ( .A(n13992), .ZN(n10912) );
  NAND2_X1 U13374 ( .A1(n13681), .A2(n14353), .ZN(n14568) );
  OAI22_X1 U13375 ( .A1(n14441), .A2(n14568), .B1(n11598), .B2(n14439), .ZN(
        n10910) );
  INV_X1 U13376 ( .A(n11591), .ZN(n14571) );
  NOR2_X1 U13377 ( .A1(n14571), .A2(n14444), .ZN(n10909) );
  AOI211_X1 U13378 ( .C1(n14441), .C2(P1_REG2_REG_10__SCAN_IN), .A(n10910), 
        .B(n10909), .ZN(n10911) );
  OAI21_X1 U13379 ( .B1(n14569), .B2(n10912), .A(n10911), .ZN(n10913) );
  AOI21_X1 U13380 ( .B1(n14575), .B2(n13953), .A(n10913), .ZN(n10914) );
  OAI21_X1 U13381 ( .B1(n14567), .B2(n13955), .A(n10914), .ZN(P1_U3283) );
  NAND2_X1 U13382 ( .A1(n10915), .A2(n13048), .ZN(n10916) );
  OAI211_X1 U13383 ( .C1(n10917), .C2(n13058), .A(n10916), .B(n12597), .ZN(
        P3_U3272) );
  XNOR2_X1 U13384 ( .A(n12406), .B(n10918), .ZN(n10925) );
  INV_X1 U13385 ( .A(n10925), .ZN(n15031) );
  INV_X1 U13386 ( .A(n12794), .ZN(n15008) );
  NAND2_X1 U13387 ( .A1(n10919), .A2(n15015), .ZN(n15028) );
  OAI22_X1 U13388 ( .A1(n14939), .A2(n15028), .B1(n10920), .B2(n14978), .ZN(
        n10927) );
  AOI22_X1 U13389 ( .A1(n14965), .A2(n12611), .B1(n12610), .B2(n14962), .ZN(
        n10924) );
  OAI211_X1 U13390 ( .C1(n10922), .C2(n12406), .A(n10921), .B(n15001), .ZN(
        n10923) );
  OAI211_X1 U13391 ( .C1(n10925), .C2(n15004), .A(n10924), .B(n10923), .ZN(
        n15029) );
  MUX2_X1 U13392 ( .A(n15029), .B(P3_REG2_REG_4__SCAN_IN), .S(n15012), .Z(
        n10926) );
  AOI211_X1 U13393 ( .C1(n15031), .C2(n15008), .A(n10927), .B(n10926), .ZN(
        n10928) );
  INV_X1 U13394 ( .A(n10928), .ZN(P3_U3229) );
  XNOR2_X1 U13395 ( .A(n10929), .B(n12563), .ZN(n15041) );
  NAND2_X1 U13396 ( .A1(n15015), .A2(n10930), .ZN(n15038) );
  OAI22_X1 U13397 ( .A1(n14939), .A2(n15038), .B1(n10931), .B2(n14978), .ZN(
        n10939) );
  OAI211_X1 U13398 ( .C1(n10934), .C2(n10933), .A(n10932), .B(n15001), .ZN(
        n10937) );
  AOI22_X1 U13399 ( .A1(n12610), .A2(n14965), .B1(n14962), .B2(n12609), .ZN(
        n10936) );
  INV_X1 U13400 ( .A(n15004), .ZN(n14985) );
  NAND2_X1 U13401 ( .A1(n15041), .A2(n14985), .ZN(n10935) );
  NAND3_X1 U13402 ( .A1(n10937), .A2(n10936), .A3(n10935), .ZN(n15039) );
  MUX2_X1 U13403 ( .A(n15039), .B(P3_REG2_REG_6__SCAN_IN), .S(n15012), .Z(
        n10938) );
  AOI211_X1 U13404 ( .C1(n15041), .C2(n15008), .A(n10939), .B(n10938), .ZN(
        n10940) );
  INV_X1 U13405 ( .A(n10940), .ZN(P3_U3227) );
  XNOR2_X1 U13406 ( .A(n12432), .B(n10097), .ZN(n11073) );
  XNOR2_X1 U13407 ( .A(n11073), .B(n14935), .ZN(n10950) );
  NAND2_X1 U13408 ( .A1(n10941), .A2(n10942), .ZN(n10945) );
  INV_X1 U13409 ( .A(n10942), .ZN(n10943) );
  NAND2_X1 U13410 ( .A1(n10945), .A2(n10944), .ZN(n12297) );
  XNOR2_X1 U13411 ( .A(n10097), .B(n15048), .ZN(n10947) );
  XNOR2_X1 U13412 ( .A(n10947), .B(n10946), .ZN(n12296) );
  OAI21_X1 U13413 ( .B1(n10950), .B2(n10949), .A(n11076), .ZN(n10951) );
  NAND2_X1 U13414 ( .A1(n10951), .A2(n12376), .ZN(n10955) );
  NOR2_X1 U13415 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10952), .ZN(n14898) );
  OAI22_X1 U13416 ( .A1(n12386), .A2(n11249), .B1(n12380), .B2(n14201), .ZN(
        n10953) );
  AOI211_X1 U13417 ( .C1(n12355), .C2(n14950), .A(n14898), .B(n10953), .ZN(
        n10954) );
  OAI211_X1 U13418 ( .C1(n11250), .C2(n10956), .A(n10955), .B(n10954), .ZN(
        P3_U3171) );
  INV_X1 U13419 ( .A(n10957), .ZN(n10958) );
  OAI21_X1 U13420 ( .B1(n10960), .B2(n10959), .A(n10958), .ZN(n10961) );
  NOR2_X1 U13421 ( .A1(n10970), .A2(n10961), .ZN(n10962) );
  XOR2_X1 U13422 ( .A(n10961), .B(n14379), .Z(n14369) );
  NOR2_X1 U13423 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14369), .ZN(n14368) );
  NOR2_X1 U13424 ( .A1(n10962), .A2(n14368), .ZN(n10966) );
  NOR2_X1 U13425 ( .A1(n13776), .A2(n10963), .ZN(n10964) );
  AOI21_X1 U13426 ( .B1(n10963), .B2(n13776), .A(n10964), .ZN(n10965) );
  NAND2_X1 U13427 ( .A1(n10965), .A2(n10966), .ZN(n13775) );
  OAI211_X1 U13428 ( .C1(n10966), .C2(n10965), .A(n13811), .B(n13775), .ZN(
        n10980) );
  OR2_X1 U13429 ( .A1(n10967), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10968) );
  XNOR2_X1 U13430 ( .A(n10971), .B(n14379), .ZN(n14374) );
  INV_X1 U13431 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14373) );
  NAND2_X1 U13432 ( .A1(n14374), .A2(n14373), .ZN(n14372) );
  OAI21_X1 U13433 ( .B1(n10971), .B2(n10970), .A(n14372), .ZN(n10974) );
  INV_X1 U13434 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11904) );
  NOR2_X1 U13435 ( .A1(n13763), .A2(n11904), .ZN(n10972) );
  AOI21_X1 U13436 ( .B1(n11904), .B2(n13763), .A(n10972), .ZN(n10973) );
  NOR2_X1 U13437 ( .A1(n10973), .A2(n10974), .ZN(n13762) );
  AOI211_X1 U13438 ( .C1(n10974), .C2(n10973), .A(n13762), .B(n13767), .ZN(
        n10978) );
  NAND2_X1 U13439 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14259)
         );
  INV_X1 U13440 ( .A(n14259), .ZN(n10975) );
  AOI21_X1 U13441 ( .B1(n13787), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10975), 
        .ZN(n10976) );
  OAI21_X1 U13442 ( .B1(n13776), .B2(n14380), .A(n10976), .ZN(n10977) );
  NOR2_X1 U13443 ( .A1(n10978), .A2(n10977), .ZN(n10979) );
  NAND2_X1 U13444 ( .A1(n10980), .A2(n10979), .ZN(P1_U3259) );
  OR2_X1 U13445 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  NAND2_X1 U13446 ( .A1(n10984), .A2(n10983), .ZN(n14703) );
  NAND2_X1 U13447 ( .A1(n14703), .A2(n14745), .ZN(n10991) );
  OAI21_X1 U13448 ( .B1(n10987), .B2(n10986), .A(n10985), .ZN(n10988) );
  NAND2_X1 U13449 ( .A1(n10988), .A2(n13541), .ZN(n10990) );
  NAND3_X1 U13450 ( .A1(n10991), .A2(n10990), .A3(n10989), .ZN(n14701) );
  MUX2_X1 U13451 ( .A(n14701), .B(P2_REG2_REG_4__SCAN_IN), .S(n13402), .Z(
        n10992) );
  INV_X1 U13452 ( .A(n10992), .ZN(n11003) );
  INV_X1 U13453 ( .A(n11364), .ZN(n13420) );
  INV_X1 U13454 ( .A(n10994), .ZN(n14700) );
  AOI21_X1 U13455 ( .B1(n10995), .B2(n10994), .A(n10230), .ZN(n10997) );
  AND2_X1 U13456 ( .A1(n10997), .A2(n10996), .ZN(n14698) );
  NAND2_X1 U13457 ( .A1(n13422), .A2(n14698), .ZN(n11000) );
  OR2_X1 U13458 ( .A1(n13414), .A2(n10998), .ZN(n10999) );
  OAI211_X1 U13459 ( .C1(n14700), .C2(n13417), .A(n11000), .B(n10999), .ZN(
        n11001) );
  AOI21_X1 U13460 ( .B1(n14703), .B2(n13420), .A(n11001), .ZN(n11002) );
  NAND2_X1 U13461 ( .A1(n11003), .A2(n11002), .ZN(P2_U3261) );
  INV_X1 U13462 ( .A(n13680), .ZN(n11589) );
  XNOR2_X1 U13463 ( .A(n11228), .B(n11227), .ZN(n11006) );
  OAI22_X1 U13464 ( .A1(n11589), .A2(n13658), .B1(n11699), .B2(n14356), .ZN(
        n14278) );
  INV_X1 U13465 ( .A(n14278), .ZN(n11005) );
  OAI21_X1 U13466 ( .B1(n11006), .B2(n14566), .A(n11005), .ZN(n14321) );
  INV_X1 U13467 ( .A(n14321), .ZN(n11015) );
  INV_X1 U13468 ( .A(n14010), .ZN(n13987) );
  XNOR2_X1 U13469 ( .A(n11234), .B(n7194), .ZN(n14323) );
  INV_X1 U13470 ( .A(n14276), .ZN(n14320) );
  NAND2_X1 U13471 ( .A1(n14320), .A2(n11009), .ZN(n11237) );
  OAI211_X1 U13472 ( .C1(n14320), .C2(n11009), .A(n14448), .B(n11237), .ZN(
        n14319) );
  OAI22_X1 U13473 ( .A1(n14010), .A2(n11010), .B1(n14281), .B2(n14439), .ZN(
        n11011) );
  AOI21_X1 U13474 ( .B1(n14276), .B2(n14396), .A(n11011), .ZN(n11012) );
  OAI21_X1 U13475 ( .B1(n14319), .B2(n13917), .A(n11012), .ZN(n11013) );
  AOI21_X1 U13476 ( .B1(n14323), .B2(n13953), .A(n11013), .ZN(n11014) );
  OAI21_X1 U13477 ( .B1(n11015), .B2(n13987), .A(n11014), .ZN(P1_U3282) );
  AOI22_X1 U13478 ( .A1(n11027), .A2(n12130), .B1(n12131), .B2(n13683), .ZN(
        n11016) );
  XNOR2_X1 U13479 ( .A(n11016), .B(n12140), .ZN(n11383) );
  NOR2_X1 U13480 ( .A1(n10373), .A2(n11017), .ZN(n11018) );
  AOI21_X1 U13481 ( .B1(n11027), .B2(n12131), .A(n11018), .ZN(n11384) );
  XNOR2_X1 U13482 ( .A(n11383), .B(n11384), .ZN(n11385) );
  INV_X1 U13483 ( .A(n11019), .ZN(n11022) );
  INV_X1 U13484 ( .A(n11020), .ZN(n11021) );
  AOI22_X2 U13485 ( .A1(n11024), .A2(n11023), .B1(n11022), .B2(n11021), .ZN(
        n11386) );
  XOR2_X1 U13486 ( .A(n11386), .B(n11385), .Z(n11031) );
  NAND2_X1 U13487 ( .A1(n13684), .A2(n14353), .ZN(n11026) );
  NAND2_X1 U13488 ( .A1(n13682), .A2(n14003), .ZN(n11025) );
  NAND2_X1 U13489 ( .A1(n11026), .A2(n11025), .ZN(n14407) );
  AND2_X1 U13490 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13750) );
  AOI21_X1 U13491 ( .B1(n14364), .B2(n14407), .A(n13750), .ZN(n11029) );
  NAND2_X1 U13492 ( .A1(n14297), .A2(n11027), .ZN(n11028) );
  OAI211_X1 U13493 ( .C1(n14367), .C2(n14409), .A(n11029), .B(n11028), .ZN(
        n11030) );
  AOI21_X1 U13494 ( .B1(n11031), .B2(n14359), .A(n11030), .ZN(n11032) );
  INV_X1 U13495 ( .A(n11032), .ZN(P1_U3213) );
  MUX2_X1 U13496 ( .A(n11034), .B(n11033), .S(n13406), .Z(n11040) );
  OAI22_X1 U13497 ( .A1(n13417), .A2(n11036), .B1(n13414), .B2(n11035), .ZN(
        n11037) );
  AOI21_X1 U13498 ( .B1(n11038), .B2(n13422), .A(n11037), .ZN(n11039) );
  OAI211_X1 U13499 ( .C1(n11041), .C2(n11364), .A(n11040), .B(n11039), .ZN(
        P2_U3260) );
  MUX2_X1 U13500 ( .A(n11043), .B(n11042), .S(n13406), .Z(n11048) );
  OAI22_X1 U13501 ( .A1(n13417), .A2(n11044), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13414), .ZN(n11045) );
  AOI21_X1 U13502 ( .B1(n11046), .B2(n13422), .A(n11045), .ZN(n11047) );
  OAI211_X1 U13503 ( .C1(n11049), .C2(n11364), .A(n11048), .B(n11047), .ZN(
        P2_U3262) );
  NAND2_X1 U13504 ( .A1(n11050), .A2(n10245), .ZN(n11051) );
  NAND2_X1 U13505 ( .A1(n11052), .A2(n13195), .ZN(n11053) );
  OAI21_X1 U13506 ( .B1(n11056), .B2(n11055), .A(n11270), .ZN(n14708) );
  OAI21_X1 U13507 ( .B1(n11060), .B2(n11059), .A(n11275), .ZN(n11062) );
  AOI21_X1 U13508 ( .B1(n11062), .B2(n13541), .A(n11061), .ZN(n14709) );
  MUX2_X1 U13509 ( .A(n11063), .B(n14709), .S(n13406), .Z(n11071) );
  INV_X1 U13510 ( .A(n11064), .ZN(n11066) );
  INV_X1 U13511 ( .A(n14706), .ZN(n11068) );
  NAND2_X1 U13512 ( .A1(n11068), .A2(n11064), .ZN(n11460) );
  INV_X1 U13513 ( .A(n11460), .ZN(n11065) );
  AOI211_X1 U13514 ( .C1(n14706), .C2(n11066), .A(n10230), .B(n11065), .ZN(
        n14705) );
  OAI22_X1 U13515 ( .A1(n11068), .A2(n13417), .B1(n13414), .B2(n11067), .ZN(
        n11069) );
  AOI21_X1 U13516 ( .B1(n14705), .B2(n13422), .A(n11069), .ZN(n11070) );
  OAI211_X1 U13517 ( .C1(n13411), .C2(n14708), .A(n11071), .B(n11070), .ZN(
        P2_U3259) );
  NAND2_X1 U13518 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  AND2_X1 U13519 ( .A1(n11076), .A2(n11074), .ZN(n11078) );
  XNOR2_X1 U13520 ( .A(n14940), .B(n10097), .ZN(n11255) );
  XNOR2_X1 U13521 ( .A(n11255), .B(n14201), .ZN(n11077) );
  AND2_X1 U13522 ( .A1(n11077), .A2(n11074), .ZN(n11075) );
  OAI211_X1 U13523 ( .C1(n11078), .C2(n11077), .A(n12376), .B(n11257), .ZN(
        n11085) );
  INV_X1 U13524 ( .A(n14936), .ZN(n11771) );
  INV_X1 U13525 ( .A(n11079), .ZN(n14941) );
  NAND2_X1 U13526 ( .A1(n12383), .A2(n14941), .ZN(n11082) );
  INV_X1 U13527 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11080) );
  NOR2_X1 U13528 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11080), .ZN(n14909) );
  AOI21_X1 U13529 ( .B1(n12355), .B2(n14935), .A(n14909), .ZN(n11081) );
  OAI211_X1 U13530 ( .C1(n11771), .C2(n12380), .A(n11082), .B(n11081), .ZN(
        n11083) );
  INV_X1 U13531 ( .A(n11083), .ZN(n11084) );
  OAI211_X1 U13532 ( .C1(n12386), .C2(n14940), .A(n11085), .B(n11084), .ZN(
        P3_U3157) );
  XNOR2_X1 U13533 ( .A(n11086), .B(n12569), .ZN(n11090) );
  INV_X1 U13534 ( .A(n11090), .ZN(n15050) );
  INV_X1 U13535 ( .A(n11087), .ZN(n11088) );
  AOI21_X1 U13536 ( .B1(n12569), .B2(n11089), .A(n11088), .ZN(n11093) );
  AOI22_X1 U13537 ( .A1(n14965), .A2(n12609), .B1(n14935), .B2(n14962), .ZN(
        n11092) );
  NAND2_X1 U13538 ( .A1(n11090), .A2(n14985), .ZN(n11091) );
  OAI211_X1 U13539 ( .C1(n11093), .C2(n14988), .A(n11092), .B(n11091), .ZN(
        n15052) );
  NAND2_X1 U13540 ( .A1(n15052), .A2(n15010), .ZN(n11097) );
  OAI22_X1 U13541 ( .A1(n15010), .A2(n11199), .B1(n11094), .B2(n14978), .ZN(
        n11095) );
  AOI21_X1 U13542 ( .B1(n12878), .B2(n12300), .A(n11095), .ZN(n11096) );
  OAI211_X1 U13543 ( .C1(n15050), .C2(n12794), .A(n11097), .B(n11096), .ZN(
        P3_U3225) );
  INV_X1 U13544 ( .A(n11098), .ZN(n11101) );
  INV_X1 U13545 ( .A(n11099), .ZN(n11100) );
  NAND2_X1 U13546 ( .A1(n11101), .A2(n11100), .ZN(n11102) );
  XNOR2_X1 U13547 ( .A(n11302), .B(n12213), .ZN(n11415) );
  NAND2_X1 U13548 ( .A1(n13189), .A2(n10230), .ZN(n11413) );
  XNOR2_X1 U13549 ( .A(n11415), .B(n11413), .ZN(n11417) );
  XNOR2_X1 U13550 ( .A(n11418), .B(n11417), .ZN(n11111) );
  NOR2_X1 U13551 ( .A1(n14243), .A2(n11288), .ZN(n11109) );
  NAND2_X1 U13552 ( .A1(n13190), .A2(n13141), .ZN(n11106) );
  NAND2_X1 U13553 ( .A1(n13188), .A2(n13139), .ZN(n11105) );
  AND2_X1 U13554 ( .A1(n11106), .A2(n11105), .ZN(n11286) );
  OAI22_X1 U13555 ( .A1(n13143), .A2(n11286), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11107), .ZN(n11108) );
  AOI211_X1 U13556 ( .C1(n11302), .C2(n14240), .A(n11109), .B(n11108), .ZN(
        n11110) );
  OAI21_X1 U13557 ( .B1(n11111), .B2(n13168), .A(n11110), .ZN(P2_U3208) );
  OAI21_X1 U13558 ( .B1(n11114), .B2(n11113), .A(n11112), .ZN(n11115) );
  NAND2_X1 U13559 ( .A1(n11124), .A2(n11115), .ZN(n11116) );
  XNOR2_X1 U13560 ( .A(n11115), .B(n14643), .ZN(n14648) );
  NAND2_X1 U13561 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14648), .ZN(n14647) );
  NAND2_X1 U13562 ( .A1(n14653), .A2(n11117), .ZN(n11118) );
  NAND2_X1 U13563 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14656), .ZN(n14654) );
  NAND2_X1 U13564 ( .A1(n11118), .A2(n14654), .ZN(n11121) );
  XOR2_X1 U13565 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11119), .Z(n11120) );
  OAI211_X1 U13566 ( .C1(n11121), .C2(n11120), .A(n14655), .B(n11324), .ZN(
        n11135) );
  NAND2_X1 U13567 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13104)
         );
  AOI21_X1 U13568 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11123), .A(n11122), 
        .ZN(n14640) );
  XNOR2_X1 U13569 ( .A(n11124), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14641) );
  OR2_X1 U13570 ( .A1(n14640), .A2(n14641), .ZN(n11125) );
  OAI21_X1 U13571 ( .B1(n11126), .B2(n14643), .A(n11125), .ZN(n11127) );
  NAND2_X1 U13572 ( .A1(n14653), .A2(n11127), .ZN(n11129) );
  XNOR2_X1 U13573 ( .A(n11128), .B(n11127), .ZN(n14659) );
  NAND2_X1 U13574 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14659), .ZN(n14657) );
  NAND2_X1 U13575 ( .A1(n11129), .A2(n14657), .ZN(n11131) );
  XNOR2_X1 U13576 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n11326), .ZN(n11130) );
  NAND2_X1 U13577 ( .A1(n11130), .A2(n11131), .ZN(n11316) );
  OAI211_X1 U13578 ( .C1(n11131), .C2(n11130), .A(n14658), .B(n11316), .ZN(
        n11132) );
  NAND2_X1 U13579 ( .A1(n13104), .A2(n11132), .ZN(n11133) );
  AOI21_X1 U13580 ( .B1(n14652), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11133), 
        .ZN(n11134) );
  OAI211_X1 U13581 ( .C1(n14644), .C2(n11326), .A(n11135), .B(n11134), .ZN(
        P2_U3230) );
  INV_X1 U13582 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14204) );
  INV_X1 U13583 ( .A(n14895), .ZN(n11205) );
  NAND2_X1 U13584 ( .A1(n11152), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U13585 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  XNOR2_X1 U13586 ( .A(n11138), .B(n11168), .ZN(n14781) );
  NAND2_X1 U13587 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n14807), .ZN(n11140) );
  OAI21_X1 U13588 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n14807), .A(n11140), .ZN(
        n14799) );
  NOR2_X1 U13589 ( .A1(n11181), .A2(n11141), .ZN(n11142) );
  XNOR2_X1 U13590 ( .A(n11141), .B(n11181), .ZN(n14818) );
  NAND2_X1 U13591 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n14842), .ZN(n11143) );
  OAI21_X1 U13592 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n14842), .A(n11143), .ZN(
        n14834) );
  INV_X1 U13593 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U13594 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n14876), .ZN(n11146) );
  OAI21_X1 U13595 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14876), .A(n11146), .ZN(
        n14869) );
  NOR2_X1 U13596 ( .A1(n11205), .A2(n11147), .ZN(n11148) );
  INV_X1 U13597 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14888) );
  XOR2_X1 U13598 ( .A(n14895), .B(n11147), .Z(n14887) );
  NAND2_X1 U13599 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11213), .ZN(n11149) );
  OAI21_X1 U13600 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11213), .A(n11149), 
        .ZN(n14919) );
  NOR2_X1 U13601 ( .A1(n14204), .A2(n11150), .ZN(n11430) );
  AOI21_X1 U13602 ( .B1(n14204), .B2(n11150), .A(n11430), .ZN(n11226) );
  NAND2_X1 U13603 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11213), .ZN(n11164) );
  INV_X1 U13604 ( .A(n11213), .ZN(n14925) );
  AOI22_X1 U13605 ( .A1(n14925), .A2(n11210), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11213), .ZN(n14908) );
  NAND2_X1 U13606 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n14876), .ZN(n11161) );
  AOI22_X1 U13607 ( .A1(n11200), .A2(n11198), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n14876), .ZN(n14880) );
  NAND2_X1 U13608 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n14842), .ZN(n11158) );
  AOI22_X1 U13609 ( .A1(n11188), .A2(n11186), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n14842), .ZN(n14846) );
  NAND2_X1 U13610 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n14807), .ZN(n11155) );
  AOI22_X1 U13611 ( .A1(n11175), .A2(n11173), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n14807), .ZN(n14811) );
  AOI21_X1 U13612 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n11152), .A(n11151), .ZN(
        n11154) );
  XNOR2_X1 U13613 ( .A(n11154), .B(n14792), .ZN(n14794) );
  NAND2_X1 U13614 ( .A1(n14794), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U13615 ( .A1(n14824), .A2(n11156), .ZN(n11157) );
  NAND2_X1 U13616 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14828), .ZN(n14827) );
  NAND2_X1 U13617 ( .A1(n14859), .A2(n11159), .ZN(n11160) );
  NAND2_X1 U13618 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14863), .ZN(n14862) );
  NAND2_X1 U13619 ( .A1(n11160), .A2(n14862), .ZN(n14881) );
  NAND2_X1 U13620 ( .A1(n14880), .A2(n14881), .ZN(n14879) );
  NAND2_X1 U13621 ( .A1(n11161), .A2(n14879), .ZN(n11162) );
  NAND2_X1 U13622 ( .A1(n14895), .A2(n11162), .ZN(n11163) );
  XNOR2_X1 U13623 ( .A(n11205), .B(n11162), .ZN(n14901) );
  NAND2_X1 U13624 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14901), .ZN(n14900) );
  NAND2_X1 U13625 ( .A1(n11163), .A2(n14900), .ZN(n14907) );
  NAND2_X1 U13626 ( .A1(n14908), .A2(n14907), .ZN(n14906) );
  NAND2_X1 U13627 ( .A1(n11164), .A2(n14906), .ZN(n11434) );
  XNOR2_X1 U13628 ( .A(n11441), .B(n11434), .ZN(n11165) );
  NAND2_X1 U13629 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11165), .ZN(n11436) );
  OAI21_X1 U13630 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11165), .A(n11436), 
        .ZN(n11224) );
  INV_X1 U13631 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11166) );
  MUX2_X1 U13632 ( .A(n11167), .B(n11166), .S(n12729), .Z(n11169) );
  NAND2_X1 U13633 ( .A1(n11169), .A2(n11168), .ZN(n11172) );
  INV_X1 U13634 ( .A(n11169), .ZN(n11170) );
  NAND2_X1 U13635 ( .A1(n11170), .A2(n14792), .ZN(n11171) );
  NAND2_X1 U13636 ( .A1(n11172), .A2(n11171), .ZN(n14786) );
  AOI21_X1 U13637 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14803) );
  INV_X1 U13638 ( .A(n11172), .ZN(n14802) );
  MUX2_X1 U13639 ( .A(n11174), .B(n11173), .S(n12729), .Z(n11176) );
  NAND2_X1 U13640 ( .A1(n11176), .A2(n11175), .ZN(n14820) );
  INV_X1 U13641 ( .A(n11176), .ZN(n11177) );
  NAND2_X1 U13642 ( .A1(n11177), .A2(n14807), .ZN(n11178) );
  AND2_X1 U13643 ( .A1(n14820), .A2(n11178), .ZN(n14801) );
  OAI21_X1 U13644 ( .B1(n14803), .B2(n14802), .A(n14801), .ZN(n14821) );
  MUX2_X1 U13645 ( .A(n11180), .B(n11179), .S(n12729), .Z(n11182) );
  NAND2_X1 U13646 ( .A1(n11182), .A2(n11181), .ZN(n11185) );
  INV_X1 U13647 ( .A(n11182), .ZN(n11183) );
  NAND2_X1 U13648 ( .A1(n11183), .A2(n14824), .ZN(n11184) );
  NAND2_X1 U13649 ( .A1(n11185), .A2(n11184), .ZN(n14819) );
  INV_X1 U13650 ( .A(n11185), .ZN(n14837) );
  MUX2_X1 U13651 ( .A(n11187), .B(n11186), .S(n12729), .Z(n11189) );
  NAND2_X1 U13652 ( .A1(n11189), .A2(n11188), .ZN(n14855) );
  INV_X1 U13653 ( .A(n11189), .ZN(n11190) );
  NAND2_X1 U13654 ( .A1(n11190), .A2(n14842), .ZN(n11191) );
  AND2_X1 U13655 ( .A1(n14855), .A2(n11191), .ZN(n14836) );
  OAI21_X1 U13656 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14856) );
  MUX2_X1 U13657 ( .A(n14958), .B(n11192), .S(n12729), .Z(n11194) );
  NAND2_X1 U13658 ( .A1(n11194), .A2(n11193), .ZN(n11197) );
  INV_X1 U13659 ( .A(n11194), .ZN(n11195) );
  NAND2_X1 U13660 ( .A1(n11195), .A2(n14859), .ZN(n11196) );
  NAND2_X1 U13661 ( .A1(n11197), .A2(n11196), .ZN(n14854) );
  AOI21_X1 U13662 ( .B1(n14856), .B2(n14855), .A(n14854), .ZN(n14872) );
  INV_X1 U13663 ( .A(n11197), .ZN(n14871) );
  MUX2_X1 U13664 ( .A(n11199), .B(n11198), .S(n12729), .Z(n11201) );
  NAND2_X1 U13665 ( .A1(n11201), .A2(n11200), .ZN(n14890) );
  INV_X1 U13666 ( .A(n11201), .ZN(n11202) );
  NAND2_X1 U13667 ( .A1(n11202), .A2(n14876), .ZN(n11203) );
  AND2_X1 U13668 ( .A1(n14890), .A2(n11203), .ZN(n14870) );
  OAI21_X1 U13669 ( .B1(n14872), .B2(n14871), .A(n14870), .ZN(n14891) );
  MUX2_X1 U13670 ( .A(n14888), .B(n11204), .S(n12729), .Z(n11206) );
  NAND2_X1 U13671 ( .A1(n11206), .A2(n11205), .ZN(n11209) );
  INV_X1 U13672 ( .A(n11206), .ZN(n11207) );
  NAND2_X1 U13673 ( .A1(n11207), .A2(n14895), .ZN(n11208) );
  NAND2_X1 U13674 ( .A1(n11209), .A2(n11208), .ZN(n14889) );
  AOI21_X1 U13675 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(n14914) );
  INV_X1 U13676 ( .A(n11209), .ZN(n14913) );
  MUX2_X1 U13677 ( .A(n11211), .B(n11210), .S(n12729), .Z(n11212) );
  NAND2_X1 U13678 ( .A1(n11212), .A2(n14925), .ZN(n11216) );
  INV_X1 U13679 ( .A(n11212), .ZN(n11214) );
  NAND2_X1 U13680 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  AND2_X1 U13681 ( .A1(n11216), .A2(n11215), .ZN(n14912) );
  OAI21_X1 U13682 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n14917) );
  NAND2_X1 U13683 ( .A1(n14917), .A2(n11216), .ZN(n11218) );
  MUX2_X1 U13684 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12729), .Z(n11440) );
  XNOR2_X1 U13685 ( .A(n11440), .B(n11441), .ZN(n11217) );
  NAND2_X1 U13686 ( .A1(n11218), .A2(n11217), .ZN(n11444) );
  OAI21_X1 U13687 ( .B1(n11218), .B2(n11217), .A(n11444), .ZN(n11219) );
  NAND2_X1 U13688 ( .A1(n11219), .A2(n14892), .ZN(n11222) );
  NOR2_X1 U13689 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11220), .ZN(n11259) );
  AOI21_X1 U13690 ( .B1(n14899), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11259), 
        .ZN(n11221) );
  OAI211_X1 U13691 ( .C1(n14896), .C2(n11435), .A(n11222), .B(n11221), .ZN(
        n11223) );
  AOI21_X1 U13692 ( .B1(n14910), .B2(n11224), .A(n11223), .ZN(n11225) );
  OAI21_X1 U13693 ( .B1(n11226), .B2(n14921), .A(n11225), .ZN(P3_U3193) );
  INV_X1 U13694 ( .A(n13679), .ZN(n11229) );
  INV_X1 U13695 ( .A(n11374), .ZN(n11366) );
  XNOR2_X1 U13696 ( .A(n11367), .B(n11366), .ZN(n11233) );
  NAND2_X1 U13697 ( .A1(n13679), .A2(n14353), .ZN(n11231) );
  NAND2_X1 U13698 ( .A1(n13677), .A2(n14003), .ZN(n11230) );
  NAND2_X1 U13699 ( .A1(n11231), .A2(n11230), .ZN(n11710) );
  INV_X1 U13700 ( .A(n11710), .ZN(n11232) );
  OAI21_X1 U13701 ( .B1(n11233), .B2(n14566), .A(n11232), .ZN(n14159) );
  INV_X1 U13702 ( .A(n14159), .ZN(n11243) );
  NAND2_X1 U13703 ( .A1(n11234), .A2(n7194), .ZN(n11236) );
  OR2_X1 U13704 ( .A1(n14276), .A2(n13679), .ZN(n11235) );
  XNOR2_X1 U13705 ( .A(n11375), .B(n11374), .ZN(n14161) );
  INV_X1 U13706 ( .A(n11237), .ZN(n11238) );
  INV_X1 U13707 ( .A(n11701), .ZN(n14158) );
  OAI211_X1 U13708 ( .C1(n11238), .C2(n14158), .A(n14448), .B(n11377), .ZN(
        n14157) );
  OAI22_X1 U13709 ( .A1(n14010), .A2(n10143), .B1(n11707), .B2(n14439), .ZN(
        n11239) );
  AOI21_X1 U13710 ( .B1(n11701), .B2(n14396), .A(n11239), .ZN(n11240) );
  OAI21_X1 U13711 ( .B1(n14157), .B2(n13917), .A(n11240), .ZN(n11241) );
  AOI21_X1 U13712 ( .B1(n14161), .B2(n13953), .A(n11241), .ZN(n11242) );
  OAI21_X1 U13713 ( .B1(n11243), .B2(n13987), .A(n11242), .ZN(P1_U3281) );
  XNOR2_X1 U13714 ( .A(n11244), .B(n12427), .ZN(n15054) );
  OAI211_X1 U13715 ( .C1(n11246), .C2(n12427), .A(n11245), .B(n15001), .ZN(
        n11248) );
  AOI22_X1 U13716 ( .A1(n14950), .A2(n14965), .B1(n14962), .B2(n12608), .ZN(
        n11247) );
  OAI211_X1 U13717 ( .C1(n15004), .C2(n15054), .A(n11248), .B(n11247), .ZN(
        n15055) );
  NAND2_X1 U13718 ( .A1(n15055), .A2(n15010), .ZN(n11254) );
  NOR2_X1 U13719 ( .A1(n11249), .A2(n15047), .ZN(n15056) );
  INV_X1 U13720 ( .A(n15056), .ZN(n11251) );
  OAI22_X1 U13721 ( .A1(n14939), .A2(n11251), .B1(n11250), .B2(n14978), .ZN(
        n11252) );
  AOI21_X1 U13722 ( .B1(n15012), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11252), .ZN(
        n11253) );
  OAI211_X1 U13723 ( .C1(n15054), .C2(n12794), .A(n11254), .B(n11253), .ZN(
        P3_U3224) );
  NAND2_X1 U13724 ( .A1(n11255), .A2(n12608), .ZN(n11256) );
  XNOR2_X1 U13725 ( .A(n11261), .B(n10097), .ZN(n11531) );
  XNOR2_X1 U13726 ( .A(n11531), .B(n11771), .ZN(n11258) );
  XNOR2_X1 U13727 ( .A(n11534), .B(n11258), .ZN(n11267) );
  AOI21_X1 U13728 ( .B1(n12365), .B2(n12607), .A(n11259), .ZN(n11265) );
  INV_X1 U13729 ( .A(n14203), .ZN(n11260) );
  NAND2_X1 U13730 ( .A1(n12383), .A2(n11260), .ZN(n11264) );
  NAND2_X1 U13731 ( .A1(n11261), .A2(n12359), .ZN(n11263) );
  NAND2_X1 U13732 ( .A1(n12355), .A2(n12608), .ZN(n11262) );
  NAND4_X1 U13733 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11266) );
  AOI21_X1 U13734 ( .B1(n11267), .B2(n12376), .A(n11266), .ZN(n11268) );
  INV_X1 U13735 ( .A(n11268), .ZN(P3_U3176) );
  NAND2_X1 U13736 ( .A1(n14706), .A2(n13194), .ZN(n11269) );
  NAND2_X1 U13737 ( .A1(n11270), .A2(n11269), .ZN(n11467) );
  INV_X1 U13738 ( .A(n11455), .ZN(n11466) );
  NAND2_X1 U13739 ( .A1(n14714), .A2(n13193), .ZN(n11271) );
  NAND2_X1 U13740 ( .A1(n14727), .A2(n13191), .ZN(n11272) );
  NAND2_X1 U13741 ( .A1(n14736), .A2(n13190), .ZN(n11273) );
  XNOR2_X1 U13742 ( .A(n11299), .B(n11300), .ZN(n14747) );
  INV_X1 U13743 ( .A(n14747), .ZN(n11293) );
  NAND2_X1 U13744 ( .A1(n11456), .A2(n11455), .ZN(n11454) );
  NAND2_X1 U13745 ( .A1(n14714), .A2(n11276), .ZN(n11277) );
  NAND2_X1 U13746 ( .A1(n11454), .A2(n11277), .ZN(n11473) );
  INV_X1 U13747 ( .A(n11477), .ZN(n11472) );
  NAND2_X1 U13748 ( .A1(n11484), .A2(n11278), .ZN(n11279) );
  OR2_X1 U13749 ( .A1(n14727), .A2(n11281), .ZN(n11280) );
  INV_X1 U13750 ( .A(n11494), .ZN(n11489) );
  NAND2_X1 U13751 ( .A1(n11490), .A2(n11489), .ZN(n11284) );
  NAND2_X1 U13752 ( .A1(n14736), .A2(n11282), .ZN(n11283) );
  NAND2_X1 U13753 ( .A1(n11284), .A2(n11283), .ZN(n11301) );
  XNOR2_X1 U13754 ( .A(n11301), .B(n11300), .ZN(n11285) );
  NAND2_X1 U13755 ( .A1(n11285), .A2(n13541), .ZN(n11287) );
  NAND2_X1 U13756 ( .A1(n11287), .A2(n11286), .ZN(n14752) );
  INV_X1 U13757 ( .A(n11302), .ZN(n14750) );
  INV_X1 U13758 ( .A(n14727), .ZN(n11340) );
  OR2_X1 U13759 ( .A1(n11460), .A2(n14714), .ZN(n11459) );
  INV_X2 U13760 ( .A(n11479), .ZN(n11339) );
  OAI211_X1 U13761 ( .C1(n14750), .C2(n6598), .A(n6486), .B(n11307), .ZN(
        n14748) );
  OAI22_X1 U13762 ( .A1(n13406), .A2(n10163), .B1(n11288), .B2(n13414), .ZN(
        n11289) );
  AOI21_X1 U13763 ( .B1(n11302), .B2(n13399), .A(n11289), .ZN(n11290) );
  OAI21_X1 U13764 ( .B1(n14748), .B2(n13398), .A(n11290), .ZN(n11291) );
  AOI21_X1 U13765 ( .B1(n14752), .B2(n13406), .A(n11291), .ZN(n11292) );
  OAI21_X1 U13766 ( .B1(n13411), .B2(n11293), .A(n11292), .ZN(P2_U3254) );
  OAI222_X1 U13767 ( .A1(n9655), .A2(P3_U3151), .B1(n13058), .B2(n11295), .C1(
        n13056), .C2(n11294), .ZN(P3_U3271) );
  INV_X1 U13768 ( .A(n11296), .ZN(n11345) );
  OAI222_X1 U13769 ( .A1(n14125), .A2(n7162), .B1(n14128), .B2(n11345), .C1(
        n11297), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13770 ( .A(n13189), .ZN(n11305) );
  NAND2_X1 U13771 ( .A1(n14750), .A2(n11305), .ZN(n11298) );
  XOR2_X1 U13772 ( .A(n11304), .B(n11514), .Z(n11569) );
  INV_X1 U13773 ( .A(n11569), .ZN(n11315) );
  NAND2_X1 U13774 ( .A1(n11302), .A2(n11305), .ZN(n11303) );
  XNOR2_X1 U13775 ( .A(n11518), .B(n11304), .ZN(n11306) );
  OAI22_X1 U13776 ( .A1(n11305), .A2(n13163), .B1(n11648), .B2(n13161), .ZN(
        n11426) );
  AOI21_X1 U13777 ( .B1(n11306), .B2(n13541), .A(n11426), .ZN(n11567) );
  INV_X1 U13778 ( .A(n11567), .ZN(n11313) );
  NAND2_X1 U13779 ( .A1(n11307), .A2(n11520), .ZN(n11308) );
  NAND3_X1 U13780 ( .A1(n11522), .A2(n6486), .A3(n11308), .ZN(n11566) );
  OAI22_X1 U13781 ( .A1(n13406), .A2(n11309), .B1(n11423), .B2(n13414), .ZN(
        n11310) );
  AOI21_X1 U13782 ( .B1(n11520), .B2(n13399), .A(n11310), .ZN(n11311) );
  OAI21_X1 U13783 ( .B1(n11566), .B2(n13398), .A(n11311), .ZN(n11312) );
  AOI21_X1 U13784 ( .B1(n11313), .B2(n13406), .A(n11312), .ZN(n11314) );
  OAI21_X1 U13785 ( .B1(n11315), .B2(n13411), .A(n11314), .ZN(P2_U3253) );
  NAND2_X1 U13786 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13114)
         );
  XNOR2_X1 U13787 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13208), .ZN(n11319) );
  OAI21_X1 U13788 ( .B1(n11326), .B2(n11317), .A(n11316), .ZN(n11318) );
  NAND2_X1 U13789 ( .A1(n11319), .A2(n11318), .ZN(n13207) );
  OAI211_X1 U13790 ( .C1(n11319), .C2(n11318), .A(n14658), .B(n13207), .ZN(
        n11320) );
  NAND2_X1 U13791 ( .A1(n13114), .A2(n11320), .ZN(n11321) );
  AOI21_X1 U13792 ( .B1(n14652), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n11321), 
        .ZN(n11330) );
  INV_X1 U13793 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11322) );
  MUX2_X1 U13794 ( .A(n11322), .B(P2_REG2_REG_17__SCAN_IN), .S(n13201), .Z(
        n11323) );
  INV_X1 U13795 ( .A(n11323), .ZN(n11328) );
  INV_X1 U13796 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U13797 ( .A1(n11328), .A2(n11327), .ZN(n13202) );
  OAI211_X1 U13798 ( .C1(n11328), .C2(n11327), .A(n14655), .B(n13202), .ZN(
        n11329) );
  OAI211_X1 U13799 ( .C1(n14644), .C2(n13208), .A(n11330), .B(n11329), .ZN(
        P2_U3231) );
  OAI21_X1 U13800 ( .B1(n11332), .B2(n11333), .A(n11331), .ZN(n14730) );
  XNOR2_X1 U13801 ( .A(n11334), .B(n11333), .ZN(n11336) );
  OAI21_X1 U13802 ( .B1(n11336), .B2(n13529), .A(n11335), .ZN(n14732) );
  NAND2_X1 U13803 ( .A1(n14732), .A2(n13406), .ZN(n11344) );
  OAI22_X1 U13804 ( .A1(n13406), .A2(n11338), .B1(n11337), .B2(n13414), .ZN(
        n11342) );
  OAI211_X1 U13805 ( .C1(n11340), .C2(n11339), .A(n6486), .B(n11498), .ZN(
        n14729) );
  NOR2_X1 U13806 ( .A1(n14729), .A2(n13398), .ZN(n11341) );
  AOI211_X1 U13807 ( .C1(n13399), .C2(n14727), .A(n11342), .B(n11341), .ZN(
        n11343) );
  OAI211_X1 U13808 ( .C1(n13411), .C2(n14730), .A(n11344), .B(n11343), .ZN(
        P2_U3256) );
  OAI222_X1 U13809 ( .A1(n13578), .A2(n7164), .B1(P2_U3088), .B2(n6472), .C1(
        n13581), .C2(n11345), .ZN(P2_U3307) );
  OAI21_X1 U13810 ( .B1(n11349), .B2(n11348), .A(n11347), .ZN(n14696) );
  INV_X1 U13811 ( .A(n14696), .ZN(n11365) );
  OAI22_X1 U13812 ( .A1(n13406), .A2(n8513), .B1(n11350), .B2(n13414), .ZN(
        n11355) );
  OAI21_X1 U13813 ( .B1(n11351), .B2(n14693), .A(n6486), .ZN(n11353) );
  OR2_X1 U13814 ( .A1(n11353), .A2(n11352), .ZN(n14692) );
  NOR2_X1 U13815 ( .A1(n13398), .A2(n14692), .ZN(n11354) );
  AOI211_X1 U13816 ( .C1(n13399), .C2(n11356), .A(n11355), .B(n11354), .ZN(
        n11363) );
  NAND2_X1 U13817 ( .A1(n11359), .A2(n13541), .ZN(n11360) );
  OAI211_X1 U13818 ( .C1(n11365), .C2(n10245), .A(n11361), .B(n11360), .ZN(
        n14694) );
  NAND2_X1 U13819 ( .A1(n14694), .A2(n13406), .ZN(n11362) );
  OAI211_X1 U13820 ( .C1(n11365), .C2(n11364), .A(n11363), .B(n11362), .ZN(
        P2_U3263) );
  OR2_X1 U13821 ( .A1(n11701), .A2(n11699), .ZN(n11368) );
  NAND2_X1 U13822 ( .A1(n11369), .A2(n11368), .ZN(n11610) );
  XNOR2_X1 U13823 ( .A(n11610), .B(n11609), .ZN(n11373) );
  NAND2_X1 U13824 ( .A1(n13676), .A2(n14003), .ZN(n11371) );
  NAND2_X1 U13825 ( .A1(n13678), .A2(n14353), .ZN(n11370) );
  NAND2_X1 U13826 ( .A1(n11371), .A2(n11370), .ZN(n11819) );
  INV_X1 U13827 ( .A(n11819), .ZN(n11372) );
  OAI21_X1 U13828 ( .B1(n11373), .B2(n14566), .A(n11372), .ZN(n14315) );
  INV_X1 U13829 ( .A(n14315), .ZN(n11382) );
  OR2_X1 U13830 ( .A1(n11701), .A2(n13678), .ZN(n11376) );
  INV_X1 U13831 ( .A(n11609), .ZN(n11603) );
  XNOR2_X1 U13832 ( .A(n11604), .B(n11603), .ZN(n14317) );
  OAI211_X1 U13833 ( .C1(n6819), .C2(n6820), .A(n14448), .B(n11607), .ZN(
        n14314) );
  OAI22_X1 U13834 ( .A1(n14010), .A2(n10388), .B1(n11822), .B2(n14439), .ZN(
        n11378) );
  AOI21_X1 U13835 ( .B1(n11824), .B2(n14396), .A(n11378), .ZN(n11379) );
  OAI21_X1 U13836 ( .B1(n14314), .B2(n13917), .A(n11379), .ZN(n11380) );
  AOI21_X1 U13837 ( .B1(n14317), .B2(n13953), .A(n11380), .ZN(n11381) );
  OAI21_X1 U13838 ( .B1(n11382), .B2(n14395), .A(n11381), .ZN(P1_U3280) );
  NAND2_X1 U13839 ( .A1(n14550), .A2(n12130), .ZN(n11388) );
  NAND2_X1 U13840 ( .A1(n12131), .A2(n13682), .ZN(n11387) );
  NAND2_X1 U13841 ( .A1(n11388), .A2(n11387), .ZN(n11389) );
  XNOR2_X1 U13842 ( .A(n11389), .B(n12039), .ZN(n11393) );
  NOR2_X1 U13843 ( .A1(n10373), .A2(n11390), .ZN(n11391) );
  AOI21_X1 U13844 ( .B1(n14550), .B2(n12131), .A(n11391), .ZN(n11392) );
  NAND2_X1 U13845 ( .A1(n11393), .A2(n11392), .ZN(n11394) );
  OAI21_X1 U13846 ( .B1(n11393), .B2(n11392), .A(n11394), .ZN(n11557) );
  AOI22_X1 U13847 ( .A1(n14557), .A2(n12131), .B1(n12135), .B2(n13681), .ZN(
        n11585) );
  NAND2_X1 U13848 ( .A1(n14557), .A2(n12130), .ZN(n11396) );
  NAND2_X1 U13849 ( .A1(n12131), .A2(n13681), .ZN(n11395) );
  NAND2_X1 U13850 ( .A1(n11396), .A2(n11395), .ZN(n11397) );
  XNOR2_X1 U13851 ( .A(n11397), .B(n12140), .ZN(n11587) );
  XOR2_X1 U13852 ( .A(n11585), .B(n11587), .Z(n11398) );
  AOI21_X1 U13853 ( .B1(n11399), .B2(n11398), .A(n11594), .ZN(n11407) );
  INV_X1 U13854 ( .A(n11400), .ZN(n14393) );
  NAND2_X1 U13855 ( .A1(n13682), .A2(n14353), .ZN(n11402) );
  NAND2_X1 U13856 ( .A1(n13680), .A2(n14003), .ZN(n11401) );
  AND2_X1 U13857 ( .A1(n11402), .A2(n11401), .ZN(n14390) );
  OAI21_X1 U13858 ( .B1(n14284), .B2(n14390), .A(n11403), .ZN(n11404) );
  AOI21_X1 U13859 ( .B1(n13653), .B2(n14393), .A(n11404), .ZN(n11406) );
  NAND2_X1 U13860 ( .A1(n14557), .A2(n14297), .ZN(n11405) );
  OAI211_X1 U13861 ( .C1(n11407), .C2(n13663), .A(n11406), .B(n11405), .ZN(
        P1_U3231) );
  XNOR2_X1 U13862 ( .A(n11520), .B(n12205), .ZN(n11408) );
  NAND2_X1 U13863 ( .A1(n13188), .A2(n10230), .ZN(n11409) );
  NAND2_X1 U13864 ( .A1(n11408), .A2(n11409), .ZN(n11545) );
  INV_X1 U13865 ( .A(n11408), .ZN(n11411) );
  INV_X1 U13866 ( .A(n11409), .ZN(n11410) );
  NAND2_X1 U13867 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  AND2_X1 U13868 ( .A1(n11545), .A2(n11412), .ZN(n11420) );
  INV_X1 U13869 ( .A(n11413), .ZN(n11414) );
  AND2_X1 U13870 ( .A1(n11415), .A2(n11414), .ZN(n11416) );
  OAI21_X1 U13871 ( .B1(n11420), .B2(n11419), .A(n11546), .ZN(n11421) );
  NAND2_X1 U13872 ( .A1(n11421), .A2(n14235), .ZN(n11428) );
  INV_X1 U13873 ( .A(n11422), .ZN(n11425) );
  NOR2_X1 U13874 ( .A1(n14243), .A2(n11423), .ZN(n11424) );
  AOI211_X1 U13875 ( .C1(n14237), .C2(n11426), .A(n11425), .B(n11424), .ZN(
        n11427) );
  OAI211_X1 U13876 ( .C1(n6823), .C2(n13149), .A(n11428), .B(n11427), .ZN(
        P2_U3196) );
  NOR2_X1 U13877 ( .A1(n11441), .A2(n11429), .ZN(n11431) );
  AOI22_X1 U13878 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11721), .B1(n11714), 
        .B2(n11773), .ZN(n11432) );
  NOR2_X1 U13879 ( .A1(n11433), .A2(n11432), .ZN(n11713) );
  AOI21_X1 U13880 ( .B1(n11433), .B2(n11432), .A(n11713), .ZN(n11453) );
  AOI22_X1 U13881 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11714), .B1(n11721), 
        .B2(n9305), .ZN(n11439) );
  NAND2_X1 U13882 ( .A1(n11435), .A2(n11434), .ZN(n11437) );
  OAI21_X1 U13883 ( .B1(n11439), .B2(n11438), .A(n11716), .ZN(n11451) );
  INV_X1 U13884 ( .A(n11440), .ZN(n11442) );
  NAND2_X1 U13885 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  AND2_X1 U13886 ( .A1(n11444), .A2(n11443), .ZN(n11446) );
  MUX2_X1 U13887 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12729), .Z(n11718) );
  XNOR2_X1 U13888 ( .A(n11718), .B(n11721), .ZN(n11445) );
  NAND3_X1 U13889 ( .A1(n11444), .A2(n11443), .A3(n11445), .ZN(n11719) );
  OAI211_X1 U13890 ( .C1(n11446), .C2(n11445), .A(n14892), .B(n11719), .ZN(
        n11449) );
  NOR2_X1 U13891 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11447), .ZN(n11538) );
  AOI21_X1 U13892 ( .B1(n14899), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11538), 
        .ZN(n11448) );
  OAI211_X1 U13893 ( .C1(n14896), .C2(n11714), .A(n11449), .B(n11448), .ZN(
        n11450) );
  AOI21_X1 U13894 ( .B1(n11451), .B2(n14910), .A(n11450), .ZN(n11452) );
  OAI21_X1 U13895 ( .B1(n11453), .B2(n14921), .A(n11452), .ZN(P3_U3194) );
  OAI21_X1 U13896 ( .B1(n11456), .B2(n11455), .A(n11454), .ZN(n11458) );
  AOI21_X1 U13897 ( .B1(n11458), .B2(n13541), .A(n11457), .ZN(n14716) );
  INV_X1 U13898 ( .A(n11459), .ZN(n11480) );
  AOI211_X1 U13899 ( .C1(n14714), .C2(n11460), .A(n10230), .B(n11480), .ZN(
        n14713) );
  INV_X1 U13900 ( .A(n11461), .ZN(n11462) );
  INV_X1 U13901 ( .A(n13414), .ZN(n13381) );
  AOI22_X1 U13902 ( .A1(n13402), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11462), 
        .B2(n13381), .ZN(n11463) );
  OAI21_X1 U13903 ( .B1(n11464), .B2(n13417), .A(n11463), .ZN(n11469) );
  OAI21_X1 U13904 ( .B1(n11467), .B2(n11466), .A(n11465), .ZN(n14717) );
  NOR2_X1 U13905 ( .A1(n14717), .A2(n13411), .ZN(n11468) );
  AOI211_X1 U13906 ( .C1(n14713), .C2(n13422), .A(n11469), .B(n11468), .ZN(
        n11470) );
  OAI21_X1 U13907 ( .B1(n13402), .B2(n14716), .A(n11470), .ZN(P2_U3258) );
  OAI21_X1 U13908 ( .B1(n11473), .B2(n11472), .A(n11471), .ZN(n11475) );
  AOI21_X1 U13909 ( .B1(n11475), .B2(n13541), .A(n11474), .ZN(n14721) );
  OAI21_X1 U13910 ( .B1(n11478), .B2(n11477), .A(n11476), .ZN(n14723) );
  INV_X1 U13911 ( .A(n14723), .ZN(n11487) );
  INV_X1 U13912 ( .A(n11484), .ZN(n14722) );
  OAI211_X1 U13913 ( .C1(n14722), .C2(n11480), .A(n6486), .B(n11479), .ZN(
        n14720) );
  OAI22_X1 U13914 ( .A1(n13406), .A2(n11482), .B1(n11481), .B2(n13414), .ZN(
        n11483) );
  AOI21_X1 U13915 ( .B1(n11484), .B2(n13399), .A(n11483), .ZN(n11485) );
  OAI21_X1 U13916 ( .B1(n14720), .B2(n13398), .A(n11485), .ZN(n11486) );
  AOI21_X1 U13917 ( .B1(n11487), .B2(n13365), .A(n11486), .ZN(n11488) );
  OAI21_X1 U13918 ( .B1(n14721), .B2(n13402), .A(n11488), .ZN(P2_U3257) );
  XNOR2_X1 U13919 ( .A(n11490), .B(n11489), .ZN(n11491) );
  NAND2_X1 U13920 ( .A1(n11491), .A2(n13541), .ZN(n11493) );
  NAND2_X1 U13921 ( .A1(n11493), .A2(n11492), .ZN(n14741) );
  INV_X1 U13922 ( .A(n14741), .ZN(n11508) );
  OR2_X1 U13923 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  NAND2_X1 U13924 ( .A1(n11497), .A2(n11496), .ZN(n14740) );
  INV_X1 U13925 ( .A(n14740), .ZN(n11506) );
  NAND2_X1 U13926 ( .A1(n11498), .A2(n14736), .ZN(n11499) );
  NAND2_X1 U13927 ( .A1(n11499), .A2(n6486), .ZN(n11500) );
  OR2_X1 U13928 ( .A1(n6598), .A2(n11500), .ZN(n14738) );
  OAI22_X1 U13929 ( .A1(n13406), .A2(n11502), .B1(n11501), .B2(n13414), .ZN(
        n11503) );
  AOI21_X1 U13930 ( .B1(n14736), .B2(n13399), .A(n11503), .ZN(n11504) );
  OAI21_X1 U13931 ( .B1(n14738), .B2(n13398), .A(n11504), .ZN(n11505) );
  AOI21_X1 U13932 ( .B1(n11506), .B2(n13365), .A(n11505), .ZN(n11507) );
  OAI21_X1 U13933 ( .B1(n11508), .B2(n13402), .A(n11507), .ZN(P2_U3255) );
  INV_X1 U13934 ( .A(n11509), .ZN(n11512) );
  OAI222_X1 U13935 ( .A1(n13578), .A2(n11510), .B1(n13581), .B2(n11512), .C1(
        n8479), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13936 ( .A1(n14125), .A2(n11513), .B1(n14128), .B2(n11512), .C1(
        P1_U3086), .C2(n11511), .ZN(P1_U3334) );
  XNOR2_X1 U13937 ( .A(n11647), .B(n11521), .ZN(n13544) );
  AND2_X1 U13938 ( .A1(n11520), .A2(n11519), .ZN(n11517) );
  XOR2_X1 U13939 ( .A(n11521), .B(n11658), .Z(n13542) );
  AND2_X1 U13940 ( .A1(n13406), .A2(n13541), .ZN(n13409) );
  INV_X1 U13941 ( .A(n11522), .ZN(n11523) );
  NOR2_X1 U13942 ( .A1(n13539), .A2(n11523), .ZN(n11524) );
  OR3_X1 U13943 ( .A1(n11653), .A2(n11524), .A3(n10230), .ZN(n13538) );
  AOI22_X1 U13944 ( .A1(n13186), .A2(n13139), .B1(n13141), .B2(n13188), .ZN(
        n13537) );
  OAI22_X1 U13945 ( .A1(n13402), .A2(n13537), .B1(n11547), .B2(n13414), .ZN(
        n11526) );
  NOR2_X1 U13946 ( .A1(n13539), .A2(n13417), .ZN(n11525) );
  AOI211_X1 U13947 ( .C1(n13402), .C2(P2_REG2_REG_13__SCAN_IN), .A(n11526), 
        .B(n11525), .ZN(n11527) );
  OAI21_X1 U13948 ( .B1(n13398), .B2(n13538), .A(n11527), .ZN(n11528) );
  AOI21_X1 U13949 ( .B1(n13542), .B2(n13409), .A(n11528), .ZN(n11529) );
  OAI21_X1 U13950 ( .B1(n13411), .B2(n13544), .A(n11529), .ZN(P2_U3252) );
  INV_X1 U13951 ( .A(n14221), .ZN(n11544) );
  XNOR2_X1 U13952 ( .A(n14221), .B(n12262), .ZN(n11530) );
  NOR2_X1 U13953 ( .A1(n11530), .A2(n12607), .ZN(n11573) );
  AOI21_X1 U13954 ( .B1(n11530), .B2(n12607), .A(n11573), .ZN(n11536) );
  NAND2_X1 U13955 ( .A1(n11531), .A2(n11771), .ZN(n11533) );
  INV_X1 U13956 ( .A(n11531), .ZN(n11532) );
  OAI21_X1 U13957 ( .B1(n11536), .B2(n11535), .A(n11575), .ZN(n11537) );
  NAND2_X1 U13958 ( .A1(n11537), .A2(n12376), .ZN(n11543) );
  INV_X1 U13959 ( .A(n11772), .ZN(n11541) );
  AOI21_X1 U13960 ( .B1(n12365), .B2(n12606), .A(n11538), .ZN(n11539) );
  OAI21_X1 U13961 ( .B1(n11771), .B2(n12379), .A(n11539), .ZN(n11540) );
  AOI21_X1 U13962 ( .B1(n11541), .B2(n12383), .A(n11540), .ZN(n11542) );
  OAI211_X1 U13963 ( .C1(n11544), .C2(n12386), .A(n11543), .B(n11542), .ZN(
        P3_U3164) );
  XNOR2_X1 U13964 ( .A(n13539), .B(n12205), .ZN(n11844) );
  NOR2_X1 U13965 ( .A1(n11648), .A2(n6486), .ZN(n11843) );
  XNOR2_X1 U13966 ( .A(n11844), .B(n11843), .ZN(n11841) );
  XNOR2_X1 U13967 ( .A(n11840), .B(n11841), .ZN(n11552) );
  NOR2_X1 U13968 ( .A1(n14243), .A2(n11547), .ZN(n11550) );
  OAI21_X1 U13969 ( .B1(n13143), .B2(n13537), .A(n11548), .ZN(n11549) );
  AOI211_X1 U13970 ( .C1(n11649), .C2(n14240), .A(n11550), .B(n11549), .ZN(
        n11551) );
  OAI21_X1 U13971 ( .B1(n11552), .B2(n13168), .A(n11551), .ZN(P2_U3206) );
  AOI21_X1 U13972 ( .B1(n14364), .B2(n14548), .A(n11553), .ZN(n11554) );
  OAI21_X1 U13973 ( .B1(n14367), .B2(n11555), .A(n11554), .ZN(n11561) );
  AOI21_X1 U13974 ( .B1(n11558), .B2(n11557), .A(n11556), .ZN(n11559) );
  NOR2_X1 U13975 ( .A1(n11559), .A2(n13663), .ZN(n11560) );
  AOI211_X1 U13976 ( .C1(n14297), .C2(n14550), .A(n11561), .B(n11560), .ZN(
        n11562) );
  INV_X1 U13977 ( .A(n11562), .ZN(P1_U3221) );
  INV_X1 U13978 ( .A(n11563), .ZN(n11564) );
  OAI222_X1 U13979 ( .A1(n13578), .A2(n11565), .B1(n13581), .B2(n11564), .C1(
        n8487), .C2(P2_U3088), .ZN(P2_U3305) );
  OAI211_X1 U13980 ( .C1(n6823), .C2(n14749), .A(n11567), .B(n11566), .ZN(
        n11568) );
  AOI21_X1 U13981 ( .B1(n11569), .B2(n13525), .A(n11568), .ZN(n11572) );
  NAND2_X1 U13982 ( .A1(n14766), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11570) );
  OAI21_X1 U13983 ( .B1(n11572), .B2(n14766), .A(n11570), .ZN(P2_U3511) );
  NAND2_X1 U13984 ( .A1(n14755), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11571) );
  OAI21_X1 U13985 ( .B1(n11572), .B2(n14755), .A(n11571), .ZN(P2_U3466) );
  INV_X1 U13986 ( .A(n11573), .ZN(n11574) );
  NAND2_X1 U13987 ( .A1(n11575), .A2(n11574), .ZN(n11635) );
  XNOR2_X1 U13988 ( .A(n14193), .B(n10097), .ZN(n11576) );
  NOR2_X1 U13989 ( .A1(n11576), .A2(n12606), .ZN(n11634) );
  INV_X1 U13990 ( .A(n11634), .ZN(n11577) );
  NAND2_X1 U13991 ( .A1(n11576), .A2(n12606), .ZN(n11633) );
  NAND2_X1 U13992 ( .A1(n11577), .A2(n11633), .ZN(n11578) );
  XNOR2_X1 U13993 ( .A(n11635), .B(n11578), .ZN(n11584) );
  AND2_X1 U13994 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11726) );
  AOI21_X1 U13995 ( .B1(n12365), .B2(n12605), .A(n11726), .ZN(n11579) );
  OAI21_X1 U13996 ( .B1(n14202), .B2(n12379), .A(n11579), .ZN(n11581) );
  NOR2_X1 U13997 ( .A1(n14193), .A2(n12386), .ZN(n11580) );
  AOI211_X1 U13998 ( .C1(n11582), .C2(n12383), .A(n11581), .B(n11580), .ZN(
        n11583) );
  OAI21_X1 U13999 ( .B1(n11584), .B2(n12371), .A(n11583), .ZN(P3_U3174) );
  INV_X1 U14000 ( .A(n11585), .ZN(n11586) );
  NOR2_X1 U14001 ( .A1(n11587), .A2(n11586), .ZN(n11593) );
  AOI22_X1 U14002 ( .A1(n11591), .A2(n12130), .B1(n12131), .B2(n13680), .ZN(
        n11588) );
  XNOR2_X1 U14003 ( .A(n11588), .B(n12140), .ZN(n11692) );
  NOR2_X1 U14004 ( .A1(n10373), .A2(n11589), .ZN(n11590) );
  AOI21_X1 U14005 ( .B1(n11591), .B2(n12131), .A(n11590), .ZN(n11691) );
  XNOR2_X1 U14006 ( .A(n11692), .B(n11691), .ZN(n11592) );
  INV_X1 U14007 ( .A(n11693), .ZN(n11596) );
  OAI21_X1 U14008 ( .B1(n11594), .B2(n11593), .A(n11592), .ZN(n11595) );
  NAND3_X1 U14009 ( .A1(n11596), .A2(n14359), .A3(n11595), .ZN(n11602) );
  AOI21_X1 U14010 ( .B1(n11597), .B2(n14568), .A(n14284), .ZN(n11600) );
  NOR2_X1 U14011 ( .A1(n14367), .A2(n11598), .ZN(n11599) );
  AOI211_X1 U14012 ( .C1(P1_REG3_REG_10__SCAN_IN), .C2(P1_U3086), .A(n11600), 
        .B(n11599), .ZN(n11601) );
  OAI211_X1 U14013 ( .C1(n14571), .C2(n14286), .A(n11602), .B(n11601), .ZN(
        P1_U3217) );
  INV_X1 U14014 ( .A(n11615), .ZN(n11606) );
  OR2_X1 U14015 ( .A1(n11824), .A2(n13677), .ZN(n11605) );
  OAI21_X1 U14016 ( .B1(n11606), .B2(n6601), .A(n11666), .ZN(n11688) );
  AOI211_X1 U14017 ( .C1(n14247), .C2(n11607), .A(n14492), .B(n6818), .ZN(
        n11685) );
  INV_X1 U14018 ( .A(n11685), .ZN(n11617) );
  INV_X1 U14019 ( .A(n14252), .ZN(n11608) );
  INV_X1 U14020 ( .A(n13677), .ZN(n11611) );
  OAI22_X1 U14021 ( .A1(n12055), .A2(n14356), .B1(n11611), .B2(n13658), .ZN(
        n14249) );
  AOI21_X1 U14022 ( .B1(n14394), .B2(n11608), .A(n14249), .ZN(n11616) );
  NAND2_X1 U14023 ( .A1(n11610), .A2(n11609), .ZN(n11613) );
  OR2_X1 U14024 ( .A1(n11824), .A2(n11611), .ZN(n11612) );
  NAND2_X1 U14025 ( .A1(n11613), .A2(n11612), .ZN(n11614) );
  NAND2_X1 U14026 ( .A1(n11615), .A2(n11614), .ZN(n11663) );
  OAI211_X1 U14027 ( .C1(n11615), .C2(n11614), .A(n11663), .B(n14522), .ZN(
        n11686) );
  OAI211_X1 U14028 ( .C1(n11617), .C2(n13964), .A(n11616), .B(n11686), .ZN(
        n11618) );
  NAND2_X1 U14029 ( .A1(n11618), .A2(n14010), .ZN(n11620) );
  AOI22_X1 U14030 ( .A1(n14247), .A2(n14396), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n13987), .ZN(n11619) );
  OAI211_X1 U14031 ( .C1(n13998), .C2(n11688), .A(n11620), .B(n11619), .ZN(
        P1_U3279) );
  INV_X1 U14032 ( .A(n11625), .ZN(n11623) );
  NAND2_X1 U14033 ( .A1(n14114), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11621) );
  OAI211_X1 U14034 ( .C1(n11623), .C2(n14128), .A(n11622), .B(n11621), .ZN(
        P1_U3332) );
  NAND2_X1 U14035 ( .A1(n11625), .A2(n11624), .ZN(n11627) );
  OAI211_X1 U14036 ( .C1(n11628), .C2(n13578), .A(n11627), .B(n11626), .ZN(
        P2_U3304) );
  INV_X1 U14037 ( .A(n11629), .ZN(n11630) );
  OAI222_X1 U14038 ( .A1(n11632), .A2(P3_U3151), .B1(n13058), .B2(n11631), 
        .C1(n13056), .C2(n11630), .ZN(P3_U3270) );
  OAI21_X1 U14039 ( .B1(n11635), .B2(n11634), .A(n11633), .ZN(n11637) );
  XNOR2_X1 U14040 ( .A(n11912), .B(n10097), .ZN(n11673) );
  XNOR2_X1 U14041 ( .A(n11673), .B(n14188), .ZN(n11636) );
  NAND2_X1 U14042 ( .A1(n11637), .A2(n11636), .ZN(n11675) );
  OAI211_X1 U14043 ( .C1(n11637), .C2(n11636), .A(n11675), .B(n12376), .ZN(
        n11642) );
  INV_X1 U14044 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11638) );
  NOR2_X1 U14045 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11638), .ZN(n12632) );
  AOI21_X1 U14046 ( .B1(n12365), .B2(n12604), .A(n12632), .ZN(n11639) );
  OAI21_X1 U14047 ( .B1(n7359), .B2(n12379), .A(n11639), .ZN(n11640) );
  AOI21_X1 U14048 ( .B1(n11832), .B2(n12383), .A(n11640), .ZN(n11641) );
  OAI211_X1 U14049 ( .C1(n12386), .C2(n11912), .A(n11642), .B(n11641), .ZN(
        P3_U3155) );
  INV_X1 U14050 ( .A(n11643), .ZN(n11644) );
  OAI222_X1 U14051 ( .A1(n11646), .A2(P3_U3151), .B1(n13058), .B2(n11645), 
        .C1(n13056), .C2(n11644), .ZN(P3_U3269) );
  XOR2_X1 U14052 ( .A(n11741), .B(n11659), .Z(n13536) );
  AOI22_X1 U14053 ( .A1(n13139), .A2(n13185), .B1(n13187), .B2(n13141), .ZN(
        n13530) );
  INV_X1 U14054 ( .A(n13530), .ZN(n14238) );
  INV_X1 U14055 ( .A(n14242), .ZN(n11650) );
  AOI22_X1 U14056 ( .A1(n14238), .A2(n13406), .B1(n11650), .B2(n13381), .ZN(
        n11651) );
  OAI21_X1 U14057 ( .B1(n11652), .B2(n13406), .A(n11651), .ZN(n11656) );
  NOR2_X1 U14058 ( .A1(n13532), .A2(n11653), .ZN(n11654) );
  OR3_X1 U14059 ( .A1(n11743), .A2(n11654), .A3(n10230), .ZN(n13531) );
  NOR2_X1 U14060 ( .A1(n13531), .A2(n13398), .ZN(n11655) );
  AOI211_X1 U14061 ( .C1(n13399), .C2(n14239), .A(n11656), .B(n11655), .ZN(
        n11661) );
  AND2_X1 U14062 ( .A1(n13539), .A2(n13187), .ZN(n11657) );
  XOR2_X1 U14063 ( .A(n11659), .B(n11740), .Z(n13534) );
  NAND2_X1 U14064 ( .A1(n13534), .A2(n13409), .ZN(n11660) );
  OAI211_X1 U14065 ( .C1(n13536), .C2(n13411), .A(n11661), .B(n11660), .ZN(
        P2_U3251) );
  NAND2_X1 U14066 ( .A1(n11663), .A2(n11662), .ZN(n11794) );
  XNOR2_X1 U14067 ( .A(n11794), .B(n11667), .ZN(n11664) );
  INV_X1 U14068 ( .A(n13674), .ZN(n11866) );
  OAI22_X1 U14069 ( .A1(n11866), .A2(n14356), .B1(n12041), .B2(n13658), .ZN(
        n14300) );
  AOI21_X1 U14070 ( .B1(n11664), .B2(n14522), .A(n14300), .ZN(n14310) );
  NAND2_X1 U14071 ( .A1(n14247), .A2(n13676), .ZN(n11665) );
  INV_X1 U14072 ( .A(n11667), .ZN(n11793) );
  XNOR2_X1 U14073 ( .A(n11792), .B(n11793), .ZN(n14313) );
  OAI211_X1 U14074 ( .C1(n6817), .C2(n6818), .A(n14448), .B(n11798), .ZN(
        n14309) );
  OAI22_X1 U14075 ( .A1(n14010), .A2(n11668), .B1(n14302), .B2(n14439), .ZN(
        n11669) );
  AOI21_X1 U14076 ( .B1(n14298), .B2(n14396), .A(n11669), .ZN(n11670) );
  OAI21_X1 U14077 ( .B1(n14309), .B2(n13917), .A(n11670), .ZN(n11671) );
  AOI21_X1 U14078 ( .B1(n14313), .B2(n13953), .A(n11671), .ZN(n11672) );
  OAI21_X1 U14079 ( .B1(n14310), .B2(n14395), .A(n11672), .ZN(P1_U3278) );
  NAND2_X1 U14080 ( .A1(n11673), .A2(n12605), .ZN(n11674) );
  NAND2_X1 U14081 ( .A1(n11675), .A2(n11674), .ZN(n11753) );
  XNOR2_X1 U14082 ( .A(n11889), .B(n10097), .ZN(n11754) );
  XNOR2_X1 U14083 ( .A(n11754), .B(n12604), .ZN(n11676) );
  XNOR2_X1 U14084 ( .A(n11753), .B(n11676), .ZN(n11682) );
  NAND2_X1 U14085 ( .A1(n12383), .A2(n11890), .ZN(n11679) );
  NOR2_X1 U14086 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11677), .ZN(n12653) );
  AOI21_X1 U14087 ( .B1(n12355), .B2(n12605), .A(n12653), .ZN(n11678) );
  OAI211_X1 U14088 ( .C1(n12229), .C2(n12380), .A(n11679), .B(n11678), .ZN(
        n11680) );
  AOI21_X1 U14089 ( .B1(n11889), .B2(n12359), .A(n11680), .ZN(n11681) );
  OAI21_X1 U14090 ( .B1(n11682), .B2(n12371), .A(n11681), .ZN(P3_U3181) );
  INV_X1 U14091 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11690) );
  AOI211_X1 U14092 ( .C1(n14549), .C2(n14247), .A(n14249), .B(n11685), .ZN(
        n11687) );
  OAI211_X1 U14093 ( .C1(n14517), .C2(n11688), .A(n11687), .B(n11686), .ZN(
        n11733) );
  NAND2_X1 U14094 ( .A1(n11733), .A2(n14578), .ZN(n11689) );
  OAI21_X1 U14095 ( .B1(n14578), .B2(n11690), .A(n11689), .ZN(P1_U3501) );
  INV_X1 U14096 ( .A(n11691), .ZN(n11695) );
  INV_X1 U14097 ( .A(n11692), .ZN(n11694) );
  AOI22_X1 U14098 ( .A1(n14276), .A2(n12131), .B1(n12135), .B2(n13679), .ZN(
        n11697) );
  AOI22_X1 U14099 ( .A1(n14276), .A2(n12130), .B1(n12131), .B2(n13679), .ZN(
        n11696) );
  XNOR2_X1 U14100 ( .A(n11696), .B(n12140), .ZN(n11698) );
  XOR2_X1 U14101 ( .A(n11697), .B(n11698), .Z(n14275) );
  NAND2_X1 U14102 ( .A1(n11698), .A2(n11697), .ZN(n11703) );
  AND2_X1 U14103 ( .A1(n14273), .A2(n11703), .ZN(n11706) );
  NOR2_X1 U14104 ( .A1(n10373), .A2(n11699), .ZN(n11700) );
  AOI21_X1 U14105 ( .B1(n11701), .B2(n12131), .A(n11700), .ZN(n11811) );
  AOI22_X1 U14106 ( .A1(n11701), .A2(n12130), .B1(n12131), .B2(n13678), .ZN(
        n11702) );
  XNOR2_X1 U14107 ( .A(n11702), .B(n12140), .ZN(n11810) );
  XOR2_X1 U14108 ( .A(n11811), .B(n11810), .Z(n11705) );
  NAND2_X1 U14109 ( .A1(n14273), .A2(n11704), .ZN(n11815) );
  OAI211_X1 U14110 ( .C1(n11706), .C2(n11705), .A(n14359), .B(n11815), .ZN(
        n11712) );
  NOR2_X1 U14111 ( .A1(n14367), .A2(n11707), .ZN(n11708) );
  AOI211_X1 U14112 ( .C1(n14364), .C2(n11710), .A(n11709), .B(n11708), .ZN(
        n11711) );
  OAI211_X1 U14113 ( .C1(n14158), .C2(n14286), .A(n11712), .B(n11711), .ZN(
        P1_U3224) );
  INV_X1 U14114 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14190) );
  INV_X1 U14115 ( .A(n12617), .ZN(n12625) );
  AOI21_X1 U14116 ( .B1(n14190), .B2(n11715), .A(n12614), .ZN(n11732) );
  NAND2_X1 U14117 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11717), .ZN(n12618) );
  OAI21_X1 U14118 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11717), .A(n12618), 
        .ZN(n11730) );
  MUX2_X1 U14119 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12729), .Z(n12622) );
  XNOR2_X1 U14120 ( .A(n12617), .B(n12622), .ZN(n11723) );
  INV_X1 U14121 ( .A(n11718), .ZN(n11720) );
  OAI21_X1 U14122 ( .B1(n11721), .B2(n11720), .A(n11719), .ZN(n11722) );
  NOR2_X1 U14123 ( .A1(n11722), .A2(n11723), .ZN(n12623) );
  AOI21_X1 U14124 ( .B1(n11723), .B2(n11722), .A(n12623), .ZN(n11728) );
  NOR2_X1 U14125 ( .A1(n14930), .A2(n11724), .ZN(n11725) );
  AOI211_X1 U14126 ( .C1(n14926), .C2(n12625), .A(n11726), .B(n11725), .ZN(
        n11727) );
  OAI21_X1 U14127 ( .B1(n11728), .B2(n14915), .A(n11727), .ZN(n11729) );
  AOI21_X1 U14128 ( .B1(n11730), .B2(n14910), .A(n11729), .ZN(n11731) );
  OAI21_X1 U14129 ( .B1(n11732), .B2(n14921), .A(n11731), .ZN(P3_U3195) );
  NAND2_X1 U14130 ( .A1(n11733), .A2(n14594), .ZN(n11734) );
  OAI21_X1 U14131 ( .B1(n14594), .B2(n8095), .A(n11734), .ZN(P1_U3542) );
  INV_X1 U14132 ( .A(n11735), .ZN(n11737) );
  OAI222_X1 U14133 ( .A1(n12729), .A2(P3_U3151), .B1(n13056), .B2(n11737), 
        .C1(n11736), .C2(n13058), .ZN(P3_U3268) );
  NOR2_X1 U14134 ( .A1(n13532), .A2(n13186), .ZN(n11739) );
  NAND2_X1 U14135 ( .A1(n13532), .A2(n13186), .ZN(n11738) );
  XNOR2_X1 U14136 ( .A(n11783), .B(n11742), .ZN(n13528) );
  INV_X1 U14137 ( .A(n11742), .ZN(n11779) );
  XNOR2_X1 U14138 ( .A(n11780), .B(n11779), .ZN(n13526) );
  OAI211_X1 U14139 ( .C1(n11743), .C2(n13523), .A(n6486), .B(n11784), .ZN(
        n13522) );
  AOI22_X1 U14140 ( .A1(n13186), .A2(n13141), .B1(n13184), .B2(n13139), .ZN(
        n13521) );
  INV_X1 U14141 ( .A(n13521), .ZN(n11744) );
  AOI22_X1 U14142 ( .A1(n11744), .A2(n13406), .B1(n11858), .B2(n13381), .ZN(
        n11745) );
  OAI21_X1 U14143 ( .B1(n11746), .B2(n13406), .A(n11745), .ZN(n11747) );
  AOI21_X1 U14144 ( .B1(n11748), .B2(n13399), .A(n11747), .ZN(n11749) );
  OAI21_X1 U14145 ( .B1(n13522), .B2(n13398), .A(n11749), .ZN(n11750) );
  AOI21_X1 U14146 ( .B1(n13526), .B2(n13365), .A(n11750), .ZN(n11751) );
  OAI21_X1 U14147 ( .B1(n13375), .B2(n13528), .A(n11751), .ZN(P2_U3250) );
  NAND2_X1 U14148 ( .A1(n11754), .A2(n12921), .ZN(n11752) );
  NAND2_X1 U14149 ( .A1(n11753), .A2(n11752), .ZN(n11757) );
  INV_X1 U14150 ( .A(n11754), .ZN(n11755) );
  XNOR2_X1 U14151 ( .A(n12925), .B(n10097), .ZN(n12230) );
  XNOR2_X1 U14152 ( .A(n12230), .B(n12229), .ZN(n11758) );
  XNOR2_X1 U14153 ( .A(n11759), .B(n11758), .ZN(n11765) );
  NOR2_X1 U14154 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11760), .ZN(n12681) );
  AOI21_X1 U14155 ( .B1(n12365), .B2(n12602), .A(n12681), .ZN(n11762) );
  NAND2_X1 U14156 ( .A1(n12383), .A2(n12926), .ZN(n11761) );
  OAI211_X1 U14157 ( .C1(n12921), .C2(n12379), .A(n11762), .B(n11761), .ZN(
        n11763) );
  AOI21_X1 U14158 ( .B1(n12925), .B2(n12359), .A(n11763), .ZN(n11764) );
  OAI21_X1 U14159 ( .B1(n11765), .B2(n12371), .A(n11764), .ZN(P3_U3166) );
  NAND2_X1 U14160 ( .A1(n15004), .A2(n11766), .ZN(n14953) );
  INV_X1 U14161 ( .A(n12930), .ZN(n14209) );
  XNOR2_X1 U14162 ( .A(n11767), .B(n11769), .ZN(n14218) );
  XNOR2_X1 U14163 ( .A(n11768), .B(n11769), .ZN(n11770) );
  OAI222_X1 U14164 ( .A1(n14996), .A2(n7359), .B1(n14998), .B2(n11771), .C1(
        n11770), .C2(n14988), .ZN(n14219) );
  NAND2_X1 U14165 ( .A1(n14219), .A2(n15010), .ZN(n11776) );
  OAI22_X1 U14166 ( .A1(n15010), .A2(n11773), .B1(n11772), .B2(n14978), .ZN(
        n11774) );
  AOI21_X1 U14167 ( .B1(n12878), .B2(n14221), .A(n11774), .ZN(n11775) );
  OAI211_X1 U14168 ( .C1(n14209), .C2(n14218), .A(n11776), .B(n11775), .ZN(
        P3_U3221) );
  INV_X1 U14169 ( .A(n11777), .ZN(n11838) );
  AOI22_X1 U14170 ( .A1(n10257), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n14114), .ZN(n11778) );
  OAI21_X1 U14171 ( .B1(n11838), .B2(n14128), .A(n11778), .ZN(P1_U3331) );
  NAND2_X1 U14172 ( .A1(n11781), .A2(n11949), .ZN(n11930) );
  OAI21_X1 U14173 ( .B1(n11781), .B2(n11949), .A(n11930), .ZN(n13520) );
  AND2_X1 U14174 ( .A1(n13523), .A2(n13185), .ZN(n11782) );
  XOR2_X1 U14175 ( .A(n11949), .B(n11950), .Z(n13518) );
  AOI21_X1 U14176 ( .B1(n11784), .B2(n12157), .A(n10230), .ZN(n11785) );
  NAND2_X1 U14177 ( .A1(n11785), .A2(n13395), .ZN(n13515) );
  AOI22_X1 U14178 ( .A1(n13183), .A2(n13139), .B1(n13185), .B2(n13141), .ZN(
        n13514) );
  OAI22_X1 U14179 ( .A1(n13514), .A2(n13402), .B1(n13103), .B2(n13414), .ZN(
        n11787) );
  NOR2_X1 U14180 ( .A1(n13516), .A2(n13417), .ZN(n11786) );
  AOI211_X1 U14181 ( .C1(n13402), .C2(P2_REG2_REG_16__SCAN_IN), .A(n11787), 
        .B(n11786), .ZN(n11788) );
  OAI21_X1 U14182 ( .B1(n13515), .B2(n13398), .A(n11788), .ZN(n11789) );
  AOI21_X1 U14183 ( .B1(n13518), .B2(n13409), .A(n11789), .ZN(n11790) );
  OAI21_X1 U14184 ( .B1(n13520), .B2(n13411), .A(n11790), .ZN(P2_U3249) );
  INV_X1 U14185 ( .A(n12055), .ZN(n13675) );
  OR2_X1 U14186 ( .A1(n14298), .A2(n13675), .ZN(n11791) );
  XNOR2_X1 U14187 ( .A(n11862), .B(n11797), .ZN(n11899) );
  NAND2_X1 U14188 ( .A1(n11794), .A2(n11793), .ZN(n11796) );
  INV_X1 U14189 ( .A(n11797), .ZN(n11861) );
  OAI21_X1 U14190 ( .B1(n7387), .B2(n11797), .A(n11868), .ZN(n11896) );
  INV_X1 U14191 ( .A(n14256), .ZN(n11807) );
  NAND2_X1 U14192 ( .A1(n11798), .A2(n14256), .ZN(n11799) );
  NAND2_X1 U14193 ( .A1(n11799), .A2(n14448), .ZN(n11800) );
  NOR2_X1 U14194 ( .A1(n11873), .A2(n11800), .ZN(n11895) );
  NAND2_X1 U14195 ( .A1(n11895), .A2(n14452), .ZN(n11806) );
  NAND2_X1 U14196 ( .A1(n14002), .A2(n14003), .ZN(n11802) );
  NAND2_X1 U14197 ( .A1(n13675), .A2(n14353), .ZN(n11801) );
  NAND2_X1 U14198 ( .A1(n11802), .A2(n11801), .ZN(n14258) );
  INV_X1 U14199 ( .A(n14258), .ZN(n11803) );
  OAI22_X1 U14200 ( .A1(n14441), .A2(n11803), .B1(n14261), .B2(n14439), .ZN(
        n11804) );
  AOI21_X1 U14201 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14395), .A(n11804), 
        .ZN(n11805) );
  OAI211_X1 U14202 ( .C1(n11807), .C2(n14444), .A(n11806), .B(n11805), .ZN(
        n11808) );
  AOI21_X1 U14203 ( .B1(n11896), .B2(n13995), .A(n11808), .ZN(n11809) );
  OAI21_X1 U14204 ( .B1(n13998), .B2(n11899), .A(n11809), .ZN(P1_U3277) );
  INV_X1 U14205 ( .A(n11810), .ZN(n11813) );
  INV_X1 U14206 ( .A(n11811), .ZN(n11812) );
  NAND2_X1 U14207 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NAND2_X1 U14208 ( .A1(n11815), .A2(n11814), .ZN(n12036) );
  NAND2_X1 U14209 ( .A1(n11824), .A2(n12130), .ZN(n11817) );
  NAND2_X1 U14210 ( .A1(n12131), .A2(n13677), .ZN(n11816) );
  NAND2_X1 U14211 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  XNOR2_X1 U14212 ( .A(n11818), .B(n12140), .ZN(n12033) );
  AOI22_X1 U14213 ( .A1(n11824), .A2(n12131), .B1(n12135), .B2(n13677), .ZN(
        n12032) );
  XNOR2_X1 U14214 ( .A(n12033), .B(n12032), .ZN(n12035) );
  XNOR2_X1 U14215 ( .A(n12036), .B(n12035), .ZN(n11826) );
  NAND2_X1 U14216 ( .A1(n14364), .A2(n11819), .ZN(n11820) );
  OAI211_X1 U14217 ( .C1(n14367), .C2(n11822), .A(n11821), .B(n11820), .ZN(
        n11823) );
  AOI21_X1 U14218 ( .B1(n11824), .B2(n14297), .A(n11823), .ZN(n11825) );
  OAI21_X1 U14219 ( .B1(n11826), .B2(n13663), .A(n11825), .ZN(P1_U3234) );
  OAI211_X1 U14220 ( .C1(n11828), .C2(n9353), .A(n15001), .B(n11827), .ZN(
        n11830) );
  AOI22_X1 U14221 ( .A1(n12604), .A2(n14962), .B1(n14965), .B2(n12606), .ZN(
        n11829) );
  NAND2_X1 U14222 ( .A1(n11830), .A2(n11829), .ZN(n11905) );
  INV_X1 U14223 ( .A(n11905), .ZN(n11836) );
  XNOR2_X1 U14224 ( .A(n11831), .B(n9353), .ZN(n11906) );
  AOI22_X1 U14225 ( .A1(n15012), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15007), 
        .B2(n11832), .ZN(n11833) );
  OAI21_X1 U14226 ( .B1(n11912), .B2(n12928), .A(n11833), .ZN(n11834) );
  AOI21_X1 U14227 ( .B1(n11906), .B2(n12930), .A(n11834), .ZN(n11835) );
  OAI21_X1 U14228 ( .B1(n11836), .B2(n15012), .A(n11835), .ZN(P3_U3219) );
  OAI222_X1 U14229 ( .A1(n13578), .A2(n11839), .B1(n13581), .B2(n11838), .C1(
        P2_U3088), .C2(n11837), .ZN(P2_U3303) );
  INV_X1 U14230 ( .A(n11841), .ZN(n11842) );
  NAND2_X1 U14231 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  XNOR2_X1 U14232 ( .A(n13532), .B(n12213), .ZN(n11847) );
  OR2_X1 U14233 ( .A1(n11846), .A2(n6486), .ZN(n11848) );
  NAND2_X1 U14234 ( .A1(n11847), .A2(n11848), .ZN(n11853) );
  INV_X1 U14235 ( .A(n11847), .ZN(n11850) );
  INV_X1 U14236 ( .A(n11848), .ZN(n11849) );
  NAND2_X1 U14237 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U14238 ( .A1(n11853), .A2(n11851), .ZN(n14231) );
  XNOR2_X1 U14239 ( .A(n13523), .B(n12205), .ZN(n12151) );
  XNOR2_X2 U14240 ( .A(n12153), .B(n12151), .ZN(n12156) );
  NOR2_X1 U14241 ( .A1(n11854), .A2(n6486), .ZN(n12155) );
  XNOR2_X1 U14242 ( .A(n12156), .B(n12155), .ZN(n11860) );
  INV_X1 U14243 ( .A(n14243), .ZN(n13145) );
  OAI22_X1 U14244 ( .A1(n13143), .A2(n13521), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11855), .ZN(n11857) );
  NOR2_X1 U14245 ( .A1(n13523), .A2(n13149), .ZN(n11856) );
  AOI211_X1 U14246 ( .C1(n13145), .C2(n11858), .A(n11857), .B(n11856), .ZN(
        n11859) );
  OAI21_X1 U14247 ( .B1(n11860), .B2(n13168), .A(n11859), .ZN(P2_U3213) );
  NAND2_X1 U14248 ( .A1(n11862), .A2(n11861), .ZN(n11864) );
  OR2_X1 U14249 ( .A1(n14256), .A2(n13674), .ZN(n11863) );
  XNOR2_X1 U14250 ( .A(n12007), .B(n11869), .ZN(n14303) );
  INV_X1 U14251 ( .A(n14303), .ZN(n11879) );
  NAND2_X1 U14252 ( .A1(n14256), .A2(n11866), .ZN(n11867) );
  NAND2_X1 U14253 ( .A1(n11870), .A2(n11869), .ZN(n11871) );
  NAND3_X1 U14254 ( .A1(n11989), .A2(n14522), .A3(n11871), .ZN(n11872) );
  AOI22_X1 U14255 ( .A1(n13673), .A2(n14003), .B1(n14353), .B2(n13674), .ZN(
        n14267) );
  NAND2_X1 U14256 ( .A1(n11872), .A2(n14267), .ZN(n14307) );
  NAND2_X1 U14257 ( .A1(n11873), .A2(n14305), .ZN(n14007) );
  OAI211_X1 U14258 ( .C1(n11873), .C2(n14305), .A(n14007), .B(n14448), .ZN(
        n14304) );
  INV_X1 U14259 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11874) );
  OAI22_X1 U14260 ( .A1(n14010), .A2(n11874), .B1(n14272), .B2(n14439), .ZN(
        n11875) );
  AOI21_X1 U14261 ( .B1(n12068), .B2(n14396), .A(n11875), .ZN(n11876) );
  OAI21_X1 U14262 ( .B1(n14304), .B2(n13917), .A(n11876), .ZN(n11877) );
  AOI21_X1 U14263 ( .B1(n14307), .B2(n14010), .A(n11877), .ZN(n11878) );
  OAI21_X1 U14264 ( .B1(n13998), .B2(n11879), .A(n11878), .ZN(P1_U3276) );
  INV_X1 U14265 ( .A(n11880), .ZN(n11986) );
  OAI222_X1 U14266 ( .A1(n13578), .A2(n11882), .B1(n13581), .B2(n11986), .C1(
        P2_U3088), .C2(n11881), .ZN(P2_U3302) );
  OAI211_X1 U14267 ( .C1(n11884), .C2(n12575), .A(n11883), .B(n15001), .ZN(
        n11886) );
  AOI22_X1 U14268 ( .A1(n12909), .A2(n14962), .B1(n14965), .B2(n12605), .ZN(
        n11885) );
  NAND2_X1 U14269 ( .A1(n11886), .A2(n11885), .ZN(n11913) );
  INV_X1 U14270 ( .A(n11913), .ZN(n11894) );
  OAI21_X1 U14271 ( .B1(n11888), .B2(n12460), .A(n11887), .ZN(n11914) );
  INV_X1 U14272 ( .A(n11889), .ZN(n11920) );
  AOI22_X1 U14273 ( .A1(n15012), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15007), 
        .B2(n11890), .ZN(n11891) );
  OAI21_X1 U14274 ( .B1(n11920), .B2(n12928), .A(n11891), .ZN(n11892) );
  AOI21_X1 U14275 ( .B1(n11914), .B2(n12930), .A(n11892), .ZN(n11893) );
  OAI21_X1 U14276 ( .B1(n11894), .B2(n15012), .A(n11893), .ZN(P3_U3218) );
  INV_X1 U14277 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11901) );
  AOI211_X1 U14278 ( .C1(n14549), .C2(n14256), .A(n14258), .B(n11895), .ZN(
        n11898) );
  NAND2_X1 U14279 ( .A1(n11896), .A2(n14522), .ZN(n11897) );
  OAI211_X1 U14280 ( .C1(n14517), .C2(n11899), .A(n11898), .B(n11897), .ZN(
        n11902) );
  NAND2_X1 U14281 ( .A1(n11902), .A2(n14578), .ZN(n11900) );
  OAI21_X1 U14282 ( .B1(n14578), .B2(n11901), .A(n11900), .ZN(P1_U3507) );
  NAND2_X1 U14283 ( .A1(n11902), .A2(n14594), .ZN(n11903) );
  OAI21_X1 U14284 ( .B1(n14594), .B2(n11904), .A(n11903), .ZN(P1_U3544) );
  INV_X1 U14285 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11907) );
  AOI21_X1 U14286 ( .B1(n15063), .B2(n11906), .A(n11905), .ZN(n11909) );
  MUX2_X1 U14287 ( .A(n11907), .B(n11909), .S(n15079), .Z(n11908) );
  OAI21_X1 U14288 ( .B1(n12996), .B2(n11912), .A(n11908), .ZN(P3_U3473) );
  INV_X1 U14289 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11910) );
  MUX2_X1 U14290 ( .A(n11910), .B(n11909), .S(n15066), .Z(n11911) );
  OAI21_X1 U14291 ( .B1(n13043), .B2(n11912), .A(n11911), .ZN(P3_U3432) );
  INV_X1 U14292 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11915) );
  AOI21_X1 U14293 ( .B1(n15063), .B2(n11914), .A(n11913), .ZN(n11917) );
  MUX2_X1 U14294 ( .A(n11915), .B(n11917), .S(n15066), .Z(n11916) );
  OAI21_X1 U14295 ( .B1(n11920), .B2(n13043), .A(n11916), .ZN(P3_U3435) );
  MUX2_X1 U14296 ( .A(n11918), .B(n11917), .S(n15079), .Z(n11919) );
  OAI21_X1 U14297 ( .B1(n11920), .B2(n12996), .A(n11919), .ZN(P3_U3474) );
  OAI222_X1 U14298 ( .A1(n12393), .A2(P3_U3151), .B1(n13058), .B2(n11922), 
        .C1(n13056), .C2(n11921), .ZN(P3_U3274) );
  INV_X1 U14299 ( .A(n11923), .ZN(n11926) );
  OAI222_X1 U14300 ( .A1(n13056), .A2(n11926), .B1(n11925), .B2(P3_U3151), 
        .C1(n11924), .C2(n13058), .ZN(P3_U3267) );
  INV_X1 U14301 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11929) );
  INV_X1 U14302 ( .A(n11927), .ZN(n13574) );
  OAI222_X1 U14303 ( .A1(n14125), .A2(n11929), .B1(n14128), .B2(n13574), .C1(
        P1_U3086), .C2(n11928), .ZN(P1_U3327) );
  INV_X1 U14304 ( .A(n13474), .ZN(n13150) );
  INV_X1 U14305 ( .A(n13182), .ZN(n13076) );
  INV_X1 U14306 ( .A(n13503), .ZN(n13384) );
  OAI21_X1 U14307 ( .B1(n13516), .B2(n11947), .A(n11930), .ZN(n13392) );
  NAND2_X1 U14308 ( .A1(n13391), .A2(n11931), .ZN(n13386) );
  INV_X1 U14309 ( .A(n13498), .ZN(n13371) );
  INV_X1 U14310 ( .A(n13181), .ZN(n13154) );
  NAND2_X1 U14311 ( .A1(n13371), .A2(n13154), .ZN(n11932) );
  OAI21_X1 U14312 ( .B1(n13180), .B2(n12181), .A(n11933), .ZN(n13339) );
  INV_X1 U14313 ( .A(n13179), .ZN(n11960) );
  INV_X1 U14314 ( .A(n13177), .ZN(n13121) );
  NOR2_X1 U14315 ( .A1(n13311), .A2(n13121), .ZN(n11935) );
  INV_X1 U14316 ( .A(n11935), .ZN(n11936) );
  INV_X1 U14317 ( .A(n13292), .ZN(n13296) );
  NAND2_X1 U14318 ( .A1(n13274), .A2(n13174), .ZN(n11939) );
  AOI21_X1 U14319 ( .B1(n13265), .B2(n11939), .A(n11938), .ZN(n13257) );
  INV_X1 U14320 ( .A(n11971), .ZN(n11941) );
  NAND2_X1 U14321 ( .A1(n13240), .A2(n13255), .ZN(n13238) );
  NOR2_X2 U14322 ( .A1(n13432), .A2(n13238), .ZN(n13231) );
  INV_X1 U14323 ( .A(n11942), .ZN(n11943) );
  AOI22_X1 U14324 ( .A1(n13402), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n11943), 
        .B2(n13381), .ZN(n11944) );
  OAI21_X1 U14325 ( .B1(n11945), .B2(n13417), .A(n11944), .ZN(n11946) );
  AOI21_X1 U14326 ( .B1(n13431), .B2(n13422), .A(n11946), .ZN(n11979) );
  OR2_X1 U14327 ( .A1(n12157), .A2(n11947), .ZN(n11948) );
  NAND2_X1 U14328 ( .A1(n13400), .A2(n13153), .ZN(n11951) );
  OR2_X1 U14329 ( .A1(n13400), .A2(n13153), .ZN(n11952) );
  NAND2_X1 U14330 ( .A1(n11953), .A2(n11952), .ZN(n13376) );
  NOR2_X1 U14331 ( .A1(n13503), .A2(n13076), .ZN(n11954) );
  NAND2_X1 U14332 ( .A1(n13503), .A2(n13076), .ZN(n11955) );
  NAND2_X1 U14333 ( .A1(n12181), .A2(n13077), .ZN(n11958) );
  AND2_X1 U14334 ( .A1(n13346), .A2(n11960), .ZN(n11962) );
  OR2_X1 U14335 ( .A1(n13346), .A2(n11960), .ZN(n11961) );
  INV_X1 U14336 ( .A(n13332), .ZN(n13321) );
  INV_X1 U14337 ( .A(n13176), .ZN(n13094) );
  INV_X1 U14338 ( .A(n13457), .ZN(n13289) );
  INV_X1 U14339 ( .A(n11967), .ZN(n11968) );
  XNOR2_X1 U14340 ( .A(n11972), .B(n11971), .ZN(n11976) );
  AOI21_X1 U14341 ( .B1(n11973), .B2(P2_B_REG_SCAN_IN), .A(n13161), .ZN(n13225) );
  AND2_X1 U14342 ( .A1(n13170), .A2(n13225), .ZN(n11974) );
  INV_X1 U14343 ( .A(n13433), .ZN(n11977) );
  NAND2_X1 U14344 ( .A1(n11977), .A2(n13406), .ZN(n11978) );
  OAI211_X1 U14345 ( .C1(n13434), .C2(n13411), .A(n11979), .B(n11978), .ZN(
        P2_U3236) );
  AOI22_X1 U14346 ( .A1(n12744), .A2(n15007), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15012), .ZN(n11981) );
  OAI21_X1 U14347 ( .B1(n11982), .B2(n12928), .A(n11981), .ZN(n11983) );
  AOI21_X1 U14348 ( .B1(n11984), .B2(n12930), .A(n11983), .ZN(n11985) );
  OAI21_X1 U14349 ( .B1(n11980), .B2(n15012), .A(n11985), .ZN(P3_U3204) );
  OAI222_X1 U14350 ( .A1(n14125), .A2(n11987), .B1(n14128), .B2(n11986), .C1(
        P1_U3086), .C2(n10256), .ZN(P1_U3330) );
  INV_X1 U14351 ( .A(n14002), .ZN(n11988) );
  NAND2_X1 U14352 ( .A1(n14001), .A2(n14000), .ZN(n11991) );
  OR2_X1 U14353 ( .A1(n14092), .A2(n13600), .ZN(n11990) );
  NAND2_X1 U14354 ( .A1(n11991), .A2(n11990), .ZN(n13993) );
  INV_X1 U14355 ( .A(n13982), .ZN(n13994) );
  NAND2_X1 U14356 ( .A1(n14085), .A2(n11992), .ZN(n11993) );
  INV_X1 U14357 ( .A(n13961), .ZN(n12013) );
  NAND2_X1 U14358 ( .A1(n13960), .A2(n12013), .ZN(n11997) );
  OR2_X1 U14359 ( .A1(n14071), .A2(n11995), .ZN(n11996) );
  INV_X1 U14360 ( .A(n13670), .ZN(n13613) );
  NAND2_X1 U14361 ( .A1(n13947), .A2(n13613), .ZN(n11998) );
  INV_X1 U14362 ( .A(n13926), .ZN(n13928) );
  NAND2_X1 U14363 ( .A1(n14058), .A2(n11999), .ZN(n12000) );
  NAND2_X1 U14364 ( .A1(n13927), .A2(n12000), .ZN(n13906) );
  INV_X1 U14365 ( .A(n13920), .ZN(n14053) );
  INV_X1 U14366 ( .A(n13888), .ZN(n13893) );
  INV_X1 U14367 ( .A(n12002), .ZN(n12003) );
  AOI21_X1 U14368 ( .B1(n12004), .B2(n12006), .A(n13836), .ZN(n12005) );
  NOR2_X1 U14369 ( .A1(n12005), .A2(n14566), .ZN(n12025) );
  INV_X1 U14370 ( .A(n12006), .ZN(n12021) );
  OR2_X1 U14371 ( .A1(n14092), .A2(n13673), .ZN(n12009) );
  NOR2_X1 U14372 ( .A1(n14085), .A2(n14004), .ZN(n12011) );
  OR2_X1 U14373 ( .A1(n14077), .A2(n13614), .ZN(n12012) );
  OR2_X1 U14374 ( .A1(n14071), .A2(n13671), .ZN(n12014) );
  OR2_X1 U14375 ( .A1(n13947), .A2(n13670), .ZN(n12015) );
  NAND2_X1 U14376 ( .A1(n14058), .A2(n13669), .ZN(n12016) );
  INV_X1 U14377 ( .A(n13878), .ZN(n13873) );
  INV_X1 U14378 ( .A(n14039), .ZN(n12019) );
  NAND2_X1 U14379 ( .A1(n13666), .A2(n14353), .ZN(n12023) );
  NAND2_X1 U14380 ( .A1(n13846), .A2(n14003), .ZN(n12022) );
  NAND2_X1 U14381 ( .A1(n12023), .A2(n12022), .ZN(n13586) );
  INV_X1 U14382 ( .A(n14058), .ZN(n13938) );
  INV_X1 U14383 ( .A(n13866), .ZN(n12026) );
  AOI211_X1 U14384 ( .C1(n14033), .C2(n13882), .A(n14492), .B(n12026), .ZN(
        n14032) );
  INV_X1 U14385 ( .A(n14033), .ZN(n13835) );
  INV_X1 U14386 ( .A(n13588), .ZN(n12027) );
  AOI22_X1 U14387 ( .A1(n14395), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n12027), 
        .B2(n14394), .ZN(n12028) );
  OAI21_X1 U14388 ( .B1(n13835), .B2(n14444), .A(n12028), .ZN(n12030) );
  NOR2_X1 U14389 ( .A1(n14036), .A2(n13923), .ZN(n12029) );
  AOI211_X1 U14390 ( .C1(n14032), .C2(n14452), .A(n12030), .B(n12029), .ZN(
        n12031) );
  OAI21_X1 U14391 ( .B1(n14035), .B2(n13987), .A(n12031), .ZN(P1_U3266) );
  INV_X1 U14392 ( .A(n12032), .ZN(n12034) );
  NAND2_X1 U14393 ( .A1(n14247), .A2(n12130), .ZN(n12038) );
  NAND2_X1 U14394 ( .A1(n12131), .A2(n13676), .ZN(n12037) );
  NAND2_X1 U14395 ( .A1(n12038), .A2(n12037), .ZN(n12040) );
  XNOR2_X1 U14396 ( .A(n12040), .B(n12039), .ZN(n12044) );
  INV_X1 U14397 ( .A(n12044), .ZN(n12046) );
  NOR2_X1 U14398 ( .A1(n10373), .A2(n12041), .ZN(n12042) );
  AOI21_X1 U14399 ( .B1(n14247), .B2(n12131), .A(n12042), .ZN(n12043) );
  INV_X1 U14400 ( .A(n12043), .ZN(n12045) );
  AND2_X1 U14401 ( .A1(n12044), .A2(n12043), .ZN(n12047) );
  AOI21_X1 U14402 ( .B1(n12046), .B2(n12045), .A(n12047), .ZN(n14246) );
  INV_X1 U14403 ( .A(n12047), .ZN(n12048) );
  NAND2_X1 U14404 ( .A1(n14244), .A2(n12048), .ZN(n12053) );
  INV_X1 U14405 ( .A(n12053), .ZN(n12051) );
  OAI22_X1 U14406 ( .A1(n6817), .A2(n10731), .B1(n12055), .B2(n12139), .ZN(
        n12049) );
  XOR2_X1 U14407 ( .A(n12140), .B(n12049), .Z(n12052) );
  INV_X1 U14408 ( .A(n12052), .ZN(n12050) );
  OAI22_X1 U14409 ( .A1(n6817), .A2(n12139), .B1(n12055), .B2(n10373), .ZN(
        n14294) );
  INV_X1 U14410 ( .A(n14294), .ZN(n12056) );
  NAND2_X1 U14411 ( .A1(n14256), .A2(n12130), .ZN(n12059) );
  NAND2_X1 U14412 ( .A1(n13674), .A2(n12131), .ZN(n12058) );
  NAND2_X1 U14413 ( .A1(n12059), .A2(n12058), .ZN(n12060) );
  XNOR2_X1 U14414 ( .A(n12060), .B(n12140), .ZN(n12063) );
  AOI22_X1 U14415 ( .A1(n14256), .A2(n12131), .B1(n12135), .B2(n13674), .ZN(
        n12061) );
  XNOR2_X1 U14416 ( .A(n12063), .B(n12061), .ZN(n14255) );
  INV_X1 U14417 ( .A(n12061), .ZN(n12062) );
  NAND2_X1 U14418 ( .A1(n12068), .A2(n12130), .ZN(n12066) );
  NAND2_X1 U14419 ( .A1(n14002), .A2(n12131), .ZN(n12065) );
  NAND2_X1 U14420 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  XNOR2_X1 U14421 ( .A(n12067), .B(n12140), .ZN(n12072) );
  NAND2_X1 U14422 ( .A1(n12068), .A2(n12131), .ZN(n12070) );
  NAND2_X1 U14423 ( .A1(n14002), .A2(n12135), .ZN(n12069) );
  NAND2_X1 U14424 ( .A1(n12070), .A2(n12069), .ZN(n12071) );
  NAND2_X1 U14425 ( .A1(n12072), .A2(n12071), .ZN(n14262) );
  NOR2_X1 U14426 ( .A1(n12072), .A2(n12071), .ZN(n14264) );
  AOI22_X1 U14427 ( .A1(n14092), .A2(n12131), .B1(n12135), .B2(n13673), .ZN(
        n12076) );
  NAND2_X1 U14428 ( .A1(n14092), .A2(n12130), .ZN(n12074) );
  NAND2_X1 U14429 ( .A1(n13673), .A2(n12131), .ZN(n12073) );
  NAND2_X1 U14430 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  XNOR2_X1 U14431 ( .A(n12075), .B(n12140), .ZN(n12078) );
  XOR2_X1 U14432 ( .A(n12076), .B(n12078), .Z(n14282) );
  INV_X1 U14433 ( .A(n12076), .ZN(n12077) );
  AND2_X1 U14434 ( .A1(n14004), .A2(n12135), .ZN(n12079) );
  AOI21_X1 U14435 ( .B1(n14085), .B2(n12131), .A(n12079), .ZN(n12085) );
  NAND2_X1 U14436 ( .A1(n14085), .A2(n12130), .ZN(n12081) );
  NAND2_X1 U14437 ( .A1(n14004), .A2(n12131), .ZN(n12080) );
  NAND2_X1 U14438 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  XNOR2_X1 U14439 ( .A(n12082), .B(n12140), .ZN(n12084) );
  XOR2_X1 U14440 ( .A(n12085), .B(n12084), .Z(n13605) );
  INV_X1 U14441 ( .A(n12085), .ZN(n12086) );
  OR2_X1 U14442 ( .A1(n14077), .A2(n12139), .ZN(n12089) );
  NAND2_X1 U14443 ( .A1(n13672), .A2(n12135), .ZN(n12088) );
  NAND2_X1 U14444 ( .A1(n12089), .A2(n12088), .ZN(n12091) );
  OAI22_X1 U14445 ( .A1(n14077), .A2(n10731), .B1(n13614), .B2(n12139), .ZN(
        n12090) );
  XNOR2_X1 U14446 ( .A(n12090), .B(n12140), .ZN(n12092) );
  XOR2_X1 U14447 ( .A(n12091), .B(n12092), .Z(n13636) );
  NAND2_X1 U14448 ( .A1(n12092), .A2(n12091), .ZN(n12093) );
  AOI22_X1 U14449 ( .A1(n14071), .A2(n12130), .B1(n12131), .B2(n13671), .ZN(
        n12094) );
  XNOR2_X1 U14450 ( .A(n12094), .B(n12140), .ZN(n12096) );
  AOI22_X1 U14451 ( .A1(n14071), .A2(n12131), .B1(n12135), .B2(n13671), .ZN(
        n12095) );
  XNOR2_X1 U14452 ( .A(n12096), .B(n12095), .ZN(n13612) );
  NAND2_X1 U14453 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  NOR2_X1 U14454 ( .A1(n10373), .A2(n13613), .ZN(n12098) );
  AOI21_X1 U14455 ( .B1(n13947), .B2(n12131), .A(n12098), .ZN(n12100) );
  AOI22_X1 U14456 ( .A1(n13947), .A2(n12130), .B1(n12131), .B2(n13670), .ZN(
        n12099) );
  XNOR2_X1 U14457 ( .A(n12099), .B(n12140), .ZN(n12101) );
  XOR2_X1 U14458 ( .A(n12100), .B(n12101), .Z(n13646) );
  NAND2_X1 U14459 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  NAND2_X1 U14460 ( .A1(n14058), .A2(n12130), .ZN(n12104) );
  NAND2_X1 U14461 ( .A1(n12131), .A2(n13669), .ZN(n12103) );
  NAND2_X1 U14462 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  XNOR2_X1 U14463 ( .A(n12105), .B(n12140), .ZN(n12106) );
  AOI22_X1 U14464 ( .A1(n14058), .A2(n12131), .B1(n12135), .B2(n13669), .ZN(
        n12107) );
  XNOR2_X1 U14465 ( .A(n12106), .B(n12107), .ZN(n13593) );
  INV_X1 U14466 ( .A(n12106), .ZN(n12108) );
  NAND2_X1 U14467 ( .A1(n13920), .A2(n12130), .ZN(n12110) );
  NAND2_X1 U14468 ( .A1(n12131), .A2(n13668), .ZN(n12109) );
  NAND2_X1 U14469 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  XNOR2_X1 U14470 ( .A(n12111), .B(n12140), .ZN(n12112) );
  AOI22_X1 U14471 ( .A1(n13920), .A2(n12131), .B1(n12135), .B2(n13668), .ZN(
        n12113) );
  XNOR2_X1 U14472 ( .A(n12112), .B(n12113), .ZN(n13628) );
  NAND2_X1 U14473 ( .A1(n13627), .A2(n13628), .ZN(n12116) );
  INV_X1 U14474 ( .A(n12112), .ZN(n12114) );
  NAND2_X1 U14475 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U14476 ( .A1(n14045), .A2(n12130), .ZN(n12118) );
  NAND2_X1 U14477 ( .A1(n12131), .A2(n13667), .ZN(n12117) );
  NAND2_X1 U14478 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  XNOR2_X1 U14479 ( .A(n12119), .B(n12140), .ZN(n12120) );
  AOI22_X1 U14480 ( .A1(n14045), .A2(n12131), .B1(n12135), .B2(n13667), .ZN(
        n12121) );
  XNOR2_X1 U14481 ( .A(n12120), .B(n12121), .ZN(n13620) );
  INV_X1 U14482 ( .A(n12120), .ZN(n12122) );
  NAND2_X1 U14483 ( .A1(n12122), .A2(n12121), .ZN(n12123) );
  NAND2_X1 U14484 ( .A1(n14039), .A2(n12130), .ZN(n12125) );
  NAND2_X1 U14485 ( .A1(n12131), .A2(n13666), .ZN(n12124) );
  NAND2_X1 U14486 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  XNOR2_X1 U14487 ( .A(n12126), .B(n12140), .ZN(n12127) );
  AOI22_X1 U14488 ( .A1(n14039), .A2(n12131), .B1(n12135), .B2(n13666), .ZN(
        n12128) );
  XNOR2_X1 U14489 ( .A(n12127), .B(n12128), .ZN(n13657) );
  INV_X1 U14490 ( .A(n12127), .ZN(n12129) );
  NAND2_X1 U14491 ( .A1(n14033), .A2(n12130), .ZN(n12133) );
  NAND2_X1 U14492 ( .A1(n12131), .A2(n13834), .ZN(n12132) );
  NAND2_X1 U14493 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  XNOR2_X1 U14494 ( .A(n12134), .B(n12140), .ZN(n12136) );
  AOI22_X1 U14495 ( .A1(n14033), .A2(n12131), .B1(n12135), .B2(n13834), .ZN(
        n12137) );
  XNOR2_X1 U14496 ( .A(n12136), .B(n12137), .ZN(n13585) );
  INV_X1 U14497 ( .A(n12136), .ZN(n12138) );
  OAI22_X1 U14498 ( .A1(n13832), .A2(n10731), .B1(n13831), .B2(n12139), .ZN(
        n12143) );
  OAI22_X1 U14499 ( .A1(n13832), .A2(n12139), .B1(n13831), .B2(n10373), .ZN(
        n12141) );
  XNOR2_X1 U14500 ( .A(n12141), .B(n12140), .ZN(n12142) );
  XOR2_X1 U14501 ( .A(n12143), .B(n12142), .Z(n12144) );
  XNOR2_X1 U14502 ( .A(n12145), .B(n12144), .ZN(n12150) );
  NOR2_X1 U14503 ( .A1(n14367), .A2(n13864), .ZN(n12148) );
  AOI22_X1 U14504 ( .A1(n13665), .A2(n14003), .B1(n14353), .B2(n13834), .ZN(
        n13858) );
  OAI22_X1 U14505 ( .A1(n14284), .A2(n13858), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12146), .ZN(n12147) );
  AOI211_X1 U14506 ( .C1(n14028), .C2(n14297), .A(n12148), .B(n12147), .ZN(
        n12149) );
  OAI21_X1 U14507 ( .B1(n12150), .B2(n13663), .A(n12149), .ZN(P1_U3220) );
  INV_X1 U14508 ( .A(n12151), .ZN(n12152) );
  NOR2_X1 U14509 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  AOI21_X2 U14510 ( .B1(n12156), .B2(n12155), .A(n12154), .ZN(n13100) );
  XNOR2_X1 U14511 ( .A(n12157), .B(n12205), .ZN(n12158) );
  NAND2_X1 U14512 ( .A1(n13184), .A2(n10230), .ZN(n12159) );
  NAND2_X1 U14513 ( .A1(n12158), .A2(n12159), .ZN(n12163) );
  INV_X1 U14514 ( .A(n12158), .ZN(n12161) );
  INV_X1 U14515 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U14516 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  AND2_X1 U14517 ( .A1(n12163), .A2(n12162), .ZN(n13101) );
  XNOR2_X1 U14518 ( .A(n13400), .B(n12205), .ZN(n12164) );
  NAND2_X1 U14519 ( .A1(n13183), .A2(n10230), .ZN(n12165) );
  NAND2_X1 U14520 ( .A1(n12164), .A2(n12165), .ZN(n12169) );
  INV_X1 U14521 ( .A(n12164), .ZN(n12167) );
  INV_X1 U14522 ( .A(n12165), .ZN(n12166) );
  NAND2_X1 U14523 ( .A1(n12167), .A2(n12166), .ZN(n12168) );
  AND2_X1 U14524 ( .A1(n12169), .A2(n12168), .ZN(n13111) );
  XNOR2_X1 U14525 ( .A(n13503), .B(n12205), .ZN(n12170) );
  NAND2_X1 U14526 ( .A1(n13182), .A2(n10230), .ZN(n12171) );
  XNOR2_X1 U14527 ( .A(n12170), .B(n12171), .ZN(n13151) );
  INV_X1 U14528 ( .A(n12170), .ZN(n12173) );
  INV_X1 U14529 ( .A(n12171), .ZN(n12172) );
  NAND2_X1 U14530 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  XNOR2_X1 U14531 ( .A(n13498), .B(n12205), .ZN(n12175) );
  NAND2_X1 U14532 ( .A1(n13181), .A2(n10230), .ZN(n12176) );
  NAND2_X1 U14533 ( .A1(n12175), .A2(n12176), .ZN(n12180) );
  INV_X1 U14534 ( .A(n12175), .ZN(n12178) );
  INV_X1 U14535 ( .A(n12176), .ZN(n12177) );
  NAND2_X1 U14536 ( .A1(n12178), .A2(n12177), .ZN(n12179) );
  NAND2_X1 U14537 ( .A1(n12180), .A2(n12179), .ZN(n13074) );
  XNOR2_X1 U14538 ( .A(n12181), .B(n12205), .ZN(n12182) );
  NAND2_X1 U14539 ( .A1(n13180), .A2(n10230), .ZN(n12183) );
  NAND2_X1 U14540 ( .A1(n12182), .A2(n12183), .ZN(n12187) );
  INV_X1 U14541 ( .A(n12182), .ZN(n12185) );
  INV_X1 U14542 ( .A(n12183), .ZN(n12184) );
  NAND2_X1 U14543 ( .A1(n12185), .A2(n12184), .ZN(n12186) );
  AND2_X1 U14544 ( .A1(n12187), .A2(n12186), .ZN(n13128) );
  XNOR2_X1 U14545 ( .A(n13346), .B(n12205), .ZN(n12188) );
  NAND2_X1 U14546 ( .A1(n13179), .A2(n10230), .ZN(n12189) );
  XNOR2_X1 U14547 ( .A(n12188), .B(n12189), .ZN(n13083) );
  INV_X1 U14548 ( .A(n12188), .ZN(n12191) );
  INV_X1 U14549 ( .A(n12189), .ZN(n12190) );
  NAND2_X1 U14550 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  XOR2_X1 U14551 ( .A(n12213), .B(n13474), .Z(n12193) );
  XNOR2_X1 U14552 ( .A(n12194), .B(n12193), .ZN(n13137) );
  NAND2_X1 U14553 ( .A1(n13178), .A2(n10230), .ZN(n13136) );
  NAND2_X1 U14554 ( .A1(n13137), .A2(n13136), .ZN(n13135) );
  INV_X1 U14555 ( .A(n12193), .ZN(n12195) );
  OR2_X1 U14556 ( .A1(n12195), .A2(n12194), .ZN(n12196) );
  NAND2_X1 U14557 ( .A1(n13135), .A2(n12196), .ZN(n12197) );
  NAND2_X1 U14558 ( .A1(n13177), .A2(n10230), .ZN(n13067) );
  OAI22_X1 U14559 ( .A1(n13066), .A2(n13067), .B1(n6588), .B2(n12197), .ZN(
        n13119) );
  XNOR2_X1 U14560 ( .A(n13462), .B(n12213), .ZN(n12200) );
  NAND2_X1 U14561 ( .A1(n13176), .A2(n10230), .ZN(n12198) );
  XNOR2_X1 U14562 ( .A(n12200), .B(n12198), .ZN(n13120) );
  INV_X1 U14563 ( .A(n12198), .ZN(n12199) );
  AOI21_X2 U14564 ( .B1(n13119), .B2(n13120), .A(n12201), .ZN(n13092) );
  NAND2_X1 U14565 ( .A1(n13175), .A2(n10230), .ZN(n12203) );
  XNOR2_X1 U14566 ( .A(n13457), .B(n12213), .ZN(n12202) );
  XOR2_X1 U14567 ( .A(n12203), .B(n12202), .Z(n13091) );
  INV_X1 U14568 ( .A(n12202), .ZN(n12204) );
  XNOR2_X1 U14569 ( .A(n13274), .B(n12205), .ZN(n12207) );
  NAND2_X1 U14570 ( .A1(n13174), .A2(n10230), .ZN(n12206) );
  NAND2_X1 U14571 ( .A1(n12207), .A2(n12206), .ZN(n12208) );
  OAI21_X1 U14572 ( .B1(n12207), .B2(n12206), .A(n12208), .ZN(n13159) );
  XNOR2_X1 U14573 ( .A(n13442), .B(n12213), .ZN(n12211) );
  NAND2_X1 U14574 ( .A1(n13173), .A2(n10230), .ZN(n12209) );
  XNOR2_X1 U14575 ( .A(n12211), .B(n12209), .ZN(n13059) );
  INV_X1 U14576 ( .A(n12209), .ZN(n12210) );
  AOI21_X2 U14577 ( .B1(n13060), .B2(n13059), .A(n12212), .ZN(n12217) );
  NAND2_X1 U14578 ( .A1(n13172), .A2(n10230), .ZN(n12214) );
  XNOR2_X1 U14579 ( .A(n12214), .B(n12213), .ZN(n12215) );
  XNOR2_X1 U14580 ( .A(n13240), .B(n12215), .ZN(n12216) );
  XNOR2_X1 U14581 ( .A(n12217), .B(n12216), .ZN(n12222) );
  OAI22_X1 U14582 ( .A1(n13162), .A2(n13163), .B1(n12218), .B2(n13161), .ZN(
        n13245) );
  AOI22_X1 U14583 ( .A1(n14237), .A2(n13245), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12219) );
  OAI21_X1 U14584 ( .B1(n13247), .B2(n14243), .A(n12219), .ZN(n12220) );
  AOI21_X1 U14585 ( .B1(n13436), .B2(n14240), .A(n12220), .ZN(n12221) );
  OAI21_X1 U14586 ( .B1(n12222), .B2(n13168), .A(n12221), .ZN(P2_U3192) );
  INV_X1 U14587 ( .A(n12223), .ZN(n12224) );
  XNOR2_X1 U14588 ( .A(n12533), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12226) );
  XNOR2_X1 U14589 ( .A(n12534), .B(n12226), .ZN(n12527) );
  INV_X1 U14590 ( .A(n12527), .ZN(n12227) );
  INV_X1 U14591 ( .A(n12230), .ZN(n12231) );
  OAI22_X2 U14592 ( .A1(n12233), .A2(n12232), .B1(n12231), .B2(n12909), .ZN(
        n12328) );
  XNOR2_X1 U14593 ( .A(n12988), .B(n10097), .ZN(n12234) );
  XNOR2_X1 U14594 ( .A(n12234), .B(n12922), .ZN(n12329) );
  INV_X1 U14595 ( .A(n12234), .ZN(n12235) );
  XNOR2_X1 U14596 ( .A(n12367), .B(n10097), .ZN(n12362) );
  XNOR2_X1 U14597 ( .A(n12561), .B(n10097), .ZN(n12236) );
  XNOR2_X1 U14598 ( .A(n12236), .B(n12899), .ZN(n12289) );
  XNOR2_X1 U14599 ( .A(n12976), .B(n10097), .ZN(n12237) );
  XNOR2_X1 U14600 ( .A(n12237), .B(n12601), .ZN(n12347) );
  NAND2_X1 U14601 ( .A1(n12239), .A2(n12238), .ZN(n12306) );
  XNOR2_X1 U14602 ( .A(n12860), .B(n10097), .ZN(n12240) );
  NAND2_X1 U14603 ( .A1(n12240), .A2(n12846), .ZN(n12241) );
  OAI21_X1 U14604 ( .B1(n12240), .B2(n12846), .A(n12241), .ZN(n12309) );
  NAND2_X1 U14605 ( .A1(n12307), .A2(n12241), .ZN(n12243) );
  XNOR2_X1 U14606 ( .A(n12849), .B(n10097), .ZN(n12242) );
  XNOR2_X1 U14607 ( .A(n12963), .B(n10097), .ZN(n12247) );
  INV_X1 U14608 ( .A(n12247), .ZN(n12245) );
  NAND2_X1 U14609 ( .A1(n12246), .A2(n12245), .ZN(n12249) );
  XNOR2_X1 U14610 ( .A(n12346), .B(n12262), .ZN(n12250) );
  NAND2_X1 U14611 ( .A1(n12250), .A2(n7179), .ZN(n12317) );
  INV_X1 U14612 ( .A(n12250), .ZN(n12251) );
  NAND2_X1 U14613 ( .A1(n12251), .A2(n12832), .ZN(n12252) );
  NAND2_X1 U14614 ( .A1(n12253), .A2(n12336), .ZN(n12316) );
  NAND2_X1 U14615 ( .A1(n12316), .A2(n12317), .ZN(n12257) );
  XNOR2_X1 U14616 ( .A(n12315), .B(n10097), .ZN(n12254) );
  NAND2_X1 U14617 ( .A1(n12254), .A2(n12821), .ZN(n12258) );
  INV_X1 U14618 ( .A(n12254), .ZN(n12255) );
  NAND2_X1 U14619 ( .A1(n12255), .A2(n12600), .ZN(n12256) );
  NAND2_X1 U14620 ( .A1(n12257), .A2(n12318), .ZN(n12320) );
  NAND2_X1 U14621 ( .A1(n12320), .A2(n12258), .ZN(n12373) );
  XNOR2_X1 U14622 ( .A(n12791), .B(n12262), .ZN(n12259) );
  NOR2_X1 U14623 ( .A1(n12259), .A2(n12802), .ZN(n12260) );
  AOI21_X1 U14624 ( .B1(n12259), .B2(n12802), .A(n12260), .ZN(n12375) );
  NAND2_X1 U14625 ( .A1(n12373), .A2(n12375), .ZN(n12374) );
  INV_X1 U14626 ( .A(n12260), .ZN(n12261) );
  XNOR2_X1 U14627 ( .A(n12778), .B(n12262), .ZN(n12263) );
  NOR2_X1 U14628 ( .A1(n12263), .A2(n12758), .ZN(n12264) );
  AOI21_X1 U14629 ( .B1(n12263), .B2(n12758), .A(n12264), .ZN(n12276) );
  XNOR2_X1 U14630 ( .A(n9586), .B(n10097), .ZN(n12265) );
  AOI22_X1 U14631 ( .A1(n12761), .A2(n12383), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12266) );
  OAI21_X1 U14632 ( .B1(n12267), .B2(n12380), .A(n12266), .ZN(n12270) );
  NOR2_X1 U14633 ( .A1(n13007), .A2(n12386), .ZN(n12269) );
  AOI211_X1 U14634 ( .C1(n12355), .C2(n12758), .A(n12270), .B(n12269), .ZN(
        n12271) );
  OAI21_X1 U14635 ( .B1(n12272), .B2(n12371), .A(n12271), .ZN(P3_U3160) );
  INV_X1 U14636 ( .A(n12273), .ZN(n14118) );
  OAI222_X1 U14637 ( .A1(n13581), .A2(n14118), .B1(P2_U3088), .B2(n8453), .C1(
        n12533), .C2(n13578), .ZN(P2_U3297) );
  OAI21_X1 U14638 ( .B1(n12276), .B2(n12275), .A(n12274), .ZN(n12277) );
  NAND2_X1 U14639 ( .A1(n12277), .A2(n12376), .ZN(n12281) );
  AOI22_X1 U14640 ( .A1(n12777), .A2(n12383), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12278) );
  OAI21_X1 U14641 ( .B1(n12773), .B2(n12380), .A(n12278), .ZN(n12279) );
  AOI21_X1 U14642 ( .B1(n12355), .B2(n12802), .A(n12279), .ZN(n12280) );
  OAI211_X1 U14643 ( .C1(n13011), .C2(n12386), .A(n12281), .B(n12280), .ZN(
        P3_U3154) );
  AOI21_X1 U14644 ( .B1(n12818), .B2(n12282), .A(n12338), .ZN(n12288) );
  AOI22_X1 U14645 ( .A1(n12831), .A2(n12355), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12285) );
  NAND2_X1 U14646 ( .A1(n12835), .A2(n12383), .ZN(n12284) );
  OAI211_X1 U14647 ( .C1(n7179), .C2(n12380), .A(n12285), .B(n12284), .ZN(
        n12286) );
  AOI21_X1 U14648 ( .B1(n12963), .B2(n12359), .A(n12286), .ZN(n12287) );
  OAI21_X1 U14649 ( .B1(n12288), .B2(n12371), .A(n12287), .ZN(P3_U3156) );
  XNOR2_X1 U14650 ( .A(n12290), .B(n12289), .ZN(n12295) );
  NAND2_X1 U14651 ( .A1(n12910), .A2(n12355), .ZN(n12291) );
  NAND2_X1 U14652 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12739)
         );
  OAI211_X1 U14653 ( .C1(n12885), .C2(n12380), .A(n12291), .B(n12739), .ZN(
        n12293) );
  INV_X1 U14654 ( .A(n12561), .ZN(n13034) );
  NOR2_X1 U14655 ( .A1(n13034), .A2(n12386), .ZN(n12292) );
  AOI211_X1 U14656 ( .C1(n12889), .C2(n12383), .A(n12293), .B(n12292), .ZN(
        n12294) );
  OAI21_X1 U14657 ( .B1(n12295), .B2(n12371), .A(n12294), .ZN(P3_U3159) );
  XOR2_X1 U14658 ( .A(n12297), .B(n12296), .Z(n12298) );
  NAND2_X1 U14659 ( .A1(n12298), .A2(n12376), .ZN(n12305) );
  NOR2_X1 U14660 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12299), .ZN(n14878) );
  AOI21_X1 U14661 ( .B1(n12359), .B2(n12300), .A(n14878), .ZN(n12304) );
  AOI22_X1 U14662 ( .A1(n12365), .A2(n14935), .B1(n12355), .B2(n12609), .ZN(
        n12303) );
  NAND2_X1 U14663 ( .A1(n12383), .A2(n12301), .ZN(n12302) );
  NAND4_X1 U14664 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        P3_U3161) );
  INV_X1 U14665 ( .A(n12307), .ZN(n12308) );
  AOI21_X1 U14666 ( .B1(n12309), .B2(n12306), .A(n12308), .ZN(n12314) );
  AOI22_X1 U14667 ( .A1(n12601), .A2(n12355), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12311) );
  NAND2_X1 U14668 ( .A1(n12861), .A2(n12383), .ZN(n12310) );
  OAI211_X1 U14669 ( .C1(n12857), .C2(n12380), .A(n12311), .B(n12310), .ZN(
        n12312) );
  AOI21_X1 U14670 ( .B1(n12860), .B2(n12359), .A(n12312), .ZN(n12313) );
  OAI21_X1 U14671 ( .B1(n12314), .B2(n12371), .A(n12313), .ZN(P3_U3163) );
  INV_X1 U14672 ( .A(n12316), .ZN(n12339) );
  INV_X1 U14673 ( .A(n12317), .ZN(n12319) );
  NOR3_X1 U14674 ( .A1(n12339), .A2(n12319), .A3(n12318), .ZN(n12322) );
  INV_X1 U14675 ( .A(n12320), .ZN(n12321) );
  OAI21_X1 U14676 ( .B1(n12322), .B2(n12321), .A(n12376), .ZN(n12326) );
  AOI22_X1 U14677 ( .A1(n12805), .A2(n12383), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12323) );
  OAI21_X1 U14678 ( .B1(n7179), .B2(n12379), .A(n12323), .ZN(n12324) );
  AOI21_X1 U14679 ( .B1(n12365), .B2(n12802), .A(n12324), .ZN(n12325) );
  OAI211_X1 U14680 ( .C1(n13019), .C2(n12386), .A(n12326), .B(n12325), .ZN(
        P3_U3165) );
  INV_X1 U14681 ( .A(n12988), .ZN(n12916) );
  AOI211_X1 U14682 ( .C1(n12329), .C2(n12328), .A(n12371), .B(n12327), .ZN(
        n12330) );
  INV_X1 U14683 ( .A(n12330), .ZN(n12334) );
  NAND2_X1 U14684 ( .A1(n12355), .A2(n12909), .ZN(n12331) );
  NAND2_X1 U14685 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14174)
         );
  OAI211_X1 U14686 ( .C1(n12886), .C2(n12380), .A(n12331), .B(n14174), .ZN(
        n12332) );
  AOI21_X1 U14687 ( .B1(n12914), .B2(n12383), .A(n12332), .ZN(n12333) );
  OAI211_X1 U14688 ( .C1(n12916), .C2(n12386), .A(n12334), .B(n12333), .ZN(
        P3_U3168) );
  INV_X1 U14689 ( .A(n12335), .ZN(n12337) );
  NOR3_X1 U14690 ( .A1(n12338), .A2(n12337), .A3(n12336), .ZN(n12340) );
  OAI21_X1 U14691 ( .B1(n12340), .B2(n12339), .A(n12376), .ZN(n12345) );
  OAI22_X1 U14692 ( .A1(n12845), .A2(n12379), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12341), .ZN(n12343) );
  NOR2_X1 U14693 ( .A1(n12821), .A2(n12380), .ZN(n12342) );
  AOI211_X1 U14694 ( .C1(n12822), .C2(n12383), .A(n12343), .B(n12342), .ZN(
        n12344) );
  OAI211_X1 U14695 ( .C1(n12386), .C2(n12346), .A(n12345), .B(n12344), .ZN(
        P3_U3169) );
  XNOR2_X1 U14696 ( .A(n12348), .B(n12347), .ZN(n12353) );
  AOI22_X1 U14697 ( .A1(n12872), .A2(n12365), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12350) );
  NAND2_X1 U14698 ( .A1(n12877), .A2(n12383), .ZN(n12349) );
  OAI211_X1 U14699 ( .C1(n12899), .C2(n12379), .A(n12350), .B(n12349), .ZN(
        n12351) );
  AOI21_X1 U14700 ( .B1(n12976), .B2(n12359), .A(n12351), .ZN(n12352) );
  OAI21_X1 U14701 ( .B1(n12353), .B2(n12371), .A(n12352), .ZN(P3_U3173) );
  AOI21_X1 U14702 ( .B1(n12831), .B2(n12354), .A(n6528), .ZN(n12361) );
  AOI22_X1 U14703 ( .A1(n12872), .A2(n12355), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12357) );
  NAND2_X1 U14704 ( .A1(n12850), .A2(n12383), .ZN(n12356) );
  OAI211_X1 U14705 ( .C1(n12845), .C2(n12380), .A(n12357), .B(n12356), .ZN(
        n12358) );
  AOI21_X1 U14706 ( .B1(n12849), .B2(n12359), .A(n12358), .ZN(n12360) );
  OAI21_X1 U14707 ( .B1(n12361), .B2(n12371), .A(n12360), .ZN(P3_U3175) );
  XNOR2_X1 U14708 ( .A(n12362), .B(n12886), .ZN(n12363) );
  XNOR2_X1 U14709 ( .A(n12364), .B(n12363), .ZN(n12372) );
  NAND2_X1 U14710 ( .A1(n12866), .A2(n12365), .ZN(n12366) );
  NAND2_X1 U14711 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12704)
         );
  OAI211_X1 U14712 ( .C1(n12922), .C2(n12379), .A(n12366), .B(n12704), .ZN(
        n12369) );
  INV_X1 U14713 ( .A(n12367), .ZN(n13038) );
  NOR2_X1 U14714 ( .A1(n13038), .A2(n12386), .ZN(n12368) );
  AOI211_X1 U14715 ( .C1(n12903), .C2(n12383), .A(n12369), .B(n12368), .ZN(
        n12370) );
  OAI21_X1 U14716 ( .B1(n12372), .B2(n12371), .A(n12370), .ZN(P3_U3178) );
  OAI21_X1 U14717 ( .B1(n12375), .B2(n12373), .A(n12374), .ZN(n12377) );
  NAND2_X1 U14718 ( .A1(n12377), .A2(n12376), .ZN(n12385) );
  OAI22_X1 U14719 ( .A1(n12821), .A2(n12379), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12378), .ZN(n12382) );
  NOR2_X1 U14720 ( .A1(n12786), .A2(n12380), .ZN(n12381) );
  AOI211_X1 U14721 ( .C1(n12790), .C2(n12383), .A(n12382), .B(n12381), .ZN(
        n12384) );
  OAI211_X1 U14722 ( .C1(n13015), .C2(n12386), .A(n12385), .B(n12384), .ZN(
        P3_U3180) );
  INV_X1 U14723 ( .A(n12387), .ZN(n12519) );
  NAND2_X1 U14724 ( .A1(n12515), .A2(n12516), .ZN(n12785) );
  INV_X1 U14725 ( .A(n12785), .ZN(n12513) );
  XNOR2_X1 U14726 ( .A(n12388), .B(n12525), .ZN(n12507) );
  NAND2_X1 U14727 ( .A1(n12500), .A2(n12498), .ZN(n12847) );
  INV_X1 U14728 ( .A(n12847), .ZN(n12497) );
  NAND2_X1 U14729 ( .A1(n10094), .A2(n12389), .ZN(n12390) );
  NAND2_X1 U14730 ( .A1(n12390), .A2(n12394), .ZN(n12396) );
  OAI211_X1 U14731 ( .C1(n12396), .C2(n12392), .A(n12391), .B(n12404), .ZN(
        n12397) );
  INV_X1 U14732 ( .A(n12392), .ZN(n14982) );
  NAND3_X1 U14733 ( .A1(n14993), .A2(n12394), .A3(n12393), .ZN(n12395) );
  MUX2_X1 U14734 ( .A(n12397), .B(n7376), .S(n12514), .Z(n12398) );
  NAND2_X1 U14735 ( .A1(n12398), .A2(n12400), .ZN(n12403) );
  NAND2_X1 U14736 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NAND2_X1 U14737 ( .A1(n12401), .A2(n12514), .ZN(n12402) );
  NAND2_X1 U14738 ( .A1(n12403), .A2(n12402), .ZN(n12408) );
  NOR2_X1 U14739 ( .A1(n12404), .A2(n12525), .ZN(n12405) );
  NOR2_X1 U14740 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  NAND2_X1 U14741 ( .A1(n12408), .A2(n12407), .ZN(n12413) );
  NAND3_X1 U14742 ( .A1(n12413), .A2(n12565), .A3(n12409), .ZN(n12411) );
  NAND3_X1 U14743 ( .A1(n12411), .A2(n12410), .A3(n12415), .ZN(n12420) );
  NAND3_X1 U14744 ( .A1(n12413), .A2(n12565), .A3(n12412), .ZN(n12418) );
  AND2_X1 U14745 ( .A1(n12422), .A2(n12414), .ZN(n12417) );
  INV_X1 U14746 ( .A(n12415), .ZN(n12416) );
  AOI21_X1 U14747 ( .B1(n12418), .B2(n12417), .A(n12416), .ZN(n12419) );
  MUX2_X1 U14748 ( .A(n12420), .B(n12419), .S(n12525), .Z(n12421) );
  OAI211_X1 U14749 ( .C1(n12525), .C2(n12422), .A(n12421), .B(n14944), .ZN(
        n12426) );
  NAND2_X1 U14750 ( .A1(n12609), .A2(n14954), .ZN(n12423) );
  MUX2_X1 U14751 ( .A(n12424), .B(n12423), .S(n12514), .Z(n12425) );
  NAND3_X1 U14752 ( .A1(n12426), .A2(n12569), .A3(n12425), .ZN(n12431) );
  INV_X1 U14753 ( .A(n12427), .ZN(n12568) );
  MUX2_X1 U14754 ( .A(n12429), .B(n12428), .S(n12525), .Z(n12430) );
  NAND3_X1 U14755 ( .A1(n12431), .A2(n12568), .A3(n12430), .ZN(n12436) );
  MUX2_X1 U14756 ( .A(n14935), .B(n12432), .S(n12525), .Z(n12434) );
  NAND2_X1 U14757 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  NAND2_X1 U14758 ( .A1(n12436), .A2(n12435), .ZN(n12441) );
  MUX2_X1 U14759 ( .A(n12438), .B(n12437), .S(n12525), .Z(n12439) );
  NAND2_X1 U14760 ( .A1(n14205), .A2(n12439), .ZN(n12440) );
  AOI21_X1 U14761 ( .B1(n12441), .B2(n7348), .A(n12440), .ZN(n12451) );
  NAND2_X1 U14762 ( .A1(n12448), .A2(n12442), .ZN(n12445) );
  NAND2_X1 U14763 ( .A1(n12447), .A2(n12443), .ZN(n12444) );
  MUX2_X1 U14764 ( .A(n12445), .B(n12444), .S(n12525), .Z(n12450) );
  INV_X1 U14765 ( .A(n12446), .ZN(n12452) );
  OR2_X1 U14766 ( .A1(n12453), .A2(n12452), .ZN(n14186) );
  INV_X1 U14767 ( .A(n14186), .ZN(n14191) );
  MUX2_X1 U14768 ( .A(n12448), .B(n12447), .S(n12514), .Z(n12449) );
  OAI211_X1 U14769 ( .C1(n12451), .C2(n12450), .A(n14191), .B(n12449), .ZN(
        n12457) );
  MUX2_X1 U14770 ( .A(n12453), .B(n12452), .S(n12525), .Z(n12454) );
  INV_X1 U14771 ( .A(n12454), .ZN(n12455) );
  NAND3_X1 U14772 ( .A1(n12457), .A2(n12456), .A3(n12455), .ZN(n12458) );
  OAI21_X1 U14773 ( .B1(n12459), .B2(n12514), .A(n12458), .ZN(n12461) );
  NAND2_X1 U14774 ( .A1(n12461), .A2(n12460), .ZN(n12466) );
  OAI211_X1 U14775 ( .C1(n12575), .C2(n12463), .A(n12469), .B(n12462), .ZN(
        n12464) );
  NAND2_X1 U14776 ( .A1(n12464), .A2(n12514), .ZN(n12465) );
  AOI21_X1 U14777 ( .B1(n12466), .B2(n12465), .A(n6994), .ZN(n12471) );
  AOI21_X1 U14778 ( .B1(n12468), .B2(n12467), .A(n12514), .ZN(n12470) );
  OAI22_X1 U14779 ( .A1(n12471), .A2(n12470), .B1(n12514), .B2(n12469), .ZN(
        n12478) );
  INV_X1 U14780 ( .A(n12472), .ZN(n12477) );
  NAND2_X1 U14781 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  AOI21_X1 U14782 ( .B1(n12475), .B2(n12479), .A(n12514), .ZN(n12476) );
  NAND2_X1 U14783 ( .A1(n12476), .A2(n12485), .ZN(n12480) );
  AOI22_X1 U14784 ( .A1(n12478), .A2(n12912), .B1(n12477), .B2(n12480), .ZN(
        n12483) );
  NAND2_X1 U14785 ( .A1(n12479), .A2(n12514), .ZN(n12481) );
  OAI21_X1 U14786 ( .B1(n12484), .B2(n12481), .A(n12480), .ZN(n12482) );
  OAI21_X1 U14787 ( .B1(n12483), .B2(n9429), .A(n12482), .ZN(n12487) );
  MUX2_X1 U14788 ( .A(n12485), .B(n7014), .S(n12525), .Z(n12486) );
  NAND3_X1 U14789 ( .A1(n12487), .A2(n12873), .A3(n12486), .ZN(n12491) );
  XNOR2_X1 U14790 ( .A(n12860), .B(n12872), .ZN(n12859) );
  MUX2_X1 U14791 ( .A(n12489), .B(n12488), .S(n12525), .Z(n12490) );
  NAND3_X1 U14792 ( .A1(n12491), .A2(n12859), .A3(n12490), .ZN(n12495) );
  MUX2_X1 U14793 ( .A(n12493), .B(n12492), .S(n12525), .Z(n12494) );
  AND2_X1 U14794 ( .A1(n12495), .A2(n12494), .ZN(n12496) );
  NAND2_X1 U14795 ( .A1(n12497), .A2(n12496), .ZN(n12499) );
  AND3_X1 U14796 ( .A1(n12839), .A2(n12498), .A3(n12499), .ZN(n12504) );
  NAND3_X1 U14797 ( .A1(n12839), .A2(n12500), .A3(n12499), .ZN(n12502) );
  NAND2_X1 U14798 ( .A1(n12502), .A2(n12501), .ZN(n12503) );
  MUX2_X1 U14799 ( .A(n12504), .B(n12503), .S(n12525), .Z(n12505) );
  NAND2_X1 U14800 ( .A1(n12811), .A2(n12505), .ZN(n12506) );
  OAI211_X1 U14801 ( .C1(n12508), .C2(n12507), .A(n12797), .B(n12506), .ZN(
        n12512) );
  MUX2_X1 U14802 ( .A(n12510), .B(n12509), .S(n12525), .Z(n12511) );
  MUX2_X1 U14803 ( .A(n12516), .B(n12515), .S(n12514), .Z(n12517) );
  OAI211_X1 U14804 ( .C1(n12519), .C2(n12518), .A(n12522), .B(n12521), .ZN(
        n12520) );
  INV_X1 U14805 ( .A(n12521), .ZN(n12524) );
  OAI21_X1 U14806 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(n12526) );
  NAND2_X1 U14807 ( .A1(n12527), .A2(n12537), .ZN(n12530) );
  OR2_X1 U14808 ( .A1(n6481), .A2(n12528), .ZN(n12529) );
  NAND2_X1 U14809 ( .A1(n12530), .A2(n12529), .ZN(n13001) );
  AND2_X1 U14810 ( .A1(n13001), .A2(n12548), .ZN(n12585) );
  INV_X1 U14811 ( .A(n12585), .ZN(n12532) );
  AND2_X1 U14812 ( .A1(n12532), .A2(n12531), .ZN(n12553) );
  INV_X1 U14813 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14117) );
  XNOR2_X1 U14814 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12535) );
  INV_X1 U14815 ( .A(SI_31_), .ZN(n13053) );
  NOR2_X1 U14816 ( .A1(n6481), .A2(n13053), .ZN(n12536) );
  INV_X1 U14817 ( .A(n12749), .ZN(n12997) );
  INV_X1 U14818 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U14819 ( .A1(n12538), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12542) );
  INV_X1 U14820 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12539) );
  OR2_X1 U14821 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  OAI211_X1 U14822 ( .C1(n12544), .C2(n12543), .A(n12542), .B(n12541), .ZN(
        n12545) );
  INV_X1 U14823 ( .A(n12545), .ZN(n12546) );
  NAND2_X1 U14824 ( .A1(n12547), .A2(n12546), .ZN(n12598) );
  INV_X1 U14825 ( .A(n12598), .ZN(n12746) );
  OR2_X1 U14826 ( .A1(n13001), .A2(n12548), .ZN(n12555) );
  AND2_X1 U14827 ( .A1(n12749), .A2(n12598), .ZN(n12586) );
  AOI21_X1 U14828 ( .B1(n12549), .B2(n6582), .A(n12586), .ZN(n12591) );
  INV_X1 U14829 ( .A(n12550), .ZN(n12551) );
  INV_X1 U14830 ( .A(n13001), .ZN(n12938) );
  INV_X1 U14831 ( .A(n12586), .ZN(n12554) );
  OAI211_X1 U14832 ( .C1(n12938), .C2(n12598), .A(n12554), .B(n12553), .ZN(
        n12558) );
  INV_X1 U14833 ( .A(n12555), .ZN(n12556) );
  NOR2_X1 U14834 ( .A1(n12556), .A2(n12746), .ZN(n12557) );
  XNOR2_X1 U14835 ( .A(n12561), .B(n12899), .ZN(n12887) );
  NAND3_X1 U14836 ( .A1(n14982), .A2(n12563), .A3(n12562), .ZN(n12567) );
  INV_X1 U14837 ( .A(n10119), .ZN(n14994) );
  NAND4_X1 U14838 ( .A1(n14994), .A2(n14960), .A3(n12565), .A4(n12564), .ZN(
        n12566) );
  NOR2_X1 U14839 ( .A1(n12567), .A2(n12566), .ZN(n12570) );
  NAND4_X1 U14840 ( .A1(n12570), .A2(n12569), .A3(n14944), .A4(n12568), .ZN(
        n12571) );
  NOR2_X1 U14841 ( .A1(n12571), .A2(n14933), .ZN(n12572) );
  NAND3_X1 U14842 ( .A1(n12573), .A2(n14205), .A3(n12572), .ZN(n12574) );
  OR3_X1 U14843 ( .A1(n12575), .A2(n14186), .A3(n12574), .ZN(n12576) );
  NOR2_X1 U14844 ( .A1(n12576), .A2(n9353), .ZN(n12577) );
  NAND4_X1 U14845 ( .A1(n12897), .A2(n12923), .A3(n12912), .A4(n12577), .ZN(
        n12578) );
  NOR2_X1 U14846 ( .A1(n12887), .A2(n12578), .ZN(n12579) );
  NAND3_X1 U14847 ( .A1(n12859), .A2(n12873), .A3(n12579), .ZN(n12580) );
  NOR2_X1 U14848 ( .A1(n12847), .A2(n12580), .ZN(n12581) );
  NAND4_X1 U14849 ( .A1(n12797), .A2(n12839), .A3(n12811), .A4(n12581), .ZN(
        n12582) );
  NOR2_X1 U14850 ( .A1(n12582), .A2(n12785), .ZN(n12583) );
  OAI22_X1 U14851 ( .A1(n12589), .A2(n12588), .B1(n12591), .B2(n12587), .ZN(
        n12590) );
  NAND3_X1 U14852 ( .A1(n12593), .A2(n12592), .A3(n12729), .ZN(n12594) );
  OAI211_X1 U14853 ( .C1(n12595), .C2(n12597), .A(n12594), .B(P3_B_REG_SCAN_IN), .ZN(n12596) );
  MUX2_X1 U14854 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12598), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14855 ( .A(n12757), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12603), .Z(
        P3_U3520) );
  MUX2_X1 U14856 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12599), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14857 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12758), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14858 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12802), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14859 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12600), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14860 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12832), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14861 ( .A(n12818), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12603), .Z(
        P3_U3514) );
  MUX2_X1 U14862 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12831), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14863 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12872), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14864 ( .A(n12601), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12603), .Z(
        P3_U3511) );
  MUX2_X1 U14865 ( .A(n12866), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12603), .Z(
        P3_U3510) );
  MUX2_X1 U14866 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12910), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14867 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12602), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14868 ( .A(n12909), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12603), .Z(
        P3_U3507) );
  MUX2_X1 U14869 ( .A(n12604), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12603), .Z(
        P3_U3506) );
  MUX2_X1 U14870 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12605), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14871 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12606), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14872 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12607), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14873 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n14936), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14874 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12608), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14875 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n14935), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14876 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n14950), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14877 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12609), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14878 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n14949), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14879 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12610), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14880 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n14963), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14881 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12611), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14882 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n14964), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14883 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12612), .S(P3_U3897), .Z(
        P3_U3492) );
  NOR2_X1 U14884 ( .A1(n12625), .A2(n12613), .ZN(n12615) );
  XNOR2_X1 U14885 ( .A(n12644), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12626) );
  AOI21_X1 U14886 ( .B1(n6591), .B2(n12626), .A(n12639), .ZN(n12638) );
  NAND2_X1 U14887 ( .A1(n12617), .A2(n12616), .ZN(n12619) );
  NAND2_X1 U14888 ( .A1(n12619), .A2(n12618), .ZN(n12621) );
  NAND2_X1 U14889 ( .A1(n12644), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12645) );
  OR2_X1 U14890 ( .A1(n12644), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12620) );
  AND2_X1 U14891 ( .A1(n12645), .A2(n12620), .ZN(n12629) );
  NAND2_X1 U14892 ( .A1(n12629), .A2(n12621), .ZN(n12642) );
  OAI21_X1 U14893 ( .B1(n12621), .B2(n12629), .A(n12642), .ZN(n12636) );
  INV_X1 U14894 ( .A(n12622), .ZN(n12624) );
  AOI21_X1 U14895 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n12631) );
  INV_X1 U14896 ( .A(n12626), .ZN(n12628) );
  MUX2_X1 U14897 ( .A(n12629), .B(n12628), .S(n12627), .Z(n12630) );
  NAND2_X1 U14898 ( .A1(n12631), .A2(n12630), .ZN(n12648) );
  OAI211_X1 U14899 ( .C1(n12631), .C2(n12630), .A(n12648), .B(n14892), .ZN(
        n12634) );
  AOI21_X1 U14900 ( .B1(n14899), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12632), 
        .ZN(n12633) );
  OAI211_X1 U14901 ( .C1(n14896), .C2(n12644), .A(n12634), .B(n12633), .ZN(
        n12635) );
  AOI21_X1 U14902 ( .B1(n12636), .B2(n14910), .A(n12635), .ZN(n12637) );
  OAI21_X1 U14903 ( .B1(n12638), .B2(n14921), .A(n12637), .ZN(P3_U3196) );
  AOI21_X1 U14904 ( .B1(n12641), .B2(n12640), .A(n12662), .ZN(n12659) );
  OAI21_X1 U14905 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12643), .A(n12668), 
        .ZN(n12657) );
  MUX2_X1 U14906 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12729), .Z(n12650) );
  NAND2_X1 U14907 ( .A1(n12644), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12646) );
  MUX2_X1 U14908 ( .A(n12646), .B(n12645), .S(n12729), .Z(n12647) );
  NAND2_X1 U14909 ( .A1(n12648), .A2(n12647), .ZN(n12672) );
  XNOR2_X1 U14910 ( .A(n12672), .B(n12667), .ZN(n12649) );
  NOR2_X1 U14911 ( .A1(n12649), .A2(n12650), .ZN(n12673) );
  AOI21_X1 U14912 ( .B1(n12650), .B2(n12649), .A(n12673), .ZN(n12655) );
  NOR2_X1 U14913 ( .A1(n14930), .A2(n12651), .ZN(n12652) );
  AOI211_X1 U14914 ( .C1(n14926), .C2(n12674), .A(n12653), .B(n12652), .ZN(
        n12654) );
  OAI21_X1 U14915 ( .B1(n12655), .B2(n14915), .A(n12654), .ZN(n12656) );
  AOI21_X1 U14916 ( .B1(n14910), .B2(n12657), .A(n12656), .ZN(n12658) );
  OAI21_X1 U14917 ( .B1(n12659), .B2(n14921), .A(n12658), .ZN(P3_U3197) );
  NOR2_X1 U14918 ( .A1(n12674), .A2(n12660), .ZN(n12661) );
  NOR2_X1 U14919 ( .A1(n12662), .A2(n12661), .ZN(n12665) );
  NAND2_X1 U14920 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12706), .ZN(n12663) );
  OAI21_X1 U14921 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12706), .A(n12663), 
        .ZN(n12664) );
  AOI21_X1 U14922 ( .B1(n12665), .B2(n12664), .A(n12695), .ZN(n12688) );
  INV_X1 U14923 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U14924 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12706), .B1(n12682), 
        .B2(n12994), .ZN(n12671) );
  NAND2_X1 U14925 ( .A1(n12667), .A2(n12666), .ZN(n12669) );
  NAND2_X1 U14926 ( .A1(n12671), .A2(n12670), .ZN(n12707) );
  OAI21_X1 U14927 ( .B1(n12671), .B2(n12670), .A(n12707), .ZN(n12686) );
  INV_X1 U14928 ( .A(n12672), .ZN(n12675) );
  AOI21_X1 U14929 ( .B1(n12675), .B2(n12674), .A(n12673), .ZN(n12691) );
  MUX2_X1 U14930 ( .A(n6904), .B(n12994), .S(n12729), .Z(n12676) );
  NOR2_X1 U14931 ( .A1(n12676), .A2(n12682), .ZN(n12690) );
  NAND2_X1 U14932 ( .A1(n12676), .A2(n12682), .ZN(n12689) );
  INV_X1 U14933 ( .A(n12689), .ZN(n12677) );
  NOR2_X1 U14934 ( .A1(n12690), .A2(n12677), .ZN(n12678) );
  XNOR2_X1 U14935 ( .A(n12691), .B(n12678), .ZN(n12684) );
  NOR2_X1 U14936 ( .A1(n14930), .A2(n12679), .ZN(n12680) );
  AOI211_X1 U14937 ( .C1(n14926), .C2(n12682), .A(n12681), .B(n12680), .ZN(
        n12683) );
  OAI21_X1 U14938 ( .B1(n12684), .B2(n14915), .A(n12683), .ZN(n12685) );
  AOI21_X1 U14939 ( .B1(n14910), .B2(n12686), .A(n12685), .ZN(n12687) );
  OAI21_X1 U14940 ( .B1(n12688), .B2(n14921), .A(n12687), .ZN(P3_U3198) );
  MUX2_X1 U14941 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12729), .Z(n12694) );
  MUX2_X1 U14942 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12729), .Z(n12692) );
  OAI21_X1 U14943 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(n14178) );
  XNOR2_X1 U14944 ( .A(n12692), .B(n12709), .ZN(n14179) );
  NOR2_X1 U14945 ( .A1(n14178), .A2(n14179), .ZN(n14177) );
  AOI21_X1 U14946 ( .B1(n12692), .B2(n12709), .A(n14177), .ZN(n12727) );
  XNOR2_X1 U14947 ( .A(n12727), .B(n12726), .ZN(n12693) );
  NOR2_X1 U14948 ( .A1(n12693), .A2(n12694), .ZN(n12725) );
  AOI21_X1 U14949 ( .B1(n12694), .B2(n12693), .A(n12725), .ZN(n12719) );
  INV_X1 U14950 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14170) );
  OR2_X1 U14951 ( .A1(n12696), .A2(n14173), .ZN(n12700) );
  INV_X1 U14952 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12697) );
  OR2_X1 U14953 ( .A1(n12726), .A2(n12697), .ZN(n12720) );
  NAND2_X1 U14954 ( .A1(n12726), .A2(n12697), .ZN(n12698) );
  NAND2_X1 U14955 ( .A1(n12720), .A2(n12698), .ZN(n12699) );
  AND3_X1 U14956 ( .A1(n12701), .A2(n12700), .A3(n12699), .ZN(n12703) );
  OAI21_X1 U14957 ( .B1(n12722), .B2(n12703), .A(n12702), .ZN(n12718) );
  INV_X1 U14958 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12705) );
  OAI21_X1 U14959 ( .B1(n14930), .B2(n12705), .A(n12704), .ZN(n12716) );
  NAND2_X1 U14960 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12706), .ZN(n12708) );
  NAND2_X1 U14961 ( .A1(n12710), .A2(n12709), .ZN(n12712) );
  INV_X1 U14962 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12986) );
  XNOR2_X1 U14963 ( .A(n12726), .B(n12986), .ZN(n12711) );
  INV_X1 U14964 ( .A(n12733), .ZN(n12714) );
  NAND3_X1 U14965 ( .A1(n12712), .A2(n14171), .A3(n12711), .ZN(n12713) );
  AOI21_X1 U14966 ( .B1(n12714), .B2(n12713), .A(n14769), .ZN(n12715) );
  AOI211_X1 U14967 ( .C1(n14926), .C2(n12726), .A(n12716), .B(n12715), .ZN(
        n12717) );
  OAI211_X1 U14968 ( .C1(n12719), .C2(n14915), .A(n12718), .B(n12717), .ZN(
        P3_U3200) );
  INV_X1 U14969 ( .A(n12720), .ZN(n12721) );
  NOR2_X1 U14970 ( .A1(n12722), .A2(n12721), .ZN(n12724) );
  XNOR2_X1 U14971 ( .A(n12723), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12728) );
  XNOR2_X1 U14972 ( .A(n12724), .B(n12728), .ZN(n12743) );
  AOI21_X1 U14973 ( .B1(n12727), .B2(n12726), .A(n12725), .ZN(n12732) );
  INV_X1 U14974 ( .A(n12728), .ZN(n12730) );
  XNOR2_X1 U14975 ( .A(n12740), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12735) );
  MUX2_X1 U14976 ( .A(n12730), .B(n12735), .S(n12729), .Z(n12731) );
  XNOR2_X1 U14977 ( .A(n12732), .B(n12731), .ZN(n12742) );
  AOI21_X1 U14978 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n12734), .A(n12733), 
        .ZN(n12737) );
  INV_X1 U14979 ( .A(n12735), .ZN(n12736) );
  NAND2_X1 U14980 ( .A1(n14899), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12738) );
  OAI211_X1 U14981 ( .C1(n14896), .C2(n12740), .A(n12739), .B(n12738), .ZN(
        n12741) );
  NAND2_X1 U14982 ( .A1(n12744), .A2(n15007), .ZN(n12747) );
  OR2_X1 U14983 ( .A1(n12746), .A2(n12745), .ZN(n12933) );
  AOI21_X1 U14984 ( .B1(n12747), .B2(n12933), .A(n15012), .ZN(n12750) );
  AOI21_X1 U14985 ( .B1(n15012), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12750), 
        .ZN(n12748) );
  OAI21_X1 U14986 ( .B1(n12749), .B2(n12928), .A(n12748), .ZN(P3_U3202) );
  AOI21_X1 U14987 ( .B1(n15012), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12750), 
        .ZN(n12751) );
  OAI21_X1 U14988 ( .B1(n12938), .B2(n12928), .A(n12751), .ZN(P3_U3203) );
  NAND2_X1 U14989 ( .A1(n12768), .A2(n12752), .ZN(n12754) );
  XNOR2_X1 U14990 ( .A(n12754), .B(n12753), .ZN(n12940) );
  INV_X1 U14991 ( .A(n12940), .ZN(n12765) );
  OAI211_X1 U14992 ( .C1(n12756), .C2(n9586), .A(n15001), .B(n12755), .ZN(
        n12760) );
  AOI22_X1 U14993 ( .A1(n14965), .A2(n12758), .B1(n12757), .B2(n14962), .ZN(
        n12759) );
  NAND2_X1 U14994 ( .A1(n12760), .A2(n12759), .ZN(n12939) );
  AOI22_X1 U14995 ( .A1(n12761), .A2(n15007), .B1(n15012), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12762) );
  OAI21_X1 U14996 ( .B1(n13007), .B2(n12928), .A(n12762), .ZN(n12763) );
  AOI21_X1 U14997 ( .B1(n12939), .B2(n15010), .A(n12763), .ZN(n12764) );
  OAI21_X1 U14998 ( .B1(n12765), .B2(n14209), .A(n12764), .ZN(P3_U3205) );
  OR2_X1 U14999 ( .A1(n12766), .A2(n12769), .ZN(n12767) );
  OAI21_X1 U15000 ( .B1(n12771), .B2(n9573), .A(n12770), .ZN(n12775) );
  OAI22_X1 U15001 ( .A1(n12773), .A2(n14996), .B1(n12772), .B2(n14998), .ZN(
        n12774) );
  AOI21_X1 U15002 ( .B1(n12775), .B2(n15001), .A(n12774), .ZN(n12776) );
  OAI21_X1 U15003 ( .B1(n15004), .B2(n12943), .A(n12776), .ZN(n12944) );
  AOI22_X1 U15004 ( .A1(n12777), .A2(n15007), .B1(n15012), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U15005 ( .A1(n12778), .A2(n12878), .ZN(n12779) );
  OAI211_X1 U15006 ( .C1(n12943), .C2(n12794), .A(n12780), .B(n12779), .ZN(
        n12781) );
  AOI21_X1 U15007 ( .B1(n12944), .B2(n15010), .A(n12781), .ZN(n12782) );
  INV_X1 U15008 ( .A(n12782), .ZN(P3_U3206) );
  XNOR2_X1 U15009 ( .A(n12783), .B(n12785), .ZN(n12948) );
  XOR2_X1 U15010 ( .A(n12785), .B(n12784), .Z(n12788) );
  OAI22_X1 U15011 ( .A1(n12786), .A2(n14996), .B1(n12821), .B2(n14998), .ZN(
        n12787) );
  AOI21_X1 U15012 ( .B1(n12788), .B2(n15001), .A(n12787), .ZN(n12789) );
  OAI21_X1 U15013 ( .B1(n15004), .B2(n12948), .A(n12789), .ZN(n12949) );
  AOI22_X1 U15014 ( .A1(n12790), .A2(n15007), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n15012), .ZN(n12793) );
  NAND2_X1 U15015 ( .A1(n12791), .A2(n12878), .ZN(n12792) );
  OAI211_X1 U15016 ( .C1(n12948), .C2(n12794), .A(n12793), .B(n12792), .ZN(
        n12795) );
  AOI21_X1 U15017 ( .B1(n12949), .B2(n15010), .A(n12795), .ZN(n12796) );
  INV_X1 U15018 ( .A(n12796), .ZN(P3_U3207) );
  XNOR2_X1 U15019 ( .A(n12798), .B(n12797), .ZN(n12954) );
  INV_X1 U15020 ( .A(n12954), .ZN(n12809) );
  OAI211_X1 U15021 ( .C1(n12801), .C2(n12800), .A(n12799), .B(n15001), .ZN(
        n12804) );
  AOI22_X1 U15022 ( .A1(n12802), .A2(n14962), .B1(n14965), .B2(n12832), .ZN(
        n12803) );
  NAND2_X1 U15023 ( .A1(n12804), .A2(n12803), .ZN(n12953) );
  AOI22_X1 U15024 ( .A1(n12805), .A2(n15007), .B1(n15012), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12806) );
  OAI21_X1 U15025 ( .B1(n13019), .B2(n12928), .A(n12806), .ZN(n12807) );
  AOI21_X1 U15026 ( .B1(n12953), .B2(n15010), .A(n12807), .ZN(n12808) );
  OAI21_X1 U15027 ( .B1(n14209), .B2(n12809), .A(n12808), .ZN(P3_U3208) );
  INV_X1 U15028 ( .A(n12810), .ZN(n12814) );
  AOI21_X1 U15029 ( .B1(n12961), .B2(n12812), .A(n12811), .ZN(n12813) );
  NOR2_X1 U15030 ( .A1(n12814), .A2(n12813), .ZN(n12960) );
  OAI211_X1 U15031 ( .C1(n12817), .C2(n12816), .A(n12815), .B(n15001), .ZN(
        n12820) );
  NAND2_X1 U15032 ( .A1(n12818), .A2(n14965), .ZN(n12819) );
  OAI211_X1 U15033 ( .C1(n12821), .C2(n14996), .A(n12820), .B(n12819), .ZN(
        n12957) );
  NAND2_X1 U15034 ( .A1(n12957), .A2(n15010), .ZN(n12827) );
  INV_X1 U15035 ( .A(n12822), .ZN(n12824) );
  INV_X1 U15036 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12823) );
  OAI22_X1 U15037 ( .A1(n12824), .A2(n14978), .B1(n15010), .B2(n12823), .ZN(
        n12825) );
  AOI21_X1 U15038 ( .B1(n12958), .B2(n12878), .A(n12825), .ZN(n12826) );
  OAI211_X1 U15039 ( .C1(n12960), .C2(n14209), .A(n12827), .B(n12826), .ZN(
        P3_U3209) );
  NAND2_X1 U15040 ( .A1(n12829), .A2(n12839), .ZN(n12830) );
  NAND3_X1 U15041 ( .A1(n12828), .A2(n15001), .A3(n12830), .ZN(n12834) );
  AOI22_X1 U15042 ( .A1(n12832), .A2(n14962), .B1(n14965), .B2(n12831), .ZN(
        n12833) );
  INV_X1 U15043 ( .A(n12835), .ZN(n12837) );
  INV_X1 U15044 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12836) );
  OAI22_X1 U15045 ( .A1(n12837), .A2(n14978), .B1(n15010), .B2(n12836), .ZN(
        n12838) );
  AOI21_X1 U15046 ( .B1(n12963), .B2(n12878), .A(n12838), .ZN(n12842) );
  OR2_X1 U15047 ( .A1(n12840), .A2(n12839), .ZN(n12962) );
  NAND3_X1 U15048 ( .A1(n12962), .A2(n12961), .A3(n12930), .ZN(n12841) );
  OAI211_X1 U15049 ( .C1(n12967), .C2(n15012), .A(n12842), .B(n12841), .ZN(
        P3_U3210) );
  XNOR2_X1 U15050 ( .A(n12843), .B(n12847), .ZN(n12844) );
  OAI222_X1 U15051 ( .A1(n14998), .A2(n12846), .B1(n14996), .B2(n12845), .C1(
        n12844), .C2(n14988), .ZN(n12968) );
  INV_X1 U15052 ( .A(n12968), .ZN(n12854) );
  XNOR2_X1 U15053 ( .A(n12848), .B(n12847), .ZN(n12969) );
  INV_X1 U15054 ( .A(n12849), .ZN(n13025) );
  AOI22_X1 U15055 ( .A1(n12850), .A2(n15007), .B1(n15012), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U15056 ( .B1(n13025), .B2(n12928), .A(n12851), .ZN(n12852) );
  AOI21_X1 U15057 ( .B1(n12969), .B2(n12930), .A(n12852), .ZN(n12853) );
  OAI21_X1 U15058 ( .B1(n12854), .B2(n15012), .A(n12853), .ZN(P3_U3211) );
  XOR2_X1 U15059 ( .A(n12855), .B(n12859), .Z(n12856) );
  OAI222_X1 U15060 ( .A1(n14998), .A2(n12885), .B1(n14996), .B2(n12857), .C1(
        n14988), .C2(n12856), .ZN(n12972) );
  INV_X1 U15061 ( .A(n12972), .ZN(n12865) );
  XOR2_X1 U15062 ( .A(n12859), .B(n12858), .Z(n12973) );
  INV_X1 U15063 ( .A(n12860), .ZN(n13029) );
  AOI22_X1 U15064 ( .A1(n15012), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12861), 
        .B2(n15007), .ZN(n12862) );
  OAI21_X1 U15065 ( .B1(n13029), .B2(n12928), .A(n12862), .ZN(n12863) );
  AOI21_X1 U15066 ( .B1(n12973), .B2(n12930), .A(n12863), .ZN(n12864) );
  OAI21_X1 U15067 ( .B1(n12865), .B2(n15012), .A(n12864), .ZN(P3_U3212) );
  AND2_X1 U15068 ( .A1(n12866), .A2(n14965), .ZN(n12871) );
  INV_X1 U15069 ( .A(n12867), .ZN(n12868) );
  AOI211_X1 U15070 ( .C1(n12873), .C2(n12869), .A(n14988), .B(n12868), .ZN(
        n12870) );
  AOI211_X1 U15071 ( .C1(n14962), .C2(n12872), .A(n12871), .B(n12870), .ZN(
        n12978) );
  OR2_X1 U15072 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U15073 ( .A1(n12876), .A2(n12875), .ZN(n12979) );
  AOI22_X1 U15074 ( .A1(n15012), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15007), 
        .B2(n12877), .ZN(n12880) );
  NAND2_X1 U15075 ( .A1(n12976), .A2(n12878), .ZN(n12879) );
  OAI211_X1 U15076 ( .C1(n12979), .C2(n14209), .A(n12880), .B(n12879), .ZN(
        n12881) );
  INV_X1 U15077 ( .A(n12881), .ZN(n12882) );
  OAI21_X1 U15078 ( .B1(n12978), .B2(n15012), .A(n12882), .ZN(P3_U3213) );
  XOR2_X1 U15079 ( .A(n12887), .B(n12883), .Z(n12884) );
  OAI222_X1 U15080 ( .A1(n14998), .A2(n12886), .B1(n14996), .B2(n12885), .C1(
        n12884), .C2(n14988), .ZN(n12980) );
  INV_X1 U15081 ( .A(n12980), .ZN(n12893) );
  XOR2_X1 U15082 ( .A(n12888), .B(n12887), .Z(n12981) );
  AOI22_X1 U15083 ( .A1(n15012), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15007), 
        .B2(n12889), .ZN(n12890) );
  OAI21_X1 U15084 ( .B1(n13034), .B2(n12928), .A(n12890), .ZN(n12891) );
  AOI21_X1 U15085 ( .B1(n12981), .B2(n12930), .A(n12891), .ZN(n12892) );
  OAI21_X1 U15086 ( .B1(n12893), .B2(n15012), .A(n12892), .ZN(P3_U3214) );
  INV_X1 U15087 ( .A(n12894), .ZN(n12895) );
  AOI21_X1 U15088 ( .B1(n12897), .B2(n12896), .A(n12895), .ZN(n12898) );
  OAI222_X1 U15089 ( .A1(n14998), .A2(n12922), .B1(n14996), .B2(n12899), .C1(
        n14988), .C2(n12898), .ZN(n12984) );
  INV_X1 U15090 ( .A(n12984), .ZN(n12907) );
  INV_X1 U15091 ( .A(n12900), .ZN(n12901) );
  AOI21_X1 U15092 ( .B1(n9429), .B2(n12902), .A(n12901), .ZN(n12985) );
  AOI22_X1 U15093 ( .A1(n15012), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15007), 
        .B2(n12903), .ZN(n12904) );
  OAI21_X1 U15094 ( .B1(n13038), .B2(n12928), .A(n12904), .ZN(n12905) );
  AOI21_X1 U15095 ( .B1(n12985), .B2(n12930), .A(n12905), .ZN(n12906) );
  OAI21_X1 U15096 ( .B1(n12907), .B2(n15012), .A(n12906), .ZN(P3_U3215) );
  XNOR2_X1 U15097 ( .A(n12908), .B(n12912), .ZN(n12911) );
  AOI222_X1 U15098 ( .A1(n15001), .A2(n12911), .B1(n12910), .B2(n14962), .C1(
        n12909), .C2(n14965), .ZN(n12991) );
  XNOR2_X1 U15099 ( .A(n12913), .B(n12912), .ZN(n12989) );
  AOI22_X1 U15100 ( .A1(n15012), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15007), 
        .B2(n12914), .ZN(n12915) );
  OAI21_X1 U15101 ( .B1(n12916), .B2(n12928), .A(n12915), .ZN(n12917) );
  AOI21_X1 U15102 ( .B1(n12989), .B2(n12930), .A(n12917), .ZN(n12918) );
  OAI21_X1 U15103 ( .B1(n12991), .B2(n15012), .A(n12918), .ZN(P3_U3216) );
  XOR2_X1 U15104 ( .A(n12919), .B(n12923), .Z(n12920) );
  OAI222_X1 U15105 ( .A1(n14996), .A2(n12922), .B1(n14998), .B2(n12921), .C1(
        n12920), .C2(n14988), .ZN(n12992) );
  INV_X1 U15106 ( .A(n12992), .ZN(n12932) );
  XNOR2_X1 U15107 ( .A(n12924), .B(n12923), .ZN(n12993) );
  INV_X1 U15108 ( .A(n12925), .ZN(n13044) );
  AOI22_X1 U15109 ( .A1(n15012), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15007), 
        .B2(n12926), .ZN(n12927) );
  OAI21_X1 U15110 ( .B1(n13044), .B2(n12928), .A(n12927), .ZN(n12929) );
  AOI21_X1 U15111 ( .B1(n12993), .B2(n12930), .A(n12929), .ZN(n12931) );
  OAI21_X1 U15112 ( .B1(n12932), .B2(n15012), .A(n12931), .ZN(P3_U3217) );
  INV_X1 U15113 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U15114 ( .A1(n12997), .A2(n9689), .ZN(n12934) );
  INV_X1 U15115 ( .A(n12933), .ZN(n12998) );
  NAND2_X1 U15116 ( .A1(n12998), .A2(n15079), .ZN(n12937) );
  OAI211_X1 U15117 ( .C1(n15079), .C2(n12935), .A(n12934), .B(n12937), .ZN(
        P3_U3490) );
  NAND2_X1 U15118 ( .A1(n15077), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12936) );
  OAI211_X1 U15119 ( .C1(n12938), .C2(n12996), .A(n12937), .B(n12936), .ZN(
        P3_U3489) );
  INV_X1 U15120 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12941) );
  MUX2_X1 U15121 ( .A(n12941), .B(n13004), .S(n15079), .Z(n12942) );
  INV_X1 U15122 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12946) );
  INV_X1 U15123 ( .A(n12943), .ZN(n12945) );
  MUX2_X1 U15124 ( .A(n12946), .B(n13008), .S(n15079), .Z(n12947) );
  INV_X1 U15125 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12951) );
  INV_X1 U15126 ( .A(n12948), .ZN(n12950) );
  AOI21_X1 U15127 ( .B1(n15058), .B2(n12950), .A(n12949), .ZN(n13012) );
  MUX2_X1 U15128 ( .A(n12951), .B(n13012), .S(n15079), .Z(n12952) );
  OAI21_X1 U15129 ( .B1(n13015), .B2(n12996), .A(n12952), .ZN(P3_U3485) );
  INV_X1 U15130 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12955) );
  AOI21_X1 U15131 ( .B1(n12954), .B2(n15063), .A(n12953), .ZN(n13016) );
  MUX2_X1 U15132 ( .A(n12955), .B(n13016), .S(n15079), .Z(n12956) );
  OAI21_X1 U15133 ( .B1(n13019), .B2(n12996), .A(n12956), .ZN(P3_U3484) );
  INV_X1 U15134 ( .A(n15063), .ZN(n14217) );
  AOI21_X1 U15135 ( .B1(n15015), .B2(n12958), .A(n12957), .ZN(n12959) );
  OAI21_X1 U15136 ( .B1(n14217), .B2(n12960), .A(n12959), .ZN(n13020) );
  MUX2_X1 U15137 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13020), .S(n15079), .Z(
        P3_U3483) );
  NAND3_X1 U15138 ( .A1(n12962), .A2(n12961), .A3(n15063), .ZN(n12965) );
  NAND2_X1 U15139 ( .A1(n12963), .A2(n15015), .ZN(n12964) );
  AND2_X1 U15140 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  NAND2_X1 U15141 ( .A1(n12967), .A2(n12966), .ZN(n13021) );
  MUX2_X1 U15142 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13021), .S(n15079), .Z(
        P3_U3482) );
  INV_X1 U15143 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12970) );
  AOI21_X1 U15144 ( .B1(n15063), .B2(n12969), .A(n12968), .ZN(n13022) );
  MUX2_X1 U15145 ( .A(n12970), .B(n13022), .S(n15079), .Z(n12971) );
  OAI21_X1 U15146 ( .B1(n13025), .B2(n12996), .A(n12971), .ZN(P3_U3481) );
  INV_X1 U15147 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12974) );
  AOI21_X1 U15148 ( .B1(n12973), .B2(n15063), .A(n12972), .ZN(n13026) );
  MUX2_X1 U15149 ( .A(n12974), .B(n13026), .S(n15079), .Z(n12975) );
  OAI21_X1 U15150 ( .B1(n13029), .B2(n12996), .A(n12975), .ZN(P3_U3480) );
  NAND2_X1 U15151 ( .A1(n12976), .A2(n15015), .ZN(n12977) );
  OAI211_X1 U15152 ( .C1(n14217), .C2(n12979), .A(n12978), .B(n12977), .ZN(
        n13030) );
  MUX2_X1 U15153 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n13030), .S(n15079), .Z(
        P3_U3479) );
  INV_X1 U15154 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12982) );
  AOI21_X1 U15155 ( .B1(n12981), .B2(n15063), .A(n12980), .ZN(n13031) );
  MUX2_X1 U15156 ( .A(n12982), .B(n13031), .S(n15079), .Z(n12983) );
  OAI21_X1 U15157 ( .B1(n13034), .B2(n12996), .A(n12983), .ZN(P3_U3478) );
  AOI21_X1 U15158 ( .B1(n12985), .B2(n15063), .A(n12984), .ZN(n13035) );
  MUX2_X1 U15159 ( .A(n12986), .B(n13035), .S(n15079), .Z(n12987) );
  OAI21_X1 U15160 ( .B1(n13038), .B2(n12996), .A(n12987), .ZN(P3_U3477) );
  AOI22_X1 U15161 ( .A1(n12989), .A2(n15063), .B1(n15015), .B2(n12988), .ZN(
        n12990) );
  NAND2_X1 U15162 ( .A1(n12991), .A2(n12990), .ZN(n13039) );
  MUX2_X1 U15163 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13039), .S(n15079), .Z(
        P3_U3476) );
  AOI21_X1 U15164 ( .B1(n12993), .B2(n15063), .A(n12992), .ZN(n13040) );
  MUX2_X1 U15165 ( .A(n12994), .B(n13040), .S(n15079), .Z(n12995) );
  OAI21_X1 U15166 ( .B1(n13044), .B2(n12996), .A(n12995), .ZN(P3_U3475) );
  INV_X1 U15167 ( .A(n13043), .ZN(n13000) );
  NAND2_X1 U15168 ( .A1(n12997), .A2(n13000), .ZN(n12999) );
  NAND2_X1 U15169 ( .A1(n12998), .A2(n15066), .ZN(n13002) );
  OAI211_X1 U15170 ( .C1(n12544), .C2(n15066), .A(n12999), .B(n13002), .ZN(
        P3_U3458) );
  NAND2_X1 U15171 ( .A1(n13001), .A2(n13000), .ZN(n13003) );
  OAI211_X1 U15172 ( .C1(n9613), .C2(n15066), .A(n13003), .B(n13002), .ZN(
        P3_U3457) );
  MUX2_X1 U15173 ( .A(n13005), .B(n13004), .S(n15066), .Z(n13006) );
  MUX2_X1 U15174 ( .A(n13009), .B(n13008), .S(n15066), .Z(n13010) );
  MUX2_X1 U15175 ( .A(n13013), .B(n13012), .S(n15066), .Z(n13014) );
  OAI21_X1 U15176 ( .B1(n13015), .B2(n13043), .A(n13014), .ZN(P3_U3453) );
  MUX2_X1 U15177 ( .A(n13017), .B(n13016), .S(n15066), .Z(n13018) );
  OAI21_X1 U15178 ( .B1(n13019), .B2(n13043), .A(n13018), .ZN(P3_U3452) );
  MUX2_X1 U15179 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13020), .S(n15066), .Z(
        P3_U3451) );
  MUX2_X1 U15180 ( .A(n13021), .B(P3_REG0_REG_23__SCAN_IN), .S(n15064), .Z(
        P3_U3450) );
  MUX2_X1 U15181 ( .A(n13023), .B(n13022), .S(n15066), .Z(n13024) );
  OAI21_X1 U15182 ( .B1(n13025), .B2(n13043), .A(n13024), .ZN(P3_U3449) );
  MUX2_X1 U15183 ( .A(n13027), .B(n13026), .S(n15066), .Z(n13028) );
  OAI21_X1 U15184 ( .B1(n13029), .B2(n13043), .A(n13028), .ZN(P3_U3448) );
  MUX2_X1 U15185 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n13030), .S(n15066), .Z(
        P3_U3447) );
  INV_X1 U15186 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13032) );
  MUX2_X1 U15187 ( .A(n13032), .B(n13031), .S(n15066), .Z(n13033) );
  OAI21_X1 U15188 ( .B1(n13034), .B2(n13043), .A(n13033), .ZN(P3_U3446) );
  MUX2_X1 U15189 ( .A(n13036), .B(n13035), .S(n15066), .Z(n13037) );
  OAI21_X1 U15190 ( .B1(n13038), .B2(n13043), .A(n13037), .ZN(P3_U3444) );
  MUX2_X1 U15191 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13039), .S(n15066), .Z(
        P3_U3441) );
  MUX2_X1 U15192 ( .A(n13041), .B(n13040), .S(n15066), .Z(n13042) );
  OAI21_X1 U15193 ( .B1(n13044), .B2(n13043), .A(n13042), .ZN(P3_U3438) );
  MUX2_X1 U15194 ( .A(P3_D_REG_1__SCAN_IN), .B(n13045), .S(n13046), .Z(
        P3_U3377) );
  MUX2_X1 U15195 ( .A(P3_D_REG_0__SCAN_IN), .B(n13047), .S(n13046), .Z(
        P3_U3376) );
  NAND2_X1 U15196 ( .A1(n13049), .A2(n13048), .ZN(n13052) );
  OR4_X1 U15197 ( .A1(n13050), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n9098), .ZN(n13051) );
  OAI211_X1 U15198 ( .C1(n13053), .C2(n13058), .A(n13052), .B(n13051), .ZN(
        P3_U3264) );
  INV_X1 U15199 ( .A(n13054), .ZN(n13055) );
  OAI222_X1 U15200 ( .A1(n13058), .A2(n13057), .B1(n13056), .B2(n13055), .C1(
        P3_U3151), .C2(n9089), .ZN(P3_U3266) );
  XNOR2_X1 U15201 ( .A(n13060), .B(n13059), .ZN(n13065) );
  OAI22_X1 U15202 ( .A1(n13093), .A2(n13163), .B1(n13061), .B2(n13161), .ZN(
        n13252) );
  AOI22_X1 U15203 ( .A1(n14237), .A2(n13252), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13062) );
  OAI21_X1 U15204 ( .B1(n13258), .B2(n14243), .A(n13062), .ZN(n13063) );
  AOI21_X1 U15205 ( .B1(n13442), .B2(n14240), .A(n13063), .ZN(n13064) );
  OAI21_X1 U15206 ( .B1(n13065), .B2(n13168), .A(n13064), .ZN(P2_U3186) );
  XNOR2_X1 U15207 ( .A(n13066), .B(n13067), .ZN(n13073) );
  NAND2_X1 U15208 ( .A1(n13178), .A2(n13141), .ZN(n13069) );
  NAND2_X1 U15209 ( .A1(n13176), .A2(n13139), .ZN(n13068) );
  NAND2_X1 U15210 ( .A1(n13069), .A2(n13068), .ZN(n13467) );
  AOI22_X1 U15211 ( .A1(n14237), .A2(n13467), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13070) );
  OAI21_X1 U15212 ( .B1(n13308), .B2(n14243), .A(n13070), .ZN(n13071) );
  AOI21_X1 U15213 ( .B1(n13468), .B2(n14240), .A(n13071), .ZN(n13072) );
  OAI21_X1 U15214 ( .B1(n13073), .B2(n13168), .A(n13072), .ZN(P2_U3188) );
  AOI21_X1 U15215 ( .B1(n13075), .B2(n13074), .A(n6590), .ZN(n13082) );
  OAI22_X1 U15216 ( .A1(n13077), .A2(n13161), .B1(n13076), .B2(n13163), .ZN(
        n13497) );
  NOR2_X1 U15217 ( .A1(n13078), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13220) );
  AOI21_X1 U15218 ( .B1(n13497), .B2(n14237), .A(n13220), .ZN(n13079) );
  OAI21_X1 U15219 ( .B1(n13367), .B2(n14243), .A(n13079), .ZN(n13080) );
  AOI21_X1 U15220 ( .B1(n13498), .B2(n14240), .A(n13080), .ZN(n13081) );
  OAI21_X1 U15221 ( .B1(n13082), .B2(n13168), .A(n13081), .ZN(P2_U3191) );
  XNOR2_X1 U15222 ( .A(n13084), .B(n13083), .ZN(n13090) );
  AND2_X1 U15223 ( .A1(n13178), .A2(n13139), .ZN(n13085) );
  AOI21_X1 U15224 ( .B1(n13180), .B2(n13141), .A(n13085), .ZN(n13482) );
  INV_X1 U15225 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13086) );
  OAI22_X1 U15226 ( .A1(n13482), .A2(n13143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13086), .ZN(n13088) );
  NOR2_X1 U15227 ( .A1(n6836), .A2(n13149), .ZN(n13087) );
  AOI211_X1 U15228 ( .C1(n13145), .C2(n13342), .A(n13088), .B(n13087), .ZN(
        n13089) );
  OAI21_X1 U15229 ( .B1(n13090), .B2(n13168), .A(n13089), .ZN(P2_U3195) );
  XNOR2_X1 U15230 ( .A(n13092), .B(n13091), .ZN(n13098) );
  OAI22_X1 U15231 ( .A1(n13094), .A2(n13163), .B1(n13093), .B2(n13161), .ZN(
        n13456) );
  AOI22_X1 U15232 ( .A1(n14237), .A2(n13456), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13095) );
  OAI21_X1 U15233 ( .B1(n13284), .B2(n14243), .A(n13095), .ZN(n13096) );
  AOI21_X1 U15234 ( .B1(n13457), .B2(n14240), .A(n13096), .ZN(n13097) );
  OAI21_X1 U15235 ( .B1(n13098), .B2(n13168), .A(n13097), .ZN(P2_U3197) );
  OAI21_X1 U15236 ( .B1(n13101), .B2(n13100), .A(n13099), .ZN(n13102) );
  NAND2_X1 U15237 ( .A1(n13102), .A2(n14235), .ZN(n13108) );
  INV_X1 U15238 ( .A(n13103), .ZN(n13106) );
  OAI21_X1 U15239 ( .B1(n13143), .B2(n13514), .A(n13104), .ZN(n13105) );
  AOI21_X1 U15240 ( .B1(n13106), .B2(n13145), .A(n13105), .ZN(n13107) );
  OAI211_X1 U15241 ( .C1(n13516), .C2(n13149), .A(n13108), .B(n13107), .ZN(
        P2_U3198) );
  INV_X1 U15242 ( .A(n13400), .ZN(n13509) );
  OAI21_X1 U15243 ( .B1(n13111), .B2(n13110), .A(n13109), .ZN(n13112) );
  NAND2_X1 U15244 ( .A1(n13112), .A2(n14235), .ZN(n13118) );
  INV_X1 U15245 ( .A(n13401), .ZN(n13116) );
  AND2_X1 U15246 ( .A1(n13184), .A2(n13141), .ZN(n13113) );
  AOI21_X1 U15247 ( .B1(n13182), .B2(n13139), .A(n13113), .ZN(n13507) );
  OAI21_X1 U15248 ( .B1(n13507), .B2(n13143), .A(n13114), .ZN(n13115) );
  AOI21_X1 U15249 ( .B1(n13116), .B2(n13145), .A(n13115), .ZN(n13117) );
  OAI211_X1 U15250 ( .C1(n13509), .C2(n13149), .A(n13118), .B(n13117), .ZN(
        P2_U3200) );
  XNOR2_X1 U15251 ( .A(n13119), .B(n13120), .ZN(n13125) );
  OAI22_X1 U15252 ( .A1(n13121), .A2(n13163), .B1(n13164), .B2(n13161), .ZN(
        n13294) );
  AOI22_X1 U15253 ( .A1(n14237), .A2(n13294), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13122) );
  OAI21_X1 U15254 ( .B1(n13298), .B2(n14243), .A(n13122), .ZN(n13123) );
  AOI21_X1 U15255 ( .B1(n13462), .B2(n14240), .A(n13123), .ZN(n13124) );
  OAI21_X1 U15256 ( .B1(n13125), .B2(n13168), .A(n13124), .ZN(P2_U3201) );
  OAI21_X1 U15257 ( .B1(n13128), .B2(n13127), .A(n13126), .ZN(n13129) );
  NAND2_X1 U15258 ( .A1(n13129), .A2(n14235), .ZN(n13134) );
  INV_X1 U15259 ( .A(n13353), .ZN(n13132) );
  AOI22_X1 U15260 ( .A1(n13179), .A2(n13139), .B1(n13141), .B2(n13181), .ZN(
        n13488) );
  INV_X1 U15261 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13130) );
  OAI22_X1 U15262 ( .A1(n13488), .A2(n13143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13130), .ZN(n13131) );
  AOI21_X1 U15263 ( .B1(n13132), .B2(n13145), .A(n13131), .ZN(n13133) );
  OAI211_X1 U15264 ( .C1(n13490), .C2(n13149), .A(n13134), .B(n13133), .ZN(
        P2_U3205) );
  OAI21_X1 U15265 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(n13138) );
  NAND2_X1 U15266 ( .A1(n13138), .A2(n14235), .ZN(n13148) );
  INV_X1 U15267 ( .A(n13326), .ZN(n13146) );
  AND2_X1 U15268 ( .A1(n13177), .A2(n13139), .ZN(n13140) );
  AOI21_X1 U15269 ( .B1(n13179), .B2(n13141), .A(n13140), .ZN(n13475) );
  INV_X1 U15270 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13142) );
  OAI22_X1 U15271 ( .A1(n13475), .A2(n13143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13142), .ZN(n13144) );
  AOI21_X1 U15272 ( .B1(n13146), .B2(n13145), .A(n13144), .ZN(n13147) );
  OAI211_X1 U15273 ( .C1(n13150), .C2(n13149), .A(n13148), .B(n13147), .ZN(
        P2_U3207) );
  XNOR2_X1 U15274 ( .A(n13152), .B(n13151), .ZN(n13158) );
  OAI22_X1 U15275 ( .A1(n13154), .A2(n13161), .B1(n13153), .B2(n13163), .ZN(
        n13377) );
  NAND2_X1 U15276 ( .A1(n13377), .A2(n14237), .ZN(n13155) );
  NAND2_X1 U15277 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14675)
         );
  OAI211_X1 U15278 ( .C1(n14243), .C2(n13380), .A(n13155), .B(n14675), .ZN(
        n13156) );
  AOI21_X1 U15279 ( .B1(n13503), .B2(n14240), .A(n13156), .ZN(n13157) );
  OAI21_X1 U15280 ( .B1(n13158), .B2(n13168), .A(n13157), .ZN(P2_U3210) );
  OAI22_X1 U15281 ( .A1(n13164), .A2(n13163), .B1(n13162), .B2(n13161), .ZN(
        n13270) );
  AOI22_X1 U15282 ( .A1(n14237), .A2(n13270), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13165) );
  OAI21_X1 U15283 ( .B1(n13271), .B2(n14243), .A(n13165), .ZN(n13166) );
  AOI21_X1 U15284 ( .B1(n13274), .B2(n14240), .A(n13166), .ZN(n13167) );
  OAI21_X1 U15285 ( .B1(n13169), .B2(n13168), .A(n13167), .ZN(P2_U3212) );
  MUX2_X1 U15286 ( .A(n13226), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13199), .Z(
        P2_U3562) );
  MUX2_X1 U15287 ( .A(n13170), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13199), .Z(
        P2_U3561) );
  MUX2_X1 U15288 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13171), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15289 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13172), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15290 ( .A(n13173), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13199), .Z(
        P2_U3558) );
  MUX2_X1 U15291 ( .A(n13174), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13199), .Z(
        P2_U3557) );
  MUX2_X1 U15292 ( .A(n13175), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13199), .Z(
        P2_U3556) );
  MUX2_X1 U15293 ( .A(n13176), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13199), .Z(
        P2_U3555) );
  MUX2_X1 U15294 ( .A(n13177), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13199), .Z(
        P2_U3554) );
  MUX2_X1 U15295 ( .A(n13178), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13199), .Z(
        P2_U3553) );
  MUX2_X1 U15296 ( .A(n13179), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13199), .Z(
        P2_U3552) );
  MUX2_X1 U15297 ( .A(n13180), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13199), .Z(
        P2_U3551) );
  MUX2_X1 U15298 ( .A(n13181), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13199), .Z(
        P2_U3550) );
  MUX2_X1 U15299 ( .A(n13182), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13199), .Z(
        P2_U3549) );
  MUX2_X1 U15300 ( .A(n13183), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13199), .Z(
        P2_U3548) );
  MUX2_X1 U15301 ( .A(n13184), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13199), .Z(
        P2_U3547) );
  MUX2_X1 U15302 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13185), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15303 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13186), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U15304 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13187), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U15305 ( .A(n13188), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13199), .Z(
        P2_U3543) );
  MUX2_X1 U15306 ( .A(n13189), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13199), .Z(
        P2_U3542) );
  MUX2_X1 U15307 ( .A(n13190), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13199), .Z(
        P2_U3541) );
  MUX2_X1 U15308 ( .A(n13191), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13199), .Z(
        P2_U3540) );
  MUX2_X1 U15309 ( .A(n13192), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13199), .Z(
        P2_U3539) );
  MUX2_X1 U15310 ( .A(n13193), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13199), .Z(
        P2_U3538) );
  MUX2_X1 U15311 ( .A(n13194), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13199), .Z(
        P2_U3537) );
  MUX2_X1 U15312 ( .A(n13195), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13199), .Z(
        P2_U3536) );
  MUX2_X1 U15313 ( .A(n13196), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13199), .Z(
        P2_U3535) );
  MUX2_X1 U15314 ( .A(n13197), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13199), .Z(
        P2_U3534) );
  MUX2_X1 U15315 ( .A(n13198), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13199), .Z(
        P2_U3533) );
  MUX2_X1 U15316 ( .A(n13200), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13199), .Z(
        P2_U3532) );
  NAND2_X1 U15317 ( .A1(n13201), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U15318 ( .A1(n13203), .A2(n13202), .ZN(n13204) );
  XNOR2_X1 U15319 ( .A(n14674), .B(n13204), .ZN(n14665) );
  NOR2_X1 U15320 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14665), .ZN(n14664) );
  NOR2_X1 U15321 ( .A1(n14674), .A2(n13204), .ZN(n13205) );
  NOR2_X1 U15322 ( .A1(n14664), .A2(n13205), .ZN(n13206) );
  INV_X1 U15323 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13209) );
  OAI21_X1 U15324 ( .B1(n13209), .B2(n13208), .A(n13207), .ZN(n13210) );
  XOR2_X1 U15325 ( .A(n14674), .B(n13210), .Z(n14667) );
  NAND2_X1 U15326 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14667), .ZN(n14666) );
  NAND2_X1 U15327 ( .A1(n14674), .A2(n13210), .ZN(n13211) );
  NAND2_X1 U15328 ( .A1(n14666), .A2(n13211), .ZN(n13212) );
  XOR2_X1 U15329 ( .A(n13212), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13215) );
  NOR2_X1 U15330 ( .A1(n13215), .A2(n14668), .ZN(n13213) );
  AOI211_X1 U15331 ( .C1(n13214), .C2(n14655), .A(n14673), .B(n13213), .ZN(
        n13219) );
  AOI22_X1 U15332 ( .A1(n13216), .A2(n14655), .B1(n14658), .B2(n13215), .ZN(
        n13218) );
  MUX2_X1 U15333 ( .A(n13219), .B(n13218), .S(n13217), .Z(n13222) );
  INV_X1 U15334 ( .A(n13220), .ZN(n13221) );
  OAI211_X1 U15335 ( .C1(n7694), .C2(n14677), .A(n13222), .B(n13221), .ZN(
        P2_U3233) );
  NAND2_X1 U15336 ( .A1(n13231), .A2(n13430), .ZN(n13230) );
  NAND2_X1 U15337 ( .A1(n13226), .A2(n13225), .ZN(n13428) );
  NOR2_X1 U15338 ( .A1(n13402), .A2(n13428), .ZN(n13233) );
  NOR2_X1 U15339 ( .A1(n13223), .A2(n13417), .ZN(n13228) );
  AOI211_X1 U15340 ( .C1(n13402), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13233), 
        .B(n13228), .ZN(n13229) );
  OAI21_X1 U15341 ( .B1(n13427), .B2(n13398), .A(n13229), .ZN(P2_U3234) );
  OAI211_X1 U15342 ( .C1(n13231), .C2(n13430), .A(n6486), .B(n13230), .ZN(
        n13429) );
  NOR2_X1 U15343 ( .A1(n13430), .A2(n13417), .ZN(n13232) );
  AOI211_X1 U15344 ( .C1(n13402), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13233), 
        .B(n13232), .ZN(n13234) );
  OAI21_X1 U15345 ( .B1(n13398), .B2(n13429), .A(n13234), .ZN(P2_U3235) );
  OAI21_X1 U15346 ( .B1(n13236), .B2(n13244), .A(n13235), .ZN(n13439) );
  OR2_X1 U15347 ( .A1(n13240), .A2(n13255), .ZN(n13237) );
  AND3_X1 U15348 ( .A1(n13238), .A2(n13237), .A3(n6486), .ZN(n13435) );
  INV_X1 U15349 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13239) );
  OAI22_X1 U15350 ( .A1(n13240), .A2(n13417), .B1(n13406), .B2(n13239), .ZN(
        n13241) );
  AOI21_X1 U15351 ( .B1(n13435), .B2(n13422), .A(n13241), .ZN(n13250) );
  AOI211_X1 U15352 ( .C1(n13244), .C2(n13243), .A(n13529), .B(n13242), .ZN(
        n13246) );
  NOR2_X1 U15353 ( .A1(n13246), .A2(n13245), .ZN(n13438) );
  OAI21_X1 U15354 ( .B1(n13247), .B2(n13414), .A(n13438), .ZN(n13248) );
  NAND2_X1 U15355 ( .A1(n13248), .A2(n13406), .ZN(n13249) );
  OAI211_X1 U15356 ( .C1(n13439), .C2(n13411), .A(n13250), .B(n13249), .ZN(
        P2_U3237) );
  XNOR2_X1 U15357 ( .A(n13251), .B(n13256), .ZN(n13253) );
  AOI21_X1 U15358 ( .B1(n13253), .B2(n13541), .A(n13252), .ZN(n13445) );
  AND2_X1 U15359 ( .A1(n13442), .A2(n13268), .ZN(n13254) );
  OR3_X1 U15360 ( .A1(n13255), .A2(n13254), .A3(n10230), .ZN(n13444) );
  OR2_X1 U15361 ( .A1(n13257), .A2(n13256), .ZN(n13441) );
  NAND3_X1 U15362 ( .A1(n13441), .A2(n13440), .A3(n13365), .ZN(n13262) );
  OAI22_X1 U15363 ( .A1(n13406), .A2(n13259), .B1(n13258), .B2(n13414), .ZN(
        n13260) );
  AOI21_X1 U15364 ( .B1(n13442), .B2(n13399), .A(n13260), .ZN(n13261) );
  OAI211_X1 U15365 ( .C1(n13444), .C2(n13398), .A(n13262), .B(n13261), .ZN(
        n13263) );
  INV_X1 U15366 ( .A(n13263), .ZN(n13264) );
  OAI21_X1 U15367 ( .B1(n13402), .B2(n13445), .A(n13264), .ZN(P2_U3238) );
  XNOR2_X1 U15368 ( .A(n13265), .B(n13266), .ZN(n13453) );
  XNOR2_X1 U15369 ( .A(n13267), .B(n13266), .ZN(n13451) );
  OAI211_X1 U15370 ( .C1(n13449), .C2(n6516), .A(n6486), .B(n13268), .ZN(
        n13448) );
  NOR2_X1 U15371 ( .A1(n13406), .A2(n13269), .ZN(n13273) );
  INV_X1 U15372 ( .A(n13270), .ZN(n13447) );
  OAI22_X1 U15373 ( .A1(n13447), .A2(n13402), .B1(n13271), .B2(n13414), .ZN(
        n13272) );
  AOI211_X1 U15374 ( .C1(n13274), .C2(n13399), .A(n13273), .B(n13272), .ZN(
        n13275) );
  OAI21_X1 U15375 ( .B1(n13448), .B2(n13398), .A(n13275), .ZN(n13276) );
  AOI21_X1 U15376 ( .B1(n13451), .B2(n13409), .A(n13276), .ZN(n13277) );
  OAI21_X1 U15377 ( .B1(n13453), .B2(n13411), .A(n13277), .ZN(P2_U3239) );
  XOR2_X1 U15378 ( .A(n13280), .B(n13278), .Z(n13460) );
  OAI21_X1 U15379 ( .B1(n13281), .B2(n13280), .A(n13279), .ZN(n13454) );
  NAND2_X1 U15380 ( .A1(n13457), .A2(n13301), .ZN(n13282) );
  NAND2_X1 U15381 ( .A1(n13282), .A2(n6486), .ZN(n13283) );
  NOR2_X1 U15382 ( .A1(n6516), .A2(n13283), .ZN(n13455) );
  NAND2_X1 U15383 ( .A1(n13455), .A2(n13422), .ZN(n13288) );
  INV_X1 U15384 ( .A(n13456), .ZN(n13285) );
  OAI22_X1 U15385 ( .A1(n13285), .A2(n13402), .B1(n13284), .B2(n13414), .ZN(
        n13286) );
  AOI21_X1 U15386 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(n13402), .A(n13286), 
        .ZN(n13287) );
  OAI211_X1 U15387 ( .C1(n13289), .C2(n13417), .A(n13288), .B(n13287), .ZN(
        n13290) );
  AOI21_X1 U15388 ( .B1(n13454), .B2(n13365), .A(n13290), .ZN(n13291) );
  OAI21_X1 U15389 ( .B1(n13460), .B2(n13375), .A(n13291), .ZN(P2_U3240) );
  XNOR2_X1 U15390 ( .A(n13293), .B(n13292), .ZN(n13295) );
  AOI21_X1 U15391 ( .B1(n13295), .B2(n13541), .A(n13294), .ZN(n13464) );
  XNOR2_X1 U15392 ( .A(n13297), .B(n13296), .ZN(n13465) );
  OAI22_X1 U15393 ( .A1(n13406), .A2(n13299), .B1(n13298), .B2(n13414), .ZN(
        n13300) );
  AOI21_X1 U15394 ( .B1(n13462), .B2(n13399), .A(n13300), .ZN(n13304) );
  AOI21_X1 U15395 ( .B1(n13462), .B2(n13310), .A(n10230), .ZN(n13302) );
  AND2_X1 U15396 ( .A1(n13302), .A2(n13301), .ZN(n13461) );
  NAND2_X1 U15397 ( .A1(n13461), .A2(n13422), .ZN(n13303) );
  OAI211_X1 U15398 ( .C1(n13465), .C2(n13411), .A(n13304), .B(n13303), .ZN(
        n13305) );
  INV_X1 U15399 ( .A(n13305), .ZN(n13306) );
  OAI21_X1 U15400 ( .B1(n13402), .B2(n13464), .A(n13306), .ZN(P2_U3241) );
  XNOR2_X1 U15401 ( .A(n13307), .B(n13314), .ZN(n13466) );
  INV_X1 U15402 ( .A(n13466), .ZN(n13320) );
  OAI22_X1 U15403 ( .A1(n13406), .A2(n13309), .B1(n13308), .B2(n13414), .ZN(
        n13313) );
  OAI211_X1 U15404 ( .C1(n13325), .C2(n13311), .A(n6486), .B(n13310), .ZN(
        n13469) );
  NOR2_X1 U15405 ( .A1(n13469), .A2(n13398), .ZN(n13312) );
  AOI211_X1 U15406 ( .C1(n13399), .C2(n13468), .A(n13313), .B(n13312), .ZN(
        n13319) );
  XNOR2_X1 U15407 ( .A(n13315), .B(n13314), .ZN(n13316) );
  NAND2_X1 U15408 ( .A1(n13316), .A2(n13541), .ZN(n13470) );
  INV_X1 U15409 ( .A(n13470), .ZN(n13317) );
  OAI21_X1 U15410 ( .B1(n13317), .B2(n13467), .A(n13406), .ZN(n13318) );
  OAI211_X1 U15411 ( .C1(n13320), .C2(n13411), .A(n13319), .B(n13318), .ZN(
        P2_U3242) );
  XNOR2_X1 U15412 ( .A(n13322), .B(n13321), .ZN(n13481) );
  NAND2_X1 U15413 ( .A1(n13341), .A2(n13474), .ZN(n13323) );
  NAND2_X1 U15414 ( .A1(n13323), .A2(n6486), .ZN(n13324) );
  NOR2_X1 U15415 ( .A1(n13325), .A2(n13324), .ZN(n13478) );
  NAND2_X1 U15416 ( .A1(n13474), .A2(n13399), .ZN(n13329) );
  OAI22_X1 U15417 ( .A1(n13475), .A2(n13402), .B1(n13326), .B2(n13414), .ZN(
        n13327) );
  INV_X1 U15418 ( .A(n13327), .ZN(n13328) );
  OAI211_X1 U15419 ( .C1(n13406), .C2(n13330), .A(n13329), .B(n13328), .ZN(
        n13335) );
  OAI21_X1 U15420 ( .B1(n13333), .B2(n13332), .A(n13331), .ZN(n13473) );
  NOR2_X1 U15421 ( .A1(n13473), .A2(n13411), .ZN(n13334) );
  AOI211_X1 U15422 ( .C1(n13478), .C2(n13422), .A(n13335), .B(n13334), .ZN(
        n13336) );
  OAI21_X1 U15423 ( .B1(n13375), .B2(n13481), .A(n13336), .ZN(P2_U3243) );
  XNOR2_X1 U15424 ( .A(n13337), .B(n13338), .ZN(n13487) );
  XNOR2_X1 U15425 ( .A(n13339), .B(n13338), .ZN(n13485) );
  NAND2_X1 U15426 ( .A1(n13346), .A2(n13352), .ZN(n13340) );
  NAND3_X1 U15427 ( .A1(n13341), .A2(n6486), .A3(n13340), .ZN(n13483) );
  NAND2_X1 U15428 ( .A1(n13342), .A2(n13381), .ZN(n13344) );
  NAND2_X1 U15429 ( .A1(n13402), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13343) );
  OAI211_X1 U15430 ( .C1(n13482), .C2(n13402), .A(n13344), .B(n13343), .ZN(
        n13345) );
  AOI21_X1 U15431 ( .B1(n13346), .B2(n13399), .A(n13345), .ZN(n13347) );
  OAI21_X1 U15432 ( .B1(n13483), .B2(n13398), .A(n13347), .ZN(n13348) );
  AOI21_X1 U15433 ( .B1(n13485), .B2(n13365), .A(n13348), .ZN(n13349) );
  OAI21_X1 U15434 ( .B1(n13487), .B2(n13375), .A(n13349), .ZN(P2_U3244) );
  XNOR2_X1 U15435 ( .A(n13350), .B(n13358), .ZN(n13494) );
  INV_X1 U15436 ( .A(n13351), .ZN(n13366) );
  OAI211_X1 U15437 ( .C1(n13490), .C2(n13366), .A(n6486), .B(n13352), .ZN(
        n13489) );
  INV_X1 U15438 ( .A(n13489), .ZN(n13357) );
  OAI22_X1 U15439 ( .A1(n13488), .A2(n13402), .B1(n13353), .B2(n13414), .ZN(
        n13354) );
  AOI21_X1 U15440 ( .B1(P2_REG2_REG_20__SCAN_IN), .B2(n13402), .A(n13354), 
        .ZN(n13355) );
  OAI21_X1 U15441 ( .B1(n13490), .B2(n13417), .A(n13355), .ZN(n13356) );
  AOI21_X1 U15442 ( .B1(n13357), .B2(n13422), .A(n13356), .ZN(n13361) );
  XNOR2_X1 U15443 ( .A(n13359), .B(n13358), .ZN(n13492) );
  NAND2_X1 U15444 ( .A1(n13492), .A2(n13409), .ZN(n13360) );
  OAI211_X1 U15445 ( .C1(n13494), .C2(n13411), .A(n13361), .B(n13360), .ZN(
        P2_U3245) );
  XOR2_X1 U15446 ( .A(n13362), .B(n13363), .Z(n13501) );
  XNOR2_X1 U15447 ( .A(n13364), .B(n13363), .ZN(n13495) );
  NAND2_X1 U15448 ( .A1(n13495), .A2(n13365), .ZN(n13374) );
  AOI211_X1 U15449 ( .C1(n13498), .C2(n13379), .A(n10230), .B(n13366), .ZN(
        n13496) );
  INV_X1 U15450 ( .A(n13497), .ZN(n13368) );
  OAI22_X1 U15451 ( .A1(n13368), .A2(n13402), .B1(n13367), .B2(n13414), .ZN(
        n13369) );
  AOI21_X1 U15452 ( .B1(P2_REG2_REG_19__SCAN_IN), .B2(n13402), .A(n13369), 
        .ZN(n13370) );
  OAI21_X1 U15453 ( .B1(n13371), .B2(n13417), .A(n13370), .ZN(n13372) );
  AOI21_X1 U15454 ( .B1(n13496), .B2(n13422), .A(n13372), .ZN(n13373) );
  OAI211_X1 U15455 ( .C1(n13501), .C2(n13375), .A(n13374), .B(n13373), .ZN(
        P2_U3246) );
  XOR2_X1 U15456 ( .A(n13376), .B(n13387), .Z(n13378) );
  AOI21_X1 U15457 ( .B1(n13378), .B2(n13541), .A(n13377), .ZN(n13505) );
  AOI211_X1 U15458 ( .C1(n13503), .C2(n13396), .A(n10230), .B(n6838), .ZN(
        n13502) );
  INV_X1 U15459 ( .A(n13380), .ZN(n13382) );
  AOI22_X1 U15460 ( .A1(n13402), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13382), 
        .B2(n13381), .ZN(n13383) );
  OAI21_X1 U15461 ( .B1(n13384), .B2(n13417), .A(n13383), .ZN(n13389) );
  AOI21_X1 U15462 ( .B1(n13387), .B2(n13386), .A(n13385), .ZN(n13506) );
  NOR2_X1 U15463 ( .A1(n13506), .A2(n13411), .ZN(n13388) );
  AOI211_X1 U15464 ( .C1(n13502), .C2(n13422), .A(n13389), .B(n13388), .ZN(
        n13390) );
  OAI21_X1 U15465 ( .B1(n13402), .B2(n13505), .A(n13390), .ZN(P2_U3247) );
  OAI21_X1 U15466 ( .B1(n13392), .B2(n13393), .A(n13391), .ZN(n13513) );
  XNOR2_X1 U15467 ( .A(n13394), .B(n13393), .ZN(n13511) );
  AOI21_X1 U15468 ( .B1(n13395), .B2(n13400), .A(n10230), .ZN(n13397) );
  NAND2_X1 U15469 ( .A1(n13397), .A2(n13396), .ZN(n13508) );
  NOR2_X1 U15470 ( .A1(n13508), .A2(n13398), .ZN(n13408) );
  NAND2_X1 U15471 ( .A1(n13400), .A2(n13399), .ZN(n13405) );
  OAI22_X1 U15472 ( .A1(n13507), .A2(n13402), .B1(n13401), .B2(n13414), .ZN(
        n13403) );
  INV_X1 U15473 ( .A(n13403), .ZN(n13404) );
  OAI211_X1 U15474 ( .C1(n13406), .C2(n11322), .A(n13405), .B(n13404), .ZN(
        n13407) );
  AOI211_X1 U15475 ( .C1(n13511), .C2(n13409), .A(n13408), .B(n13407), .ZN(
        n13410) );
  OAI21_X1 U15476 ( .B1(n13513), .B2(n13411), .A(n13410), .ZN(P2_U3248) );
  MUX2_X1 U15477 ( .A(n13413), .B(n13412), .S(n13402), .Z(n13426) );
  OAI22_X1 U15478 ( .A1(n13417), .A2(n13416), .B1(n13415), .B2(n13414), .ZN(
        n13418) );
  INV_X1 U15479 ( .A(n13418), .ZN(n13425) );
  NAND2_X1 U15480 ( .A1(n13420), .A2(n13419), .ZN(n13424) );
  NAND2_X1 U15481 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  NAND4_X1 U15482 ( .A1(n13426), .A2(n13425), .A3(n13424), .A4(n13423), .ZN(
        P2_U3264) );
  OAI211_X1 U15483 ( .C1(n13223), .C2(n14749), .A(n13427), .B(n13428), .ZN(
        n13546) );
  MUX2_X1 U15484 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13546), .S(n14768), .Z(
        P2_U3530) );
  OAI211_X1 U15485 ( .C1(n13430), .C2(n14749), .A(n13429), .B(n13428), .ZN(
        n13547) );
  MUX2_X1 U15486 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13547), .S(n14768), .Z(
        P2_U3529) );
  MUX2_X1 U15487 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13548), .S(n14768), .Z(
        P2_U3528) );
  AOI21_X1 U15488 ( .B1(n14735), .B2(n13436), .A(n13435), .ZN(n13437) );
  OAI211_X1 U15489 ( .C1(n13439), .C2(n14718), .A(n13438), .B(n13437), .ZN(
        n13549) );
  MUX2_X1 U15490 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13549), .S(n14768), .Z(
        P2_U3527) );
  NAND3_X1 U15491 ( .A1(n13441), .A2(n13440), .A3(n13525), .ZN(n13446) );
  NAND2_X1 U15492 ( .A1(n13442), .A2(n14735), .ZN(n13443) );
  NAND4_X1 U15493 ( .A1(n13446), .A2(n13445), .A3(n13444), .A4(n13443), .ZN(
        n13550) );
  MUX2_X1 U15494 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13550), .S(n14768), .Z(
        P2_U3526) );
  OAI211_X1 U15495 ( .C1(n13449), .C2(n14749), .A(n13448), .B(n13447), .ZN(
        n13450) );
  AOI21_X1 U15496 ( .B1(n13451), .B2(n13541), .A(n13450), .ZN(n13452) );
  OAI21_X1 U15497 ( .B1(n13453), .B2(n14718), .A(n13452), .ZN(n13551) );
  MUX2_X1 U15498 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13551), .S(n14768), .Z(
        P2_U3525) );
  NAND2_X1 U15499 ( .A1(n13454), .A2(n13525), .ZN(n13459) );
  AOI211_X1 U15500 ( .C1(n14735), .C2(n13457), .A(n13456), .B(n13455), .ZN(
        n13458) );
  OAI211_X1 U15501 ( .C1(n13529), .C2(n13460), .A(n13459), .B(n13458), .ZN(
        n13552) );
  MUX2_X1 U15502 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13552), .S(n14768), .Z(
        P2_U3524) );
  AOI21_X1 U15503 ( .B1(n14735), .B2(n13462), .A(n13461), .ZN(n13463) );
  OAI211_X1 U15504 ( .C1(n13465), .C2(n14718), .A(n13464), .B(n13463), .ZN(
        n13553) );
  MUX2_X1 U15505 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13553), .S(n14768), .Z(
        P2_U3523) );
  NAND2_X1 U15506 ( .A1(n13466), .A2(n13525), .ZN(n13472) );
  AOI21_X1 U15507 ( .B1(n13468), .B2(n14735), .A(n13467), .ZN(n13471) );
  NAND4_X1 U15508 ( .A1(n13472), .A2(n13471), .A3(n13470), .A4(n13469), .ZN(
        n13554) );
  MUX2_X1 U15509 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13554), .S(n14768), .Z(
        P2_U3522) );
  INV_X1 U15510 ( .A(n13473), .ZN(n13479) );
  NAND2_X1 U15511 ( .A1(n13474), .A2(n14735), .ZN(n13476) );
  NAND2_X1 U15512 ( .A1(n13476), .A2(n13475), .ZN(n13477) );
  AOI211_X1 U15513 ( .C1(n13479), .C2(n13525), .A(n13478), .B(n13477), .ZN(
        n13480) );
  OAI21_X1 U15514 ( .B1(n13529), .B2(n13481), .A(n13480), .ZN(n13555) );
  MUX2_X1 U15515 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13555), .S(n14768), .Z(
        P2_U3521) );
  OAI211_X1 U15516 ( .C1(n6836), .C2(n14749), .A(n13483), .B(n13482), .ZN(
        n13484) );
  AOI21_X1 U15517 ( .B1(n13485), .B2(n13525), .A(n13484), .ZN(n13486) );
  OAI21_X1 U15518 ( .B1(n13529), .B2(n13487), .A(n13486), .ZN(n13556) );
  MUX2_X1 U15519 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13556), .S(n14768), .Z(
        P2_U3520) );
  OAI211_X1 U15520 ( .C1(n13490), .C2(n14749), .A(n13489), .B(n13488), .ZN(
        n13491) );
  AOI21_X1 U15521 ( .B1(n13492), .B2(n13541), .A(n13491), .ZN(n13493) );
  OAI21_X1 U15522 ( .B1(n13494), .B2(n14718), .A(n13493), .ZN(n13557) );
  MUX2_X1 U15523 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13557), .S(n14768), .Z(
        P2_U3519) );
  NAND2_X1 U15524 ( .A1(n13495), .A2(n13525), .ZN(n13500) );
  AOI211_X1 U15525 ( .C1(n14735), .C2(n13498), .A(n13497), .B(n13496), .ZN(
        n13499) );
  OAI211_X1 U15526 ( .C1(n13529), .C2(n13501), .A(n13500), .B(n13499), .ZN(
        n13558) );
  MUX2_X1 U15527 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13558), .S(n14768), .Z(
        P2_U3518) );
  AOI21_X1 U15528 ( .B1(n14735), .B2(n13503), .A(n13502), .ZN(n13504) );
  OAI211_X1 U15529 ( .C1(n13506), .C2(n14718), .A(n13505), .B(n13504), .ZN(
        n13559) );
  MUX2_X1 U15530 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13559), .S(n14768), .Z(
        P2_U3517) );
  OAI211_X1 U15531 ( .C1(n13509), .C2(n14749), .A(n13508), .B(n13507), .ZN(
        n13510) );
  AOI21_X1 U15532 ( .B1(n13511), .B2(n13541), .A(n13510), .ZN(n13512) );
  OAI21_X1 U15533 ( .B1(n13513), .B2(n14718), .A(n13512), .ZN(n13560) );
  MUX2_X1 U15534 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13560), .S(n14768), .Z(
        P2_U3516) );
  OAI211_X1 U15535 ( .C1(n13516), .C2(n14749), .A(n13515), .B(n13514), .ZN(
        n13517) );
  AOI21_X1 U15536 ( .B1(n13518), .B2(n13541), .A(n13517), .ZN(n13519) );
  OAI21_X1 U15537 ( .B1(n13520), .B2(n14718), .A(n13519), .ZN(n13561) );
  MUX2_X1 U15538 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13561), .S(n14768), .Z(
        P2_U3515) );
  OAI211_X1 U15539 ( .C1(n13523), .C2(n14749), .A(n13522), .B(n13521), .ZN(
        n13524) );
  AOI21_X1 U15540 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13527) );
  OAI21_X1 U15541 ( .B1(n13529), .B2(n13528), .A(n13527), .ZN(n13562) );
  MUX2_X1 U15542 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13562), .S(n14768), .Z(
        P2_U3514) );
  OAI211_X1 U15543 ( .C1(n13532), .C2(n14749), .A(n13531), .B(n13530), .ZN(
        n13533) );
  AOI21_X1 U15544 ( .B1(n13534), .B2(n13541), .A(n13533), .ZN(n13535) );
  OAI21_X1 U15545 ( .B1(n13536), .B2(n14718), .A(n13535), .ZN(n13563) );
  MUX2_X1 U15546 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13563), .S(n14768), .Z(
        P2_U3513) );
  OAI211_X1 U15547 ( .C1(n13539), .C2(n14749), .A(n13538), .B(n13537), .ZN(
        n13540) );
  AOI21_X1 U15548 ( .B1(n13542), .B2(n13541), .A(n13540), .ZN(n13543) );
  OAI21_X1 U15549 ( .B1(n13544), .B2(n14718), .A(n13543), .ZN(n13564) );
  MUX2_X1 U15550 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13564), .S(n14768), .Z(
        P2_U3512) );
  MUX2_X1 U15551 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n13545), .S(n14768), .Z(
        P2_U3500) );
  MUX2_X1 U15552 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13546), .S(n14756), .Z(
        P2_U3498) );
  MUX2_X1 U15553 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13547), .S(n14756), .Z(
        P2_U3497) );
  MUX2_X1 U15554 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13549), .S(n14756), .Z(
        P2_U3495) );
  MUX2_X1 U15555 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13550), .S(n14756), .Z(
        P2_U3494) );
  MUX2_X1 U15556 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13551), .S(n14756), .Z(
        P2_U3493) );
  MUX2_X1 U15557 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13552), .S(n14756), .Z(
        P2_U3492) );
  MUX2_X1 U15558 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13553), .S(n14756), .Z(
        P2_U3491) );
  MUX2_X1 U15559 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13554), .S(n14756), .Z(
        P2_U3490) );
  MUX2_X1 U15560 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13555), .S(n14756), .Z(
        P2_U3489) );
  MUX2_X1 U15561 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13556), .S(n14756), .Z(
        P2_U3488) );
  MUX2_X1 U15562 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13557), .S(n14756), .Z(
        P2_U3487) );
  MUX2_X1 U15563 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13558), .S(n14756), .Z(
        P2_U3486) );
  MUX2_X1 U15564 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13559), .S(n14756), .Z(
        P2_U3484) );
  MUX2_X1 U15565 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13560), .S(n14756), .Z(
        P2_U3481) );
  MUX2_X1 U15566 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13561), .S(n14756), .Z(
        P2_U3478) );
  MUX2_X1 U15567 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13562), .S(n14756), .Z(
        P2_U3475) );
  MUX2_X1 U15568 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13563), .S(n14756), .Z(
        P2_U3472) );
  MUX2_X1 U15569 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13564), .S(n14756), .Z(
        P2_U3469) );
  INV_X1 U15570 ( .A(n13565), .ZN(n14116) );
  NOR4_X1 U15571 ( .A1(n13566), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8728), .A4(
        P2_U3088), .ZN(n13567) );
  AOI21_X1 U15572 ( .B1(n13572), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13567), 
        .ZN(n13568) );
  OAI21_X1 U15573 ( .B1(n14116), .B2(n13581), .A(n13568), .ZN(P2_U3296) );
  INV_X1 U15574 ( .A(n13569), .ZN(n14121) );
  OAI222_X1 U15575 ( .A1(n13581), .A2(n14121), .B1(P2_U3088), .B2(n8455), .C1(
        n13570), .C2(n13578), .ZN(P2_U3298) );
  AOI21_X1 U15576 ( .B1(n13572), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13571), 
        .ZN(n13573) );
  OAI21_X1 U15577 ( .B1(n13574), .B2(n13581), .A(n13573), .ZN(P2_U3299) );
  INV_X1 U15578 ( .A(n13575), .ZN(n14123) );
  OAI222_X1 U15579 ( .A1(n13578), .A2(n13577), .B1(P2_U3088), .B2(n13576), 
        .C1(n13581), .C2(n14123), .ZN(P2_U3300) );
  INV_X1 U15580 ( .A(n13579), .ZN(n14127) );
  OAI222_X1 U15581 ( .A1(P2_U3088), .A2(n13582), .B1(n13581), .B2(n14127), 
        .C1(n13580), .C2(n13578), .ZN(P2_U3301) );
  MUX2_X1 U15582 ( .A(n13583), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15583 ( .A(n13585), .B(n13584), .Z(n13591) );
  AOI22_X1 U15584 ( .A1(n14364), .A2(n13586), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13587) );
  OAI21_X1 U15585 ( .B1(n14367), .B2(n13588), .A(n13587), .ZN(n13589) );
  AOI21_X1 U15586 ( .B1(n14033), .B2(n14297), .A(n13589), .ZN(n13590) );
  OAI21_X1 U15587 ( .B1(n13591), .B2(n13663), .A(n13590), .ZN(P1_U3214) );
  XOR2_X1 U15588 ( .A(n13593), .B(n13592), .Z(n13599) );
  NAND2_X1 U15589 ( .A1(n13670), .A2(n14353), .ZN(n13595) );
  NAND2_X1 U15590 ( .A1(n13668), .A2(n14003), .ZN(n13594) );
  NAND2_X1 U15591 ( .A1(n13595), .A2(n13594), .ZN(n14057) );
  AOI22_X1 U15592 ( .A1(n14364), .A2(n14057), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13596) );
  OAI21_X1 U15593 ( .B1(n14367), .B2(n13935), .A(n13596), .ZN(n13597) );
  AOI21_X1 U15594 ( .B1(n14058), .B2(n14297), .A(n13597), .ZN(n13598) );
  OAI21_X1 U15595 ( .B1(n13599), .B2(n13663), .A(n13598), .ZN(P1_U3216) );
  NAND2_X1 U15596 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13815)
         );
  OAI22_X1 U15597 ( .A1(n13614), .A2(n14356), .B1(n13600), .B2(n13658), .ZN(
        n14084) );
  NAND2_X1 U15598 ( .A1(n14084), .A2(n14364), .ZN(n13601) );
  OAI211_X1 U15599 ( .C1(n14367), .C2(n13986), .A(n13815), .B(n13601), .ZN(
        n13607) );
  INV_X1 U15600 ( .A(n13602), .ZN(n13603) );
  AOI211_X1 U15601 ( .C1(n13605), .C2(n13604), .A(n13663), .B(n13603), .ZN(
        n13606) );
  AOI211_X1 U15602 ( .C1(n14297), .C2(n14085), .A(n13607), .B(n13606), .ZN(
        n13608) );
  INV_X1 U15603 ( .A(n13608), .ZN(P1_U3219) );
  INV_X1 U15604 ( .A(n13609), .ZN(n13610) );
  AOI21_X1 U15605 ( .B1(n13612), .B2(n13611), .A(n13610), .ZN(n13618) );
  OAI22_X1 U15606 ( .A1(n13614), .A2(n13658), .B1(n13613), .B2(n14356), .ZN(
        n14070) );
  AOI22_X1 U15607 ( .A1(n14070), .A2(n14364), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13615) );
  OAI21_X1 U15608 ( .B1(n14367), .B2(n13958), .A(n13615), .ZN(n13616) );
  AOI21_X1 U15609 ( .B1(n14071), .B2(n14297), .A(n13616), .ZN(n13617) );
  OAI21_X1 U15610 ( .B1(n13618), .B2(n13663), .A(n13617), .ZN(P1_U3223) );
  XOR2_X1 U15611 ( .A(n13620), .B(n13619), .Z(n13626) );
  OAI22_X1 U15612 ( .A1(n13622), .A2(n13658), .B1(n13621), .B2(n14356), .ZN(
        n14044) );
  AOI22_X1 U15613 ( .A1(n14364), .A2(n14044), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13623) );
  OAI21_X1 U15614 ( .B1(n14367), .B2(n13895), .A(n13623), .ZN(n13624) );
  AOI21_X1 U15615 ( .B1(n14045), .B2(n14297), .A(n13624), .ZN(n13625) );
  OAI21_X1 U15616 ( .B1(n13626), .B2(n13663), .A(n13625), .ZN(P1_U3225) );
  XOR2_X1 U15617 ( .A(n13628), .B(n13627), .Z(n13634) );
  NAND2_X1 U15618 ( .A1(n13669), .A2(n14353), .ZN(n13630) );
  NAND2_X1 U15619 ( .A1(n13667), .A2(n14003), .ZN(n13629) );
  NAND2_X1 U15620 ( .A1(n13630), .A2(n13629), .ZN(n13908) );
  AOI22_X1 U15621 ( .A1(n14364), .A2(n13908), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13631) );
  OAI21_X1 U15622 ( .B1(n14367), .B2(n13913), .A(n13631), .ZN(n13632) );
  AOI21_X1 U15623 ( .B1(n13920), .B2(n14297), .A(n13632), .ZN(n13633) );
  OAI21_X1 U15624 ( .B1(n13634), .B2(n13663), .A(n13633), .ZN(P1_U3229) );
  OAI211_X1 U15625 ( .C1(n13637), .C2(n13636), .A(n13635), .B(n14359), .ZN(
        n13643) );
  INV_X1 U15626 ( .A(n13974), .ZN(n13641) );
  AND2_X1 U15627 ( .A1(n13671), .A2(n14003), .ZN(n13638) );
  AOI21_X1 U15628 ( .B1(n14004), .B2(n14353), .A(n13638), .ZN(n14076) );
  OAI22_X1 U15629 ( .A1(n14284), .A2(n14076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13639), .ZN(n13640) );
  AOI21_X1 U15630 ( .B1(n13653), .B2(n13641), .A(n13640), .ZN(n13642) );
  OAI211_X1 U15631 ( .C1(n14077), .C2(n14286), .A(n13643), .B(n13642), .ZN(
        P1_U3233) );
  OAI21_X1 U15632 ( .B1(n13646), .B2(n13645), .A(n13644), .ZN(n13647) );
  NAND2_X1 U15633 ( .A1(n13647), .A2(n14359), .ZN(n13655) );
  INV_X1 U15634 ( .A(n13948), .ZN(n13652) );
  NAND2_X1 U15635 ( .A1(n13671), .A2(n14353), .ZN(n13649) );
  NAND2_X1 U15636 ( .A1(n13669), .A2(n14003), .ZN(n13648) );
  AND2_X1 U15637 ( .A1(n13649), .A2(n13648), .ZN(n14062) );
  INV_X1 U15638 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13650) );
  OAI22_X1 U15639 ( .A1(n14284), .A2(n14062), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13650), .ZN(n13651) );
  AOI21_X1 U15640 ( .B1(n13653), .B2(n13652), .A(n13651), .ZN(n13654) );
  OAI211_X1 U15641 ( .C1(n14286), .C2(n14063), .A(n13655), .B(n13654), .ZN(
        P1_U3235) );
  XOR2_X1 U15642 ( .A(n13657), .B(n13656), .Z(n13664) );
  OAI22_X1 U15643 ( .A1(n13659), .A2(n13658), .B1(n13830), .B2(n14356), .ZN(
        n14038) );
  AOI22_X1 U15644 ( .A1(n14364), .A2(n14038), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13660) );
  OAI21_X1 U15645 ( .B1(n14367), .B2(n13875), .A(n13660), .ZN(n13661) );
  AOI21_X1 U15646 ( .B1(n14039), .B2(n14297), .A(n13661), .ZN(n13662) );
  OAI21_X1 U15647 ( .B1(n13664), .B2(n13663), .A(n13662), .ZN(P1_U3240) );
  MUX2_X1 U15648 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13821), .S(n13689), .Z(
        P1_U3591) );
  MUX2_X1 U15649 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13842), .S(n13689), .Z(
        P1_U3590) );
  MUX2_X1 U15650 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13665), .S(n13689), .Z(
        P1_U3589) );
  MUX2_X1 U15651 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13846), .S(n13689), .Z(
        P1_U3588) );
  MUX2_X1 U15652 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13834), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15653 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13666), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15654 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13667), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15655 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13668), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15656 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13669), .S(n13689), .Z(
        P1_U3583) );
  MUX2_X1 U15657 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13670), .S(n13689), .Z(
        P1_U3582) );
  MUX2_X1 U15658 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13671), .S(n13689), .Z(
        P1_U3581) );
  MUX2_X1 U15659 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13672), .S(n13689), .Z(
        P1_U3580) );
  MUX2_X1 U15660 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14004), .S(n13689), .Z(
        P1_U3579) );
  MUX2_X1 U15661 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13673), .S(n13689), .Z(
        P1_U3578) );
  MUX2_X1 U15662 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14002), .S(n13689), .Z(
        P1_U3577) );
  MUX2_X1 U15663 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13674), .S(n13689), .Z(
        P1_U3576) );
  MUX2_X1 U15664 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13675), .S(n13689), .Z(
        P1_U3575) );
  MUX2_X1 U15665 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13676), .S(n13689), .Z(
        P1_U3574) );
  MUX2_X1 U15666 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13677), .S(n13689), .Z(
        P1_U3573) );
  MUX2_X1 U15667 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13678), .S(n13689), .Z(
        P1_U3572) );
  MUX2_X1 U15668 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13679), .S(n13689), .Z(
        P1_U3571) );
  MUX2_X1 U15669 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13680), .S(n13689), .Z(
        P1_U3570) );
  MUX2_X1 U15670 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13681), .S(n13689), .Z(
        P1_U3569) );
  MUX2_X1 U15671 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13682), .S(n13689), .Z(
        P1_U3568) );
  MUX2_X1 U15672 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13683), .S(n13689), .Z(
        P1_U3567) );
  MUX2_X1 U15673 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13684), .S(n13689), .Z(
        P1_U3566) );
  MUX2_X1 U15674 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13685), .S(n13689), .Z(
        P1_U3565) );
  MUX2_X1 U15675 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13686), .S(n13689), .Z(
        P1_U3564) );
  MUX2_X1 U15676 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13687), .S(n13689), .Z(
        P1_U3563) );
  MUX2_X1 U15677 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14354), .S(n13689), .Z(
        P1_U3562) );
  MUX2_X1 U15678 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13688), .S(n13689), .Z(
        P1_U3561) );
  MUX2_X1 U15679 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13690), .S(n13689), .Z(
        P1_U3560) );
  OAI22_X1 U15680 ( .A1(n14384), .A2(n6941), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13691), .ZN(n13692) );
  AOI21_X1 U15681 ( .B1(n13693), .B2(n13718), .A(n13692), .ZN(n13702) );
  OAI211_X1 U15682 ( .C1(n9925), .C2(n13696), .A(n13811), .B(n13695), .ZN(
        n13701) );
  OAI211_X1 U15683 ( .C1(n13699), .C2(n13698), .A(n14375), .B(n13697), .ZN(
        n13700) );
  NAND3_X1 U15684 ( .A1(n13702), .A2(n13701), .A3(n13700), .ZN(P1_U3244) );
  MUX2_X1 U15685 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n13703), .S(n13711), .Z(
        n13706) );
  INV_X1 U15686 ( .A(n13704), .ZN(n13705) );
  OAI211_X1 U15687 ( .C1(n13706), .C2(n13705), .A(n13811), .B(n13726), .ZN(
        n13715) );
  OAI211_X1 U15688 ( .C1(n13709), .C2(n13708), .A(n14375), .B(n13707), .ZN(
        n13714) );
  AND2_X1 U15689 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13710) );
  AOI21_X1 U15690 ( .B1(n13787), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13710), .ZN(
        n13713) );
  NAND2_X1 U15691 ( .A1(n13718), .A2(n13711), .ZN(n13712) );
  NAND4_X1 U15692 ( .A1(n13715), .A2(n13714), .A3(n13713), .A4(n13712), .ZN(
        P1_U3246) );
  OAI21_X1 U15693 ( .B1(n14384), .B2(n6939), .A(n13716), .ZN(n13717) );
  AOI21_X1 U15694 ( .B1(n13719), .B2(n13718), .A(n13717), .ZN(n13731) );
  OAI211_X1 U15695 ( .C1(n13722), .C2(n13721), .A(n14375), .B(n13720), .ZN(
        n13730) );
  INV_X1 U15696 ( .A(n13723), .ZN(n13728) );
  NAND3_X1 U15697 ( .A1(n13726), .A2(n13725), .A3(n13724), .ZN(n13727) );
  NAND3_X1 U15698 ( .A1(n13811), .A2(n13728), .A3(n13727), .ZN(n13729) );
  NAND4_X1 U15699 ( .A1(n13732), .A2(n13731), .A3(n13730), .A4(n13729), .ZN(
        P1_U3247) );
  NOR2_X1 U15700 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13733), .ZN(n13736) );
  NOR2_X1 U15701 ( .A1(n14380), .A2(n13734), .ZN(n13735) );
  AOI211_X1 U15702 ( .C1(n13787), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13736), .B(
        n13735), .ZN(n13747) );
  INV_X1 U15703 ( .A(n13756), .ZN(n13741) );
  NAND3_X1 U15704 ( .A1(n13739), .A2(n13738), .A3(n13737), .ZN(n13740) );
  NAND3_X1 U15705 ( .A1(n13811), .A2(n13741), .A3(n13740), .ZN(n13746) );
  OAI211_X1 U15706 ( .C1(n13744), .C2(n13743), .A(n14375), .B(n13742), .ZN(
        n13745) );
  NAND3_X1 U15707 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(P1_U3249) );
  NOR2_X1 U15708 ( .A1(n14380), .A2(n13748), .ZN(n13749) );
  AOI211_X1 U15709 ( .C1(n13787), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n13750), .B(
        n13749), .ZN(n13761) );
  OAI211_X1 U15710 ( .C1(n13753), .C2(n13752), .A(n14375), .B(n13751), .ZN(
        n13760) );
  OR3_X1 U15711 ( .A1(n13756), .A2(n13755), .A3(n13754), .ZN(n13757) );
  NAND3_X1 U15712 ( .A1(n13811), .A2(n13758), .A3(n13757), .ZN(n13759) );
  NAND3_X1 U15713 ( .A1(n13761), .A2(n13760), .A3(n13759), .ZN(P1_U3250) );
  AOI21_X1 U15714 ( .B1(n13763), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13762), 
        .ZN(n13769) );
  INV_X1 U15715 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13764) );
  OR2_X1 U15716 ( .A1(n13789), .A2(n13764), .ZN(n13766) );
  NAND2_X1 U15717 ( .A1(n13789), .A2(n13764), .ZN(n13765) );
  AND2_X1 U15718 ( .A1(n13766), .A2(n13765), .ZN(n13768) );
  NOR2_X1 U15719 ( .A1(n13769), .A2(n13768), .ZN(n13788) );
  AOI211_X1 U15720 ( .C1(n13769), .C2(n13768), .A(n13788), .B(n13767), .ZN(
        n13770) );
  INV_X1 U15721 ( .A(n13770), .ZN(n13781) );
  NAND2_X1 U15722 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14270)
         );
  INV_X1 U15723 ( .A(n14270), .ZN(n13773) );
  NOR2_X1 U15724 ( .A1(n14380), .A2(n13771), .ZN(n13772) );
  AOI211_X1 U15725 ( .C1(n13787), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13773), 
        .B(n13772), .ZN(n13780) );
  OR2_X1 U15726 ( .A1(n13789), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13774) );
  NAND2_X1 U15727 ( .A1(n13789), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13783) );
  AND2_X1 U15728 ( .A1(n13774), .A2(n13783), .ZN(n13778) );
  OAI21_X1 U15729 ( .B1(n13776), .B2(n10963), .A(n13775), .ZN(n13777) );
  NAND2_X1 U15730 ( .A1(n13778), .A2(n13777), .ZN(n13782) );
  OAI211_X1 U15731 ( .C1(n13778), .C2(n13777), .A(n13811), .B(n13782), .ZN(
        n13779) );
  NAND3_X1 U15732 ( .A1(n13781), .A2(n13780), .A3(n13779), .ZN(P1_U3260) );
  NAND2_X1 U15733 ( .A1(n13783), .A2(n13782), .ZN(n13803) );
  XNOR2_X1 U15734 ( .A(n13803), .B(n13797), .ZN(n13784) );
  NAND2_X1 U15735 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13784), .ZN(n13805) );
  OAI211_X1 U15736 ( .C1(n13784), .C2(P1_REG2_REG_18__SCAN_IN), .A(n13811), 
        .B(n13805), .ZN(n13796) );
  NAND2_X1 U15737 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n14290)
         );
  INV_X1 U15738 ( .A(n14290), .ZN(n13786) );
  NOR2_X1 U15739 ( .A1(n14380), .A2(n13797), .ZN(n13785) );
  AOI211_X1 U15740 ( .C1(n13787), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n13786), 
        .B(n13785), .ZN(n13795) );
  AOI21_X1 U15741 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13789), .A(n13788), 
        .ZN(n13798) );
  XNOR2_X1 U15742 ( .A(n13797), .B(n13798), .ZN(n13790) );
  INV_X1 U15743 ( .A(n13790), .ZN(n13793) );
  NOR2_X1 U15744 ( .A1(n13791), .A2(n13790), .ZN(n13799) );
  INV_X1 U15745 ( .A(n13799), .ZN(n13792) );
  OAI211_X1 U15746 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13793), .A(n14375), 
        .B(n13792), .ZN(n13794) );
  NAND3_X1 U15747 ( .A1(n13796), .A2(n13795), .A3(n13794), .ZN(P1_U3261) );
  NOR2_X1 U15748 ( .A1(n13798), .A2(n13797), .ZN(n13800) );
  NOR2_X1 U15749 ( .A1(n13800), .A2(n13799), .ZN(n13802) );
  XOR2_X1 U15750 ( .A(n13802), .B(n13801), .Z(n13812) );
  INV_X1 U15751 ( .A(n13812), .ZN(n13809) );
  NAND2_X1 U15752 ( .A1(n13804), .A2(n13803), .ZN(n13806) );
  NAND2_X1 U15753 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  XOR2_X1 U15754 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13807), .Z(n13810) );
  OAI21_X1 U15755 ( .B1(n13810), .B2(n14370), .A(n14380), .ZN(n13808) );
  AOI21_X1 U15756 ( .B1(n13809), .B2(n14375), .A(n13808), .ZN(n13814) );
  AOI22_X1 U15757 ( .A1(n13812), .A2(n14375), .B1(n13811), .B2(n13810), .ZN(
        n13813) );
  MUX2_X1 U15758 ( .A(n13814), .B(n13813), .S(n13897), .Z(n13816) );
  OAI211_X1 U15759 ( .C1(n6901), .C2(n14384), .A(n13816), .B(n13815), .ZN(
        P1_U3262) );
  OR2_X2 U15760 ( .A1(n13866), .A2(n14028), .ZN(n13868) );
  NAND2_X1 U15761 ( .A1(n13840), .A2(n14019), .ZN(n13817) );
  XNOR2_X1 U15762 ( .A(n14016), .B(n13817), .ZN(n13818) );
  NAND2_X1 U15763 ( .A1(n13818), .A2(n14448), .ZN(n14015) );
  INV_X1 U15764 ( .A(P1_B_REG_SCAN_IN), .ZN(n13819) );
  NOR2_X1 U15765 ( .A1(n14122), .A2(n13819), .ZN(n13820) );
  NOR2_X1 U15766 ( .A1(n14356), .A2(n13820), .ZN(n13843) );
  NAND2_X1 U15767 ( .A1(n13843), .A2(n13821), .ZN(n14017) );
  NOR2_X1 U15768 ( .A1(n14395), .A2(n14017), .ZN(n13827) );
  NOR2_X1 U15769 ( .A1(n14016), .A2(n14444), .ZN(n13822) );
  AOI211_X1 U15770 ( .C1(n14441), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13827), 
        .B(n13822), .ZN(n13823) );
  OAI21_X1 U15771 ( .B1(n14015), .B2(n13917), .A(n13823), .ZN(P1_U3263) );
  XNOR2_X1 U15772 ( .A(n13840), .B(n13824), .ZN(n13825) );
  NAND2_X1 U15773 ( .A1(n13825), .A2(n14448), .ZN(n14018) );
  NOR2_X1 U15774 ( .A1(n14019), .A2(n14444), .ZN(n13826) );
  AOI211_X1 U15775 ( .C1(n14441), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13827), 
        .B(n13826), .ZN(n13828) );
  OAI21_X1 U15776 ( .B1(n13917), .B2(n14018), .A(n13828), .ZN(P1_U3264) );
  NAND2_X1 U15777 ( .A1(n13862), .A2(n13861), .ZN(n13860) );
  OAI21_X1 U15778 ( .B1(n13832), .B2(n13831), .A(n13860), .ZN(n13833) );
  NOR2_X1 U15779 ( .A1(n13835), .A2(n13834), .ZN(n13854) );
  INV_X1 U15780 ( .A(n13861), .ZN(n13855) );
  NAND2_X1 U15781 ( .A1(n13853), .A2(n13837), .ZN(n13839) );
  XNOR2_X1 U15782 ( .A(n13839), .B(n6737), .ZN(n14025) );
  NAND2_X1 U15783 ( .A1(n14024), .A2(n14452), .ZN(n13850) );
  NAND2_X1 U15784 ( .A1(n13843), .A2(n13842), .ZN(n14021) );
  OAI22_X1 U15785 ( .A1(n13845), .A2(n14021), .B1(n13844), .B2(n14439), .ZN(
        n13848) );
  NAND2_X1 U15786 ( .A1(n13846), .A2(n14353), .ZN(n14020) );
  NOR2_X1 U15787 ( .A1(n14395), .A2(n14020), .ZN(n13847) );
  AOI211_X1 U15788 ( .C1(n14441), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13848), 
        .B(n13847), .ZN(n13849) );
  OAI211_X1 U15789 ( .C1(n14022), .C2(n14444), .A(n13850), .B(n13849), .ZN(
        n13851) );
  AOI21_X1 U15790 ( .B1(n14025), .B2(n13995), .A(n13851), .ZN(n13852) );
  OAI21_X1 U15791 ( .B1(n14026), .B2(n13998), .A(n13852), .ZN(P1_U3356) );
  INV_X1 U15792 ( .A(n13853), .ZN(n13857) );
  NOR3_X1 U15793 ( .A1(n13836), .A2(n13855), .A3(n13854), .ZN(n13856) );
  OAI21_X1 U15794 ( .B1(n13857), .B2(n13856), .A(n14522), .ZN(n13859) );
  OAI21_X1 U15795 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n14031) );
  NAND2_X1 U15796 ( .A1(n14395), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13863) );
  OAI21_X1 U15797 ( .B1(n14439), .B2(n13864), .A(n13863), .ZN(n13865) );
  AOI21_X1 U15798 ( .B1(n14028), .B2(n14396), .A(n13865), .ZN(n13870) );
  AOI21_X1 U15799 ( .B1(n14028), .B2(n13866), .A(n14492), .ZN(n13867) );
  AND2_X1 U15800 ( .A1(n13868), .A2(n13867), .ZN(n14027) );
  NAND2_X1 U15801 ( .A1(n14027), .A2(n13992), .ZN(n13869) );
  OAI211_X1 U15802 ( .C1(n14031), .C2(n13998), .A(n13870), .B(n13869), .ZN(
        n13871) );
  INV_X1 U15803 ( .A(n13871), .ZN(n13872) );
  OAI21_X1 U15804 ( .B1(n14030), .B2(n13987), .A(n13872), .ZN(P1_U3265) );
  XNOR2_X1 U15805 ( .A(n13874), .B(n13873), .ZN(n14042) );
  INV_X1 U15806 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13876) );
  OAI22_X1 U15807 ( .A1(n14010), .A2(n13876), .B1(n13875), .B2(n14439), .ZN(
        n13886) );
  AOI21_X1 U15808 ( .B1(n13879), .B2(n13878), .A(n13877), .ZN(n13880) );
  OR2_X1 U15809 ( .A1(n13880), .A2(n14566), .ZN(n14041) );
  AOI21_X1 U15810 ( .B1(n14039), .B2(n13894), .A(n14492), .ZN(n13883) );
  AND2_X1 U15811 ( .A1(n13883), .A2(n13882), .ZN(n14037) );
  AOI21_X1 U15812 ( .B1(n14037), .B2(n13897), .A(n14038), .ZN(n13884) );
  AOI21_X1 U15813 ( .B1(n14041), .B2(n13884), .A(n14395), .ZN(n13885) );
  AOI211_X1 U15814 ( .C1(n14396), .C2(n14039), .A(n13886), .B(n13885), .ZN(
        n13887) );
  OAI21_X1 U15815 ( .B1(n13998), .B2(n14042), .A(n13887), .ZN(P1_U3267) );
  XNOR2_X1 U15816 ( .A(n13889), .B(n13888), .ZN(n14049) );
  INV_X1 U15817 ( .A(n13890), .ZN(n13891) );
  AOI21_X1 U15818 ( .B1(n13893), .B2(n13892), .A(n13891), .ZN(n14046) );
  AOI211_X1 U15819 ( .C1(n14045), .C2(n13915), .A(n14492), .B(n13881), .ZN(
        n14043) );
  NOR2_X1 U15820 ( .A1(n14439), .A2(n13895), .ZN(n13896) );
  AOI211_X1 U15821 ( .C1(n14043), .C2(n13897), .A(n13896), .B(n14044), .ZN(
        n13899) );
  AOI22_X1 U15822 ( .A1(n14045), .A2(n14396), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n13987), .ZN(n13898) );
  OAI21_X1 U15823 ( .B1(n13899), .B2(n13987), .A(n13898), .ZN(n13900) );
  AOI21_X1 U15824 ( .B1(n14046), .B2(n13953), .A(n13900), .ZN(n13901) );
  OAI21_X1 U15825 ( .B1(n13955), .B2(n14049), .A(n13901), .ZN(P1_U3268) );
  NAND2_X1 U15826 ( .A1(n13902), .A2(n7205), .ZN(n13903) );
  NAND2_X1 U15827 ( .A1(n13904), .A2(n13903), .ZN(n14050) );
  INV_X1 U15828 ( .A(n14050), .ZN(n13924) );
  NAND2_X1 U15829 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  NAND2_X1 U15830 ( .A1(n13907), .A2(n14522), .ZN(n13911) );
  NAND2_X1 U15831 ( .A1(n14050), .A2(n14531), .ZN(n13910) );
  INV_X1 U15832 ( .A(n13908), .ZN(n13909) );
  OAI211_X1 U15833 ( .C1(n13912), .C2(n13911), .A(n13910), .B(n13909), .ZN(
        n14055) );
  NAND2_X1 U15834 ( .A1(n14055), .A2(n14010), .ZN(n13922) );
  INV_X1 U15835 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13914) );
  OAI22_X1 U15836 ( .A1(n14010), .A2(n13914), .B1(n13913), .B2(n14439), .ZN(
        n13919) );
  AOI21_X1 U15837 ( .B1(n13920), .B2(n13932), .A(n14492), .ZN(n13916) );
  NAND2_X1 U15838 ( .A1(n13916), .A2(n13915), .ZN(n14051) );
  NOR2_X1 U15839 ( .A1(n14051), .A2(n13917), .ZN(n13918) );
  AOI211_X1 U15840 ( .C1(n14396), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        n13921) );
  OAI211_X1 U15841 ( .C1(n13924), .C2(n13923), .A(n13922), .B(n13921), .ZN(
        P1_U3269) );
  OAI21_X1 U15842 ( .B1(n7389), .B2(n13926), .A(n13925), .ZN(n14061) );
  OAI21_X1 U15843 ( .B1(n13929), .B2(n13928), .A(n13927), .ZN(n13930) );
  NAND2_X1 U15844 ( .A1(n13930), .A2(n14522), .ZN(n14059) );
  INV_X1 U15845 ( .A(n14059), .ZN(n13931) );
  OAI21_X1 U15846 ( .B1(n13931), .B2(n14057), .A(n14010), .ZN(n13941) );
  INV_X1 U15847 ( .A(n13946), .ZN(n13934) );
  INV_X1 U15848 ( .A(n13932), .ZN(n13933) );
  AOI211_X1 U15849 ( .C1(n14058), .C2(n13934), .A(n14492), .B(n13933), .ZN(
        n14056) );
  INV_X1 U15850 ( .A(n13935), .ZN(n13936) );
  AOI22_X1 U15851 ( .A1(n14395), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13936), 
        .B2(n14394), .ZN(n13937) );
  OAI21_X1 U15852 ( .B1(n13938), .B2(n14444), .A(n13937), .ZN(n13939) );
  AOI21_X1 U15853 ( .B1(n14056), .B2(n14452), .A(n13939), .ZN(n13940) );
  OAI211_X1 U15854 ( .C1(n13998), .C2(n14061), .A(n13941), .B(n13940), .ZN(
        P1_U3270) );
  XOR2_X1 U15855 ( .A(n13942), .B(n13944), .Z(n14068) );
  OAI21_X1 U15856 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n14066) );
  AOI211_X1 U15857 ( .C1(n13947), .C2(n6525), .A(n14492), .B(n13946), .ZN(
        n14064) );
  NAND2_X1 U15858 ( .A1(n14064), .A2(n14452), .ZN(n13951) );
  OAI22_X1 U15859 ( .A1(n14441), .A2(n14062), .B1(n13948), .B2(n14439), .ZN(
        n13949) );
  AOI21_X1 U15860 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n14395), .A(n13949), 
        .ZN(n13950) );
  OAI211_X1 U15861 ( .C1(n14444), .C2(n14063), .A(n13951), .B(n13950), .ZN(
        n13952) );
  AOI21_X1 U15862 ( .B1(n13953), .B2(n14066), .A(n13952), .ZN(n13954) );
  OAI21_X1 U15863 ( .B1(n14068), .B2(n13955), .A(n13954), .ZN(P1_U3271) );
  XNOR2_X1 U15864 ( .A(n13956), .B(n13961), .ZN(n14074) );
  INV_X1 U15865 ( .A(n6525), .ZN(n13957) );
  AOI211_X1 U15866 ( .C1(n14071), .C2(n6597), .A(n14492), .B(n13957), .ZN(
        n14069) );
  INV_X1 U15867 ( .A(n14069), .ZN(n13965) );
  INV_X1 U15868 ( .A(n13958), .ZN(n13959) );
  AOI21_X1 U15869 ( .B1(n13959), .B2(n14394), .A(n14070), .ZN(n13963) );
  XNOR2_X1 U15870 ( .A(n13960), .B(n13961), .ZN(n13962) );
  NAND2_X1 U15871 ( .A1(n13962), .A2(n14522), .ZN(n14072) );
  OAI211_X1 U15872 ( .C1(n13965), .C2(n13964), .A(n13963), .B(n14072), .ZN(
        n13966) );
  NAND2_X1 U15873 ( .A1(n13966), .A2(n14010), .ZN(n13968) );
  AOI22_X1 U15874 ( .A1(n14071), .A2(n14396), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n13987), .ZN(n13967) );
  OAI211_X1 U15875 ( .C1(n13998), .C2(n14074), .A(n13968), .B(n13967), .ZN(
        P1_U3272) );
  OAI21_X1 U15876 ( .B1(n13970), .B2(n13972), .A(n13969), .ZN(n14082) );
  AOI21_X1 U15877 ( .B1(n13972), .B2(n13971), .A(n6589), .ZN(n14075) );
  NAND2_X1 U15878 ( .A1(n14075), .A2(n13995), .ZN(n13981) );
  OR2_X1 U15879 ( .A1(n14077), .A2(n13984), .ZN(n13973) );
  AND2_X1 U15880 ( .A1(n6597), .A2(n13973), .ZN(n14079) );
  OAI22_X1 U15881 ( .A1(n14441), .A2(n14076), .B1(n13974), .B2(n14439), .ZN(
        n13975) );
  INV_X1 U15882 ( .A(n13975), .ZN(n13977) );
  NAND2_X1 U15883 ( .A1(n14441), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n13976) );
  OAI211_X1 U15884 ( .C1(n14077), .C2(n14444), .A(n13977), .B(n13976), .ZN(
        n13978) );
  AOI21_X1 U15885 ( .B1(n14079), .B2(n13979), .A(n13978), .ZN(n13980) );
  OAI211_X1 U15886 ( .C1(n13998), .C2(n14082), .A(n13981), .B(n13980), .ZN(
        P1_U3273) );
  XNOR2_X1 U15887 ( .A(n13983), .B(n13982), .ZN(n14089) );
  AOI211_X1 U15888 ( .C1(n14085), .C2(n13985), .A(n14492), .B(n13984), .ZN(
        n14083) );
  INV_X1 U15889 ( .A(n14084), .ZN(n13988) );
  OAI22_X1 U15890 ( .A1(n13988), .A2(n13987), .B1(n13986), .B2(n14439), .ZN(
        n13989) );
  AOI21_X1 U15891 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n14395), .A(n13989), 
        .ZN(n13990) );
  OAI21_X1 U15892 ( .B1(n6815), .B2(n14444), .A(n13990), .ZN(n13991) );
  AOI21_X1 U15893 ( .B1(n14083), .B2(n13992), .A(n13991), .ZN(n13997) );
  XNOR2_X1 U15894 ( .A(n13993), .B(n13994), .ZN(n14086) );
  NAND2_X1 U15895 ( .A1(n14086), .A2(n13995), .ZN(n13996) );
  OAI211_X1 U15896 ( .C1(n13998), .C2(n14089), .A(n13997), .B(n13996), .ZN(
        P1_U3274) );
  XNOR2_X1 U15897 ( .A(n13999), .B(n14000), .ZN(n14090) );
  XNOR2_X1 U15898 ( .A(n14001), .B(n14000), .ZN(n14005) );
  AOI22_X1 U15899 ( .A1(n14004), .A2(n14003), .B1(n14353), .B2(n14002), .ZN(
        n14285) );
  OAI21_X1 U15900 ( .B1(n14005), .B2(n14566), .A(n14285), .ZN(n14006) );
  AOI21_X1 U15901 ( .B1(n14531), .B2(n14090), .A(n14006), .ZN(n14094) );
  XNOR2_X1 U15902 ( .A(n14007), .B(n14092), .ZN(n14008) );
  NOR2_X1 U15903 ( .A1(n14008), .A2(n14492), .ZN(n14091) );
  OAI22_X1 U15904 ( .A1(n14010), .A2(n14009), .B1(n14292), .B2(n14439), .ZN(
        n14012) );
  INV_X1 U15905 ( .A(n14092), .ZN(n14287) );
  NOR2_X1 U15906 ( .A1(n14287), .A2(n14444), .ZN(n14011) );
  AOI211_X1 U15907 ( .C1(n14091), .C2(n14452), .A(n14012), .B(n14011), .ZN(
        n14014) );
  NAND2_X1 U15908 ( .A1(n14090), .A2(n14453), .ZN(n14013) );
  OAI211_X1 U15909 ( .C1(n14094), .C2(n14395), .A(n14014), .B(n14013), .ZN(
        P1_U3275) );
  MUX2_X1 U15910 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14097), .S(n14594), .Z(
        P1_U3559) );
  OAI211_X1 U15911 ( .C1(n14019), .C2(n14570), .A(n14018), .B(n14017), .ZN(
        n14098) );
  MUX2_X1 U15912 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14098), .S(n14594), .Z(
        P1_U3558) );
  OAI211_X1 U15913 ( .C1(n14022), .C2(n14570), .A(n14021), .B(n14020), .ZN(
        n14023) );
  MUX2_X1 U15914 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14099), .S(n14594), .Z(
        P1_U3557) );
  AOI21_X1 U15915 ( .B1(n14549), .B2(n14028), .A(n14027), .ZN(n14029) );
  OAI211_X1 U15916 ( .C1(n14517), .C2(n14031), .A(n14030), .B(n14029), .ZN(
        n14100) );
  MUX2_X1 U15917 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14100), .S(n14594), .Z(
        P1_U3556) );
  AOI21_X1 U15918 ( .B1(n14549), .B2(n14033), .A(n14032), .ZN(n14034) );
  MUX2_X1 U15919 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14101), .S(n14594), .Z(
        P1_U3555) );
  AOI211_X1 U15920 ( .C1(n14549), .C2(n14039), .A(n14038), .B(n14037), .ZN(
        n14040) );
  OAI211_X1 U15921 ( .C1(n14517), .C2(n14042), .A(n14041), .B(n14040), .ZN(
        n14102) );
  MUX2_X1 U15922 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14102), .S(n14594), .Z(
        P1_U3554) );
  AOI211_X1 U15923 ( .C1(n14549), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14048) );
  NAND2_X1 U15924 ( .A1(n14046), .A2(n14574), .ZN(n14047) );
  OAI211_X1 U15925 ( .C1(n14566), .C2(n14049), .A(n14048), .B(n14047), .ZN(
        n14103) );
  MUX2_X1 U15926 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14103), .S(n14594), .Z(
        P1_U3553) );
  INV_X1 U15927 ( .A(n14095), .ZN(n14564) );
  NAND2_X1 U15928 ( .A1(n14050), .A2(n14564), .ZN(n14052) );
  OAI211_X1 U15929 ( .C1(n14053), .C2(n14570), .A(n14052), .B(n14051), .ZN(
        n14054) );
  OR2_X1 U15930 ( .A1(n14055), .A2(n14054), .ZN(n14104) );
  MUX2_X1 U15931 ( .A(n14104), .B(P1_REG1_REG_24__SCAN_IN), .S(n14591), .Z(
        P1_U3552) );
  AOI211_X1 U15932 ( .C1(n14549), .C2(n14058), .A(n14057), .B(n14056), .ZN(
        n14060) );
  OAI211_X1 U15933 ( .C1(n14517), .C2(n14061), .A(n14060), .B(n14059), .ZN(
        n14105) );
  MUX2_X1 U15934 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14105), .S(n14594), .Z(
        P1_U3551) );
  OAI21_X1 U15935 ( .B1(n14063), .B2(n14570), .A(n14062), .ZN(n14065) );
  AOI211_X1 U15936 ( .C1(n14574), .C2(n14066), .A(n14065), .B(n14064), .ZN(
        n14067) );
  OAI21_X1 U15937 ( .B1(n14566), .B2(n14068), .A(n14067), .ZN(n14106) );
  MUX2_X1 U15938 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14106), .S(n14594), .Z(
        P1_U3550) );
  AOI211_X1 U15939 ( .C1(n14549), .C2(n14071), .A(n14070), .B(n14069), .ZN(
        n14073) );
  OAI211_X1 U15940 ( .C1(n14517), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        n14107) );
  MUX2_X1 U15941 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14107), .S(n14594), .Z(
        P1_U3549) );
  NAND2_X1 U15942 ( .A1(n14075), .A2(n14522), .ZN(n14081) );
  OAI21_X1 U15943 ( .B1(n14077), .B2(n14570), .A(n14076), .ZN(n14078) );
  AOI21_X1 U15944 ( .B1(n14079), .B2(n14448), .A(n14078), .ZN(n14080) );
  OAI211_X1 U15945 ( .C1(n14517), .C2(n14082), .A(n14081), .B(n14080), .ZN(
        n14108) );
  MUX2_X1 U15946 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14108), .S(n14594), .Z(
        P1_U3548) );
  AOI211_X1 U15947 ( .C1(n14549), .C2(n14085), .A(n14084), .B(n14083), .ZN(
        n14088) );
  NAND2_X1 U15948 ( .A1(n14086), .A2(n14522), .ZN(n14087) );
  OAI211_X1 U15949 ( .C1(n14517), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        n14109) );
  MUX2_X1 U15950 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14109), .S(n14594), .Z(
        P1_U3547) );
  INV_X1 U15951 ( .A(n14090), .ZN(n14096) );
  AOI21_X1 U15952 ( .B1(n14549), .B2(n14092), .A(n14091), .ZN(n14093) );
  OAI211_X1 U15953 ( .C1(n14096), .C2(n14095), .A(n14094), .B(n14093), .ZN(
        n14110) );
  MUX2_X1 U15954 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14110), .S(n14594), .Z(
        P1_U3546) );
  MUX2_X1 U15955 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14098), .S(n14578), .Z(
        P1_U3526) );
  MUX2_X1 U15956 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14099), .S(n14578), .Z(
        P1_U3525) );
  MUX2_X1 U15957 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14100), .S(n14578), .Z(
        P1_U3524) );
  MUX2_X1 U15958 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14101), .S(n14578), .Z(
        P1_U3523) );
  MUX2_X1 U15959 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14102), .S(n14578), .Z(
        P1_U3522) );
  MUX2_X1 U15960 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14103), .S(n14578), .Z(
        P1_U3521) );
  MUX2_X1 U15961 ( .A(n14104), .B(P1_REG0_REG_24__SCAN_IN), .S(n14576), .Z(
        P1_U3520) );
  MUX2_X1 U15962 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14105), .S(n14578), .Z(
        P1_U3519) );
  MUX2_X1 U15963 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14106), .S(n14578), .Z(
        P1_U3518) );
  MUX2_X1 U15964 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14107), .S(n14578), .Z(
        P1_U3517) );
  MUX2_X1 U15965 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14108), .S(n14578), .Z(
        P1_U3516) );
  MUX2_X1 U15966 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14109), .S(n14578), .Z(
        P1_U3515) );
  MUX2_X1 U15967 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14110), .S(n14578), .Z(
        P1_U3513) );
  INV_X1 U15968 ( .A(n14111), .ZN(n14112) );
  NOR4_X1 U15969 ( .A1(n14112), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8135), .A4(
        P1_U3086), .ZN(n14113) );
  AOI21_X1 U15970 ( .B1(n14114), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14113), 
        .ZN(n14115) );
  OAI21_X1 U15971 ( .B1(n14116), .B2(n14128), .A(n14115), .ZN(P1_U3324) );
  OAI222_X1 U15972 ( .A1(n14119), .A2(P1_U3086), .B1(n14128), .B2(n14118), 
        .C1(n14117), .C2(n14125), .ZN(P1_U3325) );
  OAI222_X1 U15973 ( .A1(n14125), .A2(n6660), .B1(n14128), .B2(n14121), .C1(
        n14120), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U15974 ( .A1(n14125), .A2(n14124), .B1(n14128), .B2(n14123), .C1(
        n14122), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U15975 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14126) );
  OAI222_X1 U15976 ( .A1(P1_U3086), .A2(n14129), .B1(n14128), .B2(n14127), 
        .C1(n14126), .C2(n14125), .ZN(P1_U3329) );
  MUX2_X1 U15977 ( .A(n14131), .B(n14130), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U15978 ( .A(n14132), .ZN(n14133) );
  MUX2_X1 U15979 ( .A(n14133), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15980 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14678) );
  XNOR2_X1 U15981 ( .A(n14678), .B(n14137), .ZN(SUB_1596_U62) );
  AOI21_X1 U15982 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14138) );
  OAI21_X1 U15983 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14138), 
        .ZN(U28) );
  AOI21_X1 U15984 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14139) );
  OAI21_X1 U15985 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14139), 
        .ZN(U29) );
  AOI21_X1 U15986 ( .B1(n14142), .B2(n14141), .A(n14140), .ZN(n14143) );
  XOR2_X1 U15987 ( .A(n14143), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U15988 ( .A(n14145), .B(n14144), .Z(SUB_1596_U57) );
  XOR2_X1 U15989 ( .A(n14146), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  OAI21_X1 U15990 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14151) );
  XOR2_X1 U15991 ( .A(n14151), .B(n14150), .Z(SUB_1596_U54) );
  OAI21_X1 U15992 ( .B1(n14154), .B2(n14153), .A(n14152), .ZN(n14156) );
  XOR2_X1 U15993 ( .A(n14156), .B(n14155), .Z(SUB_1596_U70) );
  OAI21_X1 U15994 ( .B1(n14158), .B2(n14570), .A(n14157), .ZN(n14160) );
  AOI211_X1 U15995 ( .C1(n14161), .C2(n14574), .A(n14160), .B(n14159), .ZN(
        n14163) );
  INV_X1 U15996 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U15997 ( .A1(n14578), .A2(n14163), .B1(n14162), .B2(n14576), .ZN(
        P1_U3495) );
  AOI22_X1 U15998 ( .A1(n14594), .A2(n14163), .B1(n10149), .B2(n14591), .ZN(
        P1_U3540) );
  OAI21_X1 U15999 ( .B1(n14166), .B2(n14165), .A(n14164), .ZN(n14167) );
  XNOR2_X1 U16000 ( .A(n14167), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI21_X1 U16001 ( .B1(n14170), .B2(n14169), .A(n14168), .ZN(n14184) );
  OAI21_X1 U16002 ( .B1(n14172), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14171), 
        .ZN(n14182) );
  NAND2_X1 U16003 ( .A1(n14926), .A2(n14173), .ZN(n14175) );
  OAI211_X1 U16004 ( .C1(n14176), .C2(n14930), .A(n14175), .B(n14174), .ZN(
        n14181) );
  AOI211_X1 U16005 ( .C1(n14179), .C2(n14178), .A(n14915), .B(n14177), .ZN(
        n14180) );
  AOI211_X1 U16006 ( .C1(n14910), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14183) );
  OAI21_X1 U16007 ( .B1(n14184), .B2(n14921), .A(n14183), .ZN(P3_U3199) );
  XNOR2_X1 U16008 ( .A(n14185), .B(n14186), .ZN(n14187) );
  OAI222_X1 U16009 ( .A1(n14998), .A2(n14202), .B1(n14996), .B2(n14188), .C1(
        n14187), .C2(n14988), .ZN(n14214) );
  OAI22_X1 U16010 ( .A1(n14190), .A2(n15010), .B1(n14978), .B2(n14189), .ZN(
        n14197) );
  XNOR2_X1 U16011 ( .A(n14192), .B(n14191), .ZN(n14216) );
  INV_X1 U16012 ( .A(n14216), .ZN(n14195) );
  NOR2_X1 U16013 ( .A1(n14193), .A2(n15047), .ZN(n14215) );
  INV_X1 U16014 ( .A(n14215), .ZN(n14194) );
  OAI22_X1 U16015 ( .A1(n14195), .A2(n14209), .B1(n14939), .B2(n14194), .ZN(
        n14196) );
  AOI211_X1 U16016 ( .C1(n15010), .C2(n14214), .A(n14197), .B(n14196), .ZN(
        n14198) );
  INV_X1 U16017 ( .A(n14198), .ZN(P3_U3220) );
  XOR2_X1 U16018 ( .A(n14199), .B(n14205), .Z(n14200) );
  OAI222_X1 U16019 ( .A1(n14996), .A2(n14202), .B1(n14998), .B2(n14201), .C1(
        n14200), .C2(n14988), .ZN(n14222) );
  OAI22_X1 U16020 ( .A1(n14204), .A2(n15010), .B1(n14978), .B2(n14203), .ZN(
        n14212) );
  XNOR2_X1 U16021 ( .A(n14206), .B(n14205), .ZN(n14224) );
  INV_X1 U16022 ( .A(n14224), .ZN(n14210) );
  NOR2_X1 U16023 ( .A1(n14207), .A2(n15047), .ZN(n14223) );
  INV_X1 U16024 ( .A(n14223), .ZN(n14208) );
  OAI22_X1 U16025 ( .A1(n14210), .A2(n14209), .B1(n14939), .B2(n14208), .ZN(
        n14211) );
  AOI211_X1 U16026 ( .C1(n15010), .C2(n14222), .A(n14212), .B(n14211), .ZN(
        n14213) );
  INV_X1 U16027 ( .A(n14213), .ZN(P3_U3222) );
  AOI211_X1 U16028 ( .C1(n14216), .C2(n15063), .A(n14215), .B(n14214), .ZN(
        n14226) );
  AOI22_X1 U16029 ( .A1(n15079), .A2(n14226), .B1(n9316), .B2(n15077), .ZN(
        P3_U3472) );
  NOR2_X1 U16030 ( .A1(n14218), .A2(n14217), .ZN(n14220) );
  AOI211_X1 U16031 ( .C1(n15015), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14228) );
  AOI22_X1 U16032 ( .A1(n15079), .A2(n14228), .B1(n9305), .B2(n15077), .ZN(
        P3_U3471) );
  AOI211_X1 U16033 ( .C1(n14224), .C2(n15063), .A(n14223), .B(n14222), .ZN(
        n14230) );
  AOI22_X1 U16034 ( .A1(n15079), .A2(n14230), .B1(n9288), .B2(n15077), .ZN(
        P3_U3470) );
  INV_X1 U16035 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U16036 ( .A1(n15066), .A2(n14226), .B1(n14225), .B2(n15064), .ZN(
        P3_U3429) );
  INV_X1 U16037 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U16038 ( .A1(n15066), .A2(n14228), .B1(n14227), .B2(n15064), .ZN(
        P3_U3426) );
  INV_X1 U16039 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U16040 ( .A1(n15066), .A2(n14230), .B1(n14229), .B2(n15064), .ZN(
        P3_U3423) );
  NAND2_X1 U16041 ( .A1(n14232), .A2(n14231), .ZN(n14233) );
  NAND2_X1 U16042 ( .A1(n14234), .A2(n14233), .ZN(n14236) );
  AOI222_X1 U16043 ( .A1(n14240), .A2(n14239), .B1(n14238), .B2(n14237), .C1(
        n14236), .C2(n14235), .ZN(n14241) );
  NAND2_X1 U16044 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14642)
         );
  OAI211_X1 U16045 ( .C1(n14243), .C2(n14242), .A(n14241), .B(n14642), .ZN(
        P2_U3187) );
  OAI21_X1 U16046 ( .B1(n14246), .B2(n14245), .A(n14244), .ZN(n14248) );
  AOI222_X1 U16047 ( .A1(n14249), .A2(n14364), .B1(n14248), .B2(n14359), .C1(
        n14247), .C2(n14297), .ZN(n14251) );
  OAI211_X1 U16048 ( .C1(n14367), .C2(n14252), .A(n14251), .B(n14250), .ZN(
        P1_U3215) );
  OAI21_X1 U16049 ( .B1(n14255), .B2(n14254), .A(n14253), .ZN(n14257) );
  AOI222_X1 U16050 ( .A1(n14258), .A2(n14364), .B1(n14257), .B2(n14359), .C1(
        n14256), .C2(n14297), .ZN(n14260) );
  OAI211_X1 U16051 ( .C1(n14367), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        P1_U3226) );
  INV_X1 U16052 ( .A(n14262), .ZN(n14263) );
  NOR2_X1 U16053 ( .A1(n14264), .A2(n14263), .ZN(n14265) );
  XNOR2_X1 U16054 ( .A(n14266), .B(n14265), .ZN(n14269) );
  OAI22_X1 U16055 ( .A1(n14305), .A2(n14286), .B1(n14267), .B2(n14284), .ZN(
        n14268) );
  AOI21_X1 U16056 ( .B1(n14269), .B2(n14359), .A(n14268), .ZN(n14271) );
  OAI211_X1 U16057 ( .C1(n14367), .C2(n14272), .A(n14271), .B(n14270), .ZN(
        P1_U3228) );
  OAI21_X1 U16058 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14277) );
  AOI222_X1 U16059 ( .A1(n14278), .A2(n14364), .B1(n14277), .B2(n14359), .C1(
        n14276), .C2(n14297), .ZN(n14280) );
  OAI211_X1 U16060 ( .C1(n14367), .C2(n14281), .A(n14280), .B(n14279), .ZN(
        P1_U3236) );
  XNOR2_X1 U16061 ( .A(n14283), .B(n14282), .ZN(n14289) );
  OAI22_X1 U16062 ( .A1(n14287), .A2(n14286), .B1(n14285), .B2(n14284), .ZN(
        n14288) );
  AOI21_X1 U16063 ( .B1(n14289), .B2(n14359), .A(n14288), .ZN(n14291) );
  OAI211_X1 U16064 ( .C1(n14367), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        P1_U3238) );
  NAND2_X1 U16065 ( .A1(n14293), .A2(n14294), .ZN(n14295) );
  NAND2_X1 U16066 ( .A1(n14296), .A2(n14295), .ZN(n14299) );
  AOI222_X1 U16067 ( .A1(n14300), .A2(n14364), .B1(n14299), .B2(n14359), .C1(
        n14298), .C2(n14297), .ZN(n14301) );
  NAND2_X1 U16068 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14382)
         );
  OAI211_X1 U16069 ( .C1(n14367), .C2(n14302), .A(n14301), .B(n14382), .ZN(
        P1_U3241) );
  AND2_X1 U16070 ( .A1(n14303), .A2(n14574), .ZN(n14308) );
  OAI21_X1 U16071 ( .B1(n14305), .B2(n14570), .A(n14304), .ZN(n14306) );
  NOR3_X1 U16072 ( .A1(n14308), .A2(n14307), .A3(n14306), .ZN(n14325) );
  AOI22_X1 U16073 ( .A1(n14594), .A2(n14325), .B1(n13764), .B2(n14591), .ZN(
        P1_U3545) );
  OAI21_X1 U16074 ( .B1(n6817), .B2(n14570), .A(n14309), .ZN(n14312) );
  INV_X1 U16075 ( .A(n14310), .ZN(n14311) );
  AOI211_X1 U16076 ( .C1(n14313), .C2(n14574), .A(n14312), .B(n14311), .ZN(
        n14327) );
  AOI22_X1 U16077 ( .A1(n14594), .A2(n14327), .B1(n14373), .B2(n14591), .ZN(
        P1_U3543) );
  OAI21_X1 U16078 ( .B1(n6819), .B2(n14570), .A(n14314), .ZN(n14316) );
  AOI211_X1 U16079 ( .C1(n14317), .C2(n14574), .A(n14316), .B(n14315), .ZN(
        n14329) );
  AOI22_X1 U16080 ( .A1(n14594), .A2(n14329), .B1(n14318), .B2(n14591), .ZN(
        P1_U3541) );
  OAI21_X1 U16081 ( .B1(n14320), .B2(n14570), .A(n14319), .ZN(n14322) );
  AOI211_X1 U16082 ( .C1(n14323), .C2(n14574), .A(n14322), .B(n14321), .ZN(
        n14331) );
  AOI22_X1 U16083 ( .A1(n14594), .A2(n14331), .B1(n8027), .B2(n14591), .ZN(
        P1_U3539) );
  INV_X1 U16084 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14324) );
  AOI22_X1 U16085 ( .A1(n14578), .A2(n14325), .B1(n14324), .B2(n14576), .ZN(
        P1_U3510) );
  INV_X1 U16086 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14326) );
  AOI22_X1 U16087 ( .A1(n14578), .A2(n14327), .B1(n14326), .B2(n14576), .ZN(
        P1_U3504) );
  INV_X1 U16088 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U16089 ( .A1(n14578), .A2(n14329), .B1(n14328), .B2(n14576), .ZN(
        P1_U3498) );
  INV_X1 U16090 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U16091 ( .A1(n14578), .A2(n14331), .B1(n14330), .B2(n14576), .ZN(
        P1_U3492) );
  XNOR2_X1 U16092 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14332), .ZN(SUB_1596_U69)
         );
  XOR2_X1 U16093 ( .A(n14334), .B(n14333), .Z(SUB_1596_U68) );
  AOI21_X1 U16094 ( .B1(n14337), .B2(n14336), .A(n14335), .ZN(n14338) );
  XOR2_X1 U16095 ( .A(n14338), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16096 ( .B1(n14341), .B2(n14340), .A(n14339), .ZN(n14342) );
  XOR2_X1 U16097 ( .A(n14342), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16098 ( .B1(n14344), .B2(n6573), .A(n14343), .ZN(n14346) );
  XOR2_X1 U16099 ( .A(n14346), .B(n14345), .Z(SUB_1596_U65) );
  OAI222_X1 U16100 ( .A1(n14351), .A2(n14350), .B1(n14351), .B2(n14349), .C1(
        n14348), .C2(n14347), .ZN(SUB_1596_U64) );
  AND2_X1 U16101 ( .A1(n14447), .A2(n14549), .ZN(n14509) );
  AOI22_X1 U16102 ( .A1(n14352), .A2(n14509), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14366) );
  NAND2_X1 U16103 ( .A1(n14354), .A2(n14353), .ZN(n14355) );
  OAI21_X1 U16104 ( .B1(n14357), .B2(n14356), .A(n14355), .ZN(n14508) );
  OAI211_X1 U16105 ( .C1(n14361), .C2(n14360), .A(n14358), .B(n14359), .ZN(
        n14362) );
  INV_X1 U16106 ( .A(n14362), .ZN(n14363) );
  AOI21_X1 U16107 ( .B1(n14364), .B2(n14508), .A(n14363), .ZN(n14365) );
  OAI211_X1 U16108 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14367), .A(n14366), .B(
        n14365), .ZN(P1_U3218) );
  AOI21_X1 U16109 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14369), .A(n14368), 
        .ZN(n14371) );
  OR2_X1 U16110 ( .A1(n14371), .A2(n14370), .ZN(n14378) );
  OAI21_X1 U16111 ( .B1(n14374), .B2(n14373), .A(n14372), .ZN(n14376) );
  NAND2_X1 U16112 ( .A1(n14376), .A2(n14375), .ZN(n14377) );
  OAI211_X1 U16113 ( .C1(n14380), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        n14381) );
  INV_X1 U16114 ( .A(n14381), .ZN(n14383) );
  OAI211_X1 U16115 ( .C1(n14385), .C2(n14384), .A(n14383), .B(n14382), .ZN(
        P1_U3258) );
  XNOR2_X1 U16116 ( .A(n14387), .B(n14386), .ZN(n14563) );
  XNOR2_X1 U16117 ( .A(n14389), .B(n14388), .ZN(n14391) );
  OAI21_X1 U16118 ( .B1(n14391), .B2(n14566), .A(n14390), .ZN(n14392) );
  AOI21_X1 U16119 ( .B1(n14531), .B2(n14563), .A(n14392), .ZN(n14560) );
  AOI222_X1 U16120 ( .A1(n14557), .A2(n14396), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n14395), .C1(n14394), .C2(n14393), .ZN(n14401) );
  XOR2_X1 U16121 ( .A(n14397), .B(n14557), .Z(n14398) );
  NAND2_X1 U16122 ( .A1(n14398), .A2(n14448), .ZN(n14558) );
  INV_X1 U16123 ( .A(n14558), .ZN(n14399) );
  AOI22_X1 U16124 ( .A1(n14563), .A2(n14453), .B1(n14452), .B2(n14399), .ZN(
        n14400) );
  OAI211_X1 U16125 ( .C1(n14441), .C2(n14560), .A(n14401), .B(n14400), .ZN(
        P1_U3284) );
  OAI21_X1 U16126 ( .B1(n14403), .B2(n14405), .A(n14402), .ZN(n14408) );
  XNOR2_X1 U16127 ( .A(n14404), .B(n14405), .ZN(n14413) );
  NOR2_X1 U16128 ( .A1(n14413), .A2(n14497), .ZN(n14406) );
  AOI211_X1 U16129 ( .C1(n14522), .C2(n14408), .A(n14407), .B(n14406), .ZN(
        n14543) );
  NOR2_X1 U16130 ( .A1(n14439), .A2(n14409), .ZN(n14410) );
  AOI21_X1 U16131 ( .B1(n14441), .B2(P1_REG2_REG_7__SCAN_IN), .A(n14410), .ZN(
        n14411) );
  OAI21_X1 U16132 ( .B1(n14444), .B2(n14542), .A(n14411), .ZN(n14412) );
  INV_X1 U16133 ( .A(n14412), .ZN(n14418) );
  INV_X1 U16134 ( .A(n14413), .ZN(n14546) );
  OAI211_X1 U16135 ( .C1(n14542), .C2(n14415), .A(n14448), .B(n14414), .ZN(
        n14541) );
  INV_X1 U16136 ( .A(n14541), .ZN(n14416) );
  AOI22_X1 U16137 ( .A1(n14546), .A2(n14453), .B1(n14452), .B2(n14416), .ZN(
        n14417) );
  OAI211_X1 U16138 ( .C1(n14395), .C2(n14543), .A(n14418), .B(n14417), .ZN(
        P1_U3286) );
  XNOR2_X1 U16139 ( .A(n14419), .B(n14421), .ZN(n14529) );
  NAND3_X1 U16140 ( .A1(n14421), .A2(n14420), .A3(n10594), .ZN(n14422) );
  AOI21_X1 U16141 ( .B1(n10598), .B2(n14422), .A(n14566), .ZN(n14527) );
  AOI211_X1 U16142 ( .C1(n14531), .C2(n14529), .A(n14524), .B(n14527), .ZN(
        n14434) );
  INV_X1 U16143 ( .A(n14431), .ZN(n14426) );
  NOR2_X1 U16144 ( .A1(n14439), .A2(n14423), .ZN(n14424) );
  AOI21_X1 U16145 ( .B1(n14441), .B2(P1_REG2_REG_5__SCAN_IN), .A(n14424), .ZN(
        n14425) );
  OAI21_X1 U16146 ( .B1(n14444), .B2(n14426), .A(n14425), .ZN(n14427) );
  INV_X1 U16147 ( .A(n14427), .ZN(n14433) );
  INV_X1 U16148 ( .A(n14428), .ZN(n14429) );
  AOI211_X1 U16149 ( .C1(n14431), .C2(n14430), .A(n14492), .B(n14429), .ZN(
        n14526) );
  AOI22_X1 U16150 ( .A1(n14526), .A2(n14452), .B1(n14529), .B2(n14453), .ZN(
        n14432) );
  OAI211_X1 U16151 ( .C1(n14395), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        P1_U3288) );
  XNOR2_X1 U16152 ( .A(n14435), .B(n14437), .ZN(n14513) );
  NAND3_X1 U16153 ( .A1(n14437), .A2(n14436), .A3(n10630), .ZN(n14438) );
  AOI21_X1 U16154 ( .B1(n10584), .B2(n14438), .A(n14566), .ZN(n14511) );
  AOI211_X1 U16155 ( .C1(n14531), .C2(n14513), .A(n14508), .B(n14511), .ZN(
        n14456) );
  NOR2_X1 U16156 ( .A1(n14439), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14440) );
  AOI21_X1 U16157 ( .B1(n14441), .B2(P1_REG2_REG_3__SCAN_IN), .A(n14440), .ZN(
        n14442) );
  OAI21_X1 U16158 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14445) );
  INV_X1 U16159 ( .A(n14445), .ZN(n14455) );
  NAND2_X1 U16160 ( .A1(n14447), .A2(n14446), .ZN(n14449) );
  NAND2_X1 U16161 ( .A1(n14449), .A2(n14448), .ZN(n14450) );
  NOR2_X1 U16162 ( .A1(n14451), .A2(n14450), .ZN(n14510) );
  AOI22_X1 U16163 ( .A1(n14453), .A2(n14513), .B1(n14452), .B2(n14510), .ZN(
        n14454) );
  OAI211_X1 U16164 ( .C1(n14441), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        P1_U3290) );
  INV_X1 U16165 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14457) );
  NOR2_X1 U16166 ( .A1(n14488), .A2(n14457), .ZN(P1_U3294) );
  INV_X1 U16167 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14458) );
  NOR2_X1 U16168 ( .A1(n14488), .A2(n14458), .ZN(P1_U3295) );
  INV_X1 U16169 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14459) );
  NOR2_X1 U16170 ( .A1(n14488), .A2(n14459), .ZN(P1_U3296) );
  INV_X1 U16171 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14460) );
  NOR2_X1 U16172 ( .A1(n14472), .A2(n14460), .ZN(P1_U3297) );
  INV_X1 U16173 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14461) );
  NOR2_X1 U16174 ( .A1(n14472), .A2(n14461), .ZN(P1_U3298) );
  INV_X1 U16175 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14462) );
  NOR2_X1 U16176 ( .A1(n14472), .A2(n14462), .ZN(P1_U3299) );
  INV_X1 U16177 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14463) );
  NOR2_X1 U16178 ( .A1(n14472), .A2(n14463), .ZN(P1_U3300) );
  INV_X1 U16179 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14464) );
  NOR2_X1 U16180 ( .A1(n14472), .A2(n14464), .ZN(P1_U3301) );
  INV_X1 U16181 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14465) );
  NOR2_X1 U16182 ( .A1(n14472), .A2(n14465), .ZN(P1_U3302) );
  INV_X1 U16183 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14466) );
  NOR2_X1 U16184 ( .A1(n14472), .A2(n14466), .ZN(P1_U3303) );
  INV_X1 U16185 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14467) );
  NOR2_X1 U16186 ( .A1(n14472), .A2(n14467), .ZN(P1_U3304) );
  INV_X1 U16187 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14468) );
  NOR2_X1 U16188 ( .A1(n14472), .A2(n14468), .ZN(P1_U3305) );
  INV_X1 U16189 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14469) );
  NOR2_X1 U16190 ( .A1(n14472), .A2(n14469), .ZN(P1_U3306) );
  INV_X1 U16191 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14470) );
  NOR2_X1 U16192 ( .A1(n14472), .A2(n14470), .ZN(P1_U3307) );
  INV_X1 U16193 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14471) );
  NOR2_X1 U16194 ( .A1(n14472), .A2(n14471), .ZN(P1_U3308) );
  INV_X1 U16195 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14473) );
  NOR2_X1 U16196 ( .A1(n14488), .A2(n14473), .ZN(P1_U3309) );
  INV_X1 U16197 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14474) );
  NOR2_X1 U16198 ( .A1(n14488), .A2(n14474), .ZN(P1_U3310) );
  INV_X1 U16199 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14475) );
  NOR2_X1 U16200 ( .A1(n14488), .A2(n14475), .ZN(P1_U3311) );
  INV_X1 U16201 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14476) );
  NOR2_X1 U16202 ( .A1(n14488), .A2(n14476), .ZN(P1_U3312) );
  INV_X1 U16203 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14477) );
  NOR2_X1 U16204 ( .A1(n14488), .A2(n14477), .ZN(P1_U3313) );
  INV_X1 U16205 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14478) );
  NOR2_X1 U16206 ( .A1(n14488), .A2(n14478), .ZN(P1_U3314) );
  INV_X1 U16207 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14479) );
  NOR2_X1 U16208 ( .A1(n14488), .A2(n14479), .ZN(P1_U3315) );
  INV_X1 U16209 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14480) );
  NOR2_X1 U16210 ( .A1(n14488), .A2(n14480), .ZN(P1_U3316) );
  INV_X1 U16211 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14481) );
  NOR2_X1 U16212 ( .A1(n14488), .A2(n14481), .ZN(P1_U3317) );
  INV_X1 U16213 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14482) );
  NOR2_X1 U16214 ( .A1(n14488), .A2(n14482), .ZN(P1_U3318) );
  INV_X1 U16215 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14483) );
  NOR2_X1 U16216 ( .A1(n14488), .A2(n14483), .ZN(P1_U3319) );
  INV_X1 U16217 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14484) );
  NOR2_X1 U16218 ( .A1(n14488), .A2(n14484), .ZN(P1_U3320) );
  INV_X1 U16219 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14485) );
  NOR2_X1 U16220 ( .A1(n14488), .A2(n14485), .ZN(P1_U3321) );
  INV_X1 U16221 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14486) );
  NOR2_X1 U16222 ( .A1(n14488), .A2(n14486), .ZN(P1_U3322) );
  INV_X1 U16223 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14487) );
  NOR2_X1 U16224 ( .A1(n14488), .A2(n14487), .ZN(P1_U3323) );
  AOI22_X1 U16225 ( .A1(n14578), .A2(n14489), .B1(n7843), .B2(n14576), .ZN(
        P1_U3459) );
  INV_X1 U16226 ( .A(n14498), .ZN(n14501) );
  NOR3_X1 U16227 ( .A1(n14491), .A2(n14566), .A3(n14490), .ZN(n14500) );
  OAI22_X1 U16228 ( .A1(n14493), .A2(n14492), .B1(n6620), .B2(n14570), .ZN(
        n14494) );
  INV_X1 U16229 ( .A(n14494), .ZN(n14495) );
  OAI211_X1 U16230 ( .C1(n14498), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14499) );
  AOI211_X1 U16231 ( .C1(n14564), .C2(n14501), .A(n14500), .B(n14499), .ZN(
        n14580) );
  AOI22_X1 U16232 ( .A1(n14578), .A2(n14580), .B1(n7829), .B2(n14576), .ZN(
        P1_U3462) );
  OAI21_X1 U16233 ( .B1(n14503), .B2(n14570), .A(n14502), .ZN(n14506) );
  INV_X1 U16234 ( .A(n14504), .ZN(n14505) );
  AOI211_X1 U16235 ( .C1(n14564), .C2(n14507), .A(n14506), .B(n14505), .ZN(
        n14582) );
  AOI22_X1 U16236 ( .A1(n14578), .A2(n14582), .B1(n7856), .B2(n14576), .ZN(
        P1_U3465) );
  OR4_X1 U16237 ( .A1(n14511), .A2(n14510), .A3(n14509), .A4(n14508), .ZN(
        n14512) );
  AOI21_X1 U16238 ( .B1(n14574), .B2(n14513), .A(n14512), .ZN(n14584) );
  AOI22_X1 U16239 ( .A1(n14578), .A2(n14584), .B1(n7877), .B2(n14576), .ZN(
        P1_U3468) );
  OAI211_X1 U16240 ( .C1(n14516), .C2(n14570), .A(n14515), .B(n14514), .ZN(
        n14520) );
  NOR2_X1 U16241 ( .A1(n14518), .A2(n14517), .ZN(n14519) );
  AOI211_X1 U16242 ( .C1(n14522), .C2(n14521), .A(n14520), .B(n14519), .ZN(
        n14585) );
  INV_X1 U16243 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14523) );
  AOI22_X1 U16244 ( .A1(n14578), .A2(n14585), .B1(n14523), .B2(n14576), .ZN(
        P1_U3471) );
  OR4_X1 U16245 ( .A1(n14527), .A2(n14526), .A3(n14525), .A4(n14524), .ZN(
        n14528) );
  AOI21_X1 U16246 ( .B1(n14574), .B2(n14529), .A(n14528), .ZN(n14586) );
  INV_X1 U16247 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U16248 ( .A1(n14578), .A2(n14586), .B1(n14530), .B2(n14576), .ZN(
        P1_U3474) );
  NAND2_X1 U16249 ( .A1(n14532), .A2(n14564), .ZN(n14538) );
  NAND2_X1 U16250 ( .A1(n14532), .A2(n14531), .ZN(n14537) );
  NAND2_X1 U16251 ( .A1(n14533), .A2(n14549), .ZN(n14534) );
  AND2_X1 U16252 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  INV_X1 U16253 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U16254 ( .A1(n14578), .A2(n14587), .B1(n14540), .B2(n14576), .ZN(
        P1_U3477) );
  OAI21_X1 U16255 ( .B1(n14542), .B2(n14570), .A(n14541), .ZN(n14545) );
  INV_X1 U16256 ( .A(n14543), .ZN(n14544) );
  AOI211_X1 U16257 ( .C1(n14564), .C2(n14546), .A(n14545), .B(n14544), .ZN(
        n14588) );
  INV_X1 U16258 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14547) );
  AOI22_X1 U16259 ( .A1(n14578), .A2(n14588), .B1(n14547), .B2(n14576), .ZN(
        P1_U3480) );
  AOI21_X1 U16260 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(n14552) );
  OAI211_X1 U16261 ( .C1(n14553), .C2(n14566), .A(n14552), .B(n14551), .ZN(
        n14554) );
  AOI21_X1 U16262 ( .B1(n14555), .B2(n14574), .A(n14554), .ZN(n14589) );
  INV_X1 U16263 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14556) );
  AOI22_X1 U16264 ( .A1(n14578), .A2(n14589), .B1(n14556), .B2(n14576), .ZN(
        P1_U3483) );
  INV_X1 U16265 ( .A(n14557), .ZN(n14559) );
  OAI21_X1 U16266 ( .B1(n14559), .B2(n14570), .A(n14558), .ZN(n14562) );
  INV_X1 U16267 ( .A(n14560), .ZN(n14561) );
  AOI211_X1 U16268 ( .C1(n14564), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14590) );
  INV_X1 U16269 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14565) );
  AOI22_X1 U16270 ( .A1(n14578), .A2(n14590), .B1(n14565), .B2(n14576), .ZN(
        P1_U3486) );
  NOR2_X1 U16271 ( .A1(n14567), .A2(n14566), .ZN(n14573) );
  OAI211_X1 U16272 ( .C1(n14571), .C2(n14570), .A(n14569), .B(n14568), .ZN(
        n14572) );
  AOI211_X1 U16273 ( .C1(n14575), .C2(n14574), .A(n14573), .B(n14572), .ZN(
        n14593) );
  INV_X1 U16274 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14577) );
  AOI22_X1 U16275 ( .A1(n14578), .A2(n14593), .B1(n14577), .B2(n14576), .ZN(
        P1_U3489) );
  AOI22_X1 U16276 ( .A1(n14594), .A2(n14580), .B1(n14579), .B2(n14591), .ZN(
        P1_U3529) );
  AOI22_X1 U16277 ( .A1(n14594), .A2(n14582), .B1(n14581), .B2(n14591), .ZN(
        P1_U3530) );
  AOI22_X1 U16278 ( .A1(n14594), .A2(n14584), .B1(n14583), .B2(n14591), .ZN(
        P1_U3531) );
  AOI22_X1 U16279 ( .A1(n14594), .A2(n14585), .B1(n7890), .B2(n14591), .ZN(
        P1_U3532) );
  AOI22_X1 U16280 ( .A1(n14594), .A2(n14586), .B1(n9908), .B2(n14591), .ZN(
        P1_U3533) );
  AOI22_X1 U16281 ( .A1(n14594), .A2(n14587), .B1(n9910), .B2(n14591), .ZN(
        P1_U3534) );
  AOI22_X1 U16282 ( .A1(n14594), .A2(n14588), .B1(n9912), .B2(n14591), .ZN(
        P1_U3535) );
  AOI22_X1 U16283 ( .A1(n14594), .A2(n14589), .B1(n7963), .B2(n14591), .ZN(
        P1_U3536) );
  AOI22_X1 U16284 ( .A1(n14594), .A2(n14590), .B1(n9957), .B2(n14591), .ZN(
        P1_U3537) );
  AOI22_X1 U16285 ( .A1(n14594), .A2(n14593), .B1(n14592), .B2(n14591), .ZN(
        P1_U3538) );
  NOR2_X1 U16286 ( .A1(n14652), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16287 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n14658), .B1(n14655), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n14598) );
  AOI22_X1 U16288 ( .A1(n14652), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14597) );
  OAI22_X1 U16289 ( .A1(n14670), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14668), .ZN(n14595) );
  OAI21_X1 U16290 ( .B1(n14673), .B2(n14595), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14596) );
  OAI211_X1 U16291 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14598), .A(n14597), .B(
        n14596), .ZN(P2_U3214) );
  INV_X1 U16292 ( .A(n14599), .ZN(n14614) );
  OAI21_X1 U16293 ( .B1(n14614), .B2(n14600), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14601) );
  OAI21_X1 U16294 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14601), .ZN(n14612) );
  AOI211_X1 U16295 ( .C1(n14604), .C2(n14603), .A(n14602), .B(n14670), .ZN(
        n14605) );
  INV_X1 U16296 ( .A(n14605), .ZN(n14611) );
  NAND2_X1 U16297 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14652), .ZN(n14610) );
  NOR2_X1 U16298 ( .A1(n6761), .A2(n8456), .ZN(n14608) );
  OAI211_X1 U16299 ( .C1(n14608), .C2(n14607), .A(n14658), .B(n14606), .ZN(
        n14609) );
  NAND4_X1 U16300 ( .A1(n14612), .A2(n14611), .A3(n14610), .A4(n14609), .ZN(
        P2_U3215) );
  OAI21_X1 U16301 ( .B1(n14614), .B2(n14613), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14615) );
  OAI21_X1 U16302 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14615), .ZN(n14626) );
  OAI211_X1 U16303 ( .C1(n14618), .C2(n14617), .A(n14658), .B(n14616), .ZN(
        n14625) );
  NAND2_X1 U16304 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n14652), .ZN(n14624) );
  AOI211_X1 U16305 ( .C1(n14621), .C2(n14620), .A(n14619), .B(n14670), .ZN(
        n14622) );
  INV_X1 U16306 ( .A(n14622), .ZN(n14623) );
  NAND4_X1 U16307 ( .A1(n14626), .A2(n14625), .A3(n14624), .A4(n14623), .ZN(
        P2_U3216) );
  NOR2_X1 U16308 ( .A1(n14644), .A2(n14627), .ZN(n14628) );
  AOI211_X1 U16309 ( .C1(n14652), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n14629), .B(
        n14628), .ZN(n14639) );
  AOI21_X1 U16310 ( .B1(n14631), .B2(n14630), .A(n14670), .ZN(n14633) );
  NAND2_X1 U16311 ( .A1(n14633), .A2(n14632), .ZN(n14638) );
  OAI211_X1 U16312 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14658), .ZN(
        n14637) );
  NAND3_X1 U16313 ( .A1(n14639), .A2(n14638), .A3(n14637), .ZN(P2_U3221) );
  XOR2_X1 U16314 ( .A(n14641), .B(n14640), .Z(n14646) );
  OAI21_X1 U16315 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(n14645) );
  AOI21_X1 U16316 ( .B1(n14646), .B2(n14658), .A(n14645), .ZN(n14650) );
  OAI211_X1 U16317 ( .C1(n14648), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14655), 
        .B(n14647), .ZN(n14649) );
  OAI211_X1 U16318 ( .C1(n14677), .C2(n14651), .A(n14650), .B(n14649), .ZN(
        P2_U3228) );
  AOI22_X1 U16319 ( .A1(n14652), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14663) );
  NAND2_X1 U16320 ( .A1(n14673), .A2(n14653), .ZN(n14662) );
  OAI211_X1 U16321 ( .C1(n14656), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14655), 
        .B(n14654), .ZN(n14661) );
  OAI211_X1 U16322 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14659), .A(n14658), 
        .B(n14657), .ZN(n14660) );
  NAND4_X1 U16323 ( .A1(n14663), .A2(n14662), .A3(n14661), .A4(n14660), .ZN(
        P2_U3229) );
  AOI21_X1 U16324 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14665), .A(n14664), 
        .ZN(n14671) );
  OAI21_X1 U16325 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n14667), .A(n14666), 
        .ZN(n14669) );
  OAI22_X1 U16326 ( .A1(n14671), .A2(n14670), .B1(n14669), .B2(n14668), .ZN(
        n14672) );
  AOI21_X1 U16327 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(n14676) );
  OAI211_X1 U16328 ( .C1(n14678), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        P2_U3232) );
  AND2_X1 U16329 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14680), .ZN(P2_U3266) );
  AND2_X1 U16330 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14680), .ZN(P2_U3267) );
  AND2_X1 U16331 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14680), .ZN(P2_U3268) );
  AND2_X1 U16332 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14680), .ZN(P2_U3269) );
  AND2_X1 U16333 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14680), .ZN(P2_U3270) );
  AND2_X1 U16334 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14680), .ZN(P2_U3271) );
  AND2_X1 U16335 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14680), .ZN(P2_U3272) );
  AND2_X1 U16336 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14680), .ZN(P2_U3273) );
  AND2_X1 U16337 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14680), .ZN(P2_U3274) );
  AND2_X1 U16338 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14680), .ZN(P2_U3275) );
  AND2_X1 U16339 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14680), .ZN(P2_U3276) );
  AND2_X1 U16340 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14680), .ZN(P2_U3277) );
  AND2_X1 U16341 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14680), .ZN(P2_U3278) );
  AND2_X1 U16342 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14680), .ZN(P2_U3279) );
  AND2_X1 U16343 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14680), .ZN(P2_U3280) );
  AND2_X1 U16344 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14680), .ZN(P2_U3281) );
  AND2_X1 U16345 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14680), .ZN(P2_U3282) );
  AND2_X1 U16346 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14680), .ZN(P2_U3283) );
  AND2_X1 U16347 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14680), .ZN(P2_U3284) );
  AND2_X1 U16348 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14680), .ZN(P2_U3285) );
  AND2_X1 U16349 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14680), .ZN(P2_U3286) );
  AND2_X1 U16350 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14680), .ZN(P2_U3287) );
  AND2_X1 U16351 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14680), .ZN(P2_U3288) );
  AND2_X1 U16352 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14680), .ZN(P2_U3289) );
  AND2_X1 U16353 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14680), .ZN(P2_U3290) );
  AND2_X1 U16354 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14680), .ZN(P2_U3291) );
  AND2_X1 U16355 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14680), .ZN(P2_U3292) );
  AND2_X1 U16356 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14680), .ZN(P2_U3293) );
  AND2_X1 U16357 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14680), .ZN(P2_U3294) );
  AND2_X1 U16358 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14680), .ZN(P2_U3295) );
  OAI21_X1 U16359 ( .B1(n14686), .B2(n14682), .A(n14681), .ZN(P2_U3416) );
  AOI22_X1 U16360 ( .A1(n14686), .A2(n14685), .B1(n14684), .B2(n14683), .ZN(
        P2_U3417) );
  INV_X1 U16361 ( .A(n14687), .ZN(n14690) );
  AOI211_X1 U16362 ( .C1(n14690), .C2(n14746), .A(n14689), .B(n14688), .ZN(
        n14757) );
  INV_X1 U16363 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14691) );
  AOI22_X1 U16364 ( .A1(n14756), .A2(n14757), .B1(n14691), .B2(n14755), .ZN(
        P2_U3430) );
  OAI21_X1 U16365 ( .B1(n14693), .B2(n14749), .A(n14692), .ZN(n14695) );
  AOI211_X1 U16366 ( .C1(n14746), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        n14758) );
  INV_X1 U16367 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14697) );
  AOI22_X1 U16368 ( .A1(n14756), .A2(n14758), .B1(n14697), .B2(n14755), .ZN(
        P2_U3436) );
  INV_X1 U16369 ( .A(n14698), .ZN(n14699) );
  OAI21_X1 U16370 ( .B1(n14700), .B2(n14749), .A(n14699), .ZN(n14702) );
  AOI211_X1 U16371 ( .C1(n14746), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14759) );
  INV_X1 U16372 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14704) );
  AOI22_X1 U16373 ( .A1(n14756), .A2(n14759), .B1(n14704), .B2(n14755), .ZN(
        P2_U3442) );
  INV_X1 U16374 ( .A(n14708), .ZN(n14712) );
  AOI21_X1 U16375 ( .B1(n14735), .B2(n14706), .A(n14705), .ZN(n14707) );
  OAI21_X1 U16376 ( .B1(n14708), .B2(n14739), .A(n14707), .ZN(n14711) );
  INV_X1 U16377 ( .A(n14709), .ZN(n14710) );
  AOI211_X1 U16378 ( .C1(n14745), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        n14761) );
  AOI22_X1 U16379 ( .A1(n14756), .A2(n14761), .B1(n8581), .B2(n14755), .ZN(
        P2_U3448) );
  AOI21_X1 U16380 ( .B1(n14735), .B2(n14714), .A(n14713), .ZN(n14715) );
  OAI211_X1 U16381 ( .C1(n14718), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        n14719) );
  INV_X1 U16382 ( .A(n14719), .ZN(n14762) );
  AOI22_X1 U16383 ( .A1(n14756), .A2(n14762), .B1(n8600), .B2(n14755), .ZN(
        P2_U3451) );
  OAI211_X1 U16384 ( .C1(n14722), .C2(n14749), .A(n14721), .B(n14720), .ZN(
        n14725) );
  AOI21_X1 U16385 ( .B1(n10245), .B2(n14739), .A(n14723), .ZN(n14724) );
  NOR2_X1 U16386 ( .A1(n14725), .A2(n14724), .ZN(n14763) );
  INV_X1 U16387 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14726) );
  AOI22_X1 U16388 ( .A1(n14756), .A2(n14763), .B1(n14726), .B2(n14755), .ZN(
        P2_U3454) );
  INV_X1 U16389 ( .A(n14730), .ZN(n14733) );
  NAND2_X1 U16390 ( .A1(n14727), .A2(n14735), .ZN(n14728) );
  OAI211_X1 U16391 ( .C1(n14730), .C2(n14739), .A(n14729), .B(n14728), .ZN(
        n14731) );
  AOI211_X1 U16392 ( .C1(n14745), .C2(n14733), .A(n14732), .B(n14731), .ZN(
        n14764) );
  INV_X1 U16393 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16394 ( .A1(n14756), .A2(n14764), .B1(n14734), .B2(n14755), .ZN(
        P2_U3457) );
  NAND2_X1 U16395 ( .A1(n14736), .A2(n14735), .ZN(n14737) );
  OAI211_X1 U16396 ( .C1(n14740), .C2(n14739), .A(n14738), .B(n14737), .ZN(
        n14743) );
  NOR2_X1 U16397 ( .A1(n14740), .A2(n10245), .ZN(n14742) );
  NOR3_X1 U16398 ( .A1(n14743), .A2(n14742), .A3(n14741), .ZN(n14765) );
  INV_X1 U16399 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U16400 ( .A1(n14756), .A2(n14765), .B1(n14744), .B2(n14755), .ZN(
        P2_U3460) );
  AND2_X1 U16401 ( .A1(n14747), .A2(n14745), .ZN(n14754) );
  AND2_X1 U16402 ( .A1(n14747), .A2(n14746), .ZN(n14753) );
  OAI21_X1 U16403 ( .B1(n14750), .B2(n14749), .A(n14748), .ZN(n14751) );
  NOR4_X1 U16404 ( .A1(n14754), .A2(n14753), .A3(n14752), .A4(n14751), .ZN(
        n14767) );
  AOI22_X1 U16405 ( .A1(n14756), .A2(n14767), .B1(n8676), .B2(n14755), .ZN(
        P2_U3463) );
  AOI22_X1 U16406 ( .A1(n14768), .A2(n14757), .B1(n8456), .B2(n14766), .ZN(
        P2_U3499) );
  AOI22_X1 U16407 ( .A1(n14768), .A2(n14758), .B1(n9778), .B2(n14766), .ZN(
        P2_U3501) );
  AOI22_X1 U16408 ( .A1(n14768), .A2(n14759), .B1(n8540), .B2(n14766), .ZN(
        P2_U3503) );
  AOI22_X1 U16409 ( .A1(n14768), .A2(n14761), .B1(n14760), .B2(n14766), .ZN(
        P2_U3505) );
  AOI22_X1 U16410 ( .A1(n14768), .A2(n14762), .B1(n9842), .B2(n14766), .ZN(
        P2_U3506) );
  AOI22_X1 U16411 ( .A1(n14768), .A2(n14763), .B1(n8620), .B2(n14766), .ZN(
        P2_U3507) );
  AOI22_X1 U16412 ( .A1(n14768), .A2(n14764), .B1(n8639), .B2(n14766), .ZN(
        P2_U3508) );
  AOI22_X1 U16413 ( .A1(n14768), .A2(n14765), .B1(n10133), .B2(n14766), .ZN(
        P2_U3509) );
  AOI22_X1 U16414 ( .A1(n14768), .A2(n14767), .B1(n8673), .B2(n14766), .ZN(
        P2_U3510) );
  NOR2_X1 U16415 ( .A1(P3_U3897), .A2(n14899), .ZN(P3_U3150) );
  NAND3_X1 U16416 ( .A1(n14921), .A2(n14769), .A3(n14915), .ZN(n14774) );
  OAI21_X1 U16417 ( .B1(n14772), .B2(n14771), .A(n14770), .ZN(n14773) );
  NAND2_X1 U16418 ( .A1(n14774), .A2(n14773), .ZN(n14779) );
  OAI22_X1 U16419 ( .A1(n14896), .A2(n14776), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14775), .ZN(n14777) );
  INV_X1 U16420 ( .A(n14777), .ZN(n14778) );
  OAI211_X1 U16421 ( .C1(n14780), .C2(n14930), .A(n14779), .B(n14778), .ZN(
        P3_U3182) );
  INV_X1 U16422 ( .A(n14781), .ZN(n14782) );
  NAND2_X1 U16423 ( .A1(n14782), .A2(n11167), .ZN(n14783) );
  AND2_X1 U16424 ( .A1(n14784), .A2(n14783), .ZN(n14798) );
  AOI21_X1 U16425 ( .B1(n14899), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n14785), .ZN(
        n14791) );
  AND3_X1 U16426 ( .A1(n14788), .A2(n14787), .A3(n14786), .ZN(n14789) );
  OAI21_X1 U16427 ( .B1(n14803), .B2(n14789), .A(n14892), .ZN(n14790) );
  OAI211_X1 U16428 ( .C1(n14896), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14793) );
  INV_X1 U16429 ( .A(n14793), .ZN(n14797) );
  XNOR2_X1 U16430 ( .A(n14794), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14795) );
  NAND2_X1 U16431 ( .A1(n14910), .A2(n14795), .ZN(n14796) );
  OAI211_X1 U16432 ( .C1(n14798), .C2(n14921), .A(n14797), .B(n14796), .ZN(
        P3_U3185) );
  AOI21_X1 U16433 ( .B1(n14800), .B2(n14799), .A(n6611), .ZN(n14816) );
  INV_X1 U16434 ( .A(n14821), .ZN(n14805) );
  NOR3_X1 U16435 ( .A1(n14803), .A2(n14802), .A3(n14801), .ZN(n14804) );
  OAI21_X1 U16436 ( .B1(n14805), .B2(n14804), .A(n14892), .ZN(n14806) );
  OAI21_X1 U16437 ( .B1(n14896), .B2(n14807), .A(n14806), .ZN(n14808) );
  AOI211_X1 U16438 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14899), .A(n14809), .B(
        n14808), .ZN(n14815) );
  OAI21_X1 U16439 ( .B1(n14812), .B2(n14811), .A(n14810), .ZN(n14813) );
  NAND2_X1 U16440 ( .A1(n14910), .A2(n14813), .ZN(n14814) );
  OAI211_X1 U16441 ( .C1(n14816), .C2(n14921), .A(n14815), .B(n14814), .ZN(
        P3_U3186) );
  AOI21_X1 U16442 ( .B1(n11180), .B2(n14818), .A(n14817), .ZN(n14832) );
  AND3_X1 U16443 ( .A1(n14821), .A2(n14820), .A3(n14819), .ZN(n14822) );
  OAI21_X1 U16444 ( .B1(n14838), .B2(n14822), .A(n14892), .ZN(n14823) );
  OAI21_X1 U16445 ( .B1(n14896), .B2(n14824), .A(n14823), .ZN(n14825) );
  AOI211_X1 U16446 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14899), .A(n14826), .B(
        n14825), .ZN(n14831) );
  OAI21_X1 U16447 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14828), .A(n14827), .ZN(
        n14829) );
  NAND2_X1 U16448 ( .A1(n14910), .A2(n14829), .ZN(n14830) );
  OAI211_X1 U16449 ( .C1(n14832), .C2(n14921), .A(n14831), .B(n14830), .ZN(
        P3_U3187) );
  AOI21_X1 U16450 ( .B1(n14835), .B2(n14834), .A(n14833), .ZN(n14851) );
  INV_X1 U16451 ( .A(n14856), .ZN(n14840) );
  NOR3_X1 U16452 ( .A1(n14838), .A2(n14837), .A3(n14836), .ZN(n14839) );
  OAI21_X1 U16453 ( .B1(n14840), .B2(n14839), .A(n14892), .ZN(n14841) );
  OAI21_X1 U16454 ( .B1(n14896), .B2(n14842), .A(n14841), .ZN(n14843) );
  AOI211_X1 U16455 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14899), .A(n14844), .B(
        n14843), .ZN(n14850) );
  OAI21_X1 U16456 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(n14848) );
  NAND2_X1 U16457 ( .A1(n14848), .A2(n14910), .ZN(n14849) );
  OAI211_X1 U16458 ( .C1(n14851), .C2(n14921), .A(n14850), .B(n14849), .ZN(
        P3_U3188) );
  AOI21_X1 U16459 ( .B1(n14958), .B2(n14853), .A(n14852), .ZN(n14867) );
  AND3_X1 U16460 ( .A1(n14856), .A2(n14855), .A3(n14854), .ZN(n14857) );
  OAI21_X1 U16461 ( .B1(n14872), .B2(n14857), .A(n14892), .ZN(n14858) );
  OAI21_X1 U16462 ( .B1(n14896), .B2(n14859), .A(n14858), .ZN(n14860) );
  AOI211_X1 U16463 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14899), .A(n14861), .B(
        n14860), .ZN(n14866) );
  OAI21_X1 U16464 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14863), .A(n14862), .ZN(
        n14864) );
  NAND2_X1 U16465 ( .A1(n14864), .A2(n14910), .ZN(n14865) );
  OAI211_X1 U16466 ( .C1(n14867), .C2(n14921), .A(n14866), .B(n14865), .ZN(
        P3_U3189) );
  AOI21_X1 U16467 ( .B1(n6608), .B2(n14869), .A(n14868), .ZN(n14885) );
  INV_X1 U16468 ( .A(n14891), .ZN(n14874) );
  NOR3_X1 U16469 ( .A1(n14872), .A2(n14871), .A3(n14870), .ZN(n14873) );
  OAI21_X1 U16470 ( .B1(n14874), .B2(n14873), .A(n14892), .ZN(n14875) );
  OAI21_X1 U16471 ( .B1(n14896), .B2(n14876), .A(n14875), .ZN(n14877) );
  AOI211_X1 U16472 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14899), .A(n14878), .B(
        n14877), .ZN(n14884) );
  OAI21_X1 U16473 ( .B1(n14881), .B2(n14880), .A(n14879), .ZN(n14882) );
  NAND2_X1 U16474 ( .A1(n14882), .A2(n14910), .ZN(n14883) );
  OAI211_X1 U16475 ( .C1(n14885), .C2(n14921), .A(n14884), .B(n14883), .ZN(
        P3_U3190) );
  AOI21_X1 U16476 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n14905) );
  AND3_X1 U16477 ( .A1(n14891), .A2(n14890), .A3(n14889), .ZN(n14893) );
  OAI21_X1 U16478 ( .B1(n14914), .B2(n14893), .A(n14892), .ZN(n14894) );
  OAI21_X1 U16479 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  AOI211_X1 U16480 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14899), .A(n14898), .B(
        n14897), .ZN(n14904) );
  OAI21_X1 U16481 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14901), .A(n14900), .ZN(
        n14902) );
  NAND2_X1 U16482 ( .A1(n14902), .A2(n14910), .ZN(n14903) );
  OAI211_X1 U16483 ( .C1(n14905), .C2(n14921), .A(n14904), .B(n14903), .ZN(
        P3_U3191) );
  OAI21_X1 U16484 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n14911) );
  AOI21_X1 U16485 ( .B1(n14911), .B2(n14910), .A(n14909), .ZN(n14928) );
  OR3_X1 U16486 ( .A1(n14914), .A2(n14913), .A3(n14912), .ZN(n14916) );
  AOI21_X1 U16487 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n14924) );
  AOI21_X1 U16488 ( .B1(n14920), .B2(n14919), .A(n14918), .ZN(n14922) );
  NOR2_X1 U16489 ( .A1(n14922), .A2(n14921), .ZN(n14923) );
  AOI211_X1 U16490 ( .C1(n14926), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        n14927) );
  OAI211_X1 U16491 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        P3_U3192) );
  XNOR2_X1 U16492 ( .A(n14931), .B(n14933), .ZN(n15062) );
  OAI211_X1 U16493 ( .C1(n14934), .C2(n14933), .A(n14932), .B(n15001), .ZN(
        n14938) );
  AOI22_X1 U16494 ( .A1(n14962), .A2(n14936), .B1(n14935), .B2(n14965), .ZN(
        n14937) );
  NAND2_X1 U16495 ( .A1(n14938), .A2(n14937), .ZN(n15060) );
  AOI21_X1 U16496 ( .B1(n14953), .B2(n15062), .A(n15060), .ZN(n14943) );
  INV_X1 U16497 ( .A(n14939), .ZN(n14972) );
  NOR2_X1 U16498 ( .A1(n14940), .A2(n15047), .ZN(n15061) );
  AOI22_X1 U16499 ( .A1(n14972), .A2(n15061), .B1(n15007), .B2(n14941), .ZN(
        n14942) );
  OAI221_X1 U16500 ( .B1(n15012), .B2(n14943), .C1(n15010), .C2(n11211), .A(
        n14942), .ZN(P3_U3223) );
  XNOR2_X1 U16501 ( .A(n14945), .B(n14944), .ZN(n15045) );
  OAI211_X1 U16502 ( .C1(n14948), .C2(n14947), .A(n14946), .B(n15001), .ZN(
        n14952) );
  AOI22_X1 U16503 ( .A1(n14962), .A2(n14950), .B1(n14949), .B2(n14965), .ZN(
        n14951) );
  NAND2_X1 U16504 ( .A1(n14952), .A2(n14951), .ZN(n15043) );
  AOI21_X1 U16505 ( .B1(n15045), .B2(n14953), .A(n15043), .ZN(n14959) );
  NOR2_X1 U16506 ( .A1(n14954), .A2(n15047), .ZN(n15044) );
  INV_X1 U16507 ( .A(n14955), .ZN(n14956) );
  AOI22_X1 U16508 ( .A1(n14972), .A2(n15044), .B1(n15007), .B2(n14956), .ZN(
        n14957) );
  OAI221_X1 U16509 ( .B1(n15012), .B2(n14959), .C1(n15010), .C2(n14958), .A(
        n14957), .ZN(P3_U3226) );
  XNOR2_X1 U16510 ( .A(n14961), .B(n9154), .ZN(n14969) );
  INV_X1 U16511 ( .A(n14969), .ZN(n15027) );
  AOI22_X1 U16512 ( .A1(n14965), .A2(n14964), .B1(n14963), .B2(n14962), .ZN(
        n14968) );
  OAI211_X1 U16513 ( .C1(n6509), .C2(n9154), .A(n15001), .B(n14966), .ZN(
        n14967) );
  OAI211_X1 U16514 ( .C1(n14969), .C2(n15004), .A(n14968), .B(n14967), .ZN(
        n15025) );
  AOI21_X1 U16515 ( .B1(n14990), .B2(n15027), .A(n15025), .ZN(n14974) );
  AND2_X1 U16516 ( .A1(n14970), .A2(n15015), .ZN(n15026) );
  NOR2_X1 U16517 ( .A1(n14978), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n14971) );
  AOI21_X1 U16518 ( .B1(n14972), .B2(n15026), .A(n14971), .ZN(n14973) );
  OAI221_X1 U16519 ( .B1(n15012), .B2(n14974), .C1(n15010), .C2(n11167), .A(
        n14973), .ZN(P3_U3230) );
  OAI21_X1 U16520 ( .B1(n6970), .B2(n14982), .A(n14976), .ZN(n15023) );
  NOR2_X1 U16521 ( .A1(n14977), .A2(n15047), .ZN(n15022) );
  INV_X1 U16522 ( .A(n15022), .ZN(n14980) );
  OAI22_X1 U16523 ( .A1(n14980), .A2(n14979), .B1(n7575), .B2(n14978), .ZN(
        n14989) );
  XNOR2_X1 U16524 ( .A(n14981), .B(n14982), .ZN(n14987) );
  OAI22_X1 U16525 ( .A1(n9118), .A2(n14998), .B1(n14983), .B2(n14996), .ZN(
        n14984) );
  AOI21_X1 U16526 ( .B1(n15023), .B2(n14985), .A(n14984), .ZN(n14986) );
  OAI21_X1 U16527 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n15021) );
  AOI211_X1 U16528 ( .C1(n14990), .C2(n15023), .A(n14989), .B(n15021), .ZN(
        n14991) );
  AOI22_X1 U16529 ( .A1(n15012), .A2(n10046), .B1(n14991), .B2(n15010), .ZN(
        P3_U3231) );
  NOR2_X1 U16530 ( .A1(n14992), .A2(n15047), .ZN(n15018) );
  XNOR2_X1 U16531 ( .A(n14994), .B(n14993), .ZN(n15006) );
  XNOR2_X1 U16532 ( .A(n14995), .B(n10119), .ZN(n15002) );
  OAI22_X1 U16533 ( .A1(n14999), .A2(n14998), .B1(n14997), .B2(n14996), .ZN(
        n15000) );
  AOI21_X1 U16534 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15003) );
  OAI21_X1 U16535 ( .B1(n15006), .B2(n15004), .A(n15003), .ZN(n15017) );
  AOI21_X1 U16536 ( .B1(n15018), .B2(n15005), .A(n15017), .ZN(n15011) );
  INV_X1 U16537 ( .A(n15006), .ZN(n15019) );
  AOI22_X1 U16538 ( .A1(n15008), .A2(n15019), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15007), .ZN(n15009) );
  OAI221_X1 U16539 ( .B1(n15012), .B2(n15011), .C1(n15010), .C2(n10020), .A(
        n15009), .ZN(P3_U3232) );
  AOI21_X1 U16540 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15067) );
  INV_X1 U16541 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U16542 ( .A1(n15066), .A2(n15067), .B1(n15016), .B2(n15064), .ZN(
        P3_U3390) );
  AOI211_X1 U16543 ( .C1(n15058), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        n15068) );
  INV_X1 U16544 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16545 ( .A1(n15066), .A2(n15068), .B1(n15020), .B2(n15064), .ZN(
        P3_U3393) );
  AOI211_X1 U16546 ( .C1(n15058), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15069) );
  INV_X1 U16547 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U16548 ( .A1(n15066), .A2(n15069), .B1(n15024), .B2(n15064), .ZN(
        P3_U3396) );
  AOI211_X1 U16549 ( .C1(n15027), .C2(n15058), .A(n15026), .B(n15025), .ZN(
        n15070) );
  AOI22_X1 U16550 ( .A1(n15066), .A2(n15070), .B1(n9138), .B2(n15064), .ZN(
        P3_U3399) );
  INV_X1 U16551 ( .A(n15028), .ZN(n15030) );
  AOI211_X1 U16552 ( .C1(n15031), .C2(n15058), .A(n15030), .B(n15029), .ZN(
        n15071) );
  INV_X1 U16553 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15032) );
  AOI22_X1 U16554 ( .A1(n15066), .A2(n15071), .B1(n15032), .B2(n15064), .ZN(
        P3_U3402) );
  INV_X1 U16555 ( .A(n15033), .ZN(n15036) );
  AOI211_X1 U16556 ( .C1(n15036), .C2(n15058), .A(n15035), .B(n15034), .ZN(
        n15072) );
  INV_X1 U16557 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15037) );
  AOI22_X1 U16558 ( .A1(n15066), .A2(n15072), .B1(n15037), .B2(n15064), .ZN(
        P3_U3405) );
  INV_X1 U16559 ( .A(n15038), .ZN(n15040) );
  AOI211_X1 U16560 ( .C1(n15041), .C2(n15058), .A(n15040), .B(n15039), .ZN(
        n15073) );
  INV_X1 U16561 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15042) );
  AOI22_X1 U16562 ( .A1(n15066), .A2(n15073), .B1(n15042), .B2(n15064), .ZN(
        P3_U3408) );
  AOI211_X1 U16563 ( .C1(n15045), .C2(n15063), .A(n15044), .B(n15043), .ZN(
        n15074) );
  INV_X1 U16564 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15046) );
  AOI22_X1 U16565 ( .A1(n15066), .A2(n15074), .B1(n15046), .B2(n15064), .ZN(
        P3_U3411) );
  OAI22_X1 U16566 ( .A1(n15050), .A2(n15049), .B1(n15048), .B2(n15047), .ZN(
        n15051) );
  NOR2_X1 U16567 ( .A1(n15052), .A2(n15051), .ZN(n15075) );
  INV_X1 U16568 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15053) );
  AOI22_X1 U16569 ( .A1(n15066), .A2(n15075), .B1(n15053), .B2(n15064), .ZN(
        P3_U3414) );
  INV_X1 U16570 ( .A(n15054), .ZN(n15057) );
  AOI211_X1 U16571 ( .C1(n15058), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15076) );
  INV_X1 U16572 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U16573 ( .A1(n15066), .A2(n15076), .B1(n15059), .B2(n15064), .ZN(
        P3_U3417) );
  AOI211_X1 U16574 ( .C1(n15063), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15078) );
  INV_X1 U16575 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15065) );
  AOI22_X1 U16576 ( .A1(n15066), .A2(n15078), .B1(n15065), .B2(n15064), .ZN(
        P3_U3420) );
  AOI22_X1 U16577 ( .A1(n15079), .A2(n15067), .B1(n10019), .B2(n15077), .ZN(
        P3_U3459) );
  AOI22_X1 U16578 ( .A1(n15079), .A2(n15068), .B1(n10031), .B2(n15077), .ZN(
        P3_U3460) );
  AOI22_X1 U16579 ( .A1(n15079), .A2(n15069), .B1(n10045), .B2(n15077), .ZN(
        P3_U3461) );
  AOI22_X1 U16580 ( .A1(n15079), .A2(n15070), .B1(n11166), .B2(n15077), .ZN(
        P3_U3462) );
  AOI22_X1 U16581 ( .A1(n15079), .A2(n15071), .B1(n11173), .B2(n15077), .ZN(
        P3_U3463) );
  AOI22_X1 U16582 ( .A1(n15079), .A2(n15072), .B1(n11179), .B2(n15077), .ZN(
        P3_U3464) );
  AOI22_X1 U16583 ( .A1(n15079), .A2(n15073), .B1(n11186), .B2(n15077), .ZN(
        P3_U3465) );
  AOI22_X1 U16584 ( .A1(n15079), .A2(n15074), .B1(n11192), .B2(n15077), .ZN(
        P3_U3466) );
  AOI22_X1 U16585 ( .A1(n15079), .A2(n15075), .B1(n11198), .B2(n15077), .ZN(
        P3_U3467) );
  AOI22_X1 U16586 ( .A1(n15079), .A2(n15076), .B1(n11204), .B2(n15077), .ZN(
        P3_U3468) );
  AOI22_X1 U16587 ( .A1(n15079), .A2(n15078), .B1(n11210), .B2(n15077), .ZN(
        P3_U3469) );
  XOR2_X1 U16588 ( .A(n15081), .B(n15080), .Z(SUB_1596_U59) );
  XNOR2_X1 U16589 ( .A(n15082), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16590 ( .B1(n15084), .B2(n15083), .A(n15091), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16591 ( .A(n15086), .B(n15085), .ZN(SUB_1596_U56) );
  NOR2_X1 U16592 ( .A1(n15088), .A2(n15087), .ZN(n15089) );
  XOR2_X1 U16593 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15089), .Z(SUB_1596_U60) );
  XOR2_X1 U16594 ( .A(n15091), .B(n15090), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7229 ( .A(n8935), .Z(n6478) );
  INV_X1 U7221 ( .A(n12540), .ZN(n9610) );
  BUF_X2 U7226 ( .A(n7837), .Z(n8372) );
  CLKBUF_X1 U7230 ( .A(n10807), .Z(n12130) );
  CLKBUF_X2 U7237 ( .A(n8568), .Z(n6489) );
  CLKBUF_X1 U7240 ( .A(n8935), .Z(n6479) );
  NAND4_X1 U7244 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n14354)
         );
  CLKBUF_X1 U7253 ( .A(n11346), .Z(n6472) );
endmodule

