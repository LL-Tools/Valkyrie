

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209;

  CLKBUF_X2 U34610 ( .A(n3621), .Z(n4319) );
  NAND2_X1 U34620 ( .A1(n3699), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3726) );
  CLKBUF_X2 U34630 ( .A(n4740), .Z(n5896) );
  CLKBUF_X1 U34640 ( .A(n4274), .Z(n4299) );
  NOR2_X2 U34650 ( .A1(n5503), .A2(n3687), .ZN(n3712) );
  AND2_X1 U3466 ( .A1(n6613), .A2(n3567), .ZN(n3755) );
  AND2_X2 U3467 ( .A1(n3469), .A2(n3567), .ZN(n4274) );
  AND2_X1 U34680 ( .A1(n3567), .A2(n4738), .ZN(n3744) );
  CLKBUF_X1 U34690 ( .A(n5559), .Z(n3427) );
  AND2_X1 U34700 ( .A1(n3845), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4746) );
  AND2_X1 U34710 ( .A1(n6613), .A2(n4895), .ZN(n3643) );
  INV_X1 U34720 ( .A(n4624), .ZN(n4630) );
  AND2_X1 U34730 ( .A1(n4645), .A2(n4642), .ZN(n4709) );
  AND2_X1 U34740 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4895) );
  BUF_X1 U3475 ( .A(n4483), .Z(n6594) );
  NAND2_X1 U3476 ( .A1(n3687), .A2(n3713), .ZN(n4624) );
  OAI21_X1 U3477 ( .B1(n4673), .B2(n4530), .A(n4529), .ZN(n4645) );
  NAND2_X1 U3478 ( .A1(n6948), .A2(n5489), .ZN(n7014) );
  INV_X1 U3479 ( .A(n7017), .ZN(n7060) );
  NOR2_X1 U3481 ( .A1(n4487), .A2(n4488), .ZN(n6390) );
  NOR2_X2 U3482 ( .A1(n6850), .A2(n4649), .ZN(n6901) );
  AND2_X2 U3483 ( .A1(n3468), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3469)
         );
  OAI21_X2 U3484 ( .B1(n3726), .B2(n3561), .A(n3704), .ZN(n3768) );
  AND2_X2 U3485 ( .A1(n4910), .A2(n3865), .ZN(n4861) );
  CLKBUF_X2 U3486 ( .A(n7190), .Z(n7193) );
  NOR2_X1 U3487 ( .A1(n5012), .A2(n4870), .ZN(n5687) );
  CLKBUF_X2 U3488 ( .A(n3712), .Z(n7144) );
  AND4_X2 U3489 ( .A1(n3560), .A2(n3552), .A3(n3590), .A4(n3550), .ZN(n3635)
         );
  BUF_X2 U3490 ( .A(n3641), .Z(n3738) );
  CLKBUF_X2 U3491 ( .A(n4055), .Z(n4318) );
  BUF_X2 U3492 ( .A(n3653), .Z(n5897) );
  BUF_X2 U3493 ( .A(n3743), .Z(n5869) );
  CLKBUF_X2 U3494 ( .A(n3626), .Z(n5875) );
  CLKBUF_X2 U3495 ( .A(n5890), .Z(n4189) );
  BUF_X2 U3496 ( .A(n4146), .Z(n4190) );
  CLKBUF_X2 U3497 ( .A(n3658), .Z(n5876) );
  CLKBUF_X2 U3498 ( .A(n3744), .Z(n4191) );
  BUF_X2 U3499 ( .A(n3643), .Z(n5870) );
  CLKBUF_X2 U3500 ( .A(n3755), .Z(n5891) );
  NAND3_X1 U3501 ( .A1(n3516), .A2(n6505), .A3(n3515), .ZN(n5958) );
  NAND2_X1 U3502 ( .A1(n3517), .A2(n3519), .ZN(n3516) );
  AOI21_X1 U3503 ( .B1(n3488), .B2(n7057), .A(n3486), .ZN(n3485) );
  XNOR2_X1 U3504 ( .A(n3441), .B(n5918), .ZN(n6166) );
  OR2_X1 U3505 ( .A1(n6012), .A2(n3511), .ZN(n5986) );
  OAI21_X1 U3506 ( .B1(n4476), .B2(n3463), .A(n3461), .ZN(n3465) );
  NAND2_X1 U3507 ( .A1(n3497), .A2(n3496), .ZN(n5742) );
  AOI21_X1 U3508 ( .B1(n3532), .B2(n3530), .A(n3529), .ZN(n3528) );
  NOR2_X1 U3509 ( .A1(n3537), .A2(n3462), .ZN(n3461) );
  NOR2_X1 U3510 ( .A1(n3436), .A2(n3463), .ZN(n3462) );
  NOR2_X1 U3511 ( .A1(n6463), .A2(n4478), .ZN(n4479) );
  INV_X2 U3512 ( .A(n5957), .ZN(n6428) );
  INV_X1 U3513 ( .A(n5957), .ZN(n6463) );
  OAI21_X1 U3514 ( .B1(n4408), .B2(n4458), .A(n4407), .ZN(n4447) );
  NAND2_X1 U3515 ( .A1(n4401), .A2(n4437), .ZN(n4450) );
  NAND2_X1 U3516 ( .A1(n3875), .A2(n3874), .ZN(n4794) );
  AND2_X1 U3517 ( .A1(n3895), .A2(n4911), .ZN(n3866) );
  XNOR2_X1 U3518 ( .A(n3895), .B(n3896), .ZN(n4438) );
  INV_X1 U3519 ( .A(n3432), .ZN(n3865) );
  NAND2_X1 U3520 ( .A1(n3836), .A2(n3775), .ZN(n4910) );
  INV_X1 U3521 ( .A(n4806), .ZN(n6848) );
  INV_X2 U3523 ( .A(n7145), .ZN(n7185) );
  NAND2_X1 U3524 ( .A1(n3827), .A2(n7115), .ZN(n3818) );
  AND2_X1 U3525 ( .A1(n3634), .A2(n3633), .ZN(n4514) );
  NAND2_X1 U3526 ( .A1(n3673), .A2(n3672), .ZN(n4502) );
  NAND2_X1 U3527 ( .A1(n3813), .A2(n3772), .ZN(n4387) );
  CLKBUF_X1 U3528 ( .A(n3713), .Z(n4501) );
  INV_X1 U3529 ( .A(n3635), .ZN(n3466) );
  INV_X1 U3530 ( .A(n3635), .ZN(n3737) );
  CLKBUF_X1 U3531 ( .A(n3636), .Z(n4525) );
  NAND2_X1 U3532 ( .A1(n3609), .A2(n3442), .ZN(n3636) );
  OR2_X2 U3533 ( .A1(n3632), .A2(n3631), .ZN(n3713) );
  AND4_X1 U3534 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3609)
         );
  AND4_X1 U3535 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3619)
         );
  AND4_X1 U3536 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .ZN(n3667)
         );
  AND4_X1 U3537 ( .A1(n3589), .A2(n3588), .A3(n3587), .A4(n3586), .ZN(n3550)
         );
  AND4_X1 U3538 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3620)
         );
  AND4_X1 U3539 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3600)
         );
  CLKBUF_X3 U3540 ( .A(n3642), .Z(n4320) );
  AND2_X2 U3541 ( .A1(n4744), .A2(n3566), .ZN(n3653) );
  AND2_X2 U3542 ( .A1(n4746), .A2(n4738), .ZN(n4740) );
  AND2_X1 U3543 ( .A1(n3727), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4744)
         );
  AND2_X2 U3545 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4738) );
  NOR2_X2 U3546 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6613) );
  NOR2_X2 U3547 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3567) );
  CLKBUF_X1 U3548 ( .A(n5464), .Z(n3428) );
  CLKBUF_X1 U3549 ( .A(n4531), .Z(n3429) );
  INV_X1 U3550 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3430) );
  OAI21_X1 U3551 ( .B1(n4770), .B2(STATE2_REG_0__SCAN_IN), .A(n3751), .ZN(
        n3431) );
  NAND2_X1 U3552 ( .A1(n3671), .A2(n4515), .ZN(n4531) );
  OAI21_X1 U3553 ( .B1(n4770), .B2(STATE2_REG_0__SCAN_IN), .A(n3751), .ZN(
        n3777) );
  NAND2_X2 U3554 ( .A1(n3459), .A2(n4474), .ZN(n5598) );
  NAND2_X2 U3555 ( .A1(n5559), .A2(n5560), .ZN(n3459) );
  AND2_X1 U3556 ( .A1(n3561), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3566)
         );
  NOR2_X2 U3557 ( .A1(n3489), .A2(n4717), .ZN(n4815) );
  AND2_X1 U3558 ( .A1(n3610), .A2(n3675), .ZN(n3467) );
  NAND2_X2 U3559 ( .A1(n4482), .A2(n3458), .ZN(n6441) );
  OR2_X1 U3560 ( .A1(n5012), .A2(n3675), .ZN(n5655) );
  INV_X1 U3561 ( .A(n5655), .ZN(n3433) );
  OR2_X1 U3562 ( .A1(n5012), .A2(n3679), .ZN(n5634) );
  INV_X1 U3563 ( .A(n5634), .ZN(n3434) );
  OR2_X1 U3564 ( .A1(n5012), .A2(n3635), .ZN(n5641) );
  INV_X1 U3565 ( .A(n5641), .ZN(n3435) );
  INV_X1 U3566 ( .A(n6614), .ZN(n4512) );
  OR2_X1 U3567 ( .A1(n4501), .A2(n5503), .ZN(n4622) );
  AND2_X1 U3568 ( .A1(n6948), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5935) );
  NOR2_X2 U3569 ( .A1(n4880), .A2(n5503), .ZN(n5494) );
  AND2_X1 U3570 ( .A1(n3610), .A2(n3713), .ZN(n3693) );
  NAND2_X1 U3571 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  OR2_X1 U3572 ( .A1(n4640), .A2(n4513), .ZN(n4516) );
  NAND2_X1 U3573 ( .A1(n4338), .A2(n3512), .ZN(n3511) );
  INV_X1 U3574 ( .A(n5997), .ZN(n3512) );
  NAND2_X1 U3575 ( .A1(n3465), .A2(n3535), .ZN(n4481) );
  AOI21_X1 U3576 ( .B1(n3540), .B2(n3536), .A(n4479), .ZN(n3535) );
  OR2_X1 U3577 ( .A1(n5980), .A2(n7120), .ZN(n4673) );
  NAND2_X1 U3578 ( .A1(n3467), .A2(n3466), .ZN(n4070) );
  NAND2_X1 U3579 ( .A1(n4757), .A2(n4756), .ZN(n5476) );
  INV_X1 U3580 ( .A(n4673), .ZN(n5475) );
  NOR2_X1 U3581 ( .A1(n3511), .A2(n5987), .ZN(n3510) );
  OR2_X1 U3582 ( .A1(n4270), .A2(n6415), .ZN(n4312) );
  AND2_X1 U3583 ( .A1(n3505), .A2(n6024), .ZN(n3504) );
  INV_X1 U3584 ( .A(n5494), .ZN(n4633) );
  OAI21_X1 U3585 ( .B1(n5989), .B2(n4631), .A(n4630), .ZN(n5944) );
  OR2_X1 U3586 ( .A1(n6463), .A2(n6542), .ZN(n4485) );
  CLKBUF_X1 U3587 ( .A(n4497), .Z(n4498) );
  AND4_X1 U3588 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3670)
         );
  AND4_X1 U3589 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3668)
         );
  AND4_X1 U3590 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3669)
         );
  BUF_X1 U3591 ( .A(n4343), .Z(n4880) );
  OR2_X1 U3592 ( .A1(n6798), .A2(n5484), .ZN(n6948) );
  NAND2_X1 U3593 ( .A1(n4369), .A2(n4368), .ZN(n4376) );
  INV_X1 U3594 ( .A(n4409), .ZN(n3771) );
  NAND2_X1 U3595 ( .A1(n3938), .A2(n3553), .ZN(n4401) );
  INV_X1 U3596 ( .A(n6485), .ZN(n3538) );
  NOR2_X1 U3597 ( .A1(n6065), .A2(n3507), .ZN(n3506) );
  INV_X1 U3598 ( .A(n6130), .ZN(n3507) );
  AND2_X1 U3599 ( .A1(n3452), .A2(n6152), .ZN(n3498) );
  INV_X1 U3600 ( .A(n5770), .ZN(n3544) );
  INV_X1 U3601 ( .A(n5573), .ZN(n3497) );
  NAND2_X1 U3602 ( .A1(n3495), .A2(n4081), .ZN(n3788) );
  OR2_X1 U3603 ( .A1(n3477), .A2(n3479), .ZN(n3476) );
  NAND2_X1 U3604 ( .A1(n3478), .A2(n6015), .ZN(n3477) );
  INV_X1 U3605 ( .A(n6041), .ZN(n3478) );
  INV_X1 U3606 ( .A(n6421), .ZN(n4484) );
  INV_X1 U3607 ( .A(n6132), .ZN(n3472) );
  INV_X1 U3608 ( .A(n4607), .ZN(n4626) );
  AND2_X1 U3609 ( .A1(n5494), .A2(n4630), .ZN(n4607) );
  NAND2_X1 U3610 ( .A1(n3432), .A2(n3864), .ZN(n3895) );
  AND2_X1 U3611 ( .A1(n3731), .A2(n3730), .ZN(n3734) );
  OR2_X1 U3612 ( .A1(n3726), .A2(n3727), .ZN(n3731) );
  NAND2_X1 U3613 ( .A1(n3835), .A2(n3834), .ZN(n3525) );
  AOI22_X1 U3614 ( .A1(n4274), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3570) );
  AND2_X1 U3615 ( .A1(n4178), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4179)
         );
  NOR2_X1 U3616 ( .A1(n4676), .A2(n3707), .ZN(n5473) );
  NAND2_X1 U3617 ( .A1(n5475), .A2(n4694), .ZN(n7145) );
  OR2_X1 U3618 ( .A1(n5864), .A2(n5486), .ZN(n5913) );
  OR2_X1 U3619 ( .A1(n4317), .A2(n4316), .ZN(n5997) );
  NAND2_X1 U3620 ( .A1(n4269), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4270)
         );
  INV_X1 U3621 ( .A(n4268), .ZN(n4269) );
  AND2_X1 U3622 ( .A1(n4273), .A2(n4272), .ZN(n6024) );
  OR2_X1 U3623 ( .A1(n6443), .A2(n5910), .ZN(n4248) );
  AND2_X1 U3624 ( .A1(n6078), .A2(n3506), .ZN(n6037) );
  OR2_X1 U3625 ( .A1(n7039), .A2(n5910), .ZN(n4143) );
  NOR2_X1 U3626 ( .A1(n4101), .A2(n4100), .ZN(n4102) );
  NAND2_X1 U3627 ( .A1(n4102), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4137)
         );
  OR2_X1 U3628 ( .A1(n6463), .A2(n4477), .ZN(n6485) );
  AND4_X1 U3629 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n5453)
         );
  NAND2_X1 U3630 ( .A1(n6594), .A2(n3457), .ZN(n3522) );
  AND2_X1 U3631 ( .A1(n3458), .A2(n6595), .ZN(n6543) );
  NOR2_X1 U3632 ( .A1(n4657), .A2(n6916), .ZN(n6595) );
  NAND2_X1 U3633 ( .A1(n4476), .A2(n3436), .ZN(n3460) );
  NAND2_X1 U3634 ( .A1(n5758), .A2(n3531), .ZN(n3530) );
  INV_X1 U3635 ( .A(n3533), .ZN(n3531) );
  AOI21_X1 U3636 ( .B1(n6428), .B2(n3455), .A(n3437), .ZN(n3533) );
  NAND2_X1 U3637 ( .A1(n5758), .A2(n3438), .ZN(n3532) );
  NAND2_X1 U3638 ( .A1(n4549), .A2(n3470), .ZN(n4819) );
  NOR2_X1 U3639 ( .A1(n4797), .A2(n4721), .ZN(n3470) );
  NOR2_X1 U3640 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U3641 ( .A1(n6614), .A2(n4644), .ZN(n4761) );
  NAND2_X1 U3642 ( .A1(n5473), .A2(n5969), .ZN(n4638) );
  AND2_X2 U3643 ( .A1(n4393), .A2(n4392), .ZN(n5980) );
  OR2_X1 U3644 ( .A1(n4391), .A2(n4390), .ZN(n4392) );
  INV_X1 U3645 ( .A(n3713), .ZN(n4875) );
  NOR2_X1 U3646 ( .A1(n3585), .A2(n3584), .ZN(n3590) );
  AND2_X1 U3647 ( .A1(n5948), .A2(REIP_REG_31__SCAN_IN), .ZN(n3487) );
  NOR2_X1 U3648 ( .A1(n5920), .A2(n5488), .ZN(n5489) );
  INV_X1 U3649 ( .A(n7035), .ZN(n7050) );
  AND2_X1 U3650 ( .A1(n5935), .A2(n5495), .ZN(n7056) );
  INV_X1 U3651 ( .A(n6150), .ZN(n6159) );
  AND2_X1 U3652 ( .A1(n6150), .A2(n6162), .ZN(n6160) );
  INV_X1 U3653 ( .A(n6163), .ZN(n7206) );
  NAND2_X1 U3654 ( .A1(n3510), .A2(n5942), .ZN(n3509) );
  XNOR2_X1 U3655 ( .A(n4636), .B(n4635), .ZN(n5941) );
  INV_X1 U3656 ( .A(n4346), .ZN(n4358) );
  CLKBUF_X1 U3657 ( .A(n3688), .Z(n4345) );
  NAND2_X1 U3658 ( .A1(n5503), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3772) );
  OR2_X1 U3659 ( .A1(n3885), .A2(n3884), .ZN(n4439) );
  OR2_X1 U3660 ( .A1(n3765), .A2(n3764), .ZN(n4409) );
  NOR2_X1 U3661 ( .A1(n5503), .A2(n7115), .ZN(n4347) );
  NAND2_X1 U3662 ( .A1(n3635), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3813) );
  OR2_X1 U3663 ( .A1(n3809), .A2(n3808), .ZN(n4468) );
  INV_X1 U3664 ( .A(n4362), .ZN(n4377) );
  AND2_X1 U3665 ( .A1(n3692), .A2(n3635), .ZN(n3672) );
  OR2_X1 U3666 ( .A1(n3700), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3685)
         );
  NAND2_X1 U3667 ( .A1(n4633), .A2(n4630), .ZN(n4538) );
  AND2_X1 U3668 ( .A1(n3554), .A2(n3506), .ZN(n3505) );
  NOR2_X1 U3669 ( .A1(n4137), .A2(n6479), .ZN(n4138) );
  INV_X1 U3670 ( .A(n6103), .ZN(n3499) );
  NOR2_X1 U3671 ( .A1(n3502), .A2(n3501), .ZN(n3500) );
  INV_X1 U3672 ( .A(n5804), .ZN(n3502) );
  INV_X1 U3673 ( .A(n5809), .ZN(n3501) );
  AND2_X1 U3674 ( .A1(n4064), .A2(n4029), .ZN(n4034) );
  NAND2_X1 U3675 ( .A1(n3988), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4002)
         );
  NOR2_X1 U3676 ( .A1(n3779), .A2(n4856), .ZN(n3828) );
  OR2_X1 U3677 ( .A1(n6592), .A2(n6426), .ZN(n6429) );
  NOR2_X1 U3678 ( .A1(n6093), .A2(n6141), .ZN(n4596) );
  INV_X1 U3679 ( .A(n6154), .ZN(n3482) );
  AND2_X1 U3680 ( .A1(n3484), .A2(n5772), .ZN(n3483) );
  INV_X1 U3681 ( .A(n6106), .ZN(n3484) );
  INV_X1 U3682 ( .A(n4475), .ZN(n3464) );
  AND2_X1 U3683 ( .A1(n5494), .A2(n4624), .ZN(n4619) );
  AND2_X1 U3684 ( .A1(n4559), .A2(n4564), .ZN(n3481) );
  INV_X1 U3685 ( .A(n4450), .ZN(n4454) );
  OR2_X1 U3686 ( .A1(n3861), .A2(n3860), .ZN(n4431) );
  OR2_X1 U3687 ( .A1(n3750), .A2(n3749), .ZN(n4421) );
  AND2_X1 U3688 ( .A1(n3674), .A2(n3688), .ZN(n4411) );
  OR2_X1 U3689 ( .A1(n3799), .A2(n3798), .ZN(n4416) );
  NAND2_X1 U3690 ( .A1(n4347), .A2(n3737), .ZN(n4362) );
  NAND2_X1 U3691 ( .A1(n4386), .A2(n4385), .ZN(n4521) );
  OR2_X1 U3692 ( .A1(n4362), .A2(n4458), .ZN(n4391) );
  INV_X1 U3693 ( .A(n3687), .ZN(n4343) );
  AOI21_X1 U3694 ( .B1(n7117), .B2(n5179), .A(n4855), .ZN(n4869) );
  NAND2_X1 U3695 ( .A1(n4767), .A2(n4766), .ZN(n7077) );
  INV_X1 U3696 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7075) );
  NOR2_X1 U3697 ( .A1(n5974), .A2(n5975), .ZN(n4755) );
  INV_X1 U3698 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5708) );
  INV_X1 U3699 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U3700 ( .A1(n4819), .A2(n4818), .ZN(n5261) );
  CLKBUF_X1 U3701 ( .A(n3610), .Z(n3779) );
  AND2_X1 U3702 ( .A1(n4696), .A2(n5982), .ZN(n6635) );
  AND2_X1 U3703 ( .A1(n5962), .A2(n3781), .ZN(n5914) );
  INV_X1 U3704 ( .A(n3510), .ZN(n3508) );
  AND2_X1 U3705 ( .A1(n6078), .A2(n3505), .ZN(n6023) );
  NAND2_X1 U3706 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4246)
         );
  OR2_X1 U3707 ( .A1(n4246), .A2(n6052), .ZN(n4268) );
  OR2_X1 U3708 ( .A1(n7061), .A2(n5910), .ZN(n4183) );
  AND2_X1 U3709 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4138), .ZN(n4178)
         );
  INV_X1 U3710 ( .A(n6138), .ZN(n4145) );
  NOR2_X1 U3711 ( .A1(n6484), .A2(n3542), .ZN(n3541) );
  AND2_X1 U3712 ( .A1(n4104), .A2(n4103), .ZN(n6152) );
  NAND2_X1 U3713 ( .A1(n4069), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4101)
         );
  INV_X1 U3714 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4100) );
  AND2_X1 U3715 ( .A1(n6463), .A2(n4477), .ZN(n6484) );
  NAND2_X1 U3716 ( .A1(n3545), .A2(n3544), .ZN(n3543) );
  AND2_X1 U3717 ( .A1(n4054), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4069)
         );
  NOR2_X1 U3718 ( .A1(n4049), .A2(n5784), .ZN(n4054) );
  AND2_X1 U3719 ( .A1(n4018), .A2(n4001), .ZN(n3496) );
  AND2_X1 U3720 ( .A1(n3984), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3988)
         );
  CLKBUF_X1 U3721 ( .A(n5573), .Z(n5700) );
  AND2_X1 U3722 ( .A1(n3493), .A2(n3946), .ZN(n3492) );
  AND2_X1 U3723 ( .A1(n5258), .A2(n3494), .ZN(n3493) );
  INV_X1 U3724 ( .A(n5453), .ZN(n3494) );
  NAND2_X1 U3725 ( .A1(n3940), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3961)
         );
  NAND2_X1 U3726 ( .A1(n4916), .A2(n3491), .ZN(n5454) );
  AND2_X1 U3727 ( .A1(n3946), .A2(n5258), .ZN(n3491) );
  NOR2_X1 U3728 ( .A1(n3929), .A2(n6986), .ZN(n3940) );
  NAND2_X1 U3729 ( .A1(n3911), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3929)
         );
  AND2_X1 U3730 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3890), .ZN(n3911)
         );
  NOR2_X1 U3731 ( .A1(n3867), .A2(n6942), .ZN(n3890) );
  NAND2_X1 U3732 ( .A1(n3866), .A2(n4064), .ZN(n3875) );
  INV_X1 U3733 ( .A(n3788), .ZN(n3843) );
  NAND2_X1 U3734 ( .A1(n4682), .A2(n4681), .ZN(n4716) );
  NAND2_X1 U3735 ( .A1(n4493), .A2(n6493), .ZN(n3515) );
  OR2_X1 U3736 ( .A1(n6059), .A2(n3474), .ZN(n5989) );
  NAND2_X1 U3737 ( .A1(n3475), .A2(n3453), .ZN(n3474) );
  INV_X1 U3738 ( .A(n3476), .ZN(n3475) );
  BUF_X1 U3739 ( .A(n4486), .Z(n6397) );
  NOR3_X1 U3740 ( .A1(n6059), .A2(n3479), .A3(n6041), .ZN(n6027) );
  NAND2_X1 U3741 ( .A1(n6428), .A2(n4658), .ZN(n3521) );
  NAND2_X1 U3742 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4658) );
  NOR2_X1 U3743 ( .A1(n6059), .A2(n6041), .ZN(n6040) );
  AND2_X1 U3744 ( .A1(n4610), .A2(n4609), .ZN(n6060) );
  AND2_X1 U3745 ( .A1(n4603), .A2(n4602), .ZN(n6132) );
  NAND2_X1 U3746 ( .A1(n4596), .A2(n3473), .ZN(n6131) );
  NAND2_X1 U3747 ( .A1(n3545), .A2(n3539), .ZN(n3534) );
  AND2_X1 U3748 ( .A1(n5814), .A2(n3447), .ZN(n6157) );
  NAND2_X1 U3749 ( .A1(n5814), .A2(n3483), .ZN(n6155) );
  AND2_X1 U3750 ( .A1(n5812), .A2(n5811), .ZN(n5814) );
  NAND2_X1 U3751 ( .A1(n5814), .A2(n5772), .ZN(n6105) );
  INV_X1 U3752 ( .A(n5731), .ZN(n3529) );
  AND2_X1 U3753 ( .A1(n4579), .A2(n4578), .ZN(n5732) );
  NOR2_X1 U3754 ( .A1(n3440), .A2(n5732), .ZN(n5812) );
  NAND2_X1 U3755 ( .A1(n5261), .A2(n3480), .ZN(n5575) );
  AND2_X1 U3756 ( .A1(n3481), .A2(n4568), .ZN(n3480) );
  INV_X1 U3757 ( .A(n5570), .ZN(n4568) );
  NOR2_X1 U3758 ( .A1(n5575), .A2(n5576), .ZN(n5704) );
  NAND2_X1 U3759 ( .A1(n4430), .A2(n6742), .ZN(n4435) );
  NAND2_X1 U3760 ( .A1(n4624), .A2(n4622), .ZN(n4684) );
  CLKBUF_X1 U3761 ( .A(n4853), .Z(n4854) );
  NOR2_X1 U3762 ( .A1(n4909), .A2(n4861), .ZN(n5020) );
  NOR2_X1 U3763 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4869), .ZN(n4977) );
  NAND2_X1 U3764 ( .A1(n4514), .A2(n4515), .ZN(n5974) );
  INV_X1 U3765 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5488) );
  INV_X1 U3766 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3468) );
  AOI21_X1 U3767 ( .B1(n3706), .B2(n4525), .A(n3687), .ZN(n3648) );
  NAND2_X1 U3768 ( .A1(n3851), .A2(n3850), .ZN(n4901) );
  OR2_X1 U3769 ( .A1(n3726), .A2(n3845), .ZN(n3851) );
  INV_X1 U3770 ( .A(n3734), .ZN(n3732) );
  AND2_X1 U3771 ( .A1(n4978), .A2(n4909), .ZN(n5236) );
  OR2_X1 U3772 ( .A1(n4922), .A2(n4911), .ZN(n5302) );
  INV_X1 U3773 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7070) );
  INV_X1 U3774 ( .A(n4977), .ZN(n5010) );
  NOR2_X1 U3775 ( .A1(n4732), .A2(n5618), .ZN(n5511) );
  NOR2_X1 U3776 ( .A1(n5515), .A2(n5618), .ZN(n5417) );
  AOI22_X1 U3777 ( .A1(n3626), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3568) );
  AND2_X1 U3778 ( .A1(n4862), .A2(n4861), .ZN(n5043) );
  AOI21_X1 U3779 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7070), .A(n5010), .ZN(
        n5332) );
  OR3_X1 U3780 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4869), .A3(n7110), .ZN(n5012) );
  NOR2_X1 U3781 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5327) );
  INV_X1 U3782 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7097) );
  NOR2_X1 U3783 ( .A1(n5980), .A2(n4534), .ZN(n7093) );
  AND2_X1 U3784 ( .A1(n5488), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4395) );
  OR2_X1 U3785 ( .A1(n4637), .A2(n4415), .ZN(n7102) );
  INV_X1 U3786 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6787) );
  NOR2_X1 U3787 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6787), .ZN(n7129) );
  NOR2_X1 U3788 ( .A1(n6787), .A2(STATE_REG_0__SCAN_IN), .ZN(n7139) );
  INV_X1 U3789 ( .A(n7053), .ZN(n7025) );
  AND2_X1 U3790 ( .A1(n6948), .A2(n5499), .ZN(n7017) );
  AND2_X1 U3791 ( .A1(n6948), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7035) );
  INV_X1 U3792 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5696) );
  INV_X1 U3793 ( .A(n7034), .ZN(n7023) );
  CLKBUF_X1 U3794 ( .A(n4731), .Z(n4732) );
  AND2_X1 U3795 ( .A1(n5490), .A2(n7014), .ZN(n6979) );
  NAND2_X1 U3796 ( .A1(n4680), .A2(n4679), .ZN(n6150) );
  INV_X1 U3797 ( .A(n6160), .ZN(n6148) );
  AND2_X1 U3798 ( .A1(n5836), .A2(n5480), .ZN(n7204) );
  NAND2_X1 U3799 ( .A1(n5476), .A2(n5984), .ZN(n5477) );
  INV_X1 U3800 ( .A(n7204), .ZN(n6387) );
  NAND2_X1 U3801 ( .A1(n5836), .A2(n3673), .ZN(n5839) );
  AND3_X1 U3802 ( .A1(n4498), .A2(n5494), .A3(n7143), .ZN(n5474) );
  XNOR2_X1 U3803 ( .A(n5487), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5920)
         );
  NOR2_X1 U3804 ( .A1(n5913), .A2(n5964), .ZN(n5487) );
  XNOR2_X1 U3805 ( .A(n5985), .B(n5943), .ZN(n5968) );
  INV_X1 U3806 ( .A(n5942), .ZN(n5943) );
  NOR2_X1 U3807 ( .A1(n5999), .A2(n5998), .ZN(n6404) );
  AND2_X1 U3808 ( .A1(n4312), .A2(n4271), .ZN(n6417) );
  OR2_X1 U3809 ( .A1(n6051), .A2(n6050), .ZN(n6447) );
  INV_X1 U3810 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U3811 ( .A1(n6753), .A2(n4689), .ZN(n6778) );
  INV_X1 U3812 ( .A(n6748), .ZN(n6773) );
  INV_X1 U3813 ( .A(n6753), .ZN(n6772) );
  INV_X1 U3814 ( .A(n7062), .ZN(n6774) );
  AND2_X1 U3815 ( .A1(n6543), .A2(n4659), .ZN(n6535) );
  CLKBUF_X1 U3816 ( .A(n6418), .Z(n6419) );
  OAI21_X1 U3817 ( .B1(n6441), .B2(n4658), .A(n6428), .ZN(n3523) );
  OR2_X1 U3818 ( .A1(n5598), .A2(n3532), .ZN(n3527) );
  CLKBUF_X1 U3819 ( .A(n5465), .Z(n5466) );
  CLKBUF_X1 U3820 ( .A(n6762), .Z(n6763) );
  NAND2_X1 U3821 ( .A1(n3471), .A2(n4797), .ZN(n4798) );
  OR2_X1 U3822 ( .A1(n6783), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U3823 ( .A1(n6848), .A2(n4965), .ZN(n6816) );
  AND2_X1 U3824 ( .A1(n4645), .A2(n7071), .ZN(n6818) );
  AND2_X1 U3825 ( .A1(n4645), .A2(n4537), .ZN(n6920) );
  INV_X1 U3826 ( .A(n5925), .ZN(n5187) );
  CLKBUF_X1 U3827 ( .A(n4770), .Z(n4771) );
  NOR2_X1 U3828 ( .A1(n7110), .A2(n5980), .ZN(n4855) );
  AOI21_X1 U3829 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7115), .A(n7066), .ZN(
        n6627) );
  INV_X1 U3830 ( .A(n5253), .ZN(n5129) );
  AND2_X1 U3831 ( .A1(n5236), .A2(n4863), .ZN(n5512) );
  INV_X1 U3832 ( .A(n5512), .ZN(n5552) );
  INV_X1 U3833 ( .A(n5337), .ZN(n5402) );
  INV_X1 U3834 ( .A(n5290), .ZN(n5085) );
  NOR2_X1 U3835 ( .A1(n5273), .A2(n5272), .ZN(n5616) );
  NAND2_X1 U3836 ( .A1(n4947), .A2(n5272), .ZN(n5623) );
  NAND2_X1 U3837 ( .A1(n4947), .A2(n4863), .ZN(n5136) );
  INV_X1 U3838 ( .A(n5360), .ZN(n5137) );
  NOR2_X1 U3839 ( .A1(n7148), .A2(n5010), .ZN(n5398) );
  NOR2_X1 U3840 ( .A1(n7154), .A2(n5010), .ZN(n5384) );
  NOR2_X1 U3841 ( .A1(n7157), .A2(n5010), .ZN(n5375) );
  NOR2_X1 U3842 ( .A1(n7160), .A2(n5010), .ZN(n5390) );
  NOR2_X1 U3843 ( .A1(n7166), .A2(n5010), .ZN(n5380) );
  NOR2_X1 U3844 ( .A1(n4923), .A2(n5272), .ZN(n5361) );
  NOR2_X1 U3845 ( .A1(n7169), .A2(n5010), .ZN(n5357) );
  INV_X1 U3846 ( .A(n5361), .ZN(n5118) );
  NOR2_X1 U3847 ( .A1(n5012), .A2(n5503), .ZN(n5648) );
  NOR2_X1 U3848 ( .A1(n5012), .A2(n4880), .ZN(n5662) );
  INV_X1 U3849 ( .A(n5366), .ZN(n5664) );
  INV_X1 U3850 ( .A(n5384), .ZN(n5689) );
  NOR2_X1 U3851 ( .A1(n5012), .A2(n4875), .ZN(n5676) );
  INV_X1 U3852 ( .A(n5375), .ZN(n5678) );
  INV_X1 U3853 ( .A(n5371), .ZN(n5636) );
  INV_X1 U3854 ( .A(n5380), .ZN(n5657) );
  NAND2_X1 U3855 ( .A1(n5043), .A2(n4863), .ZN(n5128) );
  NAND2_X1 U3856 ( .A1(n5043), .A2(n5272), .ZN(n5117) );
  NOR2_X1 U3857 ( .A1(n5012), .A2(n6162), .ZN(n5669) );
  INV_X1 U3858 ( .A(n5357), .ZN(n5671) );
  INV_X1 U3859 ( .A(n6794), .ZN(n7117) );
  OR2_X1 U3860 ( .A1(n7128), .A2(STATE_REG_0__SCAN_IN), .ZN(n6791) );
  OAI21_X1 U3861 ( .B1(n5941), .B2(n7028), .A(n3485), .ZN(U2796) );
  OR2_X1 U3862 ( .A1(n5939), .A2(n3487), .ZN(n3486) );
  INV_X1 U3863 ( .A(n6166), .ZN(n3488) );
  NAND2_X1 U3864 ( .A1(n5810), .A2(n3500), .ZN(n5803) );
  INV_X1 U3865 ( .A(n3866), .ZN(n4909) );
  NAND2_X1 U3866 ( .A1(n6078), .A2(n6130), .ZN(n6063) );
  NOR2_X1 U3867 ( .A1(n5827), .A2(n3464), .ZN(n3436) );
  AND2_X1 U3868 ( .A1(n5810), .A2(n3452), .ZN(n6102) );
  AND2_X1 U3869 ( .A1(n6474), .A2(n5760), .ZN(n3437) );
  OR2_X1 U3870 ( .A1(n6428), .A2(n3456), .ZN(n3438) );
  NAND2_X1 U3871 ( .A1(n4514), .A2(n3648), .ZN(n3705) );
  NAND2_X1 U3872 ( .A1(n4916), .A2(n5258), .ZN(n5257) );
  NAND2_X1 U3873 ( .A1(n4796), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U3874 ( .A1(n4345), .A2(n3687), .ZN(n4458) );
  INV_X1 U3875 ( .A(n4458), .ZN(n4437) );
  INV_X1 U3876 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3727) );
  AND2_X1 U3877 ( .A1(n3473), .A2(n3472), .ZN(n3439) );
  OR2_X1 U3878 ( .A1(n5744), .A2(n5743), .ZN(n3440) );
  OR2_X1 U3879 ( .A1(n6012), .A2(n3509), .ZN(n3441) );
  NAND2_X1 U3880 ( .A1(n3534), .A2(n3536), .ZN(n6473) );
  AND2_X1 U3881 ( .A1(n5810), .A2(n5809), .ZN(n5802) );
  AND4_X1 U3882 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3442)
         );
  OAI21_X1 U3883 ( .B1(n4726), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4727), 
        .ZN(n4426) );
  OR2_X1 U3884 ( .A1(n6463), .A2(n4571), .ZN(n5758) );
  NAND2_X1 U3885 ( .A1(n3543), .A2(n5769), .ZN(n6483) );
  NAND2_X1 U3886 ( .A1(n3688), .A2(n3675), .ZN(n3694) );
  NAND2_X1 U3887 ( .A1(n3543), .A2(n3541), .ZN(n6472) );
  AND2_X1 U3888 ( .A1(n3525), .A2(n3836), .ZN(n3443) );
  NAND2_X1 U3889 ( .A1(n3523), .A2(n3522), .ZN(n6420) );
  INV_X1 U3890 ( .A(n3537), .ZN(n3536) );
  NOR2_X1 U3891 ( .A1(n3541), .A2(n3538), .ZN(n3537) );
  INV_X1 U3892 ( .A(n3540), .ZN(n3539) );
  NAND2_X1 U3893 ( .A1(n6485), .A2(n3544), .ZN(n3540) );
  NAND2_X1 U3894 ( .A1(n3635), .A2(n3688), .ZN(n3706) );
  INV_X1 U3895 ( .A(n3706), .ZN(n3503) );
  AND2_X1 U3896 ( .A1(n4484), .A2(n3521), .ZN(n3444) );
  INV_X1 U3897 ( .A(n6428), .ZN(n3519) );
  NAND2_X2 U3898 ( .A1(n3824), .A2(n3823), .ZN(n4863) );
  INV_X1 U3899 ( .A(n3675), .ZN(n3778) );
  AND2_X1 U3900 ( .A1(n3497), .A2(n4001), .ZN(n3445) );
  AND2_X1 U3901 ( .A1(n4596), .A2(n3439), .ZN(n3446) );
  AND2_X1 U3902 ( .A1(n4815), .A2(n4917), .ZN(n4916) );
  NOR2_X1 U3903 ( .A1(n6058), .A2(n6060), .ZN(n4611) );
  AND2_X1 U3904 ( .A1(n4916), .A2(n3492), .ZN(n5455) );
  NAND2_X1 U3905 ( .A1(n3460), .A2(n5826), .ZN(n5768) );
  NAND2_X1 U3906 ( .A1(n4476), .A2(n4475), .ZN(n5825) );
  NAND2_X1 U3907 ( .A1(n3527), .A2(n3530), .ZN(n5730) );
  AND2_X1 U3908 ( .A1(n3483), .A2(n3482), .ZN(n3447) );
  OR2_X1 U3909 ( .A1(n6059), .A2(n3476), .ZN(n3448) );
  OR2_X1 U3910 ( .A1(n6463), .A2(n6802), .ZN(n5826) );
  INV_X1 U3911 ( .A(n5826), .ZN(n3463) );
  AND2_X1 U3912 ( .A1(n4434), .A2(n7144), .ZN(n3449) );
  AND2_X1 U3913 ( .A1(n5455), .A2(n5561), .ZN(n5562) );
  AND2_X1 U3914 ( .A1(n3447), .A2(n6094), .ZN(n3450) );
  INV_X1 U3915 ( .A(n3780), .ZN(n5910) );
  NOR2_X1 U3916 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3780) );
  NAND2_X1 U3917 ( .A1(n5261), .A2(n3481), .ZN(n5457) );
  AND2_X1 U3918 ( .A1(n5261), .A2(n4559), .ZN(n3451) );
  INV_X1 U3919 ( .A(n5769), .ZN(n3542) );
  AND2_X1 U3920 ( .A1(n3500), .A2(n3499), .ZN(n3452) );
  AND2_X1 U3921 ( .A1(n5847), .A2(n6000), .ZN(n3453) );
  INV_X1 U3922 ( .A(n4722), .ZN(n4549) );
  NAND2_X1 U3923 ( .A1(n3844), .A2(n4719), .ZN(n4717) );
  AND2_X1 U3924 ( .A1(n3439), .A2(n6066), .ZN(n3454) );
  NAND2_X1 U3925 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3455) );
  NOR2_X1 U3926 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3456) );
  AND3_X1 U3927 ( .A1(n6581), .A2(n6545), .A3(n6564), .ZN(n3457) );
  AND2_X1 U3928 ( .A1(n6562), .A2(n6563), .ZN(n3458) );
  OAI21_X1 U3929 ( .B1(n3427), .B2(n5560), .A(n3459), .ZN(n6880) );
  AOI21_X1 U3930 ( .B1(n3866), .B2(n4437), .A(n3449), .ZN(n4804) );
  NAND3_X1 U3931 ( .A1(n3467), .A2(n3466), .A3(n4870), .ZN(n3717) );
  NAND2_X2 U3932 ( .A1(n3599), .A2(n3600), .ZN(n3610) );
  AND2_X2 U3933 ( .A1(n4744), .A2(n3469), .ZN(n3626) );
  NAND3_X1 U3934 ( .A1(n3516), .A2(n6474), .A3(n3515), .ZN(n5959) );
  AND2_X4 U3935 ( .A1(n3469), .A2(n4895), .ZN(n4038) );
  AND2_X2 U3936 ( .A1(n3469), .A2(n4746), .ZN(n4055) );
  INV_X1 U3937 ( .A(n4720), .ZN(n3471) );
  NAND2_X1 U3938 ( .A1(n4596), .A2(n3454), .ZN(n6058) );
  INV_X1 U3939 ( .A(n4596), .ZN(n6143) );
  INV_X1 U3940 ( .A(n6080), .ZN(n3473) );
  INV_X1 U3941 ( .A(n6025), .ZN(n3479) );
  NAND2_X1 U3942 ( .A1(n5814), .A2(n3450), .ZN(n6093) );
  NAND2_X1 U3943 ( .A1(n3490), .A2(n4794), .ZN(n3489) );
  INV_X1 U3944 ( .A(n4816), .ZN(n3490) );
  NAND3_X1 U3945 ( .A1(n4910), .A2(n4064), .A3(n3865), .ZN(n3495) );
  NAND2_X1 U3946 ( .A1(n5810), .A2(n3498), .ZN(n6089) );
  NAND3_X1 U3947 ( .A1(n3687), .A2(n3713), .A3(n3503), .ZN(n4508) );
  NAND2_X1 U3948 ( .A1(n6078), .A2(n3504), .ZN(n6011) );
  NOR2_X1 U3949 ( .A1(n6012), .A2(n3508), .ZN(n5985) );
  NOR2_X1 U3950 ( .A1(n6012), .A2(n5997), .ZN(n5999) );
  NOR2_X2 U3951 ( .A1(n3514), .A2(n3513), .ZN(n3675) );
  NAND4_X1 U3952 ( .A1(n3568), .A2(n3570), .A3(n3562), .A4(n3569), .ZN(n3513)
         );
  NAND4_X1 U3953 ( .A1(n3565), .A2(n3563), .A3(n3571), .A4(n3564), .ZN(n3514)
         );
  NAND2_X1 U3954 ( .A1(n4492), .A2(n4491), .ZN(n3517) );
  AOI21_X2 U3955 ( .B1(n5958), .B2(n3519), .A(n3518), .ZN(n4496) );
  OAI21_X1 U3956 ( .B1(n4493), .B2(n4494), .A(n3555), .ZN(n3518) );
  NAND2_X1 U3957 ( .A1(n6441), .A2(n6428), .ZN(n3520) );
  NAND3_X1 U3958 ( .A1(n3522), .A2(n3444), .A3(n3520), .ZN(n6418) );
  NAND3_X1 U3959 ( .A1(n4430), .A2(n6742), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4801) );
  NAND2_X1 U3960 ( .A1(n4801), .A2(n4804), .ZN(n4436) );
  NAND2_X1 U3961 ( .A1(n3832), .A2(n3833), .ZN(n3836) );
  NAND2_X1 U3962 ( .A1(n3524), .A2(n4414), .ZN(n4726) );
  NAND3_X1 U3963 ( .A1(n3525), .A2(n4437), .A3(n3836), .ZN(n3524) );
  NAND2_X1 U3964 ( .A1(n3526), .A2(n3528), .ZN(n4476) );
  NAND2_X1 U3965 ( .A1(n5598), .A2(n3530), .ZN(n3526) );
  INV_X1 U3966 ( .A(n5768), .ZN(n3545) );
  OR2_X1 U3967 ( .A1(n6517), .A2(n7062), .ZN(n4489) );
  NAND2_X1 U3968 ( .A1(n6091), .A2(n4145), .ZN(n6140) );
  OAI21_X1 U3969 ( .B1(n6390), .B2(n3547), .A(n6389), .ZN(n6391) );
  XNOR2_X1 U3970 ( .A(n6391), .B(n6505), .ZN(n6510) );
  XNOR2_X1 U3971 ( .A(n5961), .B(n4494), .ZN(n6499) );
  NAND2_X2 U3972 ( .A1(n3733), .A2(n3732), .ZN(n4900) );
  OR2_X1 U3973 ( .A1(n4338), .A2(n5999), .ZN(n4339) );
  INV_X1 U3974 ( .A(n3443), .ZN(n5295) );
  OR2_X1 U3975 ( .A1(n4070), .A2(n3679), .ZN(n6614) );
  AOI22_X1 U3976 ( .A1(n4411), .A2(n4070), .B1(n3713), .B2(n3694), .ZN(n3633)
         );
  NOR2_X2 U3977 ( .A1(n6398), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4492)
         );
  INV_X1 U3978 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7110) );
  INV_X1 U3979 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5908) );
  INV_X1 U3980 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U3981 ( .A1(n3694), .A2(n3737), .ZN(n3546) );
  AND2_X1 U3982 ( .A1(n6474), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3547)
         );
  INV_X1 U3983 ( .A(n6474), .ZN(n5957) );
  INV_X1 U3984 ( .A(n3946), .ZN(n5451) );
  OAI21_X1 U3985 ( .B1(n4459), .B2(n4053), .A(n3945), .ZN(n3946) );
  INV_X1 U3986 ( .A(n6037), .ZN(n6064) );
  OR2_X1 U3987 ( .A1(n5845), .A2(n6748), .ZN(n3548) );
  AND3_X1 U3988 ( .A1(n3721), .A2(n3720), .A3(n4772), .ZN(n3549) );
  AND4_X1 U3989 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3551)
         );
  AND4_X1 U3990 ( .A1(n3579), .A2(n3578), .A3(n3577), .A4(n3576), .ZN(n3552)
         );
  INV_X1 U3991 ( .A(n3712), .ZN(n4415) );
  AND2_X1 U3992 ( .A1(n3908), .A2(n3937), .ZN(n3553) );
  NOR2_X1 U3993 ( .A1(n4250), .A2(n6049), .ZN(n3554) );
  OR2_X1 U3994 ( .A1(n3519), .A2(n4495), .ZN(n3555) );
  INV_X1 U3995 ( .A(n5741), .ZN(n4018) );
  OR2_X1 U3996 ( .A1(n5908), .A2(n4698), .ZN(n7099) );
  OR2_X1 U3997 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3556)
         );
  OR2_X1 U3998 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3557)
         );
  OR2_X1 U3999 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3558)
         );
  AND4_X1 U4000 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3559)
         );
  INV_X1 U4001 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4494) );
  INV_X1 U4002 ( .A(n3828), .ZN(n4309) );
  NAND2_X1 U4003 ( .A1(n5465), .A2(n4473), .ZN(n5559) );
  INV_X1 U4004 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3845) );
  INV_X1 U4005 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7083) );
  AND4_X1 U4006 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3560)
         );
  AOI21_X1 U4007 ( .B1(n3689), .B2(n3679), .A(n4525), .ZN(n3690) );
  NOR2_X1 U4008 ( .A1(n3845), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4374)
         );
  OR2_X1 U4009 ( .A1(n3924), .A2(n3923), .ZN(n4461) );
  AOI21_X1 U4010 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n4383) );
  AND2_X1 U4011 ( .A1(n3674), .A2(n3713), .ZN(n4511) );
  OR2_X1 U4012 ( .A1(n3907), .A2(n3906), .ZN(n4405) );
  AND4_X1 U4013 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  INV_X1 U4014 ( .A(n3936), .ZN(n3908) );
  INV_X1 U4015 ( .A(n6092), .ZN(n4121) );
  NAND2_X1 U4016 ( .A1(n4457), .A2(n6755), .ZN(n6761) );
  OR2_X1 U4017 ( .A1(n4382), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4522)
         );
  NAND2_X1 U4018 ( .A1(n3778), .A2(n3610), .ZN(n3680) );
  INV_X1 U4019 ( .A(n5885), .ZN(n5906) );
  NAND2_X1 U4020 ( .A1(n4030), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4049)
         );
  AND2_X1 U4021 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5853), .ZN(n6030) );
  NOR2_X1 U4022 ( .A1(n3961), .A2(n5696), .ZN(n3984) );
  INV_X1 U4023 ( .A(n7102), .ZN(n4694) );
  OR2_X1 U4024 ( .A1(n4314), .A2(n6005), .ZN(n5864) );
  NAND2_X1 U4025 ( .A1(n4512), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5885) );
  NOR2_X1 U4026 ( .A1(n4002), .A2(n5708), .ZN(n4030) );
  NAND2_X1 U4027 ( .A1(n6418), .A2(n4485), .ZN(n6407) );
  OR2_X1 U4028 ( .A1(n6818), .A2(n4709), .ZN(n4806) );
  INV_X1 U4029 ( .A(n5302), .ZN(n5296) );
  INV_X1 U4030 ( .A(n5623), .ZN(n5681) );
  AND2_X1 U4031 ( .A1(n5039), .A2(n3729), .ZN(n4857) );
  OR3_X1 U4032 ( .A1(n7064), .A2(STATE2_REG_1__SCAN_IN), .A3(n4531), .ZN(n4904) );
  INV_X1 U4033 ( .A(n4669), .ZN(n5975) );
  INV_X1 U4034 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6052) );
  INV_X1 U4035 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U4036 ( .A1(n5935), .A2(n5493), .ZN(n6958) );
  AND2_X1 U4037 ( .A1(n4589), .A2(n4588), .ZN(n6154) );
  INV_X1 U4038 ( .A(n3680), .ZN(n5969) );
  AND2_X1 U4039 ( .A1(n5908), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5917) );
  INV_X1 U4040 ( .A(n4064), .ZN(n4053) );
  INV_X1 U4041 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6986) );
  NOR2_X2 U4042 ( .A1(n3778), .A2(n4856), .ZN(n4064) );
  NAND2_X1 U4043 ( .A1(n6390), .A2(n6463), .ZN(n6389) );
  INV_X1 U4044 ( .A(n6816), .ZN(n6874) );
  NAND2_X1 U4045 ( .A1(n4645), .A2(n4761), .ZN(n4965) );
  NAND2_X1 U4046 ( .A1(n5200), .A2(n4909), .ZN(n5550) );
  INV_X1 U4047 ( .A(n5400), .ZN(n5084) );
  INV_X1 U4048 ( .A(n5616), .ZN(n5684) );
  INV_X1 U4049 ( .A(n4863), .ZN(n5272) );
  INV_X1 U4050 ( .A(n5327), .ZN(n5618) );
  INV_X1 U4051 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U4052 ( .A1(n4179), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4205)
         );
  AND2_X1 U4053 ( .A1(n7021), .A2(REIP_REG_17__SCAN_IN), .ZN(n7042) );
  INV_X1 U4054 ( .A(n7014), .ZN(n7057) );
  NOR2_X1 U4055 ( .A1(n6951), .A2(n6783), .ZN(n7034) );
  AND2_X1 U4056 ( .A1(n5935), .A2(n5505), .ZN(n7053) );
  NAND2_X1 U4057 ( .A1(n5986), .A2(n4339), .ZN(n5845) );
  INV_X1 U4058 ( .A(n6151), .ZN(n5782) );
  INV_X1 U4059 ( .A(n6370), .ZN(n7207) );
  AND2_X1 U4060 ( .A1(n4184), .A2(n4183), .ZN(n6130) );
  INV_X1 U4061 ( .A(n7120), .ZN(n5984) );
  INV_X1 U4062 ( .A(n6778), .ZN(n6477) );
  OAI21_X1 U4063 ( .B1(n5941), .B2(n6897), .A(n4664), .ZN(n4665) );
  NOR2_X1 U4064 ( .A1(n6902), .A2(n4656), .ZN(n6909) );
  INV_X1 U4065 ( .A(n4965), .ZN(n6853) );
  INV_X1 U4066 ( .A(n6897), .ZN(n6926) );
  NOR2_X1 U4067 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6619) );
  AND2_X1 U4068 ( .A1(n5236), .A2(n5272), .ZN(n5253) );
  OAI211_X1 U4069 ( .C1(n5521), .C2(n5555), .A(n5520), .B(n5519), .ZN(n5554)
         );
  INV_X1 U4070 ( .A(n5303), .ZN(n5392) );
  OAI211_X1 U4071 ( .C1(n5175), .C2(n7110), .A(n5151), .B(n5520), .ZN(n5173)
         );
  AND2_X1 U4072 ( .A1(n5145), .A2(n4863), .ZN(n5400) );
  AND2_X1 U4073 ( .A1(n4771), .A2(n6618), .ZN(n5265) );
  NOR2_X1 U4074 ( .A1(n5273), .A2(n4863), .ZN(n5290) );
  AND2_X1 U4075 ( .A1(n5516), .A2(n4732), .ZN(n5624) );
  AND2_X1 U4076 ( .A1(n4924), .A2(n5272), .ZN(n5360) );
  NOR2_X1 U4077 ( .A1(n4771), .A2(n6618), .ZN(n5329) );
  NOR2_X1 U4078 ( .A1(n7151), .A2(n5010), .ZN(n5366) );
  NOR2_X1 U4079 ( .A1(n7163), .A2(n5010), .ZN(n5371) );
  INV_X1 U4080 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7115) );
  INV_X1 U4081 ( .A(READY_N), .ZN(n7143) );
  INV_X1 U4082 ( .A(n6718), .ZN(n6704) );
  NAND2_X1 U4083 ( .A1(n4668), .A2(n5475), .ZN(n7141) );
  NAND2_X1 U4084 ( .A1(n7141), .A2(n5481), .ZN(n6798) );
  INV_X1 U4085 ( .A(n7056), .ZN(n7028) );
  OAI211_X1 U4086 ( .C1(n5479), .C2(n5478), .A(n7196), .B(n5477), .ZN(n6163)
         );
  NAND2_X1 U4087 ( .A1(n6635), .A2(n4697), .ZN(n4840) );
  INV_X1 U4088 ( .A(n6635), .ZN(n6668) );
  NAND2_X2 U4089 ( .A1(n5475), .A2(n5474), .ZN(n7196) );
  NAND2_X1 U4090 ( .A1(n7062), .A2(n4397), .ZN(n6753) );
  NAND2_X1 U4091 ( .A1(n7093), .A2(n5984), .ZN(n7062) );
  INV_X1 U4092 ( .A(n4665), .ZN(n4666) );
  AOI22_X1 U4093 ( .A1(n6853), .A2(n4655), .B1(n4654), .B2(n6842), .ZN(n6902)
         );
  INV_X1 U4094 ( .A(n6920), .ZN(n6590) );
  NAND2_X1 U4095 ( .A1(n4645), .A2(n4639), .ZN(n6897) );
  INV_X1 U4096 ( .A(n4732), .ZN(n5515) );
  AOI22_X1 U4097 ( .A1(n5628), .A2(n5624), .B1(n5621), .B2(n5620), .ZN(n5690)
         );
  INV_X1 U4098 ( .A(n5648), .ZN(n5405) );
  INV_X1 U4099 ( .A(n5676), .ZN(n5379) );
  INV_X1 U4100 ( .A(n5669), .ZN(n5365) );
  INV_X1 U4101 ( .A(n5398), .ZN(n5650) );
  INV_X1 U4102 ( .A(n5390), .ZN(n5643) );
  NAND2_X1 U4103 ( .A1(n4395), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7120) );
  OAI21_X1 U4104 ( .B1(n7129), .B2(n6786), .A(n6703), .ZN(n6631) );
  AND2_X1 U4105 ( .A1(n3678), .A2(n3677), .ZN(n7128) );
  INV_X1 U4106 ( .A(n6716), .ZN(n6706) );
  INV_X1 U4107 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3561) );
  AND2_X2 U4108 ( .A1(n3566), .A2(n4746), .ZN(n5890) );
  AOI22_X1 U4109 ( .A1(n5890), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3565) );
  AND2_X2 U4110 ( .A1(n3566), .A2(n4895), .ZN(n4146) );
  AND2_X2 U4111 ( .A1(n4744), .A2(n6613), .ZN(n3621) );
  AOI22_X1 U4112 ( .A1(n4146), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3564) );
  AND2_X2 U4113 ( .A1(n4746), .A2(n6613), .ZN(n3743) );
  AND2_X2 U4114 ( .A1(n4738), .A2(n4895), .ZN(n3658) );
  AOI22_X1 U4115 ( .A1(n3743), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4116 ( .A1(n4055), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4117 ( .A1(n3653), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3571) );
  AND2_X2 U4118 ( .A1(n4744), .A2(n4738), .ZN(n3641) );
  AND2_X2 U4119 ( .A1(n3566), .A2(n3567), .ZN(n3642) );
  AOI22_X1 U4120 ( .A1(n3642), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4121 ( .A1(n3621), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4122 ( .A1(n4146), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3574)
         );
  NAND2_X1 U4123 ( .A1(n3743), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4124 ( .A1(n3658), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3572)
         );
  NAND2_X1 U4125 ( .A1(n3653), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3579)
         );
  NAND2_X1 U4126 ( .A1(n4274), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4127 ( .A1(n3641), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3577)
         );
  NAND2_X1 U4128 ( .A1(n4740), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U4129 ( .A1(n3643), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3581)
         );
  NAND2_X1 U4130 ( .A1(n3642), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4131 ( .A1(n3581), .A2(n3580), .ZN(n3585) );
  NAND2_X1 U4132 ( .A1(n3626), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3583) );
  NAND2_X1 U4133 ( .A1(n3744), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4134 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4135 ( .A1(n5890), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4136 ( .A1(n4038), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3588)
         );
  NAND2_X1 U4137 ( .A1(n4055), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U4138 ( .A1(n3755), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4139 ( .A1(n4038), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4140 ( .A1(n3653), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4141 ( .A1(n3626), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4142 ( .A1(n4146), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4143 ( .A1(n5890), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4144 ( .A1(n3642), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4145 ( .A1(n3621), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4146 ( .A1(n4274), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4147 ( .A1(n3653), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4148 ( .A1(n4274), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4149 ( .A1(n3626), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4150 ( .A1(n3642), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4151 ( .A1(n3743), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4152 ( .A1(n5890), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4153 ( .A1(n4146), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4154 ( .A1(n4055), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3605) );
  INV_X1 U4155 ( .A(n3636), .ZN(n4870) );
  NAND2_X1 U4156 ( .A1(n3717), .A2(n3680), .ZN(n3634) );
  INV_X1 U4157 ( .A(n3636), .ZN(n3674) );
  AOI22_X1 U4158 ( .A1(n5890), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4159 ( .A1(n4146), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4160 ( .A1(n3743), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4161 ( .A1(n4055), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4162 ( .A1(n4740), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4163 ( .A1(n4274), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4164 ( .A1(n3642), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4165 ( .A1(n3626), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3615) );
  NAND2_X2 U4166 ( .A1(n3620), .A2(n3619), .ZN(n3688) );
  AOI22_X1 U4167 ( .A1(n3743), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4168 ( .A1(n4146), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4169 ( .A1(n5890), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4170 ( .A1(n4055), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4171 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3632)
         );
  AOI22_X1 U4172 ( .A1(n4274), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4173 ( .A1(n3653), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4174 ( .A1(n4320), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4175 ( .A1(n3626), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4176 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3631)
         );
  AOI22_X1 U4177 ( .A1(n4038), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4178 ( .A1(n4055), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4179 ( .A1(n4146), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4180 ( .A1(n3626), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3744), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4181 ( .A1(n4274), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4182 ( .A1(n5890), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3743), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4183 ( .A1(n3653), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3755), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4184 ( .A1(n4320), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3644) );
  NAND2_X2 U4185 ( .A1(n3559), .A2(n3551), .ZN(n3687) );
  INV_X1 U4186 ( .A(n3705), .ZN(n3671) );
  NAND2_X1 U4187 ( .A1(n4038), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3652)
         );
  NAND2_X1 U4188 ( .A1(n5890), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3651) );
  NAND2_X1 U4189 ( .A1(n4055), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4190 ( .A1(n3755), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3649) );
  NAND2_X1 U4191 ( .A1(n3653), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3657)
         );
  NAND2_X1 U4192 ( .A1(n4274), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3656) );
  NAND2_X1 U4193 ( .A1(n3641), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3655)
         );
  NAND2_X1 U4194 ( .A1(n4740), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3654) );
  NAND2_X1 U4195 ( .A1(n4146), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3662)
         );
  NAND2_X1 U4196 ( .A1(n3621), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4197 ( .A1(n3743), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U4198 ( .A1(n3658), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3659)
         );
  NAND2_X1 U4199 ( .A1(n3626), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4200 ( .A1(n4320), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4201 ( .A1(n3643), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3664)
         );
  NAND2_X1 U4202 ( .A1(n3744), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3663) );
  AND4_X4 U4203 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n5503)
         );
  AND2_X1 U4204 ( .A1(n3503), .A2(n5503), .ZN(n4515) );
  NAND2_X1 U4205 ( .A1(n3694), .A2(n3610), .ZN(n5480) );
  INV_X1 U4206 ( .A(n5480), .ZN(n3673) );
  INV_X1 U4207 ( .A(n3688), .ZN(n3679) );
  NAND2_X1 U4208 ( .A1(n3679), .A2(n3778), .ZN(n3692) );
  NAND2_X1 U4209 ( .A1(n4511), .A2(n3675), .ZN(n3676) );
  NOR2_X2 U4210 ( .A1(n4502), .A2(n3676), .ZN(n4497) );
  INV_X1 U4211 ( .A(n5503), .ZN(n4697) );
  AND2_X2 U4212 ( .A1(n4497), .A2(n4697), .ZN(n4668) );
  NAND2_X1 U4213 ( .A1(n6787), .A2(STATE_REG_2__SCAN_IN), .ZN(n3678) );
  INV_X1 U4214 ( .A(n7129), .ZN(n3677) );
  NAND2_X1 U4215 ( .A1(n4343), .A2(n7128), .ZN(n3689) );
  NAND2_X1 U4216 ( .A1(n4668), .A2(n3689), .ZN(n3681) );
  NAND3_X1 U4217 ( .A1(n3679), .A2(n4870), .A3(n4875), .ZN(n4676) );
  NAND2_X1 U4218 ( .A1(n4343), .A2(n5503), .ZN(n3707) );
  NAND3_X1 U4219 ( .A1(n4531), .A2(n3681), .A3(n4638), .ZN(n3682) );
  NAND2_X1 U4220 ( .A1(n3682), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3702) );
  INV_X1 U4221 ( .A(n3702), .ZN(n3686) );
  NAND2_X1 U4222 ( .A1(n6619), .A2(n7115), .ZN(n4396) );
  NAND2_X1 U4223 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3728) );
  OAI21_X1 U4224 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n3728), .ZN(n4920) );
  OR2_X1 U4225 ( .A1(n4396), .A2(n4920), .ZN(n3684) );
  INV_X1 U4226 ( .A(n4395), .ZN(n3848) );
  NAND2_X1 U4227 ( .A1(n3848), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4228 ( .A1(n3684), .A2(n3683), .ZN(n3700) );
  NAND2_X1 U4229 ( .A1(n3686), .A2(n3685), .ZN(n3703) );
  NAND2_X1 U4230 ( .A1(n3712), .A2(n3737), .ZN(n3691) );
  NAND3_X1 U4231 ( .A1(n4508), .A2(n3691), .A3(n3690), .ZN(n3696) );
  OAI211_X1 U4232 ( .C1(n3694), .C2(n3737), .A(n3693), .B(n3692), .ZN(n4500)
         );
  INV_X1 U4233 ( .A(n4500), .ZN(n3695) );
  NAND2_X1 U4234 ( .A1(n3695), .A2(n3546), .ZN(n3716) );
  NOR2_X1 U4235 ( .A1(n3696), .A2(n3716), .ZN(n3698) );
  NAND2_X1 U4236 ( .A1(n3705), .A2(n5503), .ZN(n3697) );
  NAND2_X1 U4237 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  INV_X1 U4238 ( .A(n3700), .ZN(n3701) );
  OAI211_X1 U4239 ( .C1(n3726), .C2(n3430), .A(n3702), .B(n3701), .ZN(n3724)
         );
  NAND2_X1 U4240 ( .A1(n3703), .A2(n3724), .ZN(n3754) );
  INV_X1 U4241 ( .A(n3754), .ZN(n3723) );
  MUX2_X1 U4242 ( .A(n4396), .B(n4395), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3704) );
  NAND2_X1 U4243 ( .A1(n3706), .A2(n5503), .ZN(n3708) );
  NAND2_X1 U4244 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  NAND2_X1 U4245 ( .A1(n3705), .A2(n3709), .ZN(n4735) );
  NAND2_X1 U4246 ( .A1(n4502), .A2(n7144), .ZN(n3711) );
  NAND2_X1 U4247 ( .A1(n4697), .A2(n4525), .ZN(n3710) );
  NAND2_X1 U4248 ( .A1(n3711), .A2(n3710), .ZN(n4506) );
  INV_X1 U4249 ( .A(n4506), .ZN(n3722) );
  NAND2_X1 U4250 ( .A1(n6619), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7104) );
  INV_X1 U4251 ( .A(n7104), .ZN(n3714) );
  OAI211_X1 U4252 ( .C1(n4415), .C2(n4501), .A(n4508), .B(n3714), .ZN(n3715)
         );
  INV_X1 U4253 ( .A(n3715), .ZN(n3721) );
  NAND2_X1 U4254 ( .A1(n3716), .A2(n3687), .ZN(n3720) );
  INV_X1 U4255 ( .A(n3717), .ZN(n3719) );
  AND2_X1 U4256 ( .A1(n4875), .A2(n5503), .ZN(n3718) );
  NAND2_X1 U4257 ( .A1(n3719), .A2(n3718), .ZN(n4772) );
  NAND3_X1 U4258 ( .A1(n4735), .A2(n3722), .A3(n3549), .ZN(n3769) );
  NAND2_X1 U4259 ( .A1(n3768), .A2(n3769), .ZN(n3752) );
  NAND2_X1 U4260 ( .A1(n3723), .A2(n3752), .ZN(n3725) );
  NAND2_X1 U4261 ( .A1(n3725), .A2(n3724), .ZN(n3735) );
  INV_X1 U4262 ( .A(n3735), .ZN(n3733) );
  INV_X1 U4263 ( .A(n3728), .ZN(n5190) );
  NAND2_X1 U4264 ( .A1(n5190), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U4265 ( .A1(n3728), .A2(n7083), .ZN(n3729) );
  INV_X1 U4266 ( .A(n4396), .ZN(n3849) );
  AOI22_X1 U4267 ( .A1(n4857), .A2(n3849), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3848), .ZN(n3730) );
  NAND2_X1 U4268 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  NAND2_X1 U4269 ( .A1(n4900), .A2(n3736), .ZN(n4770) );
  AOI22_X1 U4270 ( .A1(n4190), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4271 ( .A1(n3738), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4272 ( .A1(n4038), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4273 ( .A1(n4320), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4274 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3750)
         );
  AOI22_X1 U4275 ( .A1(n5897), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4274), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4276 ( .A1(n4189), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4277 ( .A1(n5896), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4278 ( .A1(n5875), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4279 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  AOI22_X1 U4280 ( .A1(n4377), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4387), 
        .B2(n4421), .ZN(n3751) );
  INV_X1 U4281 ( .A(n3431), .ZN(n3775) );
  INV_X1 U4282 ( .A(n3752), .ZN(n3753) );
  XNOR2_X1 U4283 ( .A(n3754), .B(n3753), .ZN(n4853) );
  NAND2_X1 U4284 ( .A1(n4853), .A2(n7115), .ZN(n3767) );
  AOI22_X1 U4285 ( .A1(n4190), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4286 ( .A1(n5897), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4287 ( .A1(n4189), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4288 ( .A1(n4320), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3756) );
  NAND4_X1 U4289 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3765)
         );
  AOI22_X1 U4290 ( .A1(n4318), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4291 ( .A1(n4299), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4292 ( .A1(n3621), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4293 ( .A1(n5875), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4294 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3764)
         );
  OR2_X1 U4295 ( .A1(n3771), .A2(n3813), .ZN(n3766) );
  NAND2_X1 U4296 ( .A1(n3767), .A2(n3766), .ZN(n3832) );
  INV_X1 U4297 ( .A(n3769), .ZN(n3770) );
  XNOR2_X2 U4298 ( .A(n3768), .B(n3770), .ZN(n3827) );
  OAI21_X1 U4299 ( .B1(n3772), .B2(n3771), .A(n3813), .ZN(n3773) );
  AOI21_X1 U4300 ( .B1(n4377), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n3773), 
        .ZN(n3774) );
  NAND2_X1 U4301 ( .A1(n3818), .A2(n3774), .ZN(n3833) );
  INV_X1 U4302 ( .A(n3836), .ZN(n3776) );
  NOR2_X1 U4303 ( .A1(n3680), .A2(n4856), .ZN(n3888) );
  NAND2_X1 U4304 ( .A1(n3888), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3786) );
  INV_X2 U4305 ( .A(n4309), .ZN(n5912) );
  INV_X1 U4306 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3783) );
  INV_X1 U4307 ( .A(n5917), .ZN(n4081) );
  INV_X1 U4308 ( .A(n5910), .ZN(n3781) );
  NAND2_X1 U4309 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3867) );
  OAI21_X1 U4310 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3867), .ZN(n6940) );
  NAND2_X1 U4311 ( .A1(n3781), .A2(n6940), .ZN(n3782) );
  OAI21_X1 U4312 ( .B1(n3783), .B2(n4081), .A(n3782), .ZN(n3784) );
  AOI21_X1 U4313 ( .B1(n5912), .B2(EAX_REG_2__SCAN_IN), .A(n3784), .ZN(n3785)
         );
  AND2_X1 U4314 ( .A1(n3786), .A2(n3785), .ZN(n3842) );
  INV_X1 U4315 ( .A(n3842), .ZN(n3787) );
  NAND2_X1 U4316 ( .A1(n3788), .A2(n3787), .ZN(n3841) );
  INV_X1 U4317 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3789) );
  OR2_X1 U4318 ( .A1(n4362), .A2(n3789), .ZN(n3812) );
  AOI22_X1 U4319 ( .A1(n4190), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4320 ( .A1(n4299), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4321 ( .A1(n4189), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4322 ( .A1(n5875), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4323 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3799)
         );
  AOI22_X1 U4324 ( .A1(n4038), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4325 ( .A1(n5897), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4326 ( .A1(n4318), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4327 ( .A1(n3738), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4328 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  AOI21_X1 U4329 ( .B1(n5503), .B2(n4416), .A(n7115), .ZN(n3810) );
  AOI22_X1 U4331 ( .A1(n3738), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4332 ( .A1(n4038), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4333 ( .A1(n4190), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4334 ( .A1(n5875), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4335 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3809)
         );
  AOI22_X1 U4336 ( .A1(n5897), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4337 ( .A1(n3621), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4338 ( .A1(n4189), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4339 ( .A1(n4274), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4340 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  NAND2_X1 U4341 ( .A1(n3635), .A2(n4468), .ZN(n4402) );
  AND2_X1 U4342 ( .A1(n3810), .A2(n4402), .ZN(n3811) );
  NAND2_X1 U4343 ( .A1(n3812), .A2(n3811), .ZN(n3819) );
  INV_X1 U4344 ( .A(n3813), .ZN(n3816) );
  INV_X1 U4345 ( .A(n4468), .ZN(n3814) );
  XNOR2_X1 U4346 ( .A(n3814), .B(n4416), .ZN(n3815) );
  NAND2_X1 U4347 ( .A1(n3816), .A2(n3815), .ZN(n3820) );
  AND2_X1 U4348 ( .A1(n3819), .A2(n3820), .ZN(n3817) );
  NAND2_X1 U4349 ( .A1(n3818), .A2(n3817), .ZN(n3824) );
  INV_X1 U4350 ( .A(n3819), .ZN(n3822) );
  INV_X1 U4351 ( .A(n3820), .ZN(n3821) );
  NAND2_X1 U4352 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  NAND2_X1 U4353 ( .A1(n3675), .A2(n3779), .ZN(n3825) );
  OR2_X1 U4354 ( .A1(n4863), .A2(n3825), .ZN(n3826) );
  NAND2_X1 U4355 ( .A1(n3826), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4688) );
  INV_X1 U4356 ( .A(n3888), .ZN(n3872) );
  AOI22_X1 U4357 ( .A1(n3828), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4856), .ZN(n3829) );
  OAI21_X1 U4358 ( .B1(n3561), .B2(n3872), .A(n3829), .ZN(n3830) );
  AOI21_X1 U4359 ( .B1(n3827), .B2(n4064), .A(n3830), .ZN(n4687) );
  MUX2_X1 U4360 ( .A(n4688), .B(n5910), .S(n4687), .Z(n3831) );
  INV_X1 U4361 ( .A(n3831), .ZN(n4682) );
  INV_X1 U4362 ( .A(n3832), .ZN(n3835) );
  INV_X1 U4363 ( .A(n3833), .ZN(n3834) );
  NAND2_X1 U4364 ( .A1(n3443), .A2(n4064), .ZN(n3840) );
  NAND2_X1 U4365 ( .A1(n3888), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4366 ( .A1(n5912), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4856), .ZN(n3837) );
  AND2_X1 U4367 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  NAND2_X1 U4368 ( .A1(n3840), .A2(n3839), .ZN(n4681) );
  NAND2_X1 U4369 ( .A1(n3841), .A2(n4716), .ZN(n3844) );
  NAND2_X1 U4370 ( .A1(n3843), .A2(n3842), .ZN(n4719) );
  INV_X1 U4371 ( .A(n5039), .ZN(n3846) );
  NAND2_X1 U4372 ( .A1(n3846), .A2(n7084), .ZN(n5406) );
  NAND2_X1 U4373 ( .A1(n5039), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3847) );
  NAND2_X1 U4374 ( .A1(n5406), .A2(n3847), .ZN(n4975) );
  AOI22_X1 U4375 ( .A1(n4975), .A2(n3849), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3848), .ZN(n3850) );
  XNOR2_X1 U4376 ( .A(n4900), .B(n4901), .ZN(n4731) );
  NAND2_X1 U4377 ( .A1(n4731), .A2(n7115), .ZN(n3863) );
  AOI22_X1 U4378 ( .A1(n4190), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4379 ( .A1(n4189), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4380 ( .A1(n5869), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4381 ( .A1(n4318), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4382 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3861)
         );
  AOI22_X1 U4383 ( .A1(n4274), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4384 ( .A1(n5897), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4385 ( .A1(n4151), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4386 ( .A1(n5875), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4387 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  AOI22_X1 U4388 ( .A1(n4377), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4387), 
        .B2(n4431), .ZN(n3862) );
  INV_X1 U4389 ( .A(n3864), .ZN(n4860) );
  NAND2_X1 U4390 ( .A1(n4860), .A2(n3865), .ZN(n4911) );
  INV_X1 U4391 ( .A(n3867), .ZN(n3869) );
  INV_X1 U4392 ( .A(n3890), .ZN(n3868) );
  OAI21_X1 U4393 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3869), .A(n3868), 
        .ZN(n6941) );
  AOI22_X1 U4394 ( .A1(n3781), .A2(n6941), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4395 ( .A1(n5912), .A2(EAX_REG_3__SCAN_IN), .ZN(n3870) );
  OAI211_X1 U4396 ( .C1(n3872), .C2(n3845), .A(n3871), .B(n3870), .ZN(n3873)
         );
  INV_X1 U4397 ( .A(n3873), .ZN(n3874) );
  NAND2_X1 U4398 ( .A1(n4377), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4399 ( .A1(n4190), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4400 ( .A1(n4189), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4401 ( .A1(n5869), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4402 ( .A1(n4318), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4403 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4404 ( .A1(n4299), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4405 ( .A1(n5897), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4406 ( .A1(n4151), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4407 ( .A1(n5875), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4408 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NAND2_X1 U4409 ( .A1(n4387), .A2(n4439), .ZN(n3886) );
  NAND2_X1 U4410 ( .A1(n3887), .A2(n3886), .ZN(n3896) );
  NAND2_X1 U4411 ( .A1(n3888), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3893) );
  INV_X1 U4412 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6962) );
  AOI21_X1 U4413 ( .B1(n6962), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3889) );
  AOI21_X1 U4414 ( .B1(n5912), .B2(EAX_REG_4__SCAN_IN), .A(n3889), .ZN(n3892)
         );
  NOR2_X1 U4415 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3890), .ZN(n3891)
         );
  NOR2_X1 U4416 ( .A1(n3911), .A2(n3891), .ZN(n6963) );
  AOI22_X1 U4417 ( .A1(n3893), .A2(n3892), .B1(n3780), .B2(n6963), .ZN(n3894)
         );
  AOI21_X1 U4418 ( .B1(n4438), .B2(n4064), .A(n3894), .ZN(n4816) );
  INV_X1 U4419 ( .A(n3895), .ZN(n3897) );
  NAND2_X1 U4420 ( .A1(n3897), .A2(n3896), .ZN(n3909) );
  INV_X1 U4421 ( .A(n3909), .ZN(n3938) );
  AOI22_X1 U4422 ( .A1(n4151), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4423 ( .A1(n4190), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4424 ( .A1(n4299), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4425 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n4189), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4426 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3907)
         );
  AOI22_X1 U4427 ( .A1(n5897), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4428 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n5875), .B1(n5869), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4429 ( .A1(n4191), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4430 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n4318), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4431 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  AOI22_X1 U4432 ( .A1(n4377), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4387), 
        .B2(n4405), .ZN(n3936) );
  NAND2_X1 U4433 ( .A1(n3938), .A2(n3908), .ZN(n3928) );
  NAND2_X1 U4434 ( .A1(n3909), .A2(n3936), .ZN(n3910) );
  NAND2_X1 U4435 ( .A1(n3928), .A2(n3910), .ZN(n4408) );
  INV_X1 U4436 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6975) );
  OAI21_X1 U4437 ( .B1(n3911), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3929), 
        .ZN(n6978) );
  NAND2_X1 U4438 ( .A1(n6978), .A2(n3780), .ZN(n3912) );
  OAI21_X1 U4439 ( .B1(n6975), .B2(n4081), .A(n3912), .ZN(n3913) );
  AOI21_X1 U4440 ( .B1(n5912), .B2(EAX_REG_5__SCAN_IN), .A(n3913), .ZN(n3914)
         );
  OAI21_X1 U4441 ( .B1(n4408), .B2(n4053), .A(n3914), .ZN(n4917) );
  NAND2_X1 U4442 ( .A1(n4377), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4443 ( .A1(n4190), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4444 ( .A1(n4189), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4445 ( .A1(n5869), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4446 ( .A1(n4318), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4447 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3924)
         );
  AOI22_X1 U4448 ( .A1(n4274), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4449 ( .A1(n5897), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4450 ( .A1(n4151), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4451 ( .A1(n5875), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4452 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3923)
         );
  NAND2_X1 U4453 ( .A1(n4387), .A2(n4461), .ZN(n3925) );
  NAND2_X1 U4454 ( .A1(n3926), .A2(n3925), .ZN(n3937) );
  INV_X1 U4455 ( .A(n3937), .ZN(n3927) );
  NAND2_X1 U4456 ( .A1(n3928), .A2(n3927), .ZN(n4453) );
  NAND2_X1 U4457 ( .A1(n4453), .A2(n4064), .ZN(n3935) );
  AND2_X1 U4458 ( .A1(n3929), .A2(n6986), .ZN(n3930) );
  OR2_X1 U4459 ( .A1(n3930), .A2(n3940), .ZN(n6987) );
  INV_X1 U4460 ( .A(n6987), .ZN(n3933) );
  NOR2_X1 U4461 ( .A1(n6986), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3931) );
  AOI21_X1 U4462 ( .B1(n5912), .B2(EAX_REG_6__SCAN_IN), .A(n3931), .ZN(n3932)
         );
  MUX2_X1 U4463 ( .A(n3933), .B(n3932), .S(n5910), .Z(n3934) );
  NAND2_X1 U4464 ( .A1(n3935), .A2(n3934), .ZN(n5258) );
  AOI22_X1 U4465 ( .A1(n4377), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4387), 
        .B2(n4468), .ZN(n3939) );
  XNOR2_X1 U4466 ( .A(n4401), .B(n3939), .ZN(n4459) );
  OR2_X1 U4467 ( .A1(n3940), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4468 ( .A1(n3961), .A2(n3941), .ZN(n6999) );
  NAND2_X1 U4469 ( .A1(n6999), .A2(n3780), .ZN(n3943) );
  NAND2_X1 U4470 ( .A1(n5917), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3942)
         );
  NAND2_X1 U4471 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  AOI21_X1 U4472 ( .B1(n5912), .B2(EAX_REG_7__SCAN_IN), .A(n3944), .ZN(n3945)
         );
  AOI22_X1 U4473 ( .A1(n4318), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4474 ( .A1(n5897), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4475 ( .A1(n4151), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4476 ( .A1(n5891), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4477 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3956)
         );
  AOI22_X1 U4478 ( .A1(n4190), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4479 ( .A1(n3738), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4480 ( .A1(n5875), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4274), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4481 ( .A1(n4038), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3951) );
  NAND4_X1 U4482 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3955)
         );
  OAI21_X1 U4483 ( .B1(n3956), .B2(n3955), .A(n4064), .ZN(n3960) );
  NAND2_X1 U4484 ( .A1(n5912), .A2(EAX_REG_8__SCAN_IN), .ZN(n3959) );
  XNOR2_X1 U4485 ( .A(n3961), .B(n5696), .ZN(n5691) );
  NAND2_X1 U4486 ( .A1(n5691), .A2(n3780), .ZN(n3958) );
  NAND2_X1 U4487 ( .A1(n5917), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3957)
         );
  XOR2_X1 U4488 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3984), .Z(n5565) );
  AOI22_X1 U4489 ( .A1(n5912), .A2(EAX_REG_9__SCAN_IN), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4490 ( .A1(n4319), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4491 ( .A1(n3738), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4492 ( .A1(n4189), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4493 ( .A1(n4299), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4494 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4495 ( .A1(n5875), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4496 ( .A1(n5896), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4497 ( .A1(n4190), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4498 ( .A1(n5897), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4499 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  OAI21_X1 U4500 ( .B1(n3971), .B2(n3970), .A(n4064), .ZN(n3972) );
  OAI211_X1 U4501 ( .C1(n5565), .C2(n5910), .A(n3973), .B(n3972), .ZN(n5561)
         );
  AOI22_X1 U4502 ( .A1(n4190), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4503 ( .A1(n5897), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4504 ( .A1(n4274), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4505 ( .A1(n5875), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4506 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3983)
         );
  AOI22_X1 U4507 ( .A1(n3738), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4508 ( .A1(n4318), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4509 ( .A1(n5869), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4510 ( .A1(n4319), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4511 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3982)
         );
  NOR2_X1 U4512 ( .A1(n3983), .A2(n3982), .ZN(n3987) );
  XNOR2_X1 U4513 ( .A(n3988), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5602)
         );
  NAND2_X1 U4514 ( .A1(n5602), .A2(n3781), .ZN(n3986) );
  AOI22_X1 U4515 ( .A1(n5912), .A2(EAX_REG_10__SCAN_IN), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3985) );
  OAI211_X1 U4516 ( .C1(n3987), .C2(n4053), .A(n3986), .B(n3985), .ZN(n5574)
         );
  NAND2_X1 U4517 ( .A1(n5562), .A2(n5574), .ZN(n5573) );
  XOR2_X1 U4518 ( .A(n5708), .B(n4002), .Z(n5723) );
  AOI22_X1 U4519 ( .A1(n5912), .A2(EAX_REG_11__SCAN_IN), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4520 ( .A1(n5897), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4521 ( .A1(n4319), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4522 ( .A1(n4038), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4523 ( .A1(n5875), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U4524 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3998)
         );
  AOI22_X1 U4525 ( .A1(n4189), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4526 ( .A1(n3738), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4527 ( .A1(n4190), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4528 ( .A1(n4299), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4529 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3997)
         );
  OAI21_X1 U4530 ( .B1(n3998), .B2(n3997), .A(n4064), .ZN(n3999) );
  OAI211_X1 U4531 ( .C1(n5723), .C2(n5910), .A(n4000), .B(n3999), .ZN(n4001)
         );
  INV_X1 U4532 ( .A(n4001), .ZN(n5701) );
  XNOR2_X1 U4533 ( .A(n4030), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5763)
         );
  INV_X1 U4534 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4003) );
  INV_X1 U4535 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5749) );
  OAI22_X1 U4536 ( .A1(n4309), .A2(n4003), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5749), .ZN(n4004) );
  NAND2_X1 U4537 ( .A1(n4004), .A2(n5910), .ZN(n4016) );
  AOI22_X1 U4538 ( .A1(n4038), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4539 ( .A1(n5897), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4540 ( .A1(n4190), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4541 ( .A1(n4151), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4542 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4543 ( .A1(n4319), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4544 ( .A1(n4299), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4545 ( .A1(n4318), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4546 ( .A1(n5875), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4547 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  OAI21_X1 U4548 ( .B1(n4014), .B2(n4013), .A(n4064), .ZN(n4015) );
  NAND2_X1 U4549 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  AOI21_X1 U4550 ( .B1(n5763), .B2(n3781), .A(n4017), .ZN(n5741) );
  AOI22_X1 U4551 ( .A1(n4190), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4552 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n4318), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4553 ( .A1(n5897), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4554 ( .A1(n4299), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U4555 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4028)
         );
  AOI22_X1 U4556 ( .A1(n3738), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4557 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n4038), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4558 ( .A1(n5875), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4559 ( .A1(n4319), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4560 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  OR2_X1 U4561 ( .A1(n4028), .A2(n4027), .ZN(n4029) );
  XNOR2_X2 U4562 ( .A(n5742), .B(n4034), .ZN(n5779) );
  NAND2_X1 U4563 ( .A1(n5912), .A2(EAX_REG_13__SCAN_IN), .ZN(n4033) );
  INV_X1 U4564 ( .A(n4049), .ZN(n4031) );
  XNOR2_X1 U4565 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4031), .ZN(n5797)
         );
  AOI22_X1 U4566 ( .A1(n3781), .A2(n5797), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4567 ( .A1(n4033), .A2(n4032), .ZN(n5780) );
  NAND2_X1 U4568 ( .A1(n5779), .A2(n5780), .ZN(n4037) );
  INV_X1 U4569 ( .A(n5742), .ZN(n4035) );
  NAND2_X1 U4570 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  NAND2_X2 U4571 ( .A1(n4037), .A2(n4036), .ZN(n5810) );
  AOI22_X1 U4572 ( .A1(n4189), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4573 ( .A1(n4299), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4574 ( .A1(n5897), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4575 ( .A1(n5875), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U4576 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4048)
         );
  AOI22_X1 U4577 ( .A1(n4190), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4578 ( .A1(n4318), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4579 ( .A1(n5869), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4580 ( .A1(n4151), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4043) );
  NAND4_X1 U4581 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(n4047)
         );
  NOR2_X1 U4582 ( .A1(n4048), .A2(n4047), .ZN(n4052) );
  XNOR2_X1 U4583 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4054), .ZN(n5830)
         );
  AOI22_X1 U4584 ( .A1(n3781), .A2(n5830), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4051) );
  NAND2_X1 U4585 ( .A1(n5912), .A2(EAX_REG_14__SCAN_IN), .ZN(n4050) );
  OAI211_X1 U4586 ( .C1(n4053), .C2(n4052), .A(n4051), .B(n4050), .ZN(n5809)
         );
  XOR2_X1 U4587 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4069), .Z(n7018) );
  AOI22_X1 U4588 ( .A1(n5912), .A2(EAX_REG_15__SCAN_IN), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4589 ( .A1(n5897), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4590 ( .A1(n4299), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4591 ( .A1(n4055), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4592 ( .A1(n4190), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U4593 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4066)
         );
  AOI22_X1 U4594 ( .A1(n4189), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U4595 ( .A1(n4319), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4596 ( .A1(n5891), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4597 ( .A1(n5875), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4060) );
  NAND4_X1 U4598 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4065)
         );
  OAI21_X1 U4599 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4067) );
  OAI211_X1 U4600 ( .C1(n7018), .C2(n5910), .A(n4068), .B(n4067), .ZN(n5804)
         );
  XNOR2_X1 U4601 ( .A(n4101), .B(n4100), .ZN(n6489) );
  AOI22_X1 U4602 ( .A1(n4190), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4603 ( .A1(n5875), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4604 ( .A1(n4318), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4605 ( .A1(n4299), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U4606 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4080)
         );
  AOI22_X1 U4607 ( .A1(n4189), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4608 ( .A1(n5897), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4609 ( .A1(n3738), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4610 ( .A1(n5869), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U4611 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NOR2_X1 U4612 ( .A1(n4080), .A2(n4079), .ZN(n4084) );
  NOR2_X1 U4613 ( .A1(n4081), .A2(n4100), .ZN(n4082) );
  AOI21_X1 U4614 ( .B1(n5912), .B2(EAX_REG_16__SCAN_IN), .A(n4082), .ZN(n4083)
         );
  OAI21_X1 U4615 ( .B1(n5885), .B2(n4084), .A(n4083), .ZN(n4085) );
  AOI21_X1 U4616 ( .B1(n6489), .B2(n3781), .A(n4085), .ZN(n6103) );
  AOI22_X1 U4617 ( .A1(n4190), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4618 ( .A1(n4299), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4619 ( .A1(n4189), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4620 ( .A1(n5875), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U4621 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4095)
         );
  AOI22_X1 U4622 ( .A1(n5897), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U4623 ( .A1(n5869), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4624 ( .A1(n4151), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4625 ( .A1(n4319), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4090) );
  NAND4_X1 U4626 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4094)
         );
  NOR2_X1 U4627 ( .A1(n4095), .A2(n4094), .ZN(n4099) );
  NAND2_X1 U4628 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4096)
         );
  NAND2_X1 U4629 ( .A1(n5910), .A2(n4096), .ZN(n4097) );
  AOI21_X1 U4630 ( .B1(n5912), .B2(EAX_REG_17__SCAN_IN), .A(n4097), .ZN(n4098)
         );
  OAI21_X1 U4631 ( .B1(n5885), .B2(n4099), .A(n4098), .ZN(n4104) );
  OAI21_X1 U4632 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4102), .A(n4137), 
        .ZN(n7033) );
  OR2_X1 U4633 ( .A1(n5910), .A2(n7033), .ZN(n4103) );
  INV_X1 U4634 ( .A(n6089), .ZN(n4122) );
  AOI22_X1 U4635 ( .A1(n4319), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4636 ( .A1(n5875), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4637 ( .A1(n4320), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U4638 ( .A1(n4299), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U4639 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4116)
         );
  AOI22_X1 U4640 ( .A1(n4740), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U4641 ( .A1(n4146), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4110) );
  NAND2_X1 U4642 ( .A1(n4191), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4109) );
  AND3_X1 U4643 ( .A1(n4110), .A2(n5910), .A3(n4109), .ZN(n4113) );
  AOI22_X1 U4644 ( .A1(n3738), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4645 ( .A1(n5897), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4646 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4115)
         );
  NAND2_X1 U4647 ( .A1(n5885), .A2(n5910), .ZN(n4198) );
  OAI21_X1 U4648 ( .B1(n4116), .B2(n4115), .A(n4198), .ZN(n4118) );
  AOI22_X1 U4649 ( .A1(n5912), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4856), .ZN(n4117) );
  NAND2_X1 U4650 ( .A1(n4118), .A2(n4117), .ZN(n4120) );
  XNOR2_X1 U4651 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4137), .ZN(n6476)
         );
  NAND2_X1 U4652 ( .A1(n3780), .A2(n6476), .ZN(n4119) );
  NAND2_X1 U4653 ( .A1(n4120), .A2(n4119), .ZN(n6092) );
  NAND2_X1 U4654 ( .A1(n4122), .A2(n4121), .ZN(n6090) );
  AOI22_X1 U4655 ( .A1(n4038), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U4656 ( .A1(n4299), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U4657 ( .A1(n4318), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U4658 ( .A1(n5875), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U4659 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4132)
         );
  AOI22_X1 U4660 ( .A1(n4190), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4661 ( .A1(n5897), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U4662 ( .A1(n4151), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U4663 ( .A1(n4189), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U4664 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4131)
         );
  NOR2_X1 U4665 ( .A1(n4132), .A2(n4131), .ZN(n4136) );
  NAND2_X1 U4666 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4133)
         );
  NAND2_X1 U4667 ( .A1(n5910), .A2(n4133), .ZN(n4134) );
  AOI21_X1 U4668 ( .B1(n5912), .B2(EAX_REG_19__SCAN_IN), .A(n4134), .ZN(n4135)
         );
  OAI21_X1 U4669 ( .B1(n5885), .B2(n4136), .A(n4135), .ZN(n4144) );
  INV_X1 U4670 ( .A(n4178), .ZN(n4142) );
  INV_X1 U4671 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4140) );
  INV_X1 U4672 ( .A(n4138), .ZN(n4139) );
  NAND2_X1 U4673 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  NAND2_X1 U4674 ( .A1(n4142), .A2(n4141), .ZN(n7039) );
  NAND2_X1 U4675 ( .A1(n4144), .A2(n4143), .ZN(n6138) );
  AOI22_X1 U4676 ( .A1(n5897), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U4677 ( .A1(n3738), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U4678 ( .A1(n5875), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4679 ( .A1(n5891), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U4680 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4159)
         );
  AOI22_X1 U4681 ( .A1(n4319), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U4682 ( .A1(n4299), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U4683 ( .A1(n4038), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U4684 ( .A1(n5869), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U4685 ( .A1(n4191), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4152) );
  AND3_X1 U4686 ( .A1(n4153), .A2(n4152), .A3(n5910), .ZN(n4154) );
  NAND4_X1 U4687 ( .A1(n4157), .A2(n4156), .A3(n4155), .A4(n4154), .ZN(n4158)
         );
  OAI21_X1 U4688 ( .B1(n4159), .B2(n4158), .A(n4198), .ZN(n4161) );
  AOI22_X1 U4689 ( .A1(n5912), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n4856), .ZN(n4160) );
  NAND2_X1 U4690 ( .A1(n4161), .A2(n4160), .ZN(n4163) );
  INV_X1 U4691 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6466) );
  XNOR2_X1 U4692 ( .A(n4178), .B(n6466), .ZN(n6470) );
  NAND2_X1 U4693 ( .A1(n6470), .A2(n3781), .ZN(n4162) );
  NAND2_X1 U4694 ( .A1(n4163), .A2(n4162), .ZN(n6077) );
  NOR2_X2 U4695 ( .A1(n6140), .A2(n6077), .ZN(n6078) );
  AOI22_X1 U4696 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4190), .B1(n3621), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U4697 ( .A1(n4038), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4698 ( .A1(n5897), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4699 ( .A1(n4151), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4164) );
  NAND4_X1 U4700 ( .A1(n4167), .A2(n4166), .A3(n4165), .A4(n4164), .ZN(n4173)
         );
  AOI22_X1 U4701 ( .A1(n4299), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U4702 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n4318), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4703 ( .A1(n5875), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4704 ( .A1(n4189), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U4705 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4172)
         );
  NOR2_X1 U4706 ( .A1(n4173), .A2(n4172), .ZN(n4177) );
  NAND2_X1 U4707 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4174)
         );
  NAND2_X1 U4708 ( .A1(n5910), .A2(n4174), .ZN(n4175) );
  AOI21_X1 U4709 ( .B1(n5912), .B2(EAX_REG_21__SCAN_IN), .A(n4175), .ZN(n4176)
         );
  OAI21_X1 U4710 ( .B1(n5885), .B2(n4177), .A(n4176), .ZN(n4184) );
  INV_X1 U4711 ( .A(n4179), .ZN(n4181) );
  INV_X1 U4712 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4180) );
  NAND2_X1 U4713 ( .A1(n4181), .A2(n4180), .ZN(n4182) );
  NAND2_X1 U4714 ( .A1(n4205), .A2(n4182), .ZN(n7061) );
  AOI22_X1 U4715 ( .A1(n5897), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5875), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4716 ( .A1(n3738), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4717 ( .A1(n4319), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4740), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U4718 ( .A1(n5869), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4185) );
  NAND4_X1 U4719 ( .A1(n4188), .A2(n4187), .A3(n4186), .A4(n4185), .ZN(n4200)
         );
  AOI22_X1 U4720 ( .A1(n4190), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U4721 ( .A1(n4299), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U4722 ( .A1(n4151), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4195) );
  AOI21_X1 U4723 ( .B1(n5876), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n3781), 
        .ZN(n4193) );
  NAND2_X1 U4724 ( .A1(n4191), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4192) );
  AND2_X1 U4725 ( .A1(n4193), .A2(n4192), .ZN(n4194) );
  NAND4_X1 U4726 ( .A1(n4197), .A2(n4196), .A3(n4195), .A4(n4194), .ZN(n4199)
         );
  OAI21_X1 U4727 ( .B1(n4200), .B2(n4199), .A(n4198), .ZN(n4202) );
  AOI22_X1 U4728 ( .A1(n5912), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n4856), .ZN(n4201) );
  NAND2_X1 U4729 ( .A1(n4202), .A2(n4201), .ZN(n4204) );
  XNOR2_X1 U4730 ( .A(n4205), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6450)
         );
  NAND2_X1 U4731 ( .A1(n6450), .A2(n3780), .ZN(n4203) );
  NAND2_X1 U4732 ( .A1(n4204), .A2(n4203), .ZN(n6065) );
  INV_X1 U4733 ( .A(n4205), .ZN(n4206) );
  XNOR2_X1 U4734 ( .A(n4268), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6045)
         );
  AOI22_X1 U4735 ( .A1(n4190), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U4736 ( .A1(n4189), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4737 ( .A1(n5869), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4738 ( .A1(n4318), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4207) );
  NAND4_X1 U4739 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4216)
         );
  AOI22_X1 U4740 ( .A1(n4274), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U4741 ( .A1(n5897), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4742 ( .A1(n4320), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U4743 ( .A1(n5875), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4211) );
  NAND4_X1 U4744 ( .A1(n4214), .A2(n4213), .A3(n4212), .A4(n4211), .ZN(n4215)
         );
  OR2_X1 U4745 ( .A1(n4216), .A2(n4215), .ZN(n4240) );
  AOI22_X1 U4746 ( .A1(n4190), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U4747 ( .A1(n4189), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U4748 ( .A1(n5869), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U4749 ( .A1(n4318), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U4750 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4226)
         );
  AOI22_X1 U4751 ( .A1(n4274), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4752 ( .A1(n5897), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U4753 ( .A1(n4320), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U4754 ( .A1(n5875), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4221) );
  NAND4_X1 U4755 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  OR2_X1 U4756 ( .A1(n4226), .A2(n4225), .ZN(n4241) );
  NAND2_X1 U4757 ( .A1(n4240), .A2(n4241), .ZN(n4262) );
  AOI22_X1 U4758 ( .A1(n4190), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U4759 ( .A1(n4038), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U4760 ( .A1(n5897), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4761 ( .A1(n4320), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U4762 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4236)
         );
  AOI22_X1 U4763 ( .A1(n4274), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U4764 ( .A1(n4189), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U4765 ( .A1(n5875), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U4766 ( .A1(n4319), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4231) );
  NAND4_X1 U4767 ( .A1(n4234), .A2(n4233), .A3(n4232), .A4(n4231), .ZN(n4235)
         );
  OR2_X1 U4768 ( .A1(n4236), .A2(n4235), .ZN(n4261) );
  XNOR2_X1 U4769 ( .A(n4262), .B(n4261), .ZN(n4237) );
  NAND2_X1 U4770 ( .A1(n5906), .A2(n4237), .ZN(n4239) );
  AOI22_X1 U4771 ( .A1(n5912), .A2(EAX_REG_24__SCAN_IN), .B1(n5917), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4238) );
  OAI211_X1 U4772 ( .C1(n6045), .C2(n5910), .A(n4239), .B(n4238), .ZN(n6038)
         );
  INV_X1 U4773 ( .A(n6038), .ZN(n4250) );
  OAI21_X1 U4774 ( .B1(n4241), .B2(n4240), .A(n4262), .ZN(n4245) );
  NAND2_X1 U4775 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4242)
         );
  NAND2_X1 U4776 ( .A1(n5910), .A2(n4242), .ZN(n4243) );
  AOI21_X1 U4777 ( .B1(n5912), .B2(EAX_REG_23__SCAN_IN), .A(n4243), .ZN(n4244)
         );
  OAI21_X1 U4778 ( .B1(n5885), .B2(n4245), .A(n4244), .ZN(n4249) );
  NAND2_X1 U4779 ( .A1(n4246), .A2(n6052), .ZN(n4247) );
  NAND2_X1 U4780 ( .A1(n4268), .A2(n4247), .ZN(n6443) );
  NAND2_X1 U4781 ( .A1(n4249), .A2(n4248), .ZN(n6049) );
  AOI22_X1 U4782 ( .A1(n4190), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U4783 ( .A1(n4189), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U4784 ( .A1(n5869), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4785 ( .A1(n4318), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4251) );
  NAND4_X1 U4786 ( .A1(n4254), .A2(n4253), .A3(n4252), .A4(n4251), .ZN(n4260)
         );
  AOI22_X1 U4787 ( .A1(n4299), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U4788 ( .A1(n5897), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U4789 ( .A1(n4320), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4790 ( .A1(n5875), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4255) );
  NAND4_X1 U4791 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4259)
         );
  OR2_X1 U4792 ( .A1(n4260), .A2(n4259), .ZN(n4285) );
  INV_X1 U4793 ( .A(n4261), .ZN(n4263) );
  NOR2_X1 U4794 ( .A1(n4263), .A2(n4262), .ZN(n4286) );
  XNOR2_X1 U4795 ( .A(n4285), .B(n4286), .ZN(n4267) );
  NAND2_X1 U4796 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4264)
         );
  NAND2_X1 U4797 ( .A1(n5910), .A2(n4264), .ZN(n4265) );
  AOI21_X1 U4798 ( .B1(n5912), .B2(EAX_REG_25__SCAN_IN), .A(n4265), .ZN(n4266)
         );
  OAI21_X1 U4799 ( .B1(n5885), .B2(n4267), .A(n4266), .ZN(n4273) );
  INV_X1 U4800 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U4801 ( .A1(n4270), .A2(n6415), .ZN(n4271) );
  NAND2_X1 U4802 ( .A1(n6417), .A2(n3780), .ZN(n4272) );
  AOI22_X1 U4803 ( .A1(n3738), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U4804 ( .A1(n4189), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4805 ( .A1(n4274), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4806 ( .A1(n4319), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4275) );
  NAND4_X1 U4807 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(n4284)
         );
  AOI22_X1 U4808 ( .A1(n4190), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U4809 ( .A1(n5897), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4810 ( .A1(n4038), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U4811 ( .A1(n5875), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4279) );
  NAND4_X1 U4812 ( .A1(n4282), .A2(n4281), .A3(n4280), .A4(n4279), .ZN(n4283)
         );
  NOR2_X1 U4813 ( .A1(n4284), .A2(n4283), .ZN(n4294) );
  NAND2_X1 U4814 ( .A1(n4286), .A2(n4285), .ZN(n4293) );
  XOR2_X1 U4815 ( .A(n4294), .B(n4293), .Z(n4287) );
  NAND2_X1 U4816 ( .A1(n4287), .A2(n5906), .ZN(n4290) );
  INV_X1 U4817 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6411) );
  OAI21_X1 U4818 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6411), .A(n5910), .ZN(
        n4288) );
  AOI21_X1 U4819 ( .B1(n5912), .B2(EAX_REG_26__SCAN_IN), .A(n4288), .ZN(n4289)
         );
  NAND2_X1 U4820 ( .A1(n4290), .A2(n4289), .ZN(n4292) );
  XNOR2_X1 U4821 ( .A(n4312), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6409)
         );
  NAND2_X1 U4822 ( .A1(n6409), .A2(n3780), .ZN(n4291) );
  NAND2_X1 U4823 ( .A1(n4292), .A2(n4291), .ZN(n6014) );
  OR2_X2 U4824 ( .A1(n6011), .A2(n6014), .ZN(n6012) );
  NOR2_X1 U4825 ( .A1(n4294), .A2(n4293), .ZN(n4332) );
  AOI22_X1 U4826 ( .A1(n4190), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4298) );
  AOI22_X1 U4827 ( .A1(n4189), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4828 ( .A1(n5869), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4829 ( .A1(n4318), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4295) );
  NAND4_X1 U4830 ( .A1(n4298), .A2(n4297), .A3(n4296), .A4(n4295), .ZN(n4305)
         );
  AOI22_X1 U4831 ( .A1(n4299), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U4832 ( .A1(n3653), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U4833 ( .A1(n4320), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U4834 ( .A1(n5875), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4300) );
  NAND4_X1 U4835 ( .A1(n4303), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(n4304)
         );
  OR2_X1 U4836 ( .A1(n4305), .A2(n4304), .ZN(n4331) );
  INV_X1 U4837 ( .A(n4331), .ZN(n4306) );
  XNOR2_X1 U4838 ( .A(n4332), .B(n4306), .ZN(n4311) );
  INV_X1 U4839 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4308) );
  NAND2_X1 U4840 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4307)
         );
  OAI211_X1 U4841 ( .C1(n4309), .C2(n4308), .A(n5910), .B(n4307), .ZN(n4310)
         );
  AOI21_X1 U4842 ( .B1(n4311), .B2(n5906), .A(n4310), .ZN(n4317) );
  INV_X1 U4843 ( .A(n4312), .ZN(n4313) );
  NAND2_X1 U4844 ( .A1(n4313), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4314)
         );
  INV_X1 U4845 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U4846 ( .A1(n4314), .A2(n6005), .ZN(n4315) );
  NAND2_X1 U4847 ( .A1(n5864), .A2(n4315), .ZN(n6402) );
  NOR2_X1 U4848 ( .A1(n6402), .A2(n5910), .ZN(n4316) );
  AOI22_X1 U4849 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4189), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U4850 ( .A1(n3653), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4274), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U4851 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4319), .B1(n5869), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U4852 ( .A1(n4320), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4321) );
  NAND4_X1 U4853 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(n4330)
         );
  AOI22_X1 U4854 ( .A1(n3738), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4855 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4038), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4856 ( .A1(n5875), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4857 ( .A1(n4190), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4325) );
  NAND4_X1 U4858 ( .A1(n4328), .A2(n4327), .A3(n4326), .A4(n4325), .ZN(n4329)
         );
  NOR2_X1 U4859 ( .A1(n4330), .A2(n4329), .ZN(n5868) );
  NAND2_X1 U4860 ( .A1(n4332), .A2(n4331), .ZN(n5867) );
  XOR2_X1 U4861 ( .A(n5868), .B(n5867), .Z(n4333) );
  NAND2_X1 U4862 ( .A1(n4333), .A2(n5906), .ZN(n4337) );
  INV_X1 U4863 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5863) );
  AOI21_X1 U4864 ( .B1(n5863), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4334) );
  AOI21_X1 U4865 ( .B1(n5912), .B2(EAX_REG_28__SCAN_IN), .A(n4334), .ZN(n4336)
         );
  INV_X1 U4866 ( .A(n5864), .ZN(n4335) );
  XOR2_X1 U4867 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(n4335), .Z(n5856) );
  AOI22_X1 U4868 ( .A1(n4337), .A2(n4336), .B1(n3780), .B2(n5856), .ZN(n4338)
         );
  NAND2_X1 U4869 ( .A1(n7115), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4698) );
  INV_X1 U4870 ( .A(n4698), .ZN(n5482) );
  NAND2_X1 U4871 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5482), .ZN(n6792) );
  INV_X1 U4872 ( .A(n6792), .ZN(n4340) );
  NAND2_X2 U4873 ( .A1(n5327), .A2(n4340), .ZN(n6748) );
  XNOR2_X1 U4874 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U4875 ( .A1(n7070), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4346) );
  XNOR2_X1 U4876 ( .A(n4359), .B(n4358), .ZN(n4519) );
  INV_X1 U4877 ( .A(n4519), .ZN(n4342) );
  INV_X1 U4878 ( .A(n4391), .ZN(n4341) );
  AOI21_X1 U4879 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n4342), .A(n4341), .ZN(
        n4357) );
  INV_X1 U4880 ( .A(n4387), .ZN(n4350) );
  OAI21_X1 U4881 ( .B1(n4350), .B2(n4880), .A(n4345), .ZN(n4344) );
  AOI21_X1 U4882 ( .B1(n4377), .B2(n4519), .A(n4344), .ZN(n4356) );
  INV_X1 U4883 ( .A(n4356), .ZN(n4354) );
  INV_X1 U4884 ( .A(n4357), .ZN(n4353) );
  INV_X1 U4885 ( .A(n3707), .ZN(n5485) );
  AOI21_X1 U4886 ( .B1(n4880), .B2(n4345), .A(n5485), .ZN(n4364) );
  OAI21_X1 U4887 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7070), .A(n4346), 
        .ZN(n4349) );
  OAI21_X1 U4888 ( .B1(n3503), .B2(n4349), .A(n4347), .ZN(n4348) );
  NAND2_X1 U4889 ( .A1(n4364), .A2(n4348), .ZN(n4352) );
  OAI21_X1 U4890 ( .B1(n4350), .B2(n4349), .A(n4391), .ZN(n4351) );
  OAI211_X1 U4891 ( .C1(n4354), .C2(n4353), .A(n4352), .B(n4351), .ZN(n4355)
         );
  OAI21_X1 U4892 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n4373) );
  NAND2_X1 U4893 ( .A1(n4359), .A2(n4358), .ZN(n4361) );
  NAND2_X1 U4894 ( .A1(n7075), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U4895 ( .A1(n4361), .A2(n4360), .ZN(n4367) );
  MUX2_X1 U4896 ( .A(n7083), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n4366) );
  XNOR2_X1 U4897 ( .A(n4367), .B(n4366), .ZN(n4518) );
  INV_X1 U4898 ( .A(n4518), .ZN(n4363) );
  NAND2_X1 U4899 ( .A1(n4387), .A2(n4363), .ZN(n4365) );
  OAI211_X1 U4900 ( .C1(n4363), .C2(n4362), .A(n4364), .B(n4365), .ZN(n4372)
         );
  INV_X1 U4901 ( .A(n4364), .ZN(n4371) );
  INV_X1 U4902 ( .A(n4365), .ZN(n4370) );
  NAND2_X1 U4903 ( .A1(n4367), .A2(n4366), .ZN(n4369) );
  NAND2_X1 U4904 ( .A1(n7083), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U4905 ( .A(n7084), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4375) );
  XNOR2_X1 U4906 ( .A(n4376), .B(n4375), .ZN(n4517) );
  AOI222_X1 U4907 ( .A1(n4373), .A2(n4372), .B1(n4371), .B2(n4370), .C1(n4517), 
        .C2(n4437), .ZN(n4380) );
  INV_X1 U4908 ( .A(n4517), .ZN(n4378) );
  NAND2_X1 U4909 ( .A1(n4383), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4382) );
  AOI21_X1 U4910 ( .B1(n4378), .B2(n4522), .A(n4377), .ZN(n4379) );
  OAI22_X1 U4911 ( .A1(n4380), .A2(n4379), .B1(n4391), .B2(n4522), .ZN(n4381)
         );
  AOI21_X1 U4912 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7115), .A(n4381), 
        .ZN(n4389) );
  NAND2_X1 U4913 ( .A1(n4382), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4386) );
  INV_X1 U4914 ( .A(n4383), .ZN(n4384) );
  NAND2_X1 U4915 ( .A1(n4384), .A2(n7097), .ZN(n4385) );
  NAND2_X1 U4916 ( .A1(n4387), .A2(n4521), .ZN(n4388) );
  NAND2_X1 U4917 ( .A1(n4389), .A2(n4388), .ZN(n4393) );
  INV_X1 U4918 ( .A(n4521), .ZN(n4390) );
  NAND3_X1 U4919 ( .A1(n4697), .A2(n4870), .A3(n4501), .ZN(n4643) );
  INV_X1 U4920 ( .A(n4643), .ZN(n4394) );
  NAND3_X1 U4921 ( .A1(n4394), .A2(n5969), .A3(n3503), .ZN(n4534) );
  NAND2_X1 U4922 ( .A1(n5618), .A2(n4396), .ZN(n6799) );
  NAND2_X1 U4923 ( .A1(n6799), .A2(n7115), .ZN(n4397) );
  NAND2_X1 U4924 ( .A1(n7115), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4399) );
  INV_X1 U4925 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5617) );
  NAND2_X1 U4926 ( .A1(n5617), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U4927 ( .A1(n4399), .A2(n4398), .ZN(n4689) );
  NAND2_X1 U4928 ( .A1(n5327), .A2(n5488), .ZN(n6783) );
  INV_X2 U4929 ( .A(n6894), .ZN(n6906) );
  NAND2_X1 U4930 ( .A1(n6906), .A2(REIP_REG_28__SCAN_IN), .ZN(n6511) );
  OAI21_X1 U4931 ( .B1(n6753), .B2(n5863), .A(n6511), .ZN(n4400) );
  AOI21_X1 U4932 ( .B1(n6477), .B2(n5856), .A(n4400), .ZN(n4490) );
  OR2_X2 U4933 ( .A1(n4450), .A2(n4402), .ZN(n6474) );
  INV_X1 U4934 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4491) );
  XNOR2_X1 U4935 ( .A(n6428), .B(n4491), .ZN(n4488) );
  NAND2_X1 U4936 ( .A1(n4409), .A2(n4416), .ZN(n4422) );
  INV_X1 U4937 ( .A(n4421), .ZN(n4403) );
  NAND2_X1 U4938 ( .A1(n4422), .A2(n4403), .ZN(n4433) );
  NAND2_X1 U4939 ( .A1(n4433), .A2(n4431), .ZN(n4440) );
  INV_X1 U4940 ( .A(n4439), .ZN(n4404) );
  NOR2_X1 U4941 ( .A1(n4440), .A2(n4404), .ZN(n4406) );
  NAND2_X1 U4942 ( .A1(n4406), .A2(n4405), .ZN(n4460) );
  OAI211_X1 U4943 ( .C1(n4406), .C2(n4405), .A(n4460), .B(n7144), .ZN(n4407)
         );
  INV_X1 U4944 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4963) );
  XNOR2_X1 U4945 ( .A(n4447), .B(n4963), .ZN(n4961) );
  INV_X1 U4946 ( .A(n4416), .ZN(n4410) );
  XNOR2_X1 U4947 ( .A(n4410), .B(n4409), .ZN(n4413) );
  INV_X1 U4948 ( .A(n4411), .ZN(n4412) );
  AOI21_X1 U4949 ( .B1(n7144), .B2(n4413), .A(n4412), .ZN(n4414) );
  NAND2_X1 U4950 ( .A1(n4863), .A2(n4437), .ZN(n4419) );
  NAND2_X1 U4951 ( .A1(n5503), .A2(n4501), .ZN(n4423) );
  OAI21_X1 U4952 ( .B1(n4415), .B2(n4416), .A(n4423), .ZN(n4417) );
  INV_X1 U4953 ( .A(n4417), .ZN(n4418) );
  NAND2_X1 U4954 ( .A1(n4419), .A2(n4418), .ZN(n4690) );
  AND2_X1 U4955 ( .A1(n4690), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4727)
         );
  NAND2_X1 U4956 ( .A1(n4726), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4428)
         );
  NAND2_X1 U4957 ( .A1(n4426), .A2(n4428), .ZN(n4420) );
  NAND2_X1 U4958 ( .A1(n4420), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6741)
         );
  XNOR2_X1 U4959 ( .A(n4422), .B(n4421), .ZN(n4424) );
  OAI21_X1 U4960 ( .B1(n4424), .B2(n4415), .A(n4423), .ZN(n4425) );
  AOI21_X2 U4961 ( .B1(n4861), .B2(n4437), .A(n4425), .ZN(n6744) );
  NAND2_X1 U4962 ( .A1(n6741), .A2(n6744), .ZN(n4430) );
  INV_X1 U4963 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4427) );
  AND2_X1 U4964 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  NAND2_X1 U4965 ( .A1(n4426), .A2(n4429), .ZN(n6742) );
  INV_X1 U4966 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4811) );
  INV_X1 U4967 ( .A(n4431), .ZN(n4432) );
  XNOR2_X1 U4968 ( .A(n4433), .B(n4432), .ZN(n4434) );
  NAND2_X1 U4969 ( .A1(n4435), .A2(n4811), .ZN(n4802) );
  NAND2_X1 U4970 ( .A1(n4436), .A2(n4802), .ZN(n4843) );
  NAND2_X1 U4971 ( .A1(n4438), .A2(n4437), .ZN(n4443) );
  XNOR2_X1 U4972 ( .A(n4440), .B(n4439), .ZN(n4441) );
  NAND2_X1 U4973 ( .A1(n4441), .A2(n7144), .ZN(n4442) );
  NAND2_X1 U4974 ( .A1(n4443), .A2(n4442), .ZN(n4444) );
  XNOR2_X1 U4975 ( .A(n4444), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4844)
         );
  INV_X1 U4976 ( .A(n4444), .ZN(n4446) );
  INV_X1 U4977 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4445) );
  OAI22_X1 U4978 ( .A1(n4843), .A2(n4844), .B1(n4446), .B2(n4445), .ZN(n4960)
         );
  NAND2_X1 U4979 ( .A1(n4961), .A2(n4960), .ZN(n4449) );
  NAND2_X1 U4980 ( .A1(n4447), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4448)
         );
  NAND2_X1 U4981 ( .A1(n4449), .A2(n4448), .ZN(n6754) );
  XNOR2_X1 U4982 ( .A(n4460), .B(n4461), .ZN(n4451) );
  AND2_X1 U4983 ( .A1(n4451), .A2(n7144), .ZN(n4452) );
  AOI21_X1 U4984 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(n4455) );
  INV_X1 U4985 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U4986 ( .A1(n4455), .A2(n6857), .ZN(n6756) );
  NAND2_X1 U4987 ( .A1(n6754), .A2(n6756), .ZN(n4457) );
  INV_X1 U4988 ( .A(n4455), .ZN(n4456) );
  NAND2_X1 U4989 ( .A1(n4456), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6755)
         );
  OR2_X1 U4990 ( .A1(n4459), .A2(n4458), .ZN(n4465) );
  INV_X1 U4991 ( .A(n4460), .ZN(n4462) );
  NAND2_X1 U4992 ( .A1(n4462), .A2(n4461), .ZN(n4470) );
  XNOR2_X1 U4993 ( .A(n4470), .B(n4468), .ZN(n4463) );
  NAND2_X1 U4994 ( .A1(n4463), .A2(n7144), .ZN(n4464) );
  NAND2_X1 U4995 ( .A1(n4465), .A2(n4464), .ZN(n4466) );
  INV_X1 U4996 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6866) );
  XNOR2_X1 U4997 ( .A(n4466), .B(n6866), .ZN(n6764) );
  NAND2_X1 U4998 ( .A1(n6761), .A2(n6764), .ZN(n6762) );
  NAND2_X1 U4999 ( .A1(n4466), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4467)
         );
  NAND2_X1 U5000 ( .A1(n6762), .A2(n4467), .ZN(n5464) );
  NAND2_X1 U5001 ( .A1(n7144), .A2(n4468), .ZN(n4469) );
  OR2_X1 U5002 ( .A1(n4470), .A2(n4469), .ZN(n4471) );
  NAND2_X1 U5003 ( .A1(n6474), .A2(n4471), .ZN(n4472) );
  INV_X1 U5004 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6862) );
  XNOR2_X1 U5005 ( .A(n4472), .B(n6862), .ZN(n5467) );
  NAND2_X1 U5006 ( .A1(n5464), .A2(n5467), .ZN(n5465) );
  NAND2_X1 U5007 ( .A1(n4472), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4473)
         );
  XNOR2_X1 U5008 ( .A(n6428), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5560)
         );
  INV_X1 U5009 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6869) );
  OR2_X1 U5010 ( .A1(n6463), .A2(n6869), .ZN(n4474) );
  INV_X1 U5011 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5760) );
  INV_X1 U5012 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4571) );
  XNOR2_X1 U5013 ( .A(n6428), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5731)
         );
  INV_X1 U5014 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5015 ( .A1(n6474), .A2(n4576), .ZN(n4475) );
  AND2_X1 U5016 ( .A1(n6463), .A2(n6802), .ZN(n5827) );
  INV_X1 U5017 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5777) );
  NOR2_X1 U5018 ( .A1(n6474), .A2(n5777), .ZN(n5770) );
  NAND2_X1 U5019 ( .A1(n6474), .A2(n5777), .ZN(n5769) );
  INV_X1 U5020 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4477) );
  NOR2_X1 U5021 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U5022 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5023 ( .A1(n6474), .A2(n4657), .ZN(n4480) );
  NAND2_X1 U5024 ( .A1(n4481), .A2(n4480), .ZN(n4483) );
  INV_X1 U5025 ( .A(n4483), .ZN(n4482) );
  AND2_X1 U5026 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6562) );
  AND2_X1 U5027 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U5028 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U5029 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6545) );
  NOR2_X1 U5030 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6564) );
  INV_X1 U5031 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6542) );
  XNOR2_X1 U5032 ( .A(n6428), .B(n6542), .ZN(n6421) );
  INV_X1 U5033 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U5034 ( .A1(n6474), .A2(n6529), .ZN(n6406) );
  NAND2_X1 U5035 ( .A1(n6407), .A2(n6406), .ZN(n4486) );
  NAND2_X1 U5036 ( .A1(n4486), .A2(n6529), .ZN(n6398) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6399) );
  OAI22_X2 U5038 ( .A1(n4492), .A2(n6428), .B1(n6399), .B2(n6397), .ZN(n4487)
         );
  AOI21_X1 U5039 ( .B1(n4488), .B2(n4487), .A(n6390), .ZN(n6517) );
  NAND3_X1 U5040 ( .A1(n3548), .A2(n4490), .A3(n4489), .ZN(U2958) );
  INV_X1 U5041 ( .A(n6397), .ZN(n4493) );
  AND2_X1 U5042 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6501) );
  AND2_X1 U5043 ( .A1(n6501), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6493)
         );
  INV_X1 U5044 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U5045 ( .A1(n6493), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4661) );
  INV_X1 U5046 ( .A(n4661), .ZN(n4495) );
  INV_X1 U5047 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4780) );
  XNOR2_X1 U5048 ( .A(n4496), .B(n4780), .ZN(n5919) );
  NAND2_X1 U5049 ( .A1(n4880), .A2(n6791), .ZN(n5491) );
  AND2_X1 U5050 ( .A1(n5491), .A2(n7143), .ZN(n4758) );
  AOI21_X1 U5051 ( .B1(n4697), .B2(n3680), .A(n4525), .ZN(n4499) );
  AOI21_X1 U5052 ( .B1(n4498), .B2(n4758), .A(n4499), .ZN(n4530) );
  NAND3_X1 U5053 ( .A1(n5980), .A2(n4512), .A3(n3687), .ZN(n4527) );
  NAND2_X1 U5054 ( .A1(n4500), .A2(n4684), .ZN(n4505) );
  NAND3_X1 U5055 ( .A1(n4502), .A2(n4697), .A3(n3694), .ZN(n4504) );
  AND2_X1 U5056 ( .A1(n5503), .A2(n3687), .ZN(n5981) );
  OAI21_X1 U5057 ( .B1(n4870), .B2(n3680), .A(n5981), .ZN(n4503) );
  NAND3_X1 U5058 ( .A1(n4505), .A2(n4504), .A3(n4503), .ZN(n4507) );
  NOR2_X1 U5059 ( .A1(n4507), .A2(n4506), .ZN(n4737) );
  INV_X1 U5060 ( .A(n4508), .ZN(n4733) );
  NAND2_X1 U5061 ( .A1(n4733), .A2(n5503), .ZN(n4509) );
  AND2_X1 U5062 ( .A1(n4772), .A2(n4509), .ZN(n4510) );
  NAND2_X1 U5063 ( .A1(n4737), .A2(n4510), .ZN(n4640) );
  NAND2_X1 U5064 ( .A1(n4512), .A2(n4511), .ZN(n4532) );
  AND2_X1 U5065 ( .A1(n4532), .A2(n4643), .ZN(n4513) );
  NAND2_X1 U5066 ( .A1(n4516), .A2(n5974), .ZN(n4762) );
  NOR3_X1 U5067 ( .A1(n4519), .A2(n4518), .A3(n4517), .ZN(n4520) );
  OR2_X1 U5068 ( .A1(n4521), .A2(n4520), .ZN(n4523) );
  NAND2_X1 U5069 ( .A1(n4523), .A2(n4522), .ZN(n4669) );
  NAND2_X1 U5070 ( .A1(n3687), .A2(n6791), .ZN(n4524) );
  NAND4_X1 U5071 ( .A1(n4669), .A2(n4525), .A3(n7143), .A4(n4524), .ZN(n4526)
         );
  NAND3_X1 U5072 ( .A1(n4527), .A2(n4762), .A3(n4526), .ZN(n4528) );
  NAND2_X1 U5073 ( .A1(n4528), .A2(n5984), .ZN(n4529) );
  INV_X1 U5074 ( .A(n4532), .ZN(n4533) );
  NAND2_X1 U5075 ( .A1(n4533), .A2(n5485), .ZN(n4754) );
  AND2_X1 U5076 ( .A1(n4754), .A2(n4534), .ZN(n5973) );
  INV_X1 U5077 ( .A(n4638), .ZN(n4535) );
  AOI22_X1 U5078 ( .A1(n5494), .A2(n4498), .B1(n4535), .B2(n3737), .ZN(n4536)
         );
  NAND3_X1 U5079 ( .A1(n3429), .A2(n5973), .A3(n4536), .ZN(n4537) );
  NAND2_X1 U5080 ( .A1(n5919), .A2(n6920), .ZN(n4667) );
  OAI21_X1 U5081 ( .B1(n4684), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4538), 
        .ZN(n4539) );
  INV_X1 U5082 ( .A(n4539), .ZN(n4542) );
  MUX2_X1 U5083 ( .A(n4619), .B(n4630), .S(EBX_REG_1__SCAN_IN), .Z(n4540) );
  INV_X1 U5084 ( .A(n4540), .ZN(n4541) );
  NAND2_X1 U5085 ( .A1(n4542), .A2(n4541), .ZN(n4544) );
  INV_X1 U5086 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4543) );
  OAI22_X1 U5087 ( .A1(n4622), .A2(n4543), .B1(n4624), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4685) );
  XNOR2_X1 U5088 ( .A(n4544), .B(n4685), .ZN(n5589) );
  NAND2_X1 U5089 ( .A1(n5589), .A2(n5494), .ZN(n4546) );
  INV_X1 U5090 ( .A(n4544), .ZN(n4545) );
  NAND2_X1 U5091 ( .A1(n4546), .A2(n4545), .ZN(n4722) );
  MUX2_X1 U5092 ( .A(n4619), .B(n4630), .S(EBX_REG_2__SCAN_IN), .Z(n4547) );
  INV_X1 U5093 ( .A(n4547), .ZN(n4548) );
  NAND2_X1 U5094 ( .A1(n4548), .A2(n3558), .ZN(n4721) );
  INV_X1 U5095 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U5096 ( .A1(n4607), .A2(n6944), .ZN(n4552) );
  NAND2_X1 U5097 ( .A1(n4622), .A2(n4811), .ZN(n4550) );
  OAI211_X1 U5098 ( .C1(n4633), .C2(EBX_REG_3__SCAN_IN), .A(n4624), .B(n4550), 
        .ZN(n4551) );
  AND2_X1 U5099 ( .A1(n4552), .A2(n4551), .ZN(n4797) );
  MUX2_X1 U5100 ( .A(n4619), .B(n4630), .S(EBX_REG_4__SCAN_IN), .Z(n4553) );
  INV_X1 U5101 ( .A(n4553), .ZN(n4554) );
  NAND2_X1 U5102 ( .A1(n4554), .A2(n3557), .ZN(n4818) );
  INV_X1 U5103 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5263) );
  MUX2_X1 U5104 ( .A(n4630), .B(n4619), .S(n5263), .Z(n4556) );
  NOR2_X1 U5105 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4555)
         );
  NOR2_X1 U5106 ( .A1(n4556), .A2(n4555), .ZN(n5259) );
  NAND2_X1 U5107 ( .A1(n4622), .A2(n4963), .ZN(n4557) );
  OAI211_X1 U5108 ( .C1(n4633), .C2(EBX_REG_5__SCAN_IN), .A(n4624), .B(n4557), 
        .ZN(n4558) );
  OAI21_X1 U5109 ( .B1(n4626), .B2(EBX_REG_5__SCAN_IN), .A(n4558), .ZN(n5260)
         );
  AND2_X1 U5110 ( .A1(n5259), .A2(n5260), .ZN(n4559) );
  INV_X1 U5111 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5463) );
  MUX2_X1 U5112 ( .A(n4630), .B(n4619), .S(n5463), .Z(n4561) );
  NOR2_X1 U5113 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4560)
         );
  NOR2_X1 U5114 ( .A1(n4561), .A2(n4560), .ZN(n5458) );
  NAND2_X1 U5115 ( .A1(n4622), .A2(n6866), .ZN(n4562) );
  OAI211_X1 U5116 ( .C1(n4633), .C2(EBX_REG_7__SCAN_IN), .A(n4624), .B(n4562), 
        .ZN(n4563) );
  OAI21_X1 U5117 ( .B1(n4626), .B2(EBX_REG_7__SCAN_IN), .A(n4563), .ZN(n5459)
         );
  AND2_X1 U5118 ( .A1(n5458), .A2(n5459), .ZN(n4564) );
  INV_X1 U5119 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U5120 ( .A1(n4607), .A2(n5609), .ZN(n4567) );
  NAND2_X1 U5121 ( .A1(n4622), .A2(n6869), .ZN(n4565) );
  OAI211_X1 U5122 ( .C1(n4633), .C2(EBX_REG_9__SCAN_IN), .A(n4624), .B(n4565), 
        .ZN(n4566) );
  AND2_X1 U5123 ( .A1(n4567), .A2(n4566), .ZN(n5570) );
  MUX2_X1 U5124 ( .A(n4619), .B(n4630), .S(EBX_REG_10__SCAN_IN), .Z(n4569) );
  INV_X1 U5125 ( .A(n4569), .ZN(n4570) );
  NAND2_X1 U5126 ( .A1(n4570), .A2(n3556), .ZN(n5576) );
  NAND2_X1 U5127 ( .A1(n4622), .A2(n4571), .ZN(n4572) );
  OAI211_X1 U5128 ( .C1(n4633), .C2(EBX_REG_11__SCAN_IN), .A(n4624), .B(n4572), 
        .ZN(n4573) );
  OAI21_X1 U5129 ( .B1(n4626), .B2(EBX_REG_11__SCAN_IN), .A(n4573), .ZN(n5703)
         );
  NAND2_X1 U5130 ( .A1(n5704), .A2(n5703), .ZN(n5744) );
  INV_X1 U5131 ( .A(n4619), .ZN(n4599) );
  NAND2_X1 U5132 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4574) );
  OAI211_X1 U5133 ( .C1(n4633), .C2(EBX_REG_12__SCAN_IN), .A(n4622), .B(n4574), 
        .ZN(n4575) );
  OAI21_X1 U5134 ( .B1(n4599), .B2(EBX_REG_12__SCAN_IN), .A(n4575), .ZN(n5743)
         );
  INV_X1 U5135 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U5136 ( .A1(n4607), .A2(n5786), .ZN(n4579) );
  NAND2_X1 U5137 ( .A1(n4622), .A2(n4576), .ZN(n4577) );
  OAI211_X1 U5138 ( .C1(n4633), .C2(EBX_REG_13__SCAN_IN), .A(n4624), .B(n4577), 
        .ZN(n4578) );
  MUX2_X1 U5139 ( .A(n4619), .B(n4630), .S(EBX_REG_14__SCAN_IN), .Z(n4581) );
  NOR2_X1 U5140 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4580)
         );
  NOR2_X1 U5141 ( .A1(n4581), .A2(n4580), .ZN(n5811) );
  NAND2_X1 U5142 ( .A1(n4622), .A2(n5777), .ZN(n4582) );
  OAI211_X1 U5143 ( .C1(n4633), .C2(EBX_REG_15__SCAN_IN), .A(n4624), .B(n4582), 
        .ZN(n4583) );
  OAI21_X1 U5144 ( .B1(n4626), .B2(EBX_REG_15__SCAN_IN), .A(n4583), .ZN(n5772)
         );
  MUX2_X1 U5145 ( .A(n4619), .B(n4630), .S(EBX_REG_16__SCAN_IN), .Z(n4584) );
  INV_X1 U5146 ( .A(n4584), .ZN(n4586) );
  INV_X1 U5147 ( .A(n4684), .ZN(n4629) );
  NAND2_X1 U5148 ( .A1(n4629), .A2(n4477), .ZN(n4585) );
  NAND2_X1 U5149 ( .A1(n4586), .A2(n4585), .ZN(n6106) );
  INV_X1 U5150 ( .A(EBX_REG_17__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U5151 ( .A1(n4607), .A2(n7024), .ZN(n4589) );
  INV_X1 U5152 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U5153 ( .A1(n4622), .A2(n6917), .ZN(n4587) );
  OAI211_X1 U5154 ( .C1(n4633), .C2(EBX_REG_17__SCAN_IN), .A(n4624), .B(n4587), 
        .ZN(n4588) );
  INV_X1 U5155 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6149) );
  MUX2_X1 U5156 ( .A(n4630), .B(n4619), .S(n6149), .Z(n4591) );
  NOR2_X1 U5157 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4590)
         );
  NOR2_X1 U5158 ( .A1(n4591), .A2(n4590), .ZN(n6094) );
  INV_X1 U5159 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U5160 ( .A1(n4607), .A2(n6145), .ZN(n4595) );
  NAND2_X1 U5161 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5162 ( .A1(n4622), .A2(n4592), .ZN(n4593) );
  OAI21_X1 U5163 ( .B1(n4633), .B2(EBX_REG_19__SCAN_IN), .A(n4593), .ZN(n4594)
         );
  AND2_X1 U5164 ( .A1(n4595), .A2(n4594), .ZN(n6141) );
  NAND2_X1 U5165 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4597) );
  OAI211_X1 U5166 ( .C1(n4633), .C2(EBX_REG_20__SCAN_IN), .A(n4622), .B(n4597), 
        .ZN(n4598) );
  OAI21_X1 U5167 ( .B1(n4599), .B2(EBX_REG_20__SCAN_IN), .A(n4598), .ZN(n6080)
         );
  INV_X1 U5168 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U5169 ( .A1(n4607), .A2(n6134), .ZN(n4603) );
  NAND2_X1 U5170 ( .A1(n4624), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U5171 ( .A1(n4622), .A2(n4600), .ZN(n4601) );
  OAI21_X1 U5172 ( .B1(n4633), .B2(EBX_REG_21__SCAN_IN), .A(n4601), .ZN(n4602)
         );
  MUX2_X1 U5173 ( .A(n4619), .B(n4630), .S(EBX_REG_22__SCAN_IN), .Z(n4605) );
  NOR2_X1 U5174 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4604)
         );
  NOR2_X1 U5175 ( .A1(n4605), .A2(n4604), .ZN(n6066) );
  INV_X1 U5176 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5177 ( .A1(n4607), .A2(n4606), .ZN(n4610) );
  INV_X1 U5178 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U5179 ( .A1(n4622), .A2(n6560), .ZN(n4608) );
  OAI211_X1 U5180 ( .C1(n4633), .C2(EBX_REG_23__SCAN_IN), .A(n4624), .B(n4608), 
        .ZN(n4609) );
  INV_X1 U5181 ( .A(n4611), .ZN(n6059) );
  MUX2_X1 U5182 ( .A(n4619), .B(n4630), .S(EBX_REG_24__SCAN_IN), .Z(n4612) );
  INV_X1 U5183 ( .A(n4612), .ZN(n4614) );
  INV_X1 U5184 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U5185 ( .A1(n4629), .A2(n6546), .ZN(n4613) );
  NAND2_X1 U5186 ( .A1(n4614), .A2(n4613), .ZN(n6041) );
  NAND2_X1 U5187 ( .A1(n4622), .A2(n6542), .ZN(n4615) );
  OAI211_X1 U5188 ( .C1(n4633), .C2(EBX_REG_25__SCAN_IN), .A(n4624), .B(n4615), 
        .ZN(n4616) );
  OAI21_X1 U5189 ( .B1(n4626), .B2(EBX_REG_25__SCAN_IN), .A(n4616), .ZN(n6025)
         );
  MUX2_X1 U5190 ( .A(n4619), .B(n4630), .S(EBX_REG_26__SCAN_IN), .Z(n4618) );
  NOR2_X1 U5191 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4617)
         );
  NOR2_X1 U5192 ( .A1(n4618), .A2(n4617), .ZN(n6015) );
  MUX2_X1 U5193 ( .A(n4619), .B(n4630), .S(EBX_REG_28__SCAN_IN), .Z(n4621) );
  NOR2_X1 U5194 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4620)
         );
  NOR2_X1 U5195 ( .A1(n4621), .A2(n4620), .ZN(n5847) );
  NAND2_X1 U5196 ( .A1(n4622), .A2(n6399), .ZN(n4623) );
  OAI211_X1 U5197 ( .C1(n4633), .C2(EBX_REG_27__SCAN_IN), .A(n4624), .B(n4623), 
        .ZN(n4625) );
  OAI21_X1 U5198 ( .B1(n4626), .B2(EBX_REG_27__SCAN_IN), .A(n4625), .ZN(n6000)
         );
  OR2_X1 U5199 ( .A1(n4633), .A2(EBX_REG_29__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5200 ( .B1(n4684), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4631), 
        .ZN(n5945) );
  MUX2_X1 U5201 ( .A(n5945), .B(n4631), .S(n4630), .Z(n4627) );
  INV_X1 U5202 ( .A(n4627), .ZN(n5988) );
  INV_X1 U5203 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5204 ( .A1(n4629), .A2(n4494), .B1(n5494), .B2(n4628), .ZN(n5947)
         );
  NAND2_X1 U5205 ( .A1(n5988), .A2(n5947), .ZN(n4632) );
  OAI21_X1 U5206 ( .B1(n5989), .B2(n4632), .A(n5944), .ZN(n4636) );
  OAI22_X1 U5207 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4684), .B1(n4633), .B2(EBX_REG_31__SCAN_IN), .ZN(n4634) );
  INV_X1 U5208 ( .A(n4634), .ZN(n4635) );
  INV_X1 U5209 ( .A(n4498), .ZN(n4637) );
  OAI21_X1 U5210 ( .B1(n4638), .B2(n3737), .A(n7102), .ZN(n4639) );
  NOR2_X1 U5211 ( .A1(n5974), .A2(n4880), .ZN(n7071) );
  INV_X1 U5212 ( .A(n4640), .ZN(n4641) );
  NAND2_X1 U5213 ( .A1(n4641), .A2(n4735), .ZN(n4642) );
  OR2_X1 U5214 ( .A1(n4643), .A2(n4880), .ZN(n4644) );
  INV_X1 U5215 ( .A(n6493), .ZN(n4652) );
  AND2_X1 U5216 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4660) );
  AOI21_X1 U5217 ( .B1(n4709), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6818), 
        .ZN(n4653) );
  NAND2_X1 U5218 ( .A1(n4653), .A2(n4965), .ZN(n6922) );
  NAND2_X1 U5219 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6908) );
  INV_X1 U5220 ( .A(n6908), .ZN(n4651) );
  NAND2_X1 U5221 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U5222 ( .A1(n4576), .A2(n6889), .ZN(n6803) );
  NAND2_X1 U5223 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6803), .ZN(n4656) );
  INV_X1 U5224 ( .A(n4656), .ZN(n4650) );
  INV_X1 U5225 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5226 ( .A1(n4709), .A2(n4781), .ZN(n4647) );
  OR2_X1 U5227 ( .A1(n4645), .A2(n6906), .ZN(n4646) );
  NAND2_X1 U5228 ( .A1(n4647), .A2(n4646), .ZN(n6850) );
  NOR2_X1 U5229 ( .A1(n6862), .A2(n6866), .ZN(n6873) );
  NAND3_X1 U5230 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6873), .ZN(n4648) );
  NAND2_X1 U5231 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6828) );
  NOR2_X1 U5232 ( .A1(n4963), .A2(n6828), .ZN(n6832) );
  NAND4_X1 U5233 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .A4(n6832), .ZN(n6847) );
  NOR2_X1 U5234 ( .A1(n4648), .A2(n6847), .ZN(n4654) );
  AOI21_X1 U5235 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6839) );
  NOR2_X1 U5236 ( .A1(n6839), .A2(n6828), .ZN(n4962) );
  NAND3_X1 U5237 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4962), .ZN(n6852) );
  NOR2_X1 U5238 ( .A1(n4648), .A2(n6852), .ZN(n4655) );
  OAI22_X1 U5239 ( .A1(n4654), .A2(n6848), .B1(n4655), .B2(n4965), .ZN(n4649)
         );
  OAI21_X1 U5240 ( .B1(n6874), .B2(n4650), .A(n6901), .ZN(n6907) );
  INV_X1 U5241 ( .A(n6907), .ZN(n5774) );
  OAI21_X1 U5242 ( .B1(n6874), .B2(n4651), .A(n5774), .ZN(n6602) );
  AOI21_X1 U5243 ( .B1(n4657), .B2(n6816), .A(n6602), .ZN(n6601) );
  OAI21_X1 U5244 ( .B1(n3458), .B2(n6874), .A(n6601), .ZN(n6552) );
  AOI21_X1 U5245 ( .B1(n4658), .B2(n6922), .A(n6552), .ZN(n6544) );
  OAI21_X1 U5246 ( .B1(n6874), .B2(n4660), .A(n6544), .ZN(n6521) );
  AOI21_X1 U5247 ( .B1(n4652), .B2(n6816), .A(n6521), .ZN(n6506) );
  OAI21_X1 U5248 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6874), .A(n6506), 
        .ZN(n4663) );
  INV_X1 U5249 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5933) );
  NOR2_X1 U5250 ( .A1(n6894), .A2(n5933), .ZN(n5922) );
  INV_X1 U5251 ( .A(n4653), .ZN(n6842) );
  NAND3_X1 U5252 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6909), .ZN(n6916) );
  INV_X1 U5253 ( .A(n4658), .ZN(n4659) );
  NAND2_X1 U5254 ( .A1(n6535), .A2(n4660), .ZN(n6518) );
  NOR3_X1 U5255 ( .A1(n6518), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4661), 
        .ZN(n4662) );
  AOI211_X1 U5256 ( .C1(n4663), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5922), .B(n4662), .ZN(n4664) );
  NAND2_X1 U5257 ( .A1(n4667), .A2(n4666), .ZN(U2987) );
  INV_X1 U5258 ( .A(n4668), .ZN(n5972) );
  INV_X1 U5259 ( .A(n4755), .ZN(n4670) );
  AOI22_X1 U5260 ( .A1(n5980), .A2(n3707), .B1(n5972), .B2(n4670), .ZN(n5983)
         );
  AND2_X1 U5261 ( .A1(n5983), .A2(n5984), .ZN(n4672) );
  INV_X1 U5262 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6319) );
  NOR2_X1 U5263 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6794) );
  NAND3_X1 U5264 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6794), .A3(n7110), .ZN(
        n4671) );
  OAI21_X1 U5265 ( .B1(n4672), .B2(n6319), .A(n4671), .ZN(U2790) );
  NAND2_X1 U5266 ( .A1(n4755), .A2(n5984), .ZN(n5481) );
  INV_X1 U5267 ( .A(n5481), .ZN(n4674) );
  INV_X1 U5268 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6175) );
  OAI211_X1 U5269 ( .C1(n4674), .C2(n6175), .A(n7141), .B(n6783), .ZN(U2788)
         );
  AND2_X1 U5270 ( .A1(n4761), .A2(n5984), .ZN(n4675) );
  NAND2_X1 U5271 ( .A1(n5980), .A2(n4675), .ZN(n4680) );
  INV_X1 U5272 ( .A(n4676), .ZN(n4678) );
  INV_X1 U5273 ( .A(n3779), .ZN(n6162) );
  NAND4_X1 U5274 ( .A1(n6162), .A2(n3635), .A3(n5984), .A4(n3778), .ZN(n5478)
         );
  INV_X1 U5275 ( .A(n5478), .ZN(n4677) );
  NAND3_X1 U5276 ( .A1(n4678), .A2(n4677), .A3(n5494), .ZN(n4679) );
  NAND2_X2 U5277 ( .A1(n6150), .A2(n3779), .ZN(n6151) );
  OAI21_X1 U5278 ( .B1(n4682), .B2(n4681), .A(n4716), .ZN(n5595) );
  XNOR2_X1 U5279 ( .A(n5589), .B(n5494), .ZN(n6813) );
  AOI22_X1 U5280 ( .A1(n6160), .A2(n6813), .B1(n6159), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4683) );
  OAI21_X1 U5281 ( .B1(n6151), .B2(n5595), .A(n4683), .ZN(U2858) );
  NOR2_X1 U5282 ( .A1(n4684), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4686)
         );
  OR2_X1 U5283 ( .A1(n4686), .A2(n4685), .ZN(n5497) );
  XNOR2_X1 U5284 ( .A(n4688), .B(n4687), .ZN(n5509) );
  OAI222_X1 U5285 ( .A1(n5497), .A2(n6148), .B1(n6150), .B2(n4543), .C1(n6151), 
        .C2(n5509), .ZN(U2859) );
  OAI21_X1 U5286 ( .B1(n6772), .B2(n4689), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4693) );
  INV_X1 U5287 ( .A(n4690), .ZN(n4691) );
  AOI21_X1 U5288 ( .B1(n4691), .B2(n4781), .A(n4727), .ZN(n4713) );
  AND2_X1 U5289 ( .A1(n6906), .A2(REIP_REG_0__SCAN_IN), .ZN(n4712) );
  AOI21_X1 U5290 ( .B1(n6774), .B2(n4713), .A(n4712), .ZN(n4692) );
  OAI211_X1 U5291 ( .C1(n5509), .C2(n6748), .A(n4693), .B(n4692), .ZN(U2986)
         );
  INV_X1 U5292 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5293 ( .A1(n5475), .A2(n7071), .ZN(n4695) );
  NAND2_X1 U5294 ( .A1(n7145), .A2(n4695), .ZN(n4696) );
  INV_X1 U5295 ( .A(n6791), .ZN(n5982) );
  INV_X2 U5296 ( .A(n7099), .ZN(n6666) );
  NOR2_X4 U5297 ( .A1(n6666), .A2(n6635), .ZN(n6648) );
  AOI22_X1 U5298 ( .A1(n6666), .A2(UWORD_REG_7__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4699) );
  OAI21_X1 U5299 ( .B1(n4700), .B2(n4840), .A(n4699), .ZN(U2900) );
  INV_X1 U5300 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5301 ( .A1(n6666), .A2(UWORD_REG_5__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4701) );
  OAI21_X1 U5302 ( .B1(n4702), .B2(n4840), .A(n4701), .ZN(U2902) );
  INV_X1 U5303 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5304 ( .A1(n6666), .A2(UWORD_REG_8__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4703) );
  OAI21_X1 U5305 ( .B1(n4704), .B2(n4840), .A(n4703), .ZN(U2899) );
  INV_X1 U5306 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5307 ( .A1(n6666), .A2(UWORD_REG_6__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4705) );
  OAI21_X1 U5308 ( .B1(n4706), .B2(n4840), .A(n4705), .ZN(U2901) );
  INV_X1 U5309 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5310 ( .A1(n6666), .A2(UWORD_REG_9__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4707) );
  OAI21_X1 U5311 ( .B1(n4708), .B2(n4840), .A(n4707), .ZN(U2898) );
  INV_X1 U5312 ( .A(n6850), .ZN(n4808) );
  OAI21_X1 U5313 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4965), .A(n4808), 
        .ZN(n6815) );
  INV_X1 U5314 ( .A(n4709), .ZN(n4710) );
  NAND3_X1 U5315 ( .A1(n4710), .A2(n4781), .A3(n4965), .ZN(n4711) );
  OAI21_X1 U5316 ( .B1(n6815), .B2(n6818), .A(n4711), .ZN(n4715) );
  AOI21_X1 U5317 ( .B1(n6920), .B2(n4713), .A(n4712), .ZN(n4714) );
  OAI211_X1 U5318 ( .C1(n5497), .C2(n6897), .A(n4715), .B(n4714), .ZN(U3018)
         );
  INV_X1 U5319 ( .A(n4716), .ZN(n4718) );
  OAI21_X1 U5320 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n6935) );
  AOI21_X1 U5321 ( .B1(n4722), .B2(n4721), .A(n4720), .ZN(n6932) );
  AOI22_X1 U5322 ( .A1(n6160), .A2(n6932), .B1(n6159), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4723) );
  OAI21_X1 U5323 ( .B1(n6935), .B2(n6151), .A(n4723), .ZN(U2857) );
  INV_X1 U5324 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4725) );
  INV_X1 U5325 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5590) );
  NOR2_X1 U5326 ( .A1(n6894), .A2(n5590), .ZN(n6812) );
  AND2_X1 U5327 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4724)
         );
  AOI211_X1 U5328 ( .C1(n4725), .C2(n6477), .A(n6812), .B(n4724), .ZN(n4730)
         );
  XNOR2_X1 U5329 ( .A(n4727), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4728)
         );
  XNOR2_X1 U5330 ( .A(n4726), .B(n4728), .ZN(n6814) );
  NAND2_X1 U5331 ( .A1(n6814), .A2(n6774), .ZN(n4729) );
  OAI211_X1 U5332 ( .C1(n5595), .C2(n6748), .A(n4730), .B(n4729), .ZN(U2985)
         );
  OR2_X1 U5333 ( .A1(n4733), .A2(n5473), .ZN(n4734) );
  NOR2_X1 U5334 ( .A1(n4498), .A2(n4734), .ZN(n4736) );
  NAND4_X1 U5335 ( .A1(n4531), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4789)
         );
  NAND2_X1 U5336 ( .A1(n4732), .A2(n4789), .ZN(n4751) );
  AOI21_X1 U5337 ( .B1(n4738), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3845), 
        .ZN(n4739) );
  NOR2_X1 U5338 ( .A1(n4740), .A2(n4739), .ZN(n4752) );
  NAND2_X1 U5339 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4741) );
  INV_X1 U5340 ( .A(n4741), .ZN(n4742) );
  MUX2_X1 U5341 ( .A(n4742), .B(n4741), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4743) );
  NAND2_X1 U5342 ( .A1(n7071), .A2(n4743), .ZN(n4748) );
  MUX2_X1 U5343 ( .A(n4744), .B(n3845), .S(n4738), .Z(n4745) );
  INV_X1 U5344 ( .A(n4761), .ZN(n5979) );
  NAND2_X1 U5345 ( .A1(n5979), .A2(n4754), .ZN(n4774) );
  OAI21_X1 U5346 ( .B1(n4746), .B2(n4745), .A(n4774), .ZN(n4747) );
  OAI211_X1 U5347 ( .C1(n4752), .C2(n4772), .A(n4748), .B(n4747), .ZN(n4749)
         );
  INV_X1 U5348 ( .A(n4749), .ZN(n4750) );
  NAND2_X1 U5349 ( .A1(n4751), .A2(n4750), .ZN(n4890) );
  INV_X1 U5350 ( .A(n4752), .ZN(n4753) );
  AOI22_X1 U5351 ( .A1(n4890), .A2(n6619), .B1(n4855), .B2(n4753), .ZN(n4769)
         );
  OR2_X1 U5352 ( .A1(n5980), .A2(n4754), .ZN(n4757) );
  NAND3_X1 U5353 ( .A1(n4755), .A2(n4880), .A3(n7143), .ZN(n4756) );
  INV_X1 U5354 ( .A(n5476), .ZN(n4767) );
  OAI21_X1 U5355 ( .B1(n4668), .B2(n5982), .A(n4758), .ZN(n4759) );
  INV_X1 U5356 ( .A(n4759), .ZN(n4760) );
  OAI21_X1 U5357 ( .B1(n7071), .B2(n4498), .A(n4760), .ZN(n4764) );
  NAND2_X1 U5358 ( .A1(n5980), .A2(n4761), .ZN(n4763) );
  OAI211_X1 U5359 ( .C1(n5980), .C2(n4764), .A(n4763), .B(n4762), .ZN(n4765)
         );
  INV_X1 U5360 ( .A(n4765), .ZN(n4766) );
  INV_X1 U5361 ( .A(n7077), .ZN(n4898) );
  INV_X1 U5362 ( .A(FLUSH_REG_SCAN_IN), .ZN(n4906) );
  NAND2_X1 U5363 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n5179) );
  NOR2_X1 U5364 ( .A1(n7115), .A2(n5179), .ZN(n4907) );
  INV_X1 U5365 ( .A(n4907), .ZN(n7109) );
  OAI22_X1 U5366 ( .A1(n4898), .A2(n7120), .B1(n4906), .B2(n7109), .ZN(n7066)
         );
  NAND2_X1 U5367 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6627), .ZN(n4768) );
  OAI21_X1 U5368 ( .B1(n4769), .B2(n6627), .A(n4768), .ZN(U3456) );
  INV_X1 U5369 ( .A(n4789), .ZN(n6617) );
  OR2_X1 U5370 ( .A1(n4771), .A2(n6617), .ZN(n4779) );
  XNOR2_X1 U5371 ( .A(n3727), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4777)
         );
  INV_X1 U5372 ( .A(n4772), .ZN(n4775) );
  XNOR2_X1 U5373 ( .A(n4738), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4773)
         );
  MUX2_X1 U5374 ( .A(n4775), .B(n4774), .S(n4773), .Z(n4776) );
  AOI21_X1 U5375 ( .B1(n7071), .B2(n4777), .A(n4776), .ZN(n4778) );
  NAND2_X1 U5376 ( .A1(n4779), .A2(n4778), .ZN(n4891) );
  INV_X1 U5377 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U5378 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4780), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6817), .ZN(n6620) );
  NOR2_X1 U5379 ( .A1(n5488), .A2(n4781), .ZN(n6621) );
  INV_X1 U5380 ( .A(n6621), .ZN(n4783) );
  NAND3_X1 U5381 ( .A1(n4738), .A2(n4855), .A3(n3727), .ZN(n4782) );
  OAI21_X1 U5382 ( .B1(n6620), .B2(n4783), .A(n4782), .ZN(n4784) );
  AOI21_X1 U5383 ( .B1(n4891), .B2(n6619), .A(n4784), .ZN(n4787) );
  INV_X1 U5384 ( .A(n4855), .ZN(n7116) );
  NOR2_X1 U5385 ( .A1(n4738), .A2(n7116), .ZN(n6623) );
  OAI21_X1 U5386 ( .B1(n6623), .B2(n6627), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4786) );
  OAI21_X1 U5387 ( .B1(n4787), .B2(n6627), .A(n4786), .ZN(U3459) );
  NOR2_X1 U5388 ( .A1(n6614), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4788)
         );
  AOI21_X1 U5389 ( .B1(n3827), .B2(n4789), .A(n4788), .ZN(n7073) );
  INV_X1 U5390 ( .A(n7073), .ZN(n4791) );
  OAI22_X1 U5391 ( .A1(n5488), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7116), .ZN(n4790) );
  AOI21_X1 U5392 ( .B1(n4791), .B2(n6619), .A(n4790), .ZN(n4793) );
  AOI21_X1 U5393 ( .B1(n7071), .B2(n6619), .A(n6627), .ZN(n4792) );
  OAI22_X1 U5394 ( .A1(n4793), .A2(n6627), .B1(n4792), .B2(n3561), .ZN(U3461)
         );
  INV_X1 U5395 ( .A(n4717), .ZN(n4796) );
  OAI21_X1 U5396 ( .B1(n4796), .B2(n4794), .A(n4795), .ZN(n6943) );
  NAND2_X1 U5397 ( .A1(n4819), .A2(n4798), .ZN(n6955) );
  INV_X1 U5398 ( .A(n6955), .ZN(n4799) );
  AOI22_X1 U5399 ( .A1(n6160), .A2(n4799), .B1(n6159), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4800) );
  OAI21_X1 U5400 ( .B1(n6943), .B2(n6151), .A(n4800), .ZN(U2856) );
  NAND2_X1 U5401 ( .A1(n4801), .A2(n4802), .ZN(n4803) );
  XNOR2_X1 U5402 ( .A(n4804), .B(n4803), .ZN(n4852) );
  NAND3_X1 U5403 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6842), .ZN(n4968) );
  OAI21_X1 U5404 ( .B1(n6839), .B2(n4965), .A(n4968), .ZN(n6831) );
  INV_X1 U5405 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6949) );
  OAI22_X1 U5406 ( .A1(n6897), .A2(n6955), .B1(n6949), .B2(n6894), .ZN(n4813)
         );
  NOR2_X1 U5407 ( .A1(n4427), .A2(n6817), .ZN(n6838) );
  INV_X1 U5408 ( .A(n6838), .ZN(n4805) );
  NAND2_X1 U5409 ( .A1(n4806), .A2(n4805), .ZN(n4807) );
  NAND2_X1 U5410 ( .A1(n4808), .A2(n4807), .ZN(n6840) );
  INV_X1 U5411 ( .A(n6839), .ZN(n4809) );
  NOR2_X1 U5412 ( .A1(n4965), .A2(n4809), .ZN(n4810) );
  NOR2_X1 U5413 ( .A1(n6840), .A2(n4810), .ZN(n6826) );
  NOR2_X1 U5414 ( .A1(n6826), .A2(n4811), .ZN(n4812) );
  AOI211_X1 U5415 ( .C1(n6831), .C2(n4811), .A(n4813), .B(n4812), .ZN(n4814)
         );
  OAI21_X1 U5416 ( .B1(n4852), .B2(n6590), .A(n4814), .ZN(U3015) );
  AOI21_X1 U5417 ( .B1(n4816), .B2(n4795), .A(n4815), .ZN(n4817) );
  INV_X1 U5418 ( .A(n4817), .ZN(n6965) );
  AND2_X1 U5419 ( .A1(n4819), .A2(n4818), .ZN(n4820) );
  NOR2_X1 U5420 ( .A1(n5261), .A2(n4820), .ZN(n6960) );
  AOI22_X1 U5421 ( .A1(n6160), .A2(n6960), .B1(n6159), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4821) );
  OAI21_X1 U5422 ( .B1(n6965), .B2(n6151), .A(n4821), .ZN(U2855) );
  INV_X1 U5423 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4823) );
  AOI22_X1 U5424 ( .A1(n6666), .A2(UWORD_REG_14__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4822) );
  OAI21_X1 U5425 ( .B1(n4823), .B2(n4840), .A(n4822), .ZN(U2893) );
  INV_X1 U5426 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5427 ( .A1(n6666), .A2(UWORD_REG_0__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4824) );
  OAI21_X1 U5428 ( .B1(n4825), .B2(n4840), .A(n4824), .ZN(U2907) );
  INV_X1 U5429 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5430 ( .A1(n6666), .A2(UWORD_REG_1__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4826) );
  OAI21_X1 U5431 ( .B1(n4827), .B2(n4840), .A(n4826), .ZN(U2906) );
  INV_X1 U5432 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5433 ( .A1(n6666), .A2(UWORD_REG_2__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4828) );
  OAI21_X1 U5434 ( .B1(n4829), .B2(n4840), .A(n4828), .ZN(U2905) );
  INV_X1 U5435 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U5436 ( .A1(n6666), .A2(UWORD_REG_3__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4830) );
  OAI21_X1 U5437 ( .B1(n4831), .B2(n4840), .A(n4830), .ZN(U2904) );
  INV_X1 U5438 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5439 ( .A1(n6666), .A2(UWORD_REG_4__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4832) );
  OAI21_X1 U5440 ( .B1(n4833), .B2(n4840), .A(n4832), .ZN(U2903) );
  INV_X1 U5441 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5442 ( .A1(n6666), .A2(UWORD_REG_10__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4834) );
  OAI21_X1 U5443 ( .B1(n4835), .B2(n4840), .A(n4834), .ZN(U2897) );
  AOI22_X1 U5444 ( .A1(n6666), .A2(UWORD_REG_11__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4836) );
  OAI21_X1 U5445 ( .B1(n4308), .B2(n4840), .A(n4836), .ZN(U2896) );
  INV_X1 U5446 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5447 ( .A1(n6666), .A2(UWORD_REG_12__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4837) );
  OAI21_X1 U5448 ( .B1(n4838), .B2(n4840), .A(n4837), .ZN(U2895) );
  INV_X1 U5449 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5450 ( .A1(n6666), .A2(UWORD_REG_13__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4839) );
  OAI21_X1 U5451 ( .B1(n4841), .B2(n4840), .A(n4839), .ZN(U2894) );
  INV_X1 U5452 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6959) );
  NOR2_X1 U5453 ( .A1(n6894), .A2(n6959), .ZN(n6823) );
  NOR2_X1 U5454 ( .A1(n6753), .A2(n6962), .ZN(n4842) );
  AOI211_X1 U5455 ( .C1(n6477), .C2(n6963), .A(n6823), .B(n4842), .ZN(n4847)
         );
  INV_X1 U5456 ( .A(n4844), .ZN(n4845) );
  XNOR2_X1 U5457 ( .A(n4843), .B(n4845), .ZN(n6822) );
  NAND2_X1 U5458 ( .A1(n6822), .A2(n6774), .ZN(n4846) );
  OAI211_X1 U5459 ( .C1(n6965), .C2(n6748), .A(n4847), .B(n4846), .ZN(U2982)
         );
  INV_X1 U5460 ( .A(n6943), .ZN(n4850) );
  AOI22_X1 U5461 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6906), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4848) );
  OAI21_X1 U5462 ( .B1(n6941), .B2(n6778), .A(n4848), .ZN(n4849) );
  AOI21_X1 U5463 ( .B1(n4850), .B2(n6773), .A(n4849), .ZN(n4851) );
  OAI21_X1 U5464 ( .B1(n4852), .B2(n7062), .A(n4851), .ZN(U2983) );
  INV_X1 U5465 ( .A(n4854), .ZN(n6618) );
  NAND2_X1 U5466 ( .A1(n4857), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4976) );
  INV_X1 U5467 ( .A(n4976), .ZN(n5408) );
  NOR2_X1 U5468 ( .A1(n4920), .A2(n7084), .ZN(n5620) );
  AOI22_X1 U5469 ( .A1(n5417), .A2(n5329), .B1(n5408), .B2(n5620), .ZN(n5123)
         );
  INV_X1 U5470 ( .A(DATAI_2_), .ZN(n7154) );
  NAND3_X1 U5471 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5044) );
  NOR2_X1 U5472 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5044), .ZN(n5120)
         );
  INV_X1 U5473 ( .A(n5120), .ZN(n4859) );
  NOR2_X1 U5474 ( .A1(n5620), .A2(n4856), .ZN(n5626) );
  INV_X1 U5475 ( .A(n4857), .ZN(n4858) );
  NAND2_X1 U5476 ( .A1(n4858), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U5477 ( .A1(n4977), .A2(n4974), .ZN(n5411) );
  AOI211_X1 U5478 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4859), .A(n5626), .B(
        n5411), .ZN(n4868) );
  NOR2_X1 U5479 ( .A1(n5329), .A2(n5618), .ZN(n5144) );
  NOR2_X1 U5480 ( .A1(n4860), .A2(n5295), .ZN(n4862) );
  INV_X1 U5481 ( .A(n5117), .ZN(n4865) );
  NOR2_X1 U5482 ( .A1(n4860), .A2(n3443), .ZN(n4864) );
  NAND2_X1 U5483 ( .A1(n4864), .A2(n4861), .ZN(n4923) );
  OAI21_X1 U5484 ( .B1(n4865), .B2(n5361), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4866) );
  OAI21_X1 U5485 ( .B1(n5511), .B2(n5144), .A(n4866), .ZN(n4867) );
  NAND2_X1 U5486 ( .A1(n4868), .A2(n4867), .ZN(n5116) );
  NAND2_X1 U5487 ( .A1(n5116), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4874)
         );
  INV_X1 U5488 ( .A(DATAI_26_), .ZN(n6276) );
  OR2_X1 U5489 ( .A1(n6748), .A2(n6276), .ZN(n5683) );
  INV_X1 U5490 ( .A(DATAI_18_), .ZN(n4871) );
  OR2_X1 U5491 ( .A1(n6748), .A2(n4871), .ZN(n5551) );
  OAI22_X1 U5492 ( .A1(n5118), .A2(n5683), .B1(n5551), .B2(n5117), .ZN(n4872)
         );
  AOI21_X1 U5493 ( .B1(n5687), .B2(n5120), .A(n4872), .ZN(n4873) );
  OAI211_X1 U5494 ( .C1(n5123), .C2(n5689), .A(n4874), .B(n4873), .ZN(U3134)
         );
  INV_X1 U5495 ( .A(DATAI_3_), .ZN(n7157) );
  NAND2_X1 U5496 ( .A1(n5116), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4879)
         );
  INV_X1 U5497 ( .A(DATAI_27_), .ZN(n6277) );
  OR2_X1 U5498 ( .A1(n6748), .A2(n6277), .ZN(n5674) );
  INV_X1 U5499 ( .A(DATAI_19_), .ZN(n4876) );
  OR2_X1 U5500 ( .A1(n6748), .A2(n4876), .ZN(n5546) );
  OAI22_X1 U5501 ( .A1(n5118), .A2(n5674), .B1(n5546), .B2(n5117), .ZN(n4877)
         );
  AOI21_X1 U5502 ( .B1(n5676), .B2(n5120), .A(n4877), .ZN(n4878) );
  OAI211_X1 U5503 ( .C1(n5123), .C2(n5678), .A(n4879), .B(n4878), .ZN(U3135)
         );
  INV_X1 U5504 ( .A(DATAI_1_), .ZN(n7151) );
  NAND2_X1 U5505 ( .A1(n5116), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4884)
         );
  INV_X1 U5506 ( .A(DATAI_25_), .ZN(n6186) );
  OR2_X1 U5507 ( .A1(n6748), .A2(n6186), .ZN(n5660) );
  INV_X1 U5508 ( .A(DATAI_17_), .ZN(n4881) );
  OR2_X1 U5509 ( .A1(n6748), .A2(n4881), .ZN(n5522) );
  OAI22_X1 U5510 ( .A1(n5118), .A2(n5660), .B1(n5522), .B2(n5117), .ZN(n4882)
         );
  AOI21_X1 U5511 ( .B1(n5662), .B2(n5120), .A(n4882), .ZN(n4883) );
  OAI211_X1 U5512 ( .C1(n5123), .C2(n5664), .A(n4884), .B(n4883), .ZN(U3133)
         );
  INV_X1 U5513 ( .A(DATAI_7_), .ZN(n7169) );
  NAND2_X1 U5514 ( .A1(n5116), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4889)
         );
  INV_X1 U5515 ( .A(DATAI_31_), .ZN(n4885) );
  OR2_X1 U5516 ( .A1(n6748), .A2(n4885), .ZN(n5667) );
  INV_X1 U5517 ( .A(DATAI_23_), .ZN(n4886) );
  OR2_X1 U5518 ( .A1(n6748), .A2(n4886), .ZN(n5530) );
  OAI22_X1 U5519 ( .A1(n5118), .A2(n5667), .B1(n5530), .B2(n5117), .ZN(n4887)
         );
  AOI21_X1 U5520 ( .B1(n5669), .B2(n5120), .A(n4887), .ZN(n4888) );
  OAI211_X1 U5521 ( .C1(n5123), .C2(n5671), .A(n4889), .B(n4888), .ZN(U3139)
         );
  MUX2_X1 U5522 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4890), .S(n7077), 
        .Z(n7085) );
  OR2_X1 U5523 ( .A1(n7077), .A2(n3727), .ZN(n4893) );
  NAND2_X1 U5524 ( .A1(n7077), .A2(n4891), .ZN(n4892) );
  NAND2_X1 U5525 ( .A1(n4893), .A2(n4892), .ZN(n7082) );
  NAND3_X1 U5526 ( .A1(n7085), .A2(n5488), .A3(n7082), .ZN(n4897) );
  NOR2_X1 U5527 ( .A1(FLUSH_REG_SCAN_IN), .A2(n5488), .ZN(n4894) );
  NAND2_X1 U5528 ( .A1(n4895), .A2(n4894), .ZN(n4896) );
  NAND2_X1 U5529 ( .A1(n4897), .A2(n4896), .ZN(n7096) );
  INV_X1 U5530 ( .A(n6613), .ZN(n6622) );
  MUX2_X1 U5531 ( .A(n4906), .B(n4898), .S(n5488), .Z(n4899) );
  NAND2_X1 U5532 ( .A1(n4899), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4905) );
  INV_X1 U5533 ( .A(n4901), .ZN(n4902) );
  NOR2_X1 U5534 ( .A1(n4900), .A2(n4902), .ZN(n4903) );
  XNOR2_X1 U5535 ( .A(n4903), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7064)
         );
  NAND2_X1 U5536 ( .A1(n4905), .A2(n4904), .ZN(n7094) );
  AOI21_X1 U5537 ( .B1(n7096), .B2(n6622), .A(n7094), .ZN(n5181) );
  NAND2_X1 U5538 ( .A1(n5181), .A2(n4906), .ZN(n4908) );
  AOI21_X1 U5539 ( .B1(n4908), .B2(n4907), .A(n4977), .ZN(n6632) );
  INV_X1 U5540 ( .A(n6632), .ZN(n5927) );
  OAI21_X1 U5541 ( .B1(n5488), .B2(STATE2_REG_3__SCAN_IN), .A(n5927), .ZN(
        n5926) );
  NOR2_X1 U5542 ( .A1(n6632), .A2(n5618), .ZN(n5184) );
  INV_X1 U5543 ( .A(n5020), .ZN(n4913) );
  OR2_X1 U5544 ( .A1(n4923), .A2(n5617), .ZN(n5310) );
  OR2_X1 U5545 ( .A1(n4909), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4912) );
  INV_X1 U5546 ( .A(n4910), .ZN(n4922) );
  NAND2_X1 U5547 ( .A1(n3443), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5925) );
  NAND2_X1 U5548 ( .A1(n5296), .A2(n5187), .ZN(n5326) );
  NAND4_X1 U5549 ( .A1(n4913), .A2(n5310), .A3(n4912), .A4(n5326), .ZN(n4914)
         );
  AOI22_X1 U5550 ( .A1(n5184), .A2(n4914), .B1(n6632), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4915) );
  OAI21_X1 U5551 ( .B1(n5515), .B2(n5926), .A(n4915), .ZN(U3462) );
  NOR2_X1 U5552 ( .A1(n4815), .A2(n4917), .ZN(n4918) );
  OR2_X1 U5553 ( .A1(n4916), .A2(n4918), .ZN(n6980) );
  XOR2_X1 U5554 ( .A(n5261), .B(n5260), .Z(n6977) );
  AOI22_X1 U5555 ( .A1(n6160), .A2(n6977), .B1(n6159), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4919) );
  OAI21_X1 U5556 ( .B1(n6980), .B2(n6151), .A(n4919), .ZN(U2854) );
  NOR2_X1 U5557 ( .A1(n4771), .A2(n4854), .ZN(n5409) );
  INV_X1 U5558 ( .A(n4975), .ZN(n4921) );
  INV_X1 U5559 ( .A(n4920), .ZN(n5143) );
  NOR2_X1 U5560 ( .A1(n4921), .A2(n5143), .ZN(n5019) );
  AOI22_X1 U5561 ( .A1(n5417), .A2(n5409), .B1(n5408), .B2(n5019), .ZN(n5142)
         );
  NOR3_X1 U5562 ( .A1(n7083), .A2(n7084), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5309) );
  NAND2_X1 U5563 ( .A1(n7070), .A2(n5309), .ZN(n4929) );
  NOR2_X1 U5564 ( .A1(n5019), .A2(n5908), .ZN(n5022) );
  AOI211_X1 U5565 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4929), .A(n5022), .B(
        n5411), .ZN(n4928) );
  NOR2_X1 U5566 ( .A1(n5409), .A2(n5618), .ZN(n5416) );
  NAND2_X1 U5567 ( .A1(n4922), .A2(n3443), .ZN(n5199) );
  NOR2_X1 U5568 ( .A1(n4909), .A2(n5199), .ZN(n4947) );
  INV_X1 U5569 ( .A(n5136), .ZN(n4925) );
  INV_X1 U5570 ( .A(n4923), .ZN(n4924) );
  OAI21_X1 U5571 ( .B1(n4925), .B2(n5360), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4926) );
  OAI21_X1 U5572 ( .B1(n5511), .B2(n5416), .A(n4926), .ZN(n4927) );
  NAND2_X1 U5573 ( .A1(n4928), .A2(n4927), .ZN(n5135) );
  NAND2_X1 U5574 ( .A1(n5135), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4932)
         );
  INV_X1 U5575 ( .A(n4929), .ZN(n5139) );
  OAI22_X1 U5576 ( .A1(n5522), .A2(n5137), .B1(n5136), .B2(n5660), .ZN(n4930)
         );
  AOI21_X1 U5577 ( .B1(n5662), .B2(n5139), .A(n4930), .ZN(n4931) );
  OAI211_X1 U5578 ( .C1(n5142), .C2(n5664), .A(n4932), .B(n4931), .ZN(U3117)
         );
  NAND2_X1 U5579 ( .A1(n5135), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4935)
         );
  OAI22_X1 U5580 ( .A1(n5530), .A2(n5137), .B1(n5136), .B2(n5667), .ZN(n4933)
         );
  AOI21_X1 U5581 ( .B1(n5669), .B2(n5139), .A(n4933), .ZN(n4934) );
  OAI211_X1 U5582 ( .C1(n5142), .C2(n5671), .A(n4935), .B(n4934), .ZN(U3123)
         );
  NAND2_X1 U5583 ( .A1(n5135), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4938)
         );
  OAI22_X1 U5584 ( .A1(n5551), .A2(n5137), .B1(n5136), .B2(n5683), .ZN(n4936)
         );
  AOI21_X1 U5585 ( .B1(n5687), .B2(n5139), .A(n4936), .ZN(n4937) );
  OAI211_X1 U5586 ( .C1(n5142), .C2(n5689), .A(n4938), .B(n4937), .ZN(U3118)
         );
  NAND2_X1 U5587 ( .A1(n5135), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4941)
         );
  OAI22_X1 U5588 ( .A1(n5546), .A2(n5137), .B1(n5136), .B2(n5674), .ZN(n4939)
         );
  AOI21_X1 U5589 ( .B1(n5676), .B2(n5139), .A(n4939), .ZN(n4940) );
  OAI211_X1 U5590 ( .C1(n5142), .C2(n5678), .A(n4941), .B(n4940), .ZN(U3119)
         );
  AOI21_X1 U5591 ( .B1(n5020), .B2(n5187), .A(n5618), .ZN(n4945) );
  AND2_X1 U5592 ( .A1(n4854), .A2(n4771), .ZN(n5516) );
  NAND3_X1 U5593 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7083), .ZN(n5622) );
  NOR2_X1 U5594 ( .A1(n7070), .A2(n5622), .ZN(n5015) );
  AOI21_X1 U5595 ( .B1(n5624), .B2(n3827), .A(n5015), .ZN(n4944) );
  INV_X1 U5596 ( .A(n4944), .ZN(n4943) );
  INV_X1 U5597 ( .A(n5622), .ZN(n4942) );
  AOI22_X1 U5598 ( .A1(n4945), .A2(n4943), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4942), .ZN(n5018) );
  AOI22_X1 U5599 ( .A1(n4945), .A2(n4944), .B1(n5622), .B2(n5618), .ZN(n4946)
         );
  NAND2_X1 U5600 ( .A1(n5332), .A2(n4946), .ZN(n5011) );
  NAND2_X1 U5601 ( .A1(n5011), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4950)
         );
  OAI22_X1 U5602 ( .A1(n5546), .A2(n5136), .B1(n5623), .B2(n5674), .ZN(n4948)
         );
  AOI21_X1 U5603 ( .B1(n5676), .B2(n5015), .A(n4948), .ZN(n4949) );
  OAI211_X1 U5604 ( .C1(n5018), .C2(n5678), .A(n4950), .B(n4949), .ZN(U3111)
         );
  NAND2_X1 U5605 ( .A1(n5011), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4953)
         );
  OAI22_X1 U5606 ( .A1(n5530), .A2(n5136), .B1(n5623), .B2(n5667), .ZN(n4951)
         );
  AOI21_X1 U5607 ( .B1(n5669), .B2(n5015), .A(n4951), .ZN(n4952) );
  OAI211_X1 U5608 ( .C1(n5018), .C2(n5671), .A(n4953), .B(n4952), .ZN(U3115)
         );
  NAND2_X1 U5609 ( .A1(n5011), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4956)
         );
  OAI22_X1 U5610 ( .A1(n5551), .A2(n5136), .B1(n5623), .B2(n5683), .ZN(n4954)
         );
  AOI21_X1 U5611 ( .B1(n5687), .B2(n5015), .A(n4954), .ZN(n4955) );
  OAI211_X1 U5612 ( .C1(n5018), .C2(n5689), .A(n4956), .B(n4955), .ZN(U3110)
         );
  NAND2_X1 U5613 ( .A1(n5011), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4959)
         );
  OAI22_X1 U5614 ( .A1(n5522), .A2(n5136), .B1(n5623), .B2(n5660), .ZN(n4957)
         );
  AOI21_X1 U5615 ( .B1(n5662), .B2(n5015), .A(n4957), .ZN(n4958) );
  OAI211_X1 U5616 ( .C1(n5018), .C2(n5664), .A(n4959), .B(n4958), .ZN(U3109)
         );
  XOR2_X1 U5617 ( .A(n4960), .B(n4961), .Z(n6750) );
  INV_X1 U5618 ( .A(n6750), .ZN(n4973) );
  OAI21_X1 U5619 ( .B1(n6874), .B2(n6832), .A(n6826), .ZN(n6834) );
  INV_X1 U5620 ( .A(n4962), .ZN(n4964) );
  OAI21_X1 U5621 ( .B1(n4965), .B2(n4964), .A(n4963), .ZN(n4971) );
  INV_X1 U5622 ( .A(n6977), .ZN(n4967) );
  INV_X1 U5623 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4966) );
  OR2_X1 U5624 ( .A1(n6894), .A2(n4966), .ZN(n6751) );
  OAI21_X1 U5625 ( .B1(n6897), .B2(n4967), .A(n6751), .ZN(n4970) );
  NOR3_X1 U5626 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6828), .A3(n4968), 
        .ZN(n4969) );
  AOI211_X1 U5627 ( .C1(n6834), .C2(n4971), .A(n4970), .B(n4969), .ZN(n4972)
         );
  OAI21_X1 U5628 ( .B1(n4973), .B2(n6590), .A(n4972), .ZN(U3013) );
  INV_X1 U5629 ( .A(n4974), .ZN(n5621) );
  NOR2_X1 U5630 ( .A1(n4975), .A2(n5143), .ZN(n5407) );
  AOI22_X1 U5631 ( .A1(n5511), .A2(n5265), .B1(n5621), .B2(n5407), .ZN(n5134)
         );
  NOR2_X1 U5632 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5228) );
  NAND3_X1 U5633 ( .A1(n7075), .A2(n7070), .A3(n5228), .ZN(n4983) );
  NOR2_X1 U5634 ( .A1(n5407), .A2(n5908), .ZN(n5412) );
  NAND2_X1 U5635 ( .A1(n4977), .A2(n4976), .ZN(n5625) );
  AOI211_X1 U5636 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4983), .A(n5412), .B(
        n5625), .ZN(n4982) );
  NOR2_X1 U5637 ( .A1(n5265), .A2(n5618), .ZN(n5025) );
  NOR2_X1 U5638 ( .A1(n4861), .A2(n3443), .ZN(n4978) );
  INV_X1 U5639 ( .A(n5128), .ZN(n4979) );
  OAI21_X1 U5640 ( .B1(n5253), .B2(n4979), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4980) );
  OAI21_X1 U5641 ( .B1(n5417), .B2(n5025), .A(n4980), .ZN(n4981) );
  NAND2_X1 U5642 ( .A1(n4982), .A2(n4981), .ZN(n5127) );
  NAND2_X1 U5643 ( .A1(n5127), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4986) );
  INV_X1 U5644 ( .A(n4983), .ZN(n5131) );
  OAI22_X1 U5645 ( .A1(n5129), .A2(n5522), .B1(n5660), .B2(n5128), .ZN(n4984)
         );
  AOI21_X1 U5646 ( .B1(n5662), .B2(n5131), .A(n4984), .ZN(n4985) );
  OAI211_X1 U5647 ( .C1(n5134), .C2(n5664), .A(n4986), .B(n4985), .ZN(U3021)
         );
  NAND2_X1 U5648 ( .A1(n5127), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4989) );
  OAI22_X1 U5649 ( .A1(n5129), .A2(n5546), .B1(n5674), .B2(n5128), .ZN(n4987)
         );
  AOI21_X1 U5650 ( .B1(n5676), .B2(n5131), .A(n4987), .ZN(n4988) );
  OAI211_X1 U5651 ( .C1(n5134), .C2(n5678), .A(n4989), .B(n4988), .ZN(U3023)
         );
  NAND2_X1 U5652 ( .A1(n5127), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4992) );
  OAI22_X1 U5653 ( .A1(n5129), .A2(n5551), .B1(n5683), .B2(n5128), .ZN(n4990)
         );
  AOI21_X1 U5654 ( .B1(n5687), .B2(n5131), .A(n4990), .ZN(n4991) );
  OAI211_X1 U5655 ( .C1(n5134), .C2(n5689), .A(n4992), .B(n4991), .ZN(U3022)
         );
  NAND2_X1 U5656 ( .A1(n5127), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4995) );
  OAI22_X1 U5657 ( .A1(n5129), .A2(n5530), .B1(n5667), .B2(n5128), .ZN(n4993)
         );
  AOI21_X1 U5658 ( .B1(n5669), .B2(n5131), .A(n4993), .ZN(n4994) );
  OAI211_X1 U5659 ( .C1(n5134), .C2(n5671), .A(n4995), .B(n4994), .ZN(U3027)
         );
  INV_X1 U5660 ( .A(DATAI_6_), .ZN(n7166) );
  NAND2_X1 U5661 ( .A1(n5011), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5000)
         );
  INV_X1 U5662 ( .A(DATAI_22_), .ZN(n4996) );
  OR2_X1 U5663 ( .A1(n6748), .A2(n4996), .ZN(n5542) );
  INV_X1 U5664 ( .A(DATAI_30_), .ZN(n4997) );
  OR2_X1 U5665 ( .A1(n6748), .A2(n4997), .ZN(n5653) );
  OAI22_X1 U5666 ( .A1(n5542), .A2(n5136), .B1(n5623), .B2(n5653), .ZN(n4998)
         );
  AOI21_X1 U5667 ( .B1(n3433), .B2(n5015), .A(n4998), .ZN(n4999) );
  OAI211_X1 U5668 ( .C1(n5018), .C2(n5657), .A(n5000), .B(n4999), .ZN(U3114)
         );
  INV_X1 U5669 ( .A(DATAI_5_), .ZN(n7163) );
  NAND2_X1 U5670 ( .A1(n5011), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5005)
         );
  INV_X1 U5671 ( .A(DATAI_21_), .ZN(n5001) );
  OR2_X1 U5672 ( .A1(n6748), .A2(n5001), .ZN(n5538) );
  INV_X1 U5673 ( .A(DATAI_29_), .ZN(n5002) );
  OR2_X1 U5674 ( .A1(n6748), .A2(n5002), .ZN(n5632) );
  OAI22_X1 U5675 ( .A1(n5538), .A2(n5136), .B1(n5623), .B2(n5632), .ZN(n5003)
         );
  AOI21_X1 U5676 ( .B1(n3434), .B2(n5015), .A(n5003), .ZN(n5004) );
  OAI211_X1 U5677 ( .C1(n5018), .C2(n5636), .A(n5005), .B(n5004), .ZN(U3113)
         );
  INV_X1 U5678 ( .A(DATAI_4_), .ZN(n7160) );
  NAND2_X1 U5679 ( .A1(n5011), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5009)
         );
  INV_X1 U5680 ( .A(DATAI_20_), .ZN(n5006) );
  OR2_X1 U5681 ( .A1(n6748), .A2(n5006), .ZN(n5534) );
  INV_X1 U5682 ( .A(DATAI_28_), .ZN(n6188) );
  OR2_X1 U5683 ( .A1(n6748), .A2(n6188), .ZN(n5639) );
  OAI22_X1 U5684 ( .A1(n5534), .A2(n5136), .B1(n5623), .B2(n5639), .ZN(n5007)
         );
  AOI21_X1 U5685 ( .B1(n3435), .B2(n5015), .A(n5007), .ZN(n5008) );
  OAI211_X1 U5686 ( .C1(n5018), .C2(n5643), .A(n5009), .B(n5008), .ZN(U3112)
         );
  INV_X1 U5687 ( .A(DATAI_0_), .ZN(n7148) );
  NAND2_X1 U5688 ( .A1(n5011), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5017)
         );
  INV_X1 U5689 ( .A(DATAI_16_), .ZN(n5013) );
  OR2_X1 U5690 ( .A1(n6748), .A2(n5013), .ZN(n5526) );
  INV_X1 U5691 ( .A(DATAI_24_), .ZN(n6284) );
  OR2_X1 U5692 ( .A1(n6748), .A2(n6284), .ZN(n5646) );
  OAI22_X1 U5693 ( .A1(n5526), .A2(n5136), .B1(n5623), .B2(n5646), .ZN(n5014)
         );
  AOI21_X1 U5694 ( .B1(n5648), .B2(n5015), .A(n5014), .ZN(n5016) );
  OAI211_X1 U5695 ( .C1(n5018), .C2(n5650), .A(n5017), .B(n5016), .ZN(U3108)
         );
  AOI22_X1 U5696 ( .A1(n5417), .A2(n5265), .B1(n5621), .B2(n5019), .ZN(n5091)
         );
  NAND3_X1 U5697 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n7083), .A3(n7075), .ZN(n5269) );
  NOR2_X1 U5698 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5269), .ZN(n5087)
         );
  NAND2_X1 U5699 ( .A1(n5020), .A2(n5295), .ZN(n5273) );
  NOR2_X1 U5700 ( .A1(n5302), .A2(n5295), .ZN(n5145) );
  OAI22_X1 U5701 ( .A1(n5085), .A2(n5530), .B1(n5667), .B2(n5084), .ZN(n5021)
         );
  AOI21_X1 U5702 ( .B1(n5669), .B2(n5087), .A(n5021), .ZN(n5029) );
  INV_X1 U5703 ( .A(n5087), .ZN(n5023) );
  AOI211_X1 U5704 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5023), .A(n5022), .B(
        n5625), .ZN(n5027) );
  OAI21_X1 U5705 ( .B1(n5290), .B2(n5400), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5024) );
  OAI21_X1 U5706 ( .B1(n5511), .B2(n5025), .A(n5024), .ZN(n5026) );
  NAND2_X1 U5707 ( .A1(n5027), .A2(n5026), .ZN(n5088) );
  NAND2_X1 U5708 ( .A1(n5088), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5028) );
  OAI211_X1 U5709 ( .C1(n5091), .C2(n5671), .A(n5029), .B(n5028), .ZN(U3091)
         );
  OAI22_X1 U5710 ( .A1(n5085), .A2(n5546), .B1(n5674), .B2(n5084), .ZN(n5030)
         );
  AOI21_X1 U5711 ( .B1(n5676), .B2(n5087), .A(n5030), .ZN(n5032) );
  NAND2_X1 U5712 ( .A1(n5088), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5031) );
  OAI211_X1 U5713 ( .C1(n5091), .C2(n5678), .A(n5032), .B(n5031), .ZN(U3087)
         );
  OAI22_X1 U5714 ( .A1(n5085), .A2(n5522), .B1(n5660), .B2(n5084), .ZN(n5033)
         );
  AOI21_X1 U5715 ( .B1(n5662), .B2(n5087), .A(n5033), .ZN(n5035) );
  NAND2_X1 U5716 ( .A1(n5088), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5034) );
  OAI211_X1 U5717 ( .C1(n5091), .C2(n5664), .A(n5035), .B(n5034), .ZN(U3085)
         );
  OAI22_X1 U5718 ( .A1(n5085), .A2(n5551), .B1(n5683), .B2(n5084), .ZN(n5036)
         );
  AOI21_X1 U5719 ( .B1(n5687), .B2(n5087), .A(n5036), .ZN(n5038) );
  NAND2_X1 U5720 ( .A1(n5088), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5037) );
  OAI211_X1 U5721 ( .C1(n5091), .C2(n5689), .A(n5038), .B(n5037), .ZN(U3086)
         );
  INV_X1 U5722 ( .A(n3827), .ZN(n5496) );
  NOR2_X1 U5723 ( .A1(n5515), .A2(n5496), .ZN(n5307) );
  NOR2_X1 U5724 ( .A1(n5039), .A2(n7084), .ZN(n5071) );
  AOI21_X1 U5725 ( .B1(n5307), .B2(n5329), .A(n5071), .ZN(n5046) );
  INV_X1 U5726 ( .A(n5046), .ZN(n5041) );
  INV_X1 U5727 ( .A(n5044), .ZN(n5040) );
  AOI22_X1 U5728 ( .A1(n5041), .A2(n5327), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5040), .ZN(n5074) );
  NOR2_X1 U5729 ( .A1(n5618), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5513) );
  INV_X1 U5730 ( .A(n5513), .ZN(n5042) );
  OAI21_X1 U5731 ( .B1(n5043), .B2(n6748), .A(n5042), .ZN(n5045) );
  AOI22_X1 U5732 ( .A1(n5046), .A2(n5045), .B1(n5618), .B2(n5044), .ZN(n5047)
         );
  NAND2_X1 U5733 ( .A1(n5332), .A2(n5047), .ZN(n5069) );
  NAND2_X1 U5734 ( .A1(n5069), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5050)
         );
  OAI22_X1 U5735 ( .A1(n5534), .A2(n5128), .B1(n5117), .B2(n5639), .ZN(n5048)
         );
  AOI21_X1 U5736 ( .B1(n3435), .B2(n5071), .A(n5048), .ZN(n5049) );
  OAI211_X1 U5737 ( .C1(n5074), .C2(n5643), .A(n5050), .B(n5049), .ZN(U3144)
         );
  NAND2_X1 U5738 ( .A1(n5069), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5053)
         );
  OAI22_X1 U5739 ( .A1(n5526), .A2(n5128), .B1(n5117), .B2(n5646), .ZN(n5051)
         );
  AOI21_X1 U5740 ( .B1(n5648), .B2(n5071), .A(n5051), .ZN(n5052) );
  OAI211_X1 U5741 ( .C1(n5074), .C2(n5650), .A(n5053), .B(n5052), .ZN(U3140)
         );
  NAND2_X1 U5742 ( .A1(n5069), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5056)
         );
  OAI22_X1 U5743 ( .A1(n5542), .A2(n5128), .B1(n5117), .B2(n5653), .ZN(n5054)
         );
  AOI21_X1 U5744 ( .B1(n3433), .B2(n5071), .A(n5054), .ZN(n5055) );
  OAI211_X1 U5745 ( .C1(n5074), .C2(n5657), .A(n5056), .B(n5055), .ZN(U3146)
         );
  NAND2_X1 U5746 ( .A1(n5069), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5059)
         );
  OAI22_X1 U5747 ( .A1(n5530), .A2(n5128), .B1(n5117), .B2(n5667), .ZN(n5057)
         );
  AOI21_X1 U5748 ( .B1(n5669), .B2(n5071), .A(n5057), .ZN(n5058) );
  OAI211_X1 U5749 ( .C1(n5074), .C2(n5671), .A(n5059), .B(n5058), .ZN(U3147)
         );
  NAND2_X1 U5750 ( .A1(n5069), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5062)
         );
  OAI22_X1 U5751 ( .A1(n5522), .A2(n5128), .B1(n5117), .B2(n5660), .ZN(n5060)
         );
  AOI21_X1 U5752 ( .B1(n5662), .B2(n5071), .A(n5060), .ZN(n5061) );
  OAI211_X1 U5753 ( .C1(n5074), .C2(n5664), .A(n5062), .B(n5061), .ZN(U3141)
         );
  NAND2_X1 U5754 ( .A1(n5069), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5065)
         );
  OAI22_X1 U5755 ( .A1(n5546), .A2(n5128), .B1(n5117), .B2(n5674), .ZN(n5063)
         );
  AOI21_X1 U5756 ( .B1(n5676), .B2(n5071), .A(n5063), .ZN(n5064) );
  OAI211_X1 U5757 ( .C1(n5074), .C2(n5678), .A(n5065), .B(n5064), .ZN(U3143)
         );
  NAND2_X1 U5758 ( .A1(n5069), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5068)
         );
  OAI22_X1 U5759 ( .A1(n5551), .A2(n5128), .B1(n5117), .B2(n5683), .ZN(n5066)
         );
  AOI21_X1 U5760 ( .B1(n5687), .B2(n5071), .A(n5066), .ZN(n5067) );
  OAI211_X1 U5761 ( .C1(n5074), .C2(n5689), .A(n5068), .B(n5067), .ZN(U3142)
         );
  NAND2_X1 U5762 ( .A1(n5069), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5073)
         );
  OAI22_X1 U5763 ( .A1(n5538), .A2(n5128), .B1(n5117), .B2(n5632), .ZN(n5070)
         );
  AOI21_X1 U5764 ( .B1(n3434), .B2(n5071), .A(n5070), .ZN(n5072) );
  OAI211_X1 U5765 ( .C1(n5074), .C2(n5636), .A(n5073), .B(n5072), .ZN(U3145)
         );
  OAI22_X1 U5766 ( .A1(n5085), .A2(n5542), .B1(n5653), .B2(n5084), .ZN(n5075)
         );
  AOI21_X1 U5767 ( .B1(n3433), .B2(n5087), .A(n5075), .ZN(n5077) );
  NAND2_X1 U5768 ( .A1(n5088), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5076) );
  OAI211_X1 U5769 ( .C1(n5091), .C2(n5657), .A(n5077), .B(n5076), .ZN(U3090)
         );
  OAI22_X1 U5770 ( .A1(n5085), .A2(n5538), .B1(n5632), .B2(n5084), .ZN(n5078)
         );
  AOI21_X1 U5771 ( .B1(n3434), .B2(n5087), .A(n5078), .ZN(n5080) );
  NAND2_X1 U5772 ( .A1(n5088), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5079) );
  OAI211_X1 U5773 ( .C1(n5091), .C2(n5636), .A(n5080), .B(n5079), .ZN(U3089)
         );
  OAI22_X1 U5774 ( .A1(n5085), .A2(n5534), .B1(n5639), .B2(n5084), .ZN(n5081)
         );
  AOI21_X1 U5775 ( .B1(n3435), .B2(n5087), .A(n5081), .ZN(n5083) );
  NAND2_X1 U5776 ( .A1(n5088), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5082) );
  OAI211_X1 U5777 ( .C1(n5091), .C2(n5643), .A(n5083), .B(n5082), .ZN(U3088)
         );
  OAI22_X1 U5778 ( .A1(n5085), .A2(n5526), .B1(n5646), .B2(n5084), .ZN(n5086)
         );
  AOI21_X1 U5779 ( .B1(n5648), .B2(n5087), .A(n5086), .ZN(n5090) );
  NAND2_X1 U5780 ( .A1(n5088), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5089) );
  OAI211_X1 U5781 ( .C1(n5091), .C2(n5650), .A(n5090), .B(n5089), .ZN(U3084)
         );
  NAND2_X1 U5782 ( .A1(n5135), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5094)
         );
  OAI22_X1 U5783 ( .A1(n5526), .A2(n5137), .B1(n5136), .B2(n5646), .ZN(n5092)
         );
  AOI21_X1 U5784 ( .B1(n5648), .B2(n5139), .A(n5092), .ZN(n5093) );
  OAI211_X1 U5785 ( .C1(n5142), .C2(n5650), .A(n5094), .B(n5093), .ZN(U3116)
         );
  NAND2_X1 U5786 ( .A1(n5116), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5097)
         );
  OAI22_X1 U5787 ( .A1(n5118), .A2(n5639), .B1(n5534), .B2(n5117), .ZN(n5095)
         );
  AOI21_X1 U5788 ( .B1(n3435), .B2(n5120), .A(n5095), .ZN(n5096) );
  OAI211_X1 U5789 ( .C1(n5123), .C2(n5643), .A(n5097), .B(n5096), .ZN(U3136)
         );
  NAND2_X1 U5790 ( .A1(n5135), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5100)
         );
  OAI22_X1 U5791 ( .A1(n5534), .A2(n5137), .B1(n5136), .B2(n5639), .ZN(n5098)
         );
  AOI21_X1 U5792 ( .B1(n3435), .B2(n5139), .A(n5098), .ZN(n5099) );
  OAI211_X1 U5793 ( .C1(n5142), .C2(n5643), .A(n5100), .B(n5099), .ZN(U3120)
         );
  NAND2_X1 U5794 ( .A1(n5127), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5103) );
  OAI22_X1 U5795 ( .A1(n5129), .A2(n5526), .B1(n5646), .B2(n5128), .ZN(n5101)
         );
  AOI21_X1 U5796 ( .B1(n5648), .B2(n5131), .A(n5101), .ZN(n5102) );
  OAI211_X1 U5797 ( .C1(n5134), .C2(n5650), .A(n5103), .B(n5102), .ZN(U3020)
         );
  NAND2_X1 U5798 ( .A1(n5127), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5106) );
  OAI22_X1 U5799 ( .A1(n5129), .A2(n5538), .B1(n5632), .B2(n5128), .ZN(n5104)
         );
  AOI21_X1 U5800 ( .B1(n3434), .B2(n5131), .A(n5104), .ZN(n5105) );
  OAI211_X1 U5801 ( .C1(n5134), .C2(n5636), .A(n5106), .B(n5105), .ZN(U3025)
         );
  NAND2_X1 U5802 ( .A1(n5116), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5109)
         );
  OAI22_X1 U5803 ( .A1(n5118), .A2(n5632), .B1(n5538), .B2(n5117), .ZN(n5107)
         );
  AOI21_X1 U5804 ( .B1(n3434), .B2(n5120), .A(n5107), .ZN(n5108) );
  OAI211_X1 U5805 ( .C1(n5123), .C2(n5636), .A(n5109), .B(n5108), .ZN(U3137)
         );
  NAND2_X1 U5806 ( .A1(n5116), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5112)
         );
  OAI22_X1 U5807 ( .A1(n5118), .A2(n5646), .B1(n5526), .B2(n5117), .ZN(n5110)
         );
  AOI21_X1 U5808 ( .B1(n5648), .B2(n5120), .A(n5110), .ZN(n5111) );
  OAI211_X1 U5809 ( .C1(n5123), .C2(n5650), .A(n5112), .B(n5111), .ZN(U3132)
         );
  NAND2_X1 U5810 ( .A1(n5135), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5115)
         );
  OAI22_X1 U5811 ( .A1(n5542), .A2(n5137), .B1(n5136), .B2(n5653), .ZN(n5113)
         );
  AOI21_X1 U5812 ( .B1(n3433), .B2(n5139), .A(n5113), .ZN(n5114) );
  OAI211_X1 U5813 ( .C1(n5142), .C2(n5657), .A(n5115), .B(n5114), .ZN(U3122)
         );
  NAND2_X1 U5814 ( .A1(n5116), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5122)
         );
  OAI22_X1 U5815 ( .A1(n5118), .A2(n5653), .B1(n5542), .B2(n5117), .ZN(n5119)
         );
  AOI21_X1 U5816 ( .B1(n3433), .B2(n5120), .A(n5119), .ZN(n5121) );
  OAI211_X1 U5817 ( .C1(n5123), .C2(n5657), .A(n5122), .B(n5121), .ZN(U3138)
         );
  NAND2_X1 U5818 ( .A1(n5127), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5126) );
  OAI22_X1 U5819 ( .A1(n5129), .A2(n5542), .B1(n5653), .B2(n5128), .ZN(n5124)
         );
  AOI21_X1 U5820 ( .B1(n3433), .B2(n5131), .A(n5124), .ZN(n5125) );
  OAI211_X1 U5821 ( .C1(n5134), .C2(n5657), .A(n5126), .B(n5125), .ZN(U3026)
         );
  NAND2_X1 U5822 ( .A1(n5127), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5133) );
  OAI22_X1 U5823 ( .A1(n5129), .A2(n5534), .B1(n5639), .B2(n5128), .ZN(n5130)
         );
  AOI21_X1 U5824 ( .B1(n3435), .B2(n5131), .A(n5130), .ZN(n5132) );
  OAI211_X1 U5825 ( .C1(n5134), .C2(n5643), .A(n5133), .B(n5132), .ZN(U3024)
         );
  NAND2_X1 U5826 ( .A1(n5135), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5141)
         );
  OAI22_X1 U5827 ( .A1(n5538), .A2(n5137), .B1(n5136), .B2(n5632), .ZN(n5138)
         );
  AOI21_X1 U5828 ( .B1(n3434), .B2(n5139), .A(n5138), .ZN(n5140) );
  OAI211_X1 U5829 ( .C1(n5142), .C2(n5636), .A(n5141), .B(n5140), .ZN(U3121)
         );
  NAND2_X1 U5830 ( .A1(n5143), .A2(n7084), .ZN(n5150) );
  INV_X1 U5831 ( .A(n5150), .ZN(n5510) );
  AOI22_X1 U5832 ( .A1(n5511), .A2(n5329), .B1(n5510), .B2(n5408), .ZN(n5178)
         );
  NAND3_X1 U5833 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7084), .ZN(n5334) );
  NOR2_X1 U5834 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5334), .ZN(n5175)
         );
  INV_X1 U5835 ( .A(n5417), .ZN(n5148) );
  INV_X1 U5836 ( .A(n5144), .ZN(n5147) );
  NAND2_X1 U5837 ( .A1(n5145), .A2(n5272), .ZN(n5337) );
  NAND3_X1 U5838 ( .A1(n5296), .A2(n5295), .A3(n4863), .ZN(n5303) );
  AOI21_X1 U5839 ( .B1(n5337), .B2(n5303), .A(n5617), .ZN(n5146) );
  AOI21_X1 U5840 ( .B1(n5148), .B2(n5147), .A(n5146), .ZN(n5149) );
  NOR2_X1 U5841 ( .A1(n5149), .A2(n5411), .ZN(n5151) );
  NAND2_X1 U5842 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5150), .ZN(n5520) );
  NAND2_X1 U5843 ( .A1(n5173), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5154) );
  OAI22_X1 U5844 ( .A1(n5337), .A2(n5530), .B1(n5303), .B2(n5667), .ZN(n5152)
         );
  AOI21_X1 U5845 ( .B1(n5669), .B2(n5175), .A(n5152), .ZN(n5153) );
  OAI211_X1 U5846 ( .C1(n5178), .C2(n5671), .A(n5154), .B(n5153), .ZN(U3075)
         );
  NAND2_X1 U5847 ( .A1(n5173), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U5848 ( .A1(n5337), .A2(n5522), .B1(n5303), .B2(n5660), .ZN(n5155)
         );
  AOI21_X1 U5849 ( .B1(n5662), .B2(n5175), .A(n5155), .ZN(n5156) );
  OAI211_X1 U5850 ( .C1(n5178), .C2(n5664), .A(n5157), .B(n5156), .ZN(U3069)
         );
  NAND2_X1 U5851 ( .A1(n5173), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5160) );
  OAI22_X1 U5852 ( .A1(n5337), .A2(n5526), .B1(n5303), .B2(n5646), .ZN(n5158)
         );
  AOI21_X1 U5853 ( .B1(n5648), .B2(n5175), .A(n5158), .ZN(n5159) );
  OAI211_X1 U5854 ( .C1(n5178), .C2(n5650), .A(n5160), .B(n5159), .ZN(U3068)
         );
  NAND2_X1 U5855 ( .A1(n5173), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5163) );
  OAI22_X1 U5856 ( .A1(n5337), .A2(n5538), .B1(n5303), .B2(n5632), .ZN(n5161)
         );
  AOI21_X1 U5857 ( .B1(n3434), .B2(n5175), .A(n5161), .ZN(n5162) );
  OAI211_X1 U5858 ( .C1(n5178), .C2(n5636), .A(n5163), .B(n5162), .ZN(U3073)
         );
  NAND2_X1 U5859 ( .A1(n5173), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5166) );
  OAI22_X1 U5860 ( .A1(n5337), .A2(n5534), .B1(n5303), .B2(n5639), .ZN(n5164)
         );
  AOI21_X1 U5861 ( .B1(n3435), .B2(n5175), .A(n5164), .ZN(n5165) );
  OAI211_X1 U5862 ( .C1(n5178), .C2(n5643), .A(n5166), .B(n5165), .ZN(U3072)
         );
  NAND2_X1 U5863 ( .A1(n5173), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5169) );
  OAI22_X1 U5864 ( .A1(n5337), .A2(n5551), .B1(n5303), .B2(n5683), .ZN(n5167)
         );
  AOI21_X1 U5865 ( .B1(n5687), .B2(n5175), .A(n5167), .ZN(n5168) );
  OAI211_X1 U5866 ( .C1(n5178), .C2(n5689), .A(n5169), .B(n5168), .ZN(U3070)
         );
  NAND2_X1 U5867 ( .A1(n5173), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5172) );
  OAI22_X1 U5868 ( .A1(n5337), .A2(n5542), .B1(n5303), .B2(n5653), .ZN(n5170)
         );
  AOI21_X1 U5869 ( .B1(n3433), .B2(n5175), .A(n5170), .ZN(n5171) );
  OAI211_X1 U5870 ( .C1(n5178), .C2(n5657), .A(n5172), .B(n5171), .ZN(U3074)
         );
  NAND2_X1 U5871 ( .A1(n5173), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5177) );
  OAI22_X1 U5872 ( .A1(n5337), .A2(n5546), .B1(n5303), .B2(n5674), .ZN(n5174)
         );
  AOI21_X1 U5873 ( .B1(n5676), .B2(n5175), .A(n5174), .ZN(n5176) );
  OAI211_X1 U5874 ( .C1(n5178), .C2(n5678), .A(n5177), .B(n5176), .ZN(U3071)
         );
  INV_X1 U5875 ( .A(n5179), .ZN(n5180) );
  AND2_X1 U5876 ( .A1(n5181), .A2(n5180), .ZN(n7113) );
  MUX2_X1 U5877 ( .A(n7113), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(n6632), 
        .Z(n5182) );
  AOI21_X1 U5878 ( .B1(n5184), .B2(n4863), .A(n5182), .ZN(n5183) );
  OAI21_X1 U5879 ( .B1(n5496), .B2(n5926), .A(n5183), .ZN(U3465) );
  INV_X1 U5880 ( .A(n5184), .ZN(n5928) );
  AOI211_X1 U5881 ( .C1(n5295), .C2(n5617), .A(n5187), .B(n5928), .ZN(n5185)
         );
  AOI21_X1 U5882 ( .B1(n6632), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5185), 
        .ZN(n5186) );
  OAI21_X1 U5883 ( .B1(n6618), .B2(n5926), .A(n5186), .ZN(U3464) );
  INV_X1 U5884 ( .A(n4861), .ZN(n5188) );
  NAND3_X1 U5885 ( .A1(n4909), .A2(n5188), .A3(n5187), .ZN(n5189) );
  NAND2_X1 U5886 ( .A1(n5189), .A2(n5327), .ZN(n5195) );
  INV_X1 U5887 ( .A(n5195), .ZN(n5193) );
  OR2_X1 U5888 ( .A1(n4732), .A2(n5496), .ZN(n5229) );
  INV_X1 U5889 ( .A(n5516), .ZN(n5191) );
  NAND2_X1 U5890 ( .A1(n5190), .A2(n5228), .ZN(n5197) );
  OAI21_X1 U5891 ( .B1(n5229), .B2(n5191), .A(n5197), .ZN(n5196) );
  NAND2_X1 U5892 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5228), .ZN(n5518) );
  INV_X1 U5893 ( .A(n5518), .ZN(n5192) );
  AOI22_X1 U5894 ( .A1(n5193), .A2(n5196), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5192), .ZN(n5227) );
  NAND2_X1 U5895 ( .A1(n5618), .A2(n5518), .ZN(n5194) );
  OAI211_X1 U5896 ( .C1(n5196), .C2(n5195), .A(n5332), .B(n5194), .ZN(n5222)
         );
  NAND2_X1 U5897 ( .A1(n5222), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5203) );
  INV_X1 U5898 ( .A(n5197), .ZN(n5224) );
  INV_X1 U5899 ( .A(n5199), .ZN(n5198) );
  NAND3_X1 U5900 ( .A1(n5198), .A2(n4863), .A3(n4909), .ZN(n5443) );
  NOR2_X1 U5901 ( .A1(n5199), .A2(n4863), .ZN(n5200) );
  OAI22_X1 U5902 ( .A1(n5542), .A2(n5443), .B1(n5550), .B2(n5653), .ZN(n5201)
         );
  AOI21_X1 U5903 ( .B1(n3433), .B2(n5224), .A(n5201), .ZN(n5202) );
  OAI211_X1 U5904 ( .C1(n5227), .C2(n5657), .A(n5203), .B(n5202), .ZN(U3050)
         );
  NAND2_X1 U5905 ( .A1(n5222), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5206) );
  OAI22_X1 U5906 ( .A1(n5538), .A2(n5443), .B1(n5550), .B2(n5632), .ZN(n5204)
         );
  AOI21_X1 U5907 ( .B1(n3434), .B2(n5224), .A(n5204), .ZN(n5205) );
  OAI211_X1 U5908 ( .C1(n5227), .C2(n5636), .A(n5206), .B(n5205), .ZN(U3049)
         );
  NAND2_X1 U5909 ( .A1(n5222), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5209) );
  OAI22_X1 U5910 ( .A1(n5522), .A2(n5443), .B1(n5550), .B2(n5660), .ZN(n5207)
         );
  AOI21_X1 U5911 ( .B1(n5662), .B2(n5224), .A(n5207), .ZN(n5208) );
  OAI211_X1 U5912 ( .C1(n5227), .C2(n5664), .A(n5209), .B(n5208), .ZN(U3045)
         );
  NAND2_X1 U5913 ( .A1(n5222), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5212) );
  OAI22_X1 U5914 ( .A1(n5551), .A2(n5443), .B1(n5550), .B2(n5683), .ZN(n5210)
         );
  AOI21_X1 U5915 ( .B1(n5687), .B2(n5224), .A(n5210), .ZN(n5211) );
  OAI211_X1 U5916 ( .C1(n5227), .C2(n5689), .A(n5212), .B(n5211), .ZN(U3046)
         );
  NAND2_X1 U5917 ( .A1(n5222), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5215) );
  OAI22_X1 U5918 ( .A1(n5530), .A2(n5443), .B1(n5550), .B2(n5667), .ZN(n5213)
         );
  AOI21_X1 U5919 ( .B1(n5669), .B2(n5224), .A(n5213), .ZN(n5214) );
  OAI211_X1 U5920 ( .C1(n5227), .C2(n5671), .A(n5215), .B(n5214), .ZN(U3051)
         );
  NAND2_X1 U5921 ( .A1(n5222), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5218) );
  OAI22_X1 U5922 ( .A1(n5546), .A2(n5443), .B1(n5550), .B2(n5674), .ZN(n5216)
         );
  AOI21_X1 U5923 ( .B1(n5676), .B2(n5224), .A(n5216), .ZN(n5217) );
  OAI211_X1 U5924 ( .C1(n5227), .C2(n5678), .A(n5218), .B(n5217), .ZN(U3047)
         );
  NAND2_X1 U5925 ( .A1(n5222), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5221) );
  OAI22_X1 U5926 ( .A1(n5534), .A2(n5443), .B1(n5550), .B2(n5639), .ZN(n5219)
         );
  AOI21_X1 U5927 ( .B1(n3435), .B2(n5224), .A(n5219), .ZN(n5220) );
  OAI211_X1 U5928 ( .C1(n5227), .C2(n5643), .A(n5221), .B(n5220), .ZN(U3048)
         );
  NAND2_X1 U5929 ( .A1(n5222), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5226) );
  OAI22_X1 U5930 ( .A1(n5526), .A2(n5443), .B1(n5550), .B2(n5646), .ZN(n5223)
         );
  AOI21_X1 U5931 ( .B1(n5648), .B2(n5224), .A(n5223), .ZN(n5225) );
  OAI211_X1 U5932 ( .C1(n5227), .C2(n5650), .A(n5226), .B(n5225), .ZN(U3044)
         );
  NAND2_X1 U5933 ( .A1(n5228), .A2(n7075), .ZN(n5233) );
  NOR2_X1 U5934 ( .A1(n7070), .A2(n5233), .ZN(n5230) );
  INV_X1 U5935 ( .A(n5230), .ZN(n5256) );
  INV_X1 U5936 ( .A(n5229), .ZN(n5330) );
  AOI21_X1 U5937 ( .B1(n5330), .B2(n5265), .A(n5230), .ZN(n5235) );
  AOI21_X1 U5938 ( .B1(n5236), .B2(STATEBS16_REG_SCAN_IN), .A(n5618), .ZN(
        n5232) );
  AOI22_X1 U5939 ( .A1(n5235), .A2(n5232), .B1(n5618), .B2(n5233), .ZN(n5231)
         );
  NAND2_X1 U5940 ( .A1(n5332), .A2(n5231), .ZN(n5252) );
  INV_X1 U5941 ( .A(n5232), .ZN(n5234) );
  OAI22_X1 U5942 ( .A1(n5235), .A2(n5234), .B1(n5908), .B2(n5233), .ZN(n5251)
         );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5252), .B1(n5375), 
        .B2(n5251), .ZN(n5238) );
  INV_X1 U5944 ( .A(n5546), .ZN(n5672) );
  INV_X1 U5945 ( .A(n5674), .ZN(n5376) );
  AOI22_X1 U5946 ( .A1(n5672), .A2(n5512), .B1(n5253), .B2(n5376), .ZN(n5237)
         );
  OAI211_X1 U5947 ( .C1(n5379), .C2(n5256), .A(n5238), .B(n5237), .ZN(U3031)
         );
  AOI22_X1 U5948 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5252), .B1(n5398), 
        .B2(n5251), .ZN(n5240) );
  INV_X1 U5949 ( .A(n5526), .ZN(n5644) );
  INV_X1 U5950 ( .A(n5646), .ZN(n5401) );
  AOI22_X1 U5951 ( .A1(n5644), .A2(n5512), .B1(n5253), .B2(n5401), .ZN(n5239)
         );
  OAI211_X1 U5952 ( .C1(n5405), .C2(n5256), .A(n5240), .B(n5239), .ZN(U3028)
         );
  INV_X1 U5953 ( .A(n5687), .ZN(n5388) );
  AOI22_X1 U5954 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5252), .B1(n5384), 
        .B2(n5251), .ZN(n5242) );
  INV_X1 U5955 ( .A(n5551), .ZN(n5680) );
  INV_X1 U5956 ( .A(n5683), .ZN(n5385) );
  AOI22_X1 U5957 ( .A1(n5680), .A2(n5512), .B1(n5253), .B2(n5385), .ZN(n5241)
         );
  OAI211_X1 U5958 ( .C1(n5388), .C2(n5256), .A(n5242), .B(n5241), .ZN(U3030)
         );
  AOI22_X1 U5959 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5252), .B1(n5357), 
        .B2(n5251), .ZN(n5244) );
  INV_X1 U5960 ( .A(n5530), .ZN(n5665) );
  INV_X1 U5961 ( .A(n5667), .ZN(n5359) );
  AOI22_X1 U5962 ( .A1(n5665), .A2(n5512), .B1(n5253), .B2(n5359), .ZN(n5243)
         );
  OAI211_X1 U5963 ( .C1(n5365), .C2(n5256), .A(n5244), .B(n5243), .ZN(U3035)
         );
  AOI22_X1 U5964 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5252), .B1(n5380), 
        .B2(n5251), .ZN(n5246) );
  INV_X1 U5965 ( .A(n5542), .ZN(n5651) );
  INV_X1 U5966 ( .A(n5653), .ZN(n5381) );
  AOI22_X1 U5967 ( .A1(n5651), .A2(n5512), .B1(n5253), .B2(n5381), .ZN(n5245)
         );
  OAI211_X1 U5968 ( .C1(n5655), .C2(n5256), .A(n5246), .B(n5245), .ZN(U3034)
         );
  AOI22_X1 U5969 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5252), .B1(n5371), 
        .B2(n5251), .ZN(n5248) );
  INV_X1 U5970 ( .A(n5538), .ZN(n5630) );
  INV_X1 U5971 ( .A(n5632), .ZN(n5372) );
  AOI22_X1 U5972 ( .A1(n5630), .A2(n5512), .B1(n5253), .B2(n5372), .ZN(n5247)
         );
  OAI211_X1 U5973 ( .C1(n5634), .C2(n5256), .A(n5248), .B(n5247), .ZN(U3033)
         );
  AOI22_X1 U5974 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5252), .B1(n5390), 
        .B2(n5251), .ZN(n5250) );
  INV_X1 U5975 ( .A(n5534), .ZN(n5637) );
  INV_X1 U5976 ( .A(n5639), .ZN(n5393) );
  AOI22_X1 U5977 ( .A1(n5637), .A2(n5512), .B1(n5253), .B2(n5393), .ZN(n5249)
         );
  OAI211_X1 U5978 ( .C1(n5641), .C2(n5256), .A(n5250), .B(n5249), .ZN(U3032)
         );
  INV_X1 U5979 ( .A(n5662), .ZN(n5370) );
  AOI22_X1 U5980 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5252), .B1(n5366), 
        .B2(n5251), .ZN(n5255) );
  INV_X1 U5981 ( .A(n5522), .ZN(n5658) );
  INV_X1 U5982 ( .A(n5660), .ZN(n5367) );
  AOI22_X1 U5983 ( .A1(n5658), .A2(n5512), .B1(n5253), .B2(n5367), .ZN(n5254)
         );
  OAI211_X1 U5984 ( .C1(n5370), .C2(n5256), .A(n5255), .B(n5254), .ZN(U3029)
         );
  OAI21_X1 U5985 ( .B1(n4916), .B2(n5258), .A(n5257), .ZN(n6988) );
  AOI21_X1 U5986 ( .B1(n5261), .B2(n5260), .A(n5259), .ZN(n5262) );
  OR2_X1 U5987 ( .A1(n3451), .A2(n5262), .ZN(n6833) );
  OAI222_X1 U5988 ( .A1(n6988), .A2(n6151), .B1(n6150), .B2(n5263), .C1(n6148), 
        .C2(n6833), .ZN(U2853) );
  NOR2_X1 U5989 ( .A1(n7070), .A2(n5269), .ZN(n5264) );
  INV_X1 U5990 ( .A(n5264), .ZN(n5293) );
  AOI21_X1 U5991 ( .B1(n5307), .B2(n5265), .A(n5264), .ZN(n5271) );
  OR2_X1 U5992 ( .A1(n5273), .A2(n5617), .ZN(n5266) );
  AND2_X1 U5993 ( .A1(n5266), .A2(n5327), .ZN(n5268) );
  AOI22_X1 U5994 ( .A1(n5271), .A2(n5268), .B1(n5618), .B2(n5269), .ZN(n5267)
         );
  NAND2_X1 U5995 ( .A1(n5332), .A2(n5267), .ZN(n5289) );
  INV_X1 U5996 ( .A(n5268), .ZN(n5270) );
  OAI22_X1 U5997 ( .A1(n5271), .A2(n5270), .B1(n5908), .B2(n5269), .ZN(n5288)
         );
  AOI22_X1 U5998 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5289), .B1(n5398), 
        .B2(n5288), .ZN(n5275) );
  AOI22_X1 U5999 ( .A1(n5616), .A2(n5644), .B1(n5290), .B2(n5401), .ZN(n5274)
         );
  OAI211_X1 U6000 ( .C1(n5293), .C2(n5405), .A(n5275), .B(n5274), .ZN(U3092)
         );
  AOI22_X1 U6001 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5289), .B1(n5384), 
        .B2(n5288), .ZN(n5277) );
  AOI22_X1 U6002 ( .A1(n5616), .A2(n5680), .B1(n5290), .B2(n5385), .ZN(n5276)
         );
  OAI211_X1 U6003 ( .C1(n5293), .C2(n5388), .A(n5277), .B(n5276), .ZN(U3094)
         );
  AOI22_X1 U6004 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5289), .B1(n5366), 
        .B2(n5288), .ZN(n5279) );
  AOI22_X1 U6005 ( .A1(n5616), .A2(n5658), .B1(n5290), .B2(n5367), .ZN(n5278)
         );
  OAI211_X1 U6006 ( .C1(n5293), .C2(n5370), .A(n5279), .B(n5278), .ZN(U3093)
         );
  AOI22_X1 U6007 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5289), .B1(n5390), 
        .B2(n5288), .ZN(n5281) );
  AOI22_X1 U6008 ( .A1(n5616), .A2(n5637), .B1(n5290), .B2(n5393), .ZN(n5280)
         );
  OAI211_X1 U6009 ( .C1(n5293), .C2(n5641), .A(n5281), .B(n5280), .ZN(U3096)
         );
  AOI22_X1 U6010 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5289), .B1(n5375), 
        .B2(n5288), .ZN(n5283) );
  AOI22_X1 U6011 ( .A1(n5616), .A2(n5672), .B1(n5290), .B2(n5376), .ZN(n5282)
         );
  OAI211_X1 U6012 ( .C1(n5293), .C2(n5379), .A(n5283), .B(n5282), .ZN(U3095)
         );
  AOI22_X1 U6013 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5289), .B1(n5380), 
        .B2(n5288), .ZN(n5285) );
  AOI22_X1 U6014 ( .A1(n5616), .A2(n5651), .B1(n5290), .B2(n5381), .ZN(n5284)
         );
  OAI211_X1 U6015 ( .C1(n5293), .C2(n5655), .A(n5285), .B(n5284), .ZN(U3098)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5289), .B1(n5357), 
        .B2(n5288), .ZN(n5287) );
  AOI22_X1 U6017 ( .A1(n5616), .A2(n5665), .B1(n5290), .B2(n5359), .ZN(n5286)
         );
  OAI211_X1 U6018 ( .C1(n5293), .C2(n5365), .A(n5287), .B(n5286), .ZN(U3099)
         );
  AOI22_X1 U6019 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5289), .B1(n5371), 
        .B2(n5288), .ZN(n5292) );
  AOI22_X1 U6020 ( .A1(n5616), .A2(n5630), .B1(n5290), .B2(n5372), .ZN(n5291)
         );
  OAI211_X1 U6021 ( .C1(n5293), .C2(n5634), .A(n5292), .B(n5291), .ZN(U3097)
         );
  NAND3_X1 U6022 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7084), .A3(n7075), .ZN(n5410) );
  NOR2_X1 U6023 ( .A1(n7070), .A2(n5410), .ZN(n5294) );
  INV_X1 U6024 ( .A(n5294), .ZN(n5396) );
  AOI21_X1 U6025 ( .B1(n5330), .B2(n5409), .A(n5294), .ZN(n5301) );
  INV_X1 U6026 ( .A(n5301), .ZN(n5299) );
  NAND3_X1 U6027 ( .A1(n5296), .A2(STATEBS16_REG_SCAN_IN), .A3(n5295), .ZN(
        n5297) );
  NAND2_X1 U6028 ( .A1(n5297), .A2(n5327), .ZN(n5300) );
  NAND2_X1 U6029 ( .A1(n5618), .A2(n5410), .ZN(n5298) );
  OAI211_X1 U6030 ( .C1(n5299), .C2(n5300), .A(n5332), .B(n5298), .ZN(n5391)
         );
  OAI22_X1 U6031 ( .A1(n5301), .A2(n5300), .B1(n5908), .B2(n5410), .ZN(n5389)
         );
  AOI22_X1 U6032 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5391), .B1(n5398), 
        .B2(n5389), .ZN(n5305) );
  NOR3_X2 U6033 ( .A1(n5302), .A2(n3443), .A3(n4863), .ZN(n5420) );
  AOI22_X1 U6034 ( .A1(n5401), .A2(n5420), .B1(n5392), .B2(n5644), .ZN(n5304)
         );
  OAI211_X1 U6035 ( .C1(n5405), .C2(n5396), .A(n5305), .B(n5304), .ZN(U3060)
         );
  INV_X1 U6036 ( .A(n5309), .ZN(n5311) );
  NOR2_X1 U6037 ( .A1(n7070), .A2(n5311), .ZN(n5306) );
  INV_X1 U6038 ( .A(n5306), .ZN(n5364) );
  AOI21_X1 U6039 ( .B1(n5307), .B2(n5409), .A(n5306), .ZN(n5313) );
  NAND3_X1 U6040 ( .A1(n5327), .A2(n5313), .A3(n5310), .ZN(n5308) );
  OAI211_X1 U6041 ( .C1(n5327), .C2(n5309), .A(n5332), .B(n5308), .ZN(n5358)
         );
  NAND2_X1 U6042 ( .A1(n5327), .A2(n5310), .ZN(n5312) );
  OAI22_X1 U6043 ( .A1(n5313), .A2(n5312), .B1(n4856), .B2(n5311), .ZN(n5356)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5358), .B1(n5398), 
        .B2(n5356), .ZN(n5315) );
  AOI22_X1 U6045 ( .A1(n5644), .A2(n5361), .B1(n5360), .B2(n5401), .ZN(n5314)
         );
  OAI211_X1 U6046 ( .C1(n5405), .C2(n5364), .A(n5315), .B(n5314), .ZN(U3124)
         );
  AOI22_X1 U6047 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5391), .B1(n5366), 
        .B2(n5389), .ZN(n5317) );
  AOI22_X1 U6048 ( .A1(n5367), .A2(n5420), .B1(n5392), .B2(n5658), .ZN(n5316)
         );
  OAI211_X1 U6049 ( .C1(n5370), .C2(n5396), .A(n5317), .B(n5316), .ZN(U3061)
         );
  AOI22_X1 U6050 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5358), .B1(n5384), 
        .B2(n5356), .ZN(n5319) );
  AOI22_X1 U6051 ( .A1(n5680), .A2(n5361), .B1(n5360), .B2(n5385), .ZN(n5318)
         );
  OAI211_X1 U6052 ( .C1(n5388), .C2(n5364), .A(n5319), .B(n5318), .ZN(U3126)
         );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5358), .B1(n5366), 
        .B2(n5356), .ZN(n5321) );
  AOI22_X1 U6054 ( .A1(n5658), .A2(n5361), .B1(n5360), .B2(n5367), .ZN(n5320)
         );
  OAI211_X1 U6055 ( .C1(n5370), .C2(n5364), .A(n5321), .B(n5320), .ZN(U3125)
         );
  AOI22_X1 U6056 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5358), .B1(n5390), 
        .B2(n5356), .ZN(n5323) );
  AOI22_X1 U6057 ( .A1(n5637), .A2(n5361), .B1(n5360), .B2(n5393), .ZN(n5322)
         );
  OAI211_X1 U6058 ( .C1(n5641), .C2(n5364), .A(n5323), .B(n5322), .ZN(U3128)
         );
  AOI22_X1 U6059 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5391), .B1(n5357), 
        .B2(n5389), .ZN(n5325) );
  AOI22_X1 U6060 ( .A1(n5359), .A2(n5420), .B1(n5392), .B2(n5665), .ZN(n5324)
         );
  OAI211_X1 U6061 ( .C1(n5365), .C2(n5396), .A(n5325), .B(n5324), .ZN(U3067)
         );
  NAND2_X1 U6062 ( .A1(n5327), .A2(n5326), .ZN(n5335) );
  INV_X1 U6063 ( .A(n5406), .ZN(n5328) );
  AOI21_X1 U6064 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(n5336) );
  INV_X1 U6065 ( .A(n5336), .ZN(n5333) );
  NAND2_X1 U6066 ( .A1(n5618), .A2(n5334), .ZN(n5331) );
  OAI211_X1 U6067 ( .C1(n5335), .C2(n5333), .A(n5332), .B(n5331), .ZN(n5399)
         );
  OAI22_X1 U6068 ( .A1(n5336), .A2(n5335), .B1(n4856), .B2(n5334), .ZN(n5397)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5399), .B1(n5380), 
        .B2(n5397), .ZN(n5339) );
  AOI22_X1 U6070 ( .A1(n5402), .A2(n5381), .B1(n5400), .B2(n5651), .ZN(n5338)
         );
  OAI211_X1 U6071 ( .C1(n5406), .C2(n5655), .A(n5339), .B(n5338), .ZN(U3082)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5399), .B1(n5357), 
        .B2(n5397), .ZN(n5341) );
  AOI22_X1 U6073 ( .A1(n5402), .A2(n5359), .B1(n5400), .B2(n5665), .ZN(n5340)
         );
  OAI211_X1 U6074 ( .C1(n5406), .C2(n5365), .A(n5341), .B(n5340), .ZN(U3083)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5358), .B1(n5380), 
        .B2(n5356), .ZN(n5343) );
  AOI22_X1 U6076 ( .A1(n5651), .A2(n5361), .B1(n5360), .B2(n5381), .ZN(n5342)
         );
  OAI211_X1 U6077 ( .C1(n5655), .C2(n5364), .A(n5343), .B(n5342), .ZN(U3130)
         );
  AOI22_X1 U6078 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5358), .B1(n5375), 
        .B2(n5356), .ZN(n5345) );
  AOI22_X1 U6079 ( .A1(n5672), .A2(n5361), .B1(n5360), .B2(n5376), .ZN(n5344)
         );
  OAI211_X1 U6080 ( .C1(n5379), .C2(n5364), .A(n5345), .B(n5344), .ZN(U3127)
         );
  AOI22_X1 U6081 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5399), .B1(n5384), 
        .B2(n5397), .ZN(n5347) );
  AOI22_X1 U6082 ( .A1(n5402), .A2(n5385), .B1(n5400), .B2(n5680), .ZN(n5346)
         );
  OAI211_X1 U6083 ( .C1(n5406), .C2(n5388), .A(n5347), .B(n5346), .ZN(U3078)
         );
  AOI22_X1 U6084 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5399), .B1(n5375), 
        .B2(n5397), .ZN(n5349) );
  AOI22_X1 U6085 ( .A1(n5402), .A2(n5376), .B1(n5400), .B2(n5672), .ZN(n5348)
         );
  OAI211_X1 U6086 ( .C1(n5406), .C2(n5379), .A(n5349), .B(n5348), .ZN(U3079)
         );
  AOI22_X1 U6087 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5399), .B1(n5390), 
        .B2(n5397), .ZN(n5351) );
  AOI22_X1 U6088 ( .A1(n5402), .A2(n5393), .B1(n5400), .B2(n5637), .ZN(n5350)
         );
  OAI211_X1 U6089 ( .C1(n5406), .C2(n5641), .A(n5351), .B(n5350), .ZN(U3080)
         );
  AOI22_X1 U6090 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5358), .B1(n5371), 
        .B2(n5356), .ZN(n5353) );
  AOI22_X1 U6091 ( .A1(n5630), .A2(n5361), .B1(n5360), .B2(n5372), .ZN(n5352)
         );
  OAI211_X1 U6092 ( .C1(n5634), .C2(n5364), .A(n5353), .B(n5352), .ZN(U3129)
         );
  AOI22_X1 U6093 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5391), .B1(n5371), 
        .B2(n5389), .ZN(n5355) );
  AOI22_X1 U6094 ( .A1(n5372), .A2(n5420), .B1(n5392), .B2(n5630), .ZN(n5354)
         );
  OAI211_X1 U6095 ( .C1(n5634), .C2(n5396), .A(n5355), .B(n5354), .ZN(U3065)
         );
  AOI22_X1 U6096 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5358), .B1(n5357), 
        .B2(n5356), .ZN(n5363) );
  AOI22_X1 U6097 ( .A1(n5665), .A2(n5361), .B1(n5360), .B2(n5359), .ZN(n5362)
         );
  OAI211_X1 U6098 ( .C1(n5365), .C2(n5364), .A(n5363), .B(n5362), .ZN(U3131)
         );
  AOI22_X1 U6099 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5399), .B1(n5366), 
        .B2(n5397), .ZN(n5369) );
  AOI22_X1 U6100 ( .A1(n5402), .A2(n5367), .B1(n5400), .B2(n5658), .ZN(n5368)
         );
  OAI211_X1 U6101 ( .C1(n5406), .C2(n5370), .A(n5369), .B(n5368), .ZN(U3077)
         );
  AOI22_X1 U6102 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5399), .B1(n5371), 
        .B2(n5397), .ZN(n5374) );
  AOI22_X1 U6103 ( .A1(n5402), .A2(n5372), .B1(n5400), .B2(n5630), .ZN(n5373)
         );
  OAI211_X1 U6104 ( .C1(n5406), .C2(n5634), .A(n5374), .B(n5373), .ZN(U3081)
         );
  AOI22_X1 U6105 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5391), .B1(n5375), 
        .B2(n5389), .ZN(n5378) );
  AOI22_X1 U6106 ( .A1(n5376), .A2(n5420), .B1(n5392), .B2(n5672), .ZN(n5377)
         );
  OAI211_X1 U6107 ( .C1(n5379), .C2(n5396), .A(n5378), .B(n5377), .ZN(U3063)
         );
  AOI22_X1 U6108 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5391), .B1(n5380), 
        .B2(n5389), .ZN(n5383) );
  AOI22_X1 U6109 ( .A1(n5381), .A2(n5420), .B1(n5392), .B2(n5651), .ZN(n5382)
         );
  OAI211_X1 U6110 ( .C1(n5655), .C2(n5396), .A(n5383), .B(n5382), .ZN(U3066)
         );
  AOI22_X1 U6111 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5391), .B1(n5384), 
        .B2(n5389), .ZN(n5387) );
  AOI22_X1 U6112 ( .A1(n5385), .A2(n5420), .B1(n5392), .B2(n5680), .ZN(n5386)
         );
  OAI211_X1 U6113 ( .C1(n5388), .C2(n5396), .A(n5387), .B(n5386), .ZN(U3062)
         );
  AOI22_X1 U6114 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5391), .B1(n5390), 
        .B2(n5389), .ZN(n5395) );
  AOI22_X1 U6115 ( .A1(n5393), .A2(n5420), .B1(n5392), .B2(n5637), .ZN(n5394)
         );
  OAI211_X1 U6116 ( .C1(n5641), .C2(n5396), .A(n5395), .B(n5394), .ZN(U3064)
         );
  AOI22_X1 U6117 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5399), .B1(n5398), 
        .B2(n5397), .ZN(n5404) );
  AOI22_X1 U6118 ( .A1(n5402), .A2(n5401), .B1(n5400), .B2(n5644), .ZN(n5403)
         );
  OAI211_X1 U6119 ( .C1(n5406), .C2(n5405), .A(n5404), .B(n5403), .ZN(U3076)
         );
  AOI22_X1 U6120 ( .A1(n5511), .A2(n5409), .B1(n5408), .B2(n5407), .ZN(n5449)
         );
  NOR2_X1 U6121 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5410), .ZN(n5446)
         );
  INV_X1 U6122 ( .A(n5446), .ZN(n5413) );
  AOI211_X1 U6123 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5413), .A(n5412), .B(
        n5411), .ZN(n5419) );
  INV_X1 U6124 ( .A(n5443), .ZN(n5414) );
  OAI21_X1 U6125 ( .B1(n5420), .B2(n5414), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5415) );
  OAI21_X1 U6126 ( .B1(n5417), .B2(n5416), .A(n5415), .ZN(n5418) );
  NAND2_X1 U6127 ( .A1(n5419), .A2(n5418), .ZN(n5442) );
  NAND2_X1 U6128 ( .A1(n5442), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5423) );
  INV_X1 U6129 ( .A(n5420), .ZN(n5444) );
  OAI22_X1 U6130 ( .A1(n5444), .A2(n5538), .B1(n5632), .B2(n5443), .ZN(n5421)
         );
  AOI21_X1 U6131 ( .B1(n3434), .B2(n5446), .A(n5421), .ZN(n5422) );
  OAI211_X1 U6132 ( .C1(n5449), .C2(n5636), .A(n5423), .B(n5422), .ZN(U3057)
         );
  NAND2_X1 U6133 ( .A1(n5442), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5426) );
  OAI22_X1 U6134 ( .A1(n5444), .A2(n5526), .B1(n5646), .B2(n5443), .ZN(n5424)
         );
  AOI21_X1 U6135 ( .B1(n5648), .B2(n5446), .A(n5424), .ZN(n5425) );
  OAI211_X1 U6136 ( .C1(n5449), .C2(n5650), .A(n5426), .B(n5425), .ZN(U3052)
         );
  NAND2_X1 U6137 ( .A1(n5442), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5429) );
  OAI22_X1 U6138 ( .A1(n5444), .A2(n5546), .B1(n5674), .B2(n5443), .ZN(n5427)
         );
  AOI21_X1 U6139 ( .B1(n5676), .B2(n5446), .A(n5427), .ZN(n5428) );
  OAI211_X1 U6140 ( .C1(n5449), .C2(n5678), .A(n5429), .B(n5428), .ZN(U3055)
         );
  NAND2_X1 U6141 ( .A1(n5442), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5432) );
  OAI22_X1 U6142 ( .A1(n5444), .A2(n5534), .B1(n5639), .B2(n5443), .ZN(n5430)
         );
  AOI21_X1 U6143 ( .B1(n3435), .B2(n5446), .A(n5430), .ZN(n5431) );
  OAI211_X1 U6144 ( .C1(n5449), .C2(n5643), .A(n5432), .B(n5431), .ZN(U3056)
         );
  NAND2_X1 U6145 ( .A1(n5442), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5435) );
  OAI22_X1 U6146 ( .A1(n5444), .A2(n5522), .B1(n5660), .B2(n5443), .ZN(n5433)
         );
  AOI21_X1 U6147 ( .B1(n5662), .B2(n5446), .A(n5433), .ZN(n5434) );
  OAI211_X1 U6148 ( .C1(n5449), .C2(n5664), .A(n5435), .B(n5434), .ZN(U3053)
         );
  NAND2_X1 U6149 ( .A1(n5442), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5438) );
  OAI22_X1 U6150 ( .A1(n5444), .A2(n5551), .B1(n5683), .B2(n5443), .ZN(n5436)
         );
  AOI21_X1 U6151 ( .B1(n5687), .B2(n5446), .A(n5436), .ZN(n5437) );
  OAI211_X1 U6152 ( .C1(n5449), .C2(n5689), .A(n5438), .B(n5437), .ZN(U3054)
         );
  NAND2_X1 U6153 ( .A1(n5442), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5441) );
  OAI22_X1 U6154 ( .A1(n5444), .A2(n5530), .B1(n5667), .B2(n5443), .ZN(n5439)
         );
  AOI21_X1 U6155 ( .B1(n5669), .B2(n5446), .A(n5439), .ZN(n5440) );
  OAI211_X1 U6156 ( .C1(n5449), .C2(n5671), .A(n5441), .B(n5440), .ZN(U3059)
         );
  NAND2_X1 U6157 ( .A1(n5442), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5448) );
  OAI22_X1 U6158 ( .A1(n5444), .A2(n5542), .B1(n5653), .B2(n5443), .ZN(n5445)
         );
  AOI21_X1 U6159 ( .B1(n3433), .B2(n5446), .A(n5445), .ZN(n5447) );
  OAI211_X1 U6160 ( .C1(n5449), .C2(n5657), .A(n5448), .B(n5447), .ZN(U3058)
         );
  INV_X1 U6161 ( .A(n5454), .ZN(n5450) );
  AOI21_X1 U6162 ( .B1(n5451), .B2(n5257), .A(n5450), .ZN(n6766) );
  INV_X1 U6163 ( .A(n6766), .ZN(n7000) );
  XOR2_X1 U6164 ( .A(n5459), .B(n3451), .Z(n6996) );
  AOI22_X1 U6165 ( .A1(n6160), .A2(n6996), .B1(n6159), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5452) );
  OAI21_X1 U6166 ( .B1(n7000), .B2(n6151), .A(n5452), .ZN(U2852) );
  AND2_X1 U6167 ( .A1(n5454), .A2(n5453), .ZN(n5456) );
  OR2_X1 U6168 ( .A1(n5456), .A2(n5455), .ZN(n5692) );
  INV_X1 U6169 ( .A(n5457), .ZN(n5461) );
  AOI21_X1 U6170 ( .B1(n3451), .B2(n5459), .A(n5458), .ZN(n5460) );
  NOR2_X1 U6171 ( .A1(n5461), .A2(n5460), .ZN(n6855) );
  INV_X1 U6172 ( .A(n6855), .ZN(n5462) );
  OAI222_X1 U6173 ( .A1(n5692), .A2(n6151), .B1(n6150), .B2(n5463), .C1(n6148), 
        .C2(n5462), .ZN(U2851) );
  OAI21_X1 U6174 ( .B1(n3428), .B2(n5467), .A(n5466), .ZN(n5468) );
  INV_X1 U6175 ( .A(n5468), .ZN(n6859) );
  NAND2_X1 U6176 ( .A1(n6859), .A2(n6774), .ZN(n5472) );
  INV_X1 U6177 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5469) );
  NOR2_X1 U6178 ( .A1(n6894), .A2(n5469), .ZN(n6854) );
  NOR2_X1 U6179 ( .A1(n6778), .A2(n5691), .ZN(n5470) );
  AOI211_X1 U6180 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6854), 
        .B(n5470), .ZN(n5471) );
  OAI211_X1 U6181 ( .C1(n6748), .C2(n5692), .A(n5472), .B(n5471), .ZN(U2978)
         );
  INV_X1 U6182 ( .A(n5473), .ZN(n5479) );
  INV_X1 U6183 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6637) );
  OAI222_X1 U6184 ( .A1(n6387), .A2(n5509), .B1(n5839), .B2(n7148), .C1(n5836), 
        .C2(n6637), .ZN(U2891) );
  AND2_X1 U6185 ( .A1(n3781), .A2(n5482), .ZN(n7105) );
  NOR3_X1 U6186 ( .A1(n7115), .A2(n7110), .A3(n7117), .ZN(n7111) );
  NOR2_X1 U6187 ( .A1(n7105), .A2(n7111), .ZN(n5483) );
  NAND2_X1 U6188 ( .A1(n5483), .A2(n6894), .ZN(n5484) );
  NAND2_X1 U6189 ( .A1(n5935), .A2(n5485), .ZN(n5490) );
  NAND2_X1 U6190 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5486) );
  INV_X1 U6191 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U6192 ( .A1(n5617), .A2(n7143), .ZN(n5501) );
  NOR2_X1 U6193 ( .A1(n5503), .A2(n5501), .ZN(n5492) );
  AND2_X1 U6194 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  NAND2_X1 U6195 ( .A1(n6958), .A2(n6948), .ZN(n6971) );
  AND3_X1 U6196 ( .A1(n5494), .A2(EBX_REG_31__SCAN_IN), .A3(n5501), .ZN(n5495)
         );
  NAND2_X1 U6197 ( .A1(n5935), .A2(n5981), .ZN(n6970) );
  OAI22_X1 U6198 ( .A1(n7028), .A2(n5497), .B1(n5496), .B2(n6970), .ZN(n5498)
         );
  AOI21_X1 U6199 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6971), .A(n5498), .ZN(n5508)
         );
  AND2_X1 U6200 ( .A1(n5920), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6201 ( .A1(n7050), .A2(n7060), .ZN(n5506) );
  INV_X1 U6202 ( .A(n5501), .ZN(n5500) );
  NAND2_X1 U6203 ( .A1(n5982), .A2(n5500), .ZN(n7103) );
  AND2_X1 U6204 ( .A1(n7144), .A2(n7103), .ZN(n5934) );
  INV_X1 U6205 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U6206 ( .A1(n5940), .A2(n5501), .ZN(n5502) );
  NOR2_X1 U6207 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  OR2_X1 U6208 ( .A1(n5934), .A2(n5504), .ZN(n5505) );
  AOI22_X1 U6209 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5506), .B1(n7053), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U6210 ( .C1(n6979), .C2(n5509), .A(n5508), .B(n5507), .ZN(U2827)
         );
  INV_X1 U6211 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6643) );
  OAI222_X1 U6212 ( .A1(n6943), .A2(n6387), .B1(n5839), .B2(n7157), .C1(n5836), 
        .C2(n6643), .ZN(U2888) );
  INV_X1 U6213 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6652) );
  OAI222_X1 U6214 ( .A1(n7000), .A2(n6387), .B1(n5839), .B2(n7169), .C1(n5836), 
        .C2(n6652), .ZN(U2884) );
  INV_X1 U6215 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6650) );
  OAI222_X1 U6216 ( .A1(n6988), .A2(n6387), .B1(n5839), .B2(n7166), .C1(n5836), 
        .C2(n6650), .ZN(U2885) );
  INV_X1 U6217 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6647) );
  OAI222_X1 U6218 ( .A1(n6980), .A2(n6387), .B1(n5839), .B2(n7163), .C1(n6163), 
        .C2(n6647), .ZN(U2886) );
  INV_X1 U6219 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6645) );
  OAI222_X1 U6220 ( .A1(n6965), .A2(n6387), .B1(n5839), .B2(n7160), .C1(n6645), 
        .C2(n5836), .ZN(U2887) );
  INV_X1 U6221 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6639) );
  OAI222_X1 U6222 ( .A1(n5595), .A2(n6387), .B1(n5839), .B2(n7151), .C1(n5836), 
        .C2(n6639), .ZN(U2890) );
  INV_X1 U6223 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6641) );
  OAI222_X1 U6224 ( .A1(n6935), .A2(n6387), .B1(n5839), .B2(n7154), .C1(n5836), 
        .C2(n6641), .ZN(U2889) );
  INV_X1 U6225 ( .A(DATAI_8_), .ZN(n7172) );
  INV_X1 U6226 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6654) );
  OAI222_X1 U6227 ( .A1(n5692), .A2(n6387), .B1(n5839), .B2(n7172), .C1(n5836), 
        .C2(n6654), .ZN(U2883) );
  AOI22_X1 U6228 ( .A1(n5511), .A2(n5516), .B1(n5510), .B2(n5621), .ZN(n5558)
         );
  AOI21_X1 U6229 ( .B1(n5552), .B2(n5550), .A(n5513), .ZN(n5514) );
  AOI21_X1 U6230 ( .B1(n5516), .B2(n5515), .A(n5514), .ZN(n5517) );
  NOR2_X1 U6231 ( .A1(n5517), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5521) );
  NOR2_X1 U6232 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5518), .ZN(n5555)
         );
  INV_X1 U6233 ( .A(n5625), .ZN(n5519) );
  OAI22_X1 U6234 ( .A1(n5552), .A2(n5660), .B1(n5522), .B2(n5550), .ZN(n5523)
         );
  AOI21_X1 U6235 ( .B1(n5554), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n5523), 
        .ZN(n5525) );
  NAND2_X1 U6236 ( .A1(n5662), .A2(n5555), .ZN(n5524) );
  OAI211_X1 U6237 ( .C1(n5558), .C2(n5664), .A(n5525), .B(n5524), .ZN(U3037)
         );
  OAI22_X1 U6238 ( .A1(n5552), .A2(n5646), .B1(n5526), .B2(n5550), .ZN(n5527)
         );
  AOI21_X1 U6239 ( .B1(n5554), .B2(INSTQUEUE_REG_2__0__SCAN_IN), .A(n5527), 
        .ZN(n5529) );
  NAND2_X1 U6240 ( .A1(n5648), .A2(n5555), .ZN(n5528) );
  OAI211_X1 U6241 ( .C1(n5558), .C2(n5650), .A(n5529), .B(n5528), .ZN(U3036)
         );
  OAI22_X1 U6242 ( .A1(n5552), .A2(n5667), .B1(n5530), .B2(n5550), .ZN(n5531)
         );
  AOI21_X1 U6243 ( .B1(n5554), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n5531), 
        .ZN(n5533) );
  NAND2_X1 U6244 ( .A1(n5669), .A2(n5555), .ZN(n5532) );
  OAI211_X1 U6245 ( .C1(n5558), .C2(n5671), .A(n5533), .B(n5532), .ZN(U3043)
         );
  OAI22_X1 U6246 ( .A1(n5552), .A2(n5639), .B1(n5534), .B2(n5550), .ZN(n5535)
         );
  AOI21_X1 U6247 ( .B1(n5554), .B2(INSTQUEUE_REG_2__4__SCAN_IN), .A(n5535), 
        .ZN(n5537) );
  NAND2_X1 U6248 ( .A1(n3435), .A2(n5555), .ZN(n5536) );
  OAI211_X1 U6249 ( .C1(n5558), .C2(n5643), .A(n5537), .B(n5536), .ZN(U3040)
         );
  OAI22_X1 U6250 ( .A1(n5552), .A2(n5632), .B1(n5538), .B2(n5550), .ZN(n5539)
         );
  AOI21_X1 U6251 ( .B1(n5554), .B2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n5539), 
        .ZN(n5541) );
  NAND2_X1 U6252 ( .A1(n3434), .A2(n5555), .ZN(n5540) );
  OAI211_X1 U6253 ( .C1(n5558), .C2(n5636), .A(n5541), .B(n5540), .ZN(U3041)
         );
  OAI22_X1 U6254 ( .A1(n5552), .A2(n5653), .B1(n5542), .B2(n5550), .ZN(n5543)
         );
  AOI21_X1 U6255 ( .B1(n5554), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n5543), 
        .ZN(n5545) );
  NAND2_X1 U6256 ( .A1(n3433), .A2(n5555), .ZN(n5544) );
  OAI211_X1 U6257 ( .C1(n5558), .C2(n5657), .A(n5545), .B(n5544), .ZN(U3042)
         );
  OAI22_X1 U6258 ( .A1(n5552), .A2(n5674), .B1(n5546), .B2(n5550), .ZN(n5547)
         );
  AOI21_X1 U6259 ( .B1(n5554), .B2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n5547), 
        .ZN(n5549) );
  NAND2_X1 U6260 ( .A1(n5676), .A2(n5555), .ZN(n5548) );
  OAI211_X1 U6261 ( .C1(n5558), .C2(n5678), .A(n5549), .B(n5548), .ZN(U3039)
         );
  OAI22_X1 U6262 ( .A1(n5552), .A2(n5683), .B1(n5551), .B2(n5550), .ZN(n5553)
         );
  AOI21_X1 U6263 ( .B1(n5554), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n5553), 
        .ZN(n5557) );
  NAND2_X1 U6264 ( .A1(n5687), .A2(n5555), .ZN(n5556) );
  OAI211_X1 U6265 ( .C1(n5558), .C2(n5689), .A(n5557), .B(n5556), .ZN(U3038)
         );
  INV_X1 U6266 ( .A(n5561), .ZN(n5564) );
  INV_X1 U6267 ( .A(n5455), .ZN(n5563) );
  AOI21_X1 U6268 ( .B1(n5564), .B2(n5563), .A(n5562), .ZN(n5569) );
  INV_X1 U6269 ( .A(n5565), .ZN(n5607) );
  AOI22_X1 U6270 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6906), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5566) );
  OAI21_X1 U6271 ( .B1(n6778), .B2(n5607), .A(n5566), .ZN(n5567) );
  AOI21_X1 U6272 ( .B1(n5569), .B2(n6773), .A(n5567), .ZN(n5568) );
  OAI21_X1 U6273 ( .B1(n6880), .B2(n7062), .A(n5568), .ZN(U2977) );
  INV_X1 U6274 ( .A(n5569), .ZN(n5608) );
  NAND2_X1 U6275 ( .A1(n5457), .A2(n5570), .ZN(n5571) );
  NAND2_X1 U6276 ( .A1(n5575), .A2(n5571), .ZN(n5613) );
  INV_X1 U6277 ( .A(n5613), .ZN(n6879) );
  AOI22_X1 U6278 ( .A1(n6160), .A2(n6879), .B1(n6159), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5572) );
  OAI21_X1 U6279 ( .B1(n5608), .B2(n6151), .A(n5572), .ZN(U2850) );
  INV_X1 U6280 ( .A(DATAI_9_), .ZN(n7175) );
  INV_X1 U6281 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6656) );
  OAI222_X1 U6282 ( .A1(n5608), .A2(n6387), .B1(n5839), .B2(n7175), .C1(n6163), 
        .C2(n6656), .ZN(U2882) );
  OAI21_X1 U6283 ( .B1(n5562), .B2(n5574), .A(n5700), .ZN(n5606) );
  AOI21_X1 U6284 ( .B1(n5576), .B2(n5575), .A(n5704), .ZN(n6871) );
  AOI22_X1 U6285 ( .A1(n6871), .A2(n6160), .B1(EBX_REG_10__SCAN_IN), .B2(n6159), .ZN(n5577) );
  OAI21_X1 U6286 ( .B1(n5606), .B2(n6151), .A(n5577), .ZN(U2849) );
  NAND2_X1 U6287 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6950) );
  NOR2_X1 U6288 ( .A1(n6950), .A2(n6949), .ZN(n6956) );
  NAND4_X1 U6289 ( .A1(n6956), .A2(REIP_REG_4__SCAN_IN), .A3(
        REIP_REG_5__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5579) );
  NOR2_X1 U6290 ( .A1(n6958), .A2(n5579), .ZN(n6995) );
  INV_X1 U6291 ( .A(n6995), .ZN(n5578) );
  INV_X1 U6292 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7006) );
  NOR3_X1 U6293 ( .A1(n5578), .A2(n5469), .A3(n7006), .ZN(n5584) );
  INV_X1 U6294 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U6295 ( .A1(n5584), .A2(n6679), .ZN(n5611) );
  NOR3_X1 U6296 ( .A1(n5579), .A2(n7006), .A3(n5469), .ZN(n5819) );
  NAND2_X1 U6297 ( .A1(n5819), .A2(n6948), .ZN(n5580) );
  NAND2_X1 U6298 ( .A1(n6971), .A2(n5580), .ZN(n5693) );
  NAND2_X1 U6299 ( .A1(n5611), .A2(n5693), .ZN(n5583) );
  INV_X1 U6300 ( .A(n6948), .ZN(n6951) );
  AOI21_X1 U6301 ( .B1(n7035), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7034), 
        .ZN(n5581) );
  OAI21_X1 U6302 ( .B1(n7060), .B2(n5602), .A(n5581), .ZN(n5582) );
  AOI21_X1 U6303 ( .B1(n5583), .B2(REIP_REG_10__SCAN_IN), .A(n5582), .ZN(n5588) );
  NAND2_X1 U6304 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5584), .ZN(n5754) );
  AOI22_X1 U6305 ( .A1(EBX_REG_10__SCAN_IN), .A2(n7053), .B1(n7056), .B2(n6871), .ZN(n5585) );
  OAI21_X1 U6306 ( .B1(REIP_REG_10__SCAN_IN), .B2(n5754), .A(n5585), .ZN(n5586) );
  INV_X1 U6307 ( .A(n5586), .ZN(n5587) );
  OAI211_X1 U6308 ( .C1(n5606), .C2(n7014), .A(n5588), .B(n5587), .ZN(U2817)
         );
  INV_X1 U6309 ( .A(n5589), .ZN(n5592) );
  INV_X1 U6310 ( .A(n6970), .ZN(n6947) );
  AOI22_X1 U6311 ( .A1(n6947), .A2(n4854), .B1(n7053), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5591) );
  INV_X1 U6312 ( .A(n6958), .ZN(n6112) );
  NAND2_X1 U6313 ( .A1(n6112), .A2(n5590), .ZN(n6930) );
  OAI211_X1 U6314 ( .C1(n5592), .C2(n7028), .A(n5591), .B(n6930), .ZN(n5597)
         );
  AOI22_X1 U6315 ( .A1(n7017), .A2(n4725), .B1(n6951), .B2(REIP_REG_1__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6316 ( .A1(n7035), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5593)
         );
  OAI211_X1 U6317 ( .C1(n6979), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5596)
         );
  OR2_X1 U6318 ( .A1(n5597), .A2(n5596), .ZN(U2826) );
  XNOR2_X1 U6319 ( .A(n6428), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5599)
         );
  NAND2_X1 U6320 ( .A1(n5598), .A2(n5599), .ZN(n5718) );
  OAI21_X1 U6321 ( .B1(n5598), .B2(n5599), .A(n5718), .ZN(n5600) );
  INV_X1 U6322 ( .A(n5600), .ZN(n6875) );
  NAND2_X1 U6323 ( .A1(n6875), .A2(n6774), .ZN(n5605) );
  INV_X1 U6324 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5601) );
  NOR2_X1 U6325 ( .A1(n6894), .A2(n5601), .ZN(n6870) );
  NOR2_X1 U6326 ( .A1(n6778), .A2(n5602), .ZN(n5603) );
  AOI211_X1 U6327 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6870), 
        .B(n5603), .ZN(n5604) );
  OAI211_X1 U6328 ( .C1(n6748), .C2(n5606), .A(n5605), .B(n5604), .ZN(U2976)
         );
  INV_X1 U6329 ( .A(DATAI_10_), .ZN(n7178) );
  INV_X1 U6330 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6658) );
  OAI222_X1 U6331 ( .A1(n5606), .A2(n6387), .B1(n5839), .B2(n7178), .C1(n5836), 
        .C2(n6658), .ZN(U2881) );
  OAI22_X1 U6332 ( .A1(n5608), .A2(n7014), .B1(n7060), .B2(n5607), .ZN(n5615)
         );
  OAI22_X1 U6333 ( .A1(n5609), .A2(n7025), .B1(n6679), .B2(n5693), .ZN(n5610)
         );
  AOI211_X1 U6334 ( .C1(n7035), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n7034), 
        .B(n5610), .ZN(n5612) );
  OAI211_X1 U6335 ( .C1(n5613), .C2(n7028), .A(n5612), .B(n5611), .ZN(n5614)
         );
  OR2_X1 U6336 ( .A1(n5615), .A2(n5614), .ZN(U2818) );
  AOI21_X1 U6337 ( .B1(n5684), .B2(n5623), .A(n5617), .ZN(n5619) );
  NOR2_X1 U6338 ( .A1(n5619), .A2(n5618), .ZN(n5628) );
  NOR2_X1 U6339 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5622), .ZN(n5686)
         );
  INV_X1 U6340 ( .A(n5624), .ZN(n5627) );
  AOI211_X1 U6341 ( .C1(n5628), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5629)
         );
  OAI21_X1 U6342 ( .B1(n5686), .B2(n7110), .A(n5629), .ZN(n5679) );
  AOI22_X1 U6343 ( .A1(n5681), .A2(n5630), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5679), .ZN(n5631) );
  OAI21_X1 U6344 ( .B1(n5684), .B2(n5632), .A(n5631), .ZN(n5633) );
  AOI21_X1 U6345 ( .B1(n3434), .B2(n5686), .A(n5633), .ZN(n5635) );
  OAI21_X1 U6346 ( .B1(n5690), .B2(n5636), .A(n5635), .ZN(U3105) );
  AOI22_X1 U6347 ( .A1(n5681), .A2(n5637), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5679), .ZN(n5638) );
  OAI21_X1 U6348 ( .B1(n5684), .B2(n5639), .A(n5638), .ZN(n5640) );
  AOI21_X1 U6349 ( .B1(n3435), .B2(n5686), .A(n5640), .ZN(n5642) );
  OAI21_X1 U6350 ( .B1(n5690), .B2(n5643), .A(n5642), .ZN(U3104) );
  AOI22_X1 U6351 ( .A1(n5681), .A2(n5644), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5679), .ZN(n5645) );
  OAI21_X1 U6352 ( .B1(n5684), .B2(n5646), .A(n5645), .ZN(n5647) );
  AOI21_X1 U6353 ( .B1(n5648), .B2(n5686), .A(n5647), .ZN(n5649) );
  OAI21_X1 U6354 ( .B1(n5690), .B2(n5650), .A(n5649), .ZN(U3100) );
  AOI22_X1 U6355 ( .A1(n5681), .A2(n5651), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5679), .ZN(n5652) );
  OAI21_X1 U6356 ( .B1(n5684), .B2(n5653), .A(n5652), .ZN(n5654) );
  AOI21_X1 U6357 ( .B1(n3433), .B2(n5686), .A(n5654), .ZN(n5656) );
  OAI21_X1 U6358 ( .B1(n5690), .B2(n5657), .A(n5656), .ZN(U3106) );
  AOI22_X1 U6359 ( .A1(n5681), .A2(n5658), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5679), .ZN(n5659) );
  OAI21_X1 U6360 ( .B1(n5684), .B2(n5660), .A(n5659), .ZN(n5661) );
  AOI21_X1 U6361 ( .B1(n5662), .B2(n5686), .A(n5661), .ZN(n5663) );
  OAI21_X1 U6362 ( .B1(n5690), .B2(n5664), .A(n5663), .ZN(U3101) );
  AOI22_X1 U6363 ( .A1(n5681), .A2(n5665), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5679), .ZN(n5666) );
  OAI21_X1 U6364 ( .B1(n5684), .B2(n5667), .A(n5666), .ZN(n5668) );
  AOI21_X1 U6365 ( .B1(n5669), .B2(n5686), .A(n5668), .ZN(n5670) );
  OAI21_X1 U6366 ( .B1(n5690), .B2(n5671), .A(n5670), .ZN(U3107) );
  AOI22_X1 U6367 ( .A1(n5681), .A2(n5672), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5679), .ZN(n5673) );
  OAI21_X1 U6368 ( .B1(n5684), .B2(n5674), .A(n5673), .ZN(n5675) );
  AOI21_X1 U6369 ( .B1(n5676), .B2(n5686), .A(n5675), .ZN(n5677) );
  OAI21_X1 U6370 ( .B1(n5690), .B2(n5678), .A(n5677), .ZN(U3103) );
  AOI22_X1 U6371 ( .A1(n5681), .A2(n5680), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5679), .ZN(n5682) );
  OAI21_X1 U6372 ( .B1(n5684), .B2(n5683), .A(n5682), .ZN(n5685) );
  AOI21_X1 U6373 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5688) );
  OAI21_X1 U6374 ( .B1(n5690), .B2(n5689), .A(n5688), .ZN(U3102) );
  OAI22_X1 U6375 ( .A1(n5692), .A2(n7014), .B1(n5691), .B2(n7060), .ZN(n5699)
         );
  NAND2_X1 U6376 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6995), .ZN(n5694) );
  AOI21_X1 U6377 ( .B1(n5469), .B2(n5694), .A(n5693), .ZN(n5698) );
  AOI22_X1 U6378 ( .A1(EBX_REG_8__SCAN_IN), .A2(n7053), .B1(n7056), .B2(n6855), 
        .ZN(n5695) );
  OAI211_X1 U6379 ( .C1(n7050), .C2(n5696), .A(n5695), .B(n7023), .ZN(n5697)
         );
  OR3_X1 U6380 ( .A1(n5699), .A2(n5698), .A3(n5697), .ZN(U2819) );
  AOI21_X1 U6381 ( .B1(n5701), .B2(n5700), .A(n3445), .ZN(n5727) );
  INV_X1 U6382 ( .A(n5727), .ZN(n5717) );
  NAND2_X1 U6383 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5755) );
  NOR2_X1 U6384 ( .A1(n5755), .A2(n6679), .ZN(n5818) );
  AND2_X1 U6385 ( .A1(n5818), .A2(n5819), .ZN(n5702) );
  OAI21_X1 U6386 ( .B1(n6958), .B2(n5702), .A(n6948), .ZN(n5789) );
  INV_X1 U6387 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5714) );
  OR2_X1 U6388 ( .A1(n5704), .A2(n5703), .ZN(n5705) );
  NAND2_X1 U6389 ( .A1(n5744), .A2(n5705), .ZN(n6896) );
  OAI22_X1 U6390 ( .A1(n5714), .A2(n7025), .B1(n7028), .B2(n6896), .ZN(n5706)
         );
  AOI21_X1 U6391 ( .B1(n7017), .B2(n5723), .A(n5706), .ZN(n5707) );
  INV_X1 U6392 ( .A(n5707), .ZN(n5710) );
  OAI21_X1 U6393 ( .B1(n7050), .B2(n5708), .A(n7023), .ZN(n5709) );
  AOI211_X1 U6394 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5789), .A(n5710), .B(n5709), .ZN(n5713) );
  NOR2_X1 U6395 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5754), .ZN(n5711) );
  NAND2_X1 U6396 ( .A1(n5711), .A2(REIP_REG_10__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U6397 ( .C1(n5717), .C2(n7014), .A(n5713), .B(n5712), .ZN(U2816)
         );
  OAI22_X1 U6398 ( .A1(n6148), .A2(n6896), .B1(n5714), .B2(n6150), .ZN(n5715)
         );
  AOI21_X1 U6399 ( .B1(n5727), .B2(n5782), .A(n5715), .ZN(n5716) );
  INV_X1 U6400 ( .A(n5716), .ZN(U2848) );
  INV_X1 U6401 ( .A(DATAI_11_), .ZN(n7181) );
  INV_X1 U6402 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6660) );
  OAI222_X1 U6403 ( .A1(n5717), .A2(n6387), .B1(n5839), .B2(n7181), .C1(n5836), 
        .C2(n6660), .ZN(U2880) );
  INV_X1 U6404 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6868) );
  OAI21_X1 U6405 ( .B1(n6868), .B2(n6428), .A(n5718), .ZN(n5719) );
  INV_X1 U6406 ( .A(n5719), .ZN(n5722) );
  OAI21_X1 U6407 ( .B1(n3519), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5758), 
        .ZN(n5721) );
  OAI211_X1 U6408 ( .C1(n3519), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5719), .B(n5758), .ZN(n5759) );
  INV_X1 U6409 ( .A(n5759), .ZN(n5720) );
  AOI21_X1 U6410 ( .B1(n5722), .B2(n5721), .A(n5720), .ZN(n6899) );
  INV_X1 U6411 ( .A(n6899), .ZN(n5729) );
  INV_X1 U6412 ( .A(n5723), .ZN(n5725) );
  AOI22_X1 U6413 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6906), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5724) );
  OAI21_X1 U6414 ( .B1(n6778), .B2(n5725), .A(n5724), .ZN(n5726) );
  AOI21_X1 U6415 ( .B1(n5727), .B2(n6773), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6416 ( .B1(n5729), .B2(n7062), .A(n5728), .ZN(U2975) );
  XOR2_X1 U6417 ( .A(n5730), .B(n5731), .Z(n5801) );
  AND2_X1 U6418 ( .A1(n3440), .A2(n5732), .ZN(n5733) );
  OR2_X1 U6419 ( .A1(n5733), .A2(n5812), .ZN(n5785) );
  INV_X1 U6420 ( .A(n5785), .ZN(n5739) );
  NAND2_X1 U6421 ( .A1(n6906), .A2(REIP_REG_13__SCAN_IN), .ZN(n5795) );
  INV_X1 U6422 ( .A(n5795), .ZN(n5738) );
  INV_X1 U6424 ( .A(n6803), .ZN(n5735) );
  INV_X1 U6425 ( .A(n6901), .ZN(n5734) );
  AOI21_X1 U6426 ( .B1(n6816), .B2(n5735), .A(n5734), .ZN(n6806) );
  OAI33_X1 U6427 ( .A1(1'b0), .A2(n6806), .A3(n4576), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6902), .B3(n6889), .ZN(n5737)
         );
  AOI211_X1 U6428 ( .C1(n6926), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5740)
         );
  OAI21_X1 U6429 ( .B1(n5801), .B2(n6590), .A(n5740), .ZN(U3005) );
  OAI21_X1 U6430 ( .B1(n3445), .B2(n4018), .A(n5742), .ZN(n5767) );
  NAND2_X1 U6431 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  NAND2_X1 U6432 ( .A1(n3440), .A2(n5745), .ZN(n6886) );
  INV_X1 U6433 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5746) );
  OAI22_X1 U6434 ( .A1(n6886), .A2(n6148), .B1(n5746), .B2(n6150), .ZN(n5747)
         );
  INV_X1 U6435 ( .A(n5747), .ZN(n5748) );
  OAI21_X1 U6436 ( .B1(n5767), .B2(n6151), .A(n5748), .ZN(U2847) );
  INV_X1 U6437 ( .A(n5763), .ZN(n5753) );
  OAI21_X1 U6438 ( .B1(n7050), .B2(n5749), .A(n7023), .ZN(n5752) );
  AOI22_X1 U6439 ( .A1(EBX_REG_12__SCAN_IN), .A2(n7053), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5789), .ZN(n5750) );
  OAI21_X1 U6440 ( .B1(n7028), .B2(n6886), .A(n5750), .ZN(n5751) );
  AOI211_X1 U6441 ( .C1(n7017), .C2(n5753), .A(n5752), .B(n5751), .ZN(n5757)
         );
  NOR2_X1 U6442 ( .A1(n5755), .A2(n5754), .ZN(n5816) );
  INV_X1 U6443 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U6444 ( .A1(n5816), .A2(n6682), .ZN(n5756) );
  OAI211_X1 U6445 ( .C1(n5767), .C2(n7014), .A(n5757), .B(n5756), .ZN(U2815)
         );
  NAND2_X1 U6446 ( .A1(n5759), .A2(n5758), .ZN(n5762) );
  XNOR2_X1 U6447 ( .A(n6428), .B(n5760), .ZN(n5761) );
  XNOR2_X1 U6448 ( .A(n5762), .B(n5761), .ZN(n6891) );
  NAND2_X1 U6449 ( .A1(n6891), .A2(n6774), .ZN(n5766) );
  NOR2_X1 U6450 ( .A1(n6894), .A2(n6682), .ZN(n6887) );
  NOR2_X1 U6451 ( .A1(n6778), .A2(n5763), .ZN(n5764) );
  AOI211_X1 U6452 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6887), 
        .B(n5764), .ZN(n5765) );
  OAI211_X1 U6453 ( .C1(n6748), .C2(n5767), .A(n5766), .B(n5765), .ZN(U2974)
         );
  INV_X1 U6454 ( .A(DATAI_12_), .ZN(n7184) );
  OAI222_X1 U6455 ( .A1(n5767), .A2(n6387), .B1(n5839), .B2(n7184), .C1(n5836), 
        .C2(n4003), .ZN(U2879) );
  NOR2_X1 U6456 ( .A1(n5770), .A2(n3542), .ZN(n5771) );
  XNOR2_X1 U6457 ( .A(n5768), .B(n5771), .ZN(n5844) );
  OR2_X1 U6458 ( .A1(n5814), .A2(n5772), .ZN(n5773) );
  NAND2_X1 U6459 ( .A1(n6105), .A2(n5773), .ZN(n7020) );
  INV_X1 U6460 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6688) );
  OAI22_X1 U6461 ( .A1(n7020), .A2(n6897), .B1(n6688), .B2(n6894), .ZN(n5776)
         );
  NOR2_X1 U6462 ( .A1(n5774), .A2(n5777), .ZN(n5775) );
  AOI211_X1 U6463 ( .C1(n6909), .C2(n5777), .A(n5776), .B(n5775), .ZN(n5778)
         );
  OAI21_X1 U6464 ( .B1(n5844), .B2(n6590), .A(n5778), .ZN(U3003) );
  XOR2_X1 U6465 ( .A(n5780), .B(n5779), .Z(n5799) );
  OAI22_X1 U6466 ( .A1(n5785), .A2(n6148), .B1(n5786), .B2(n6150), .ZN(n5781)
         );
  AOI21_X1 U6467 ( .B1(n5799), .B2(n5782), .A(n5781), .ZN(n5783) );
  INV_X1 U6468 ( .A(n5783), .ZN(U2846) );
  INV_X1 U6469 ( .A(n5799), .ZN(n5838) );
  INV_X1 U6470 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U6471 ( .A1(n6682), .A2(n6685), .ZN(n5817) );
  AOI21_X1 U6472 ( .B1(n6682), .B2(n6685), .A(n5817), .ZN(n5793) );
  OAI21_X1 U6473 ( .B1(n7050), .B2(n5784), .A(n7023), .ZN(n5792) );
  OAI22_X1 U6474 ( .A1(n5786), .A2(n7025), .B1(n7028), .B2(n5785), .ZN(n5788)
         );
  NOR2_X1 U6475 ( .A1(n7060), .A2(n5797), .ZN(n5787) );
  AOI211_X1 U6476 ( .C1(REIP_REG_13__SCAN_IN), .C2(n5789), .A(n5788), .B(n5787), .ZN(n5790) );
  INV_X1 U6477 ( .A(n5790), .ZN(n5791) );
  AOI211_X1 U6478 ( .C1(n5816), .C2(n5793), .A(n5792), .B(n5791), .ZN(n5794)
         );
  OAI21_X1 U6479 ( .B1(n5838), .B2(n7014), .A(n5794), .ZN(U2814) );
  NAND2_X1 U6480 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5796)
         );
  OAI211_X1 U6481 ( .C1(n6778), .C2(n5797), .A(n5796), .B(n5795), .ZN(n5798)
         );
  AOI21_X1 U6482 ( .B1(n5799), .B2(n6773), .A(n5798), .ZN(n5800) );
  OAI21_X1 U6483 ( .B1(n5801), .B2(n7062), .A(n5800), .ZN(U2973) );
  OAI21_X1 U6484 ( .B1(n5802), .B2(n5804), .A(n5803), .ZN(n7015) );
  INV_X1 U6485 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5805) );
  OAI22_X1 U6486 ( .A1(n7020), .A2(n6148), .B1(n5805), .B2(n6150), .ZN(n5806)
         );
  INV_X1 U6487 ( .A(n5806), .ZN(n5807) );
  OAI21_X1 U6488 ( .B1(n7015), .B2(n6151), .A(n5807), .ZN(U2844) );
  INV_X1 U6489 ( .A(n5802), .ZN(n5808) );
  OAI21_X1 U6490 ( .B1(n5810), .B2(n5809), .A(n5808), .ZN(n5837) );
  NOR2_X1 U6491 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  OR2_X1 U6492 ( .A1(n5814), .A2(n5813), .ZN(n5834) );
  INV_X1 U6493 ( .A(n5834), .ZN(n6805) );
  NAND2_X1 U6494 ( .A1(n7035), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5815)
         );
  OAI211_X1 U6495 ( .C1(n7060), .C2(n5830), .A(n7023), .B(n5815), .ZN(n5823)
         );
  NAND2_X1 U6496 ( .A1(n5817), .A2(n5816), .ZN(n5821) );
  NAND4_X1 U6497 ( .A1(n5819), .A2(n5818), .A3(n5817), .A4(
        REIP_REG_14__SCAN_IN), .ZN(n5849) );
  INV_X1 U6498 ( .A(n5849), .ZN(n6108) );
  OAI21_X1 U6499 ( .B1(n6958), .B2(n6108), .A(n6948), .ZN(n7011) );
  AOI22_X1 U6500 ( .A1(EBX_REG_14__SCAN_IN), .A2(n7053), .B1(
        REIP_REG_14__SCAN_IN), .B2(n7011), .ZN(n5820) );
  OAI21_X1 U6501 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5821), .A(n5820), .ZN(n5822) );
  AOI211_X1 U6502 ( .C1(n6805), .C2(n7056), .A(n5823), .B(n5822), .ZN(n5824)
         );
  OAI21_X1 U6503 ( .B1(n5837), .B2(n7014), .A(n5824), .ZN(U2813) );
  INV_X1 U6504 ( .A(DATAI_15_), .ZN(n7195) );
  INV_X1 U6505 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6669) );
  OAI222_X1 U6506 ( .A1(n7015), .A2(n6387), .B1(n5839), .B2(n7195), .C1(n5836), 
        .C2(n6669), .ZN(U2876) );
  NOR2_X1 U6507 ( .A1(n3463), .A2(n5827), .ZN(n5828) );
  XNOR2_X1 U6508 ( .A(n5825), .B(n5828), .ZN(n6808) );
  NAND2_X1 U6509 ( .A1(n6808), .A2(n6774), .ZN(n5833) );
  INV_X1 U6510 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5829) );
  NOR2_X1 U6511 ( .A1(n6894), .A2(n5829), .ZN(n6804) );
  NOR2_X1 U6512 ( .A1(n6778), .A2(n5830), .ZN(n5831) );
  AOI211_X1 U6513 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6804), 
        .B(n5831), .ZN(n5832) );
  OAI211_X1 U6514 ( .C1(n6748), .C2(n5837), .A(n5833), .B(n5832), .ZN(U2972)
         );
  INV_X1 U6515 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5835) );
  OAI222_X1 U6516 ( .A1(n5837), .A2(n6151), .B1(n6150), .B2(n5835), .C1(n6148), 
        .C2(n5834), .ZN(U2845) );
  INV_X1 U6517 ( .A(DATAI_14_), .ZN(n7192) );
  INV_X1 U6518 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6665) );
  OAI222_X1 U6519 ( .A1(n5837), .A2(n6387), .B1(n5839), .B2(n7192), .C1(n5836), 
        .C2(n6665), .ZN(U2877) );
  INV_X1 U6520 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6663) );
  INV_X1 U6521 ( .A(DATAI_13_), .ZN(n7188) );
  OAI222_X1 U6522 ( .A1(n6163), .A2(n6663), .B1(n5839), .B2(n7188), .C1(n6387), 
        .C2(n5838), .ZN(U2878) );
  INV_X1 U6523 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5840) );
  OAI22_X1 U6524 ( .A1(n6753), .A2(n5840), .B1(n6894), .B2(n6688), .ZN(n5841)
         );
  AOI21_X1 U6525 ( .B1(n6477), .B2(n7018), .A(n5841), .ZN(n5843) );
  OR2_X1 U6526 ( .A1(n7015), .A2(n6748), .ZN(n5842) );
  OAI211_X1 U6527 ( .C1(n5844), .C2(n7062), .A(n5843), .B(n5842), .ZN(U2971)
         );
  INV_X1 U6528 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5858) );
  INV_X1 U6529 ( .A(n6000), .ZN(n5846) );
  NOR2_X1 U6530 ( .A1(n3448), .A2(n5846), .ZN(n5848) );
  OAI21_X1 U6531 ( .B1(n5848), .B2(n5847), .A(n5989), .ZN(n6513) );
  OAI222_X1 U6532 ( .A1(n5858), .A2(n6150), .B1(n6151), .B2(n5845), .C1(n6148), 
        .C2(n6513), .ZN(U2831) );
  AND2_X1 U6533 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n6001) );
  AND2_X1 U6534 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5931) );
  INV_X1 U6535 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6702) );
  INV_X1 U6536 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7049) );
  NOR2_X1 U6537 ( .A1(n5849), .A2(n6688), .ZN(n6110) );
  NAND2_X1 U6538 ( .A1(n6110), .A2(REIP_REG_16__SCAN_IN), .ZN(n6067) );
  INV_X1 U6539 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6691) );
  NOR2_X1 U6540 ( .A1(n6067), .A2(n6691), .ZN(n6096) );
  NAND4_X1 U6541 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(n6096), .ZN(n6069) );
  NOR2_X1 U6542 ( .A1(n7049), .A2(n6069), .ZN(n5852) );
  AND3_X1 U6543 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        n5852), .ZN(n5850) );
  NAND2_X1 U6544 ( .A1(n6948), .A2(n5850), .ZN(n6042) );
  NOR2_X1 U6545 ( .A1(n6702), .A2(n6042), .ZN(n6028) );
  NAND3_X1 U6546 ( .A1(n6001), .A2(n5931), .A3(n6028), .ZN(n5851) );
  NAND2_X1 U6547 ( .A1(n6971), .A2(n5851), .ZN(n5994) );
  INV_X1 U6548 ( .A(n5994), .ZN(n5861) );
  NAND2_X1 U6549 ( .A1(n6112), .A2(n5852), .ZN(n6070) );
  INV_X1 U6550 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6353) );
  NOR2_X1 U6551 ( .A1(n6070), .A2(n6353), .ZN(n6053) );
  NAND2_X1 U6552 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6053), .ZN(n6044) );
  INV_X1 U6553 ( .A(n6044), .ZN(n5853) );
  NAND2_X1 U6554 ( .A1(n6030), .A2(n6001), .ZN(n6004) );
  INV_X1 U6555 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6709) );
  NOR3_X1 U6556 ( .A1(n6004), .A2(REIP_REG_28__SCAN_IN), .A3(n6709), .ZN(n5855) );
  NOR2_X1 U6557 ( .A1(n7050), .A2(n5863), .ZN(n5854) );
  AOI211_X1 U6558 ( .C1(n7017), .C2(n5856), .A(n5855), .B(n5854), .ZN(n5857)
         );
  OAI21_X1 U6559 ( .B1(n7025), .B2(n5858), .A(n5857), .ZN(n5860) );
  NOR2_X1 U6560 ( .A1(n6513), .A2(n7028), .ZN(n5859) );
  AOI211_X1 U6561 ( .C1(n5861), .C2(REIP_REG_28__SCAN_IN), .A(n5860), .B(n5859), .ZN(n5862) );
  OAI21_X1 U6562 ( .B1(n5845), .B2(n7014), .A(n5862), .ZN(U2799) );
  OR2_X1 U6563 ( .A1(n5864), .A2(n5863), .ZN(n5866) );
  INV_X1 U6564 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U6565 ( .A(n5866), .B(n5865), .ZN(n6393) );
  OR2_X1 U6566 ( .A1(n5868), .A2(n5867), .ZN(n5889) );
  AOI22_X1 U6567 ( .A1(n4189), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5874) );
  AOI22_X1 U6568 ( .A1(n4190), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5869), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5873) );
  AOI22_X1 U6569 ( .A1(n3738), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U6570 ( .A1(n5870), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5871) );
  NAND4_X1 U6571 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n5882)
         );
  AOI22_X1 U6572 ( .A1(n3653), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4274), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5880) );
  AOI22_X1 U6573 ( .A1(n5875), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5879) );
  AOI22_X1 U6574 ( .A1(n4318), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5878) );
  AOI22_X1 U6575 ( .A1(n4319), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5877) );
  NAND4_X1 U6576 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n5881)
         );
  NOR2_X1 U6577 ( .A1(n5882), .A2(n5881), .ZN(n5888) );
  XNOR2_X1 U6578 ( .A(n5889), .B(n5888), .ZN(n5886) );
  AOI21_X1 U6579 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5908), .A(n3780), 
        .ZN(n5884) );
  NAND2_X1 U6580 ( .A1(n5912), .A2(EAX_REG_29__SCAN_IN), .ZN(n5883) );
  OAI211_X1 U6581 ( .C1(n5886), .C2(n5885), .A(n5884), .B(n5883), .ZN(n5887)
         );
  OAI21_X1 U6582 ( .B1(n5910), .B2(n6393), .A(n5887), .ZN(n5987) );
  NOR2_X1 U6583 ( .A1(n5889), .A2(n5888), .ZN(n5905) );
  AOI22_X1 U6584 ( .A1(n4190), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3621), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5895) );
  AOI22_X1 U6585 ( .A1(n5890), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5894) );
  AOI22_X1 U6586 ( .A1(n5869), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5876), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5893) );
  AOI22_X1 U6587 ( .A1(n4318), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5891), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5892) );
  NAND4_X1 U6588 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n5903)
         );
  AOI22_X1 U6589 ( .A1(n4274), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3738), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5901) );
  AOI22_X1 U6590 ( .A1(n5897), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5896), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5900) );
  AOI22_X1 U6591 ( .A1(n4151), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5870), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5899) );
  AOI22_X1 U6592 ( .A1(n5875), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4191), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5898) );
  NAND4_X1 U6593 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5902)
         );
  NOR2_X1 U6594 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  XNOR2_X1 U6595 ( .A(n5905), .B(n5904), .ZN(n5907) );
  NAND2_X1 U6596 ( .A1(n5907), .A2(n5906), .ZN(n5916) );
  NAND2_X1 U6597 ( .A1(n5908), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5909)
         );
  NAND2_X1 U6598 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  AOI21_X1 U6599 ( .B1(n5912), .B2(EAX_REG_30__SCAN_IN), .A(n5911), .ZN(n5915)
         );
  XNOR2_X1 U6600 ( .A(n5913), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5962)
         );
  AOI21_X1 U6601 ( .B1(n5916), .B2(n5915), .A(n5914), .ZN(n5942) );
  AOI22_X1 U6602 ( .A1(n5912), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n5917), .ZN(n5918) );
  NAND2_X1 U6603 ( .A1(n5919), .A2(n6774), .ZN(n5924) );
  NOR2_X1 U6604 ( .A1(n6778), .A2(n5920), .ZN(n5921) );
  AOI211_X1 U6605 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n6772), .A(n5922), 
        .B(n5921), .ZN(n5923) );
  OAI211_X1 U6606 ( .C1(n6166), .C2(n6748), .A(n5924), .B(n5923), .ZN(U2955)
         );
  XOR2_X1 U6607 ( .A(n4861), .B(n5925), .Z(n5929) );
  OAI222_X1 U6608 ( .A1(n5929), .A2(n5928), .B1(n5927), .B2(n7083), .C1(n4771), 
        .C2(n5926), .ZN(U3463) );
  INV_X1 U6609 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6713) );
  INV_X1 U6610 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6715) );
  NOR2_X1 U6611 ( .A1(n6713), .A2(n6715), .ZN(n5930) );
  OAI21_X1 U6612 ( .B1(n5930), .B2(n6958), .A(n5994), .ZN(n5948) );
  INV_X1 U6613 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5938) );
  INV_X1 U6614 ( .A(n5931), .ZN(n5932) );
  NOR2_X1 U6615 ( .A1(n6004), .A2(n5932), .ZN(n5990) );
  NAND4_X1 U6616 ( .A1(n5990), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n5933), .ZN(n5937) );
  NAND3_X1 U6617 ( .A1(n5935), .A2(EBX_REG_31__SCAN_IN), .A3(n5934), .ZN(n5936) );
  OAI211_X1 U6618 ( .C1(n7050), .C2(n5938), .A(n5937), .B(n5936), .ZN(n5939)
         );
  OAI22_X1 U6619 ( .A1(n5941), .A2(n6148), .B1(n6150), .B2(n5940), .ZN(U2828)
         );
  INV_X1 U6620 ( .A(n5968), .ZN(n5956) );
  OAI21_X1 U6621 ( .B1(n5989), .B2(n5945), .A(n5944), .ZN(n5946) );
  XOR2_X1 U6622 ( .A(n5947), .B(n5946), .Z(n6497) );
  INV_X1 U6623 ( .A(n5948), .ZN(n5952) );
  AOI21_X1 U6624 ( .B1(n5994), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5951) );
  AOI22_X1 U6625 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7035), .B1(n7017), 
        .B2(n5962), .ZN(n5950) );
  NAND2_X1 U6626 ( .A1(n7053), .A2(EBX_REG_30__SCAN_IN), .ZN(n5949) );
  OAI211_X1 U6627 ( .C1(n5952), .C2(n5951), .A(n5950), .B(n5949), .ZN(n5953)
         );
  AOI21_X1 U6628 ( .B1(n6497), .B2(n7056), .A(n5953), .ZN(n5954) );
  OAI21_X1 U6629 ( .B1(n5956), .B2(n7014), .A(n5954), .ZN(U2797) );
  AOI22_X1 U6630 ( .A1(n6497), .A2(n6160), .B1(EBX_REG_30__SCAN_IN), .B2(n6159), .ZN(n5955) );
  OAI21_X1 U6631 ( .B1(n5956), .B2(n6151), .A(n5955), .ZN(U2829) );
  NAND2_X1 U6632 ( .A1(n5958), .A2(n5957), .ZN(n5960) );
  NAND2_X1 U6633 ( .A1(n5960), .A2(n5959), .ZN(n5961) );
  NAND2_X1 U6634 ( .A1(n6477), .A2(n5962), .ZN(n5963) );
  NAND2_X1 U6635 ( .A1(n6906), .A2(REIP_REG_30__SCAN_IN), .ZN(n6495) );
  OAI211_X1 U6636 ( .C1(n6753), .C2(n5964), .A(n5963), .B(n6495), .ZN(n5965)
         );
  AOI21_X1 U6637 ( .B1(n5968), .B2(n6773), .A(n5965), .ZN(n5966) );
  OAI21_X1 U6638 ( .B1(n6499), .B2(n7062), .A(n5966), .ZN(U2956) );
  AND2_X1 U6639 ( .A1(n3679), .A2(n3779), .ZN(n5967) );
  NAND2_X1 U6640 ( .A1(n6163), .A2(n5967), .ZN(n6370) );
  NAND2_X1 U6641 ( .A1(n5968), .A2(n7204), .ZN(n5971) );
  AND2_X1 U6642 ( .A1(n6163), .A2(n5969), .ZN(n7203) );
  AOI22_X1 U6643 ( .A1(n7203), .A2(DATAI_30_), .B1(n7206), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5970) );
  OAI211_X1 U6644 ( .C1(n6370), .C2(n7192), .A(n5971), .B(n5970), .ZN(U2861)
         );
  NAND2_X1 U6645 ( .A1(n5973), .A2(n5972), .ZN(n5977) );
  INV_X1 U6646 ( .A(n5974), .ZN(n5976) );
  AOI22_X1 U6647 ( .A1(n5980), .A2(n5977), .B1(n5976), .B2(n5975), .ZN(n5978)
         );
  OAI21_X1 U6648 ( .B1(n5980), .B2(n5979), .A(n5978), .ZN(n7091) );
  NOR2_X1 U6649 ( .A1(n7144), .A2(n5981), .ZN(n6781) );
  NOR2_X1 U6650 ( .A1(n6781), .A2(n5982), .ZN(n6796) );
  OAI21_X1 U6651 ( .B1(n6796), .B2(READY_N), .A(n5983), .ZN(n7089) );
  AND2_X1 U6652 ( .A1(n7089), .A2(n5984), .ZN(n7063) );
  MUX2_X1 U6653 ( .A(MORE_REG_SCAN_IN), .B(n7091), .S(n7063), .Z(U3471) );
  AOI21_X1 U6654 ( .B1(n5987), .B2(n5986), .A(n5985), .ZN(n6395) );
  INV_X1 U6655 ( .A(n6395), .ZN(n6120) );
  XNOR2_X1 U6656 ( .A(n5989), .B(n5988), .ZN(n6508) );
  AOI22_X1 U6657 ( .A1(n7035), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(n5990), 
        .B2(n6713), .ZN(n5991) );
  OAI21_X1 U6658 ( .B1(n7060), .B2(n6393), .A(n5991), .ZN(n5992) );
  AOI21_X1 U6659 ( .B1(n7053), .B2(EBX_REG_29__SCAN_IN), .A(n5992), .ZN(n5993)
         );
  OAI21_X1 U6660 ( .B1(n6713), .B2(n5994), .A(n5993), .ZN(n5995) );
  AOI21_X1 U6661 ( .B1(n6508), .B2(n7056), .A(n5995), .ZN(n5996) );
  OAI21_X1 U6662 ( .B1(n6120), .B2(n7014), .A(n5996), .ZN(U2798) );
  AND2_X1 U6663 ( .A1(n6012), .A2(n5997), .ZN(n5998) );
  INV_X1 U6664 ( .A(n6404), .ZN(n6122) );
  XNOR2_X1 U6665 ( .A(n3448), .B(n6000), .ZN(n6522) );
  INV_X1 U6666 ( .A(n6001), .ZN(n6003) );
  INV_X1 U6667 ( .A(n6028), .ZN(n6002) );
  OAI21_X1 U6668 ( .B1(n6003), .B2(n6002), .A(n6971), .ZN(n6016) );
  NOR2_X1 U6669 ( .A1(n7060), .A2(n6402), .ZN(n6007) );
  OAI22_X1 U6670 ( .A1(n7050), .A2(n6005), .B1(REIP_REG_27__SCAN_IN), .B2(
        n6004), .ZN(n6006) );
  AOI211_X1 U6671 ( .C1(EBX_REG_27__SCAN_IN), .C2(n7053), .A(n6007), .B(n6006), 
        .ZN(n6008) );
  OAI21_X1 U6672 ( .B1(n6709), .B2(n6016), .A(n6008), .ZN(n6009) );
  AOI21_X1 U6673 ( .B1(n6522), .B2(n7056), .A(n6009), .ZN(n6010) );
  OAI21_X1 U6674 ( .B1(n6122), .B2(n7014), .A(n6010), .ZN(U2800) );
  INV_X1 U6675 ( .A(n6012), .ZN(n6013) );
  AOI21_X1 U6676 ( .B1(n6014), .B2(n6011), .A(n6013), .ZN(n6413) );
  INV_X1 U6677 ( .A(n6413), .ZN(n6123) );
  OAI21_X1 U6678 ( .B1(n6027), .B2(n6015), .A(n3448), .ZN(n6124) );
  INV_X1 U6679 ( .A(n6124), .ZN(n6531) );
  INV_X1 U6680 ( .A(n6016), .ZN(n6017) );
  OAI221_X1 U6681 ( .B1(REIP_REG_26__SCAN_IN), .B2(REIP_REG_25__SCAN_IN), .C1(
        REIP_REG_26__SCAN_IN), .C2(n6030), .A(n6017), .ZN(n6018) );
  OAI21_X1 U6682 ( .B1(n7050), .B2(n6411), .A(n6018), .ZN(n6021) );
  INV_X1 U6683 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6125) );
  INV_X1 U6684 ( .A(n6409), .ZN(n6019) );
  OAI22_X1 U6685 ( .A1(n7025), .A2(n6125), .B1(n6019), .B2(n7060), .ZN(n6020)
         );
  AOI211_X1 U6686 ( .C1(n6531), .C2(n7056), .A(n6021), .B(n6020), .ZN(n6022)
         );
  OAI21_X1 U6687 ( .B1(n6123), .B2(n7014), .A(n6022), .ZN(U2801) );
  OAI21_X1 U6688 ( .B1(n6023), .B2(n6024), .A(n6011), .ZN(n6424) );
  NOR2_X1 U6689 ( .A1(n6040), .A2(n6025), .ZN(n6026) );
  OR2_X1 U6690 ( .A1(n6027), .A2(n6026), .ZN(n6538) );
  INV_X1 U6691 ( .A(n6538), .ZN(n6035) );
  INV_X1 U6692 ( .A(n6971), .ZN(n6029) );
  INV_X1 U6693 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6707) );
  NOR3_X1 U6694 ( .A1(n6029), .A2(n6028), .A3(n6707), .ZN(n6034) );
  INV_X1 U6695 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6126) );
  AOI22_X1 U6696 ( .A1(n7035), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6030), 
        .B2(n6707), .ZN(n6032) );
  NAND2_X1 U6697 ( .A1(n7017), .A2(n6417), .ZN(n6031) );
  OAI211_X1 U6698 ( .C1(n7025), .C2(n6126), .A(n6032), .B(n6031), .ZN(n6033)
         );
  AOI211_X1 U6699 ( .C1(n6035), .C2(n7056), .A(n6034), .B(n6033), .ZN(n6036)
         );
  OAI21_X1 U6700 ( .B1(n6424), .B2(n7014), .A(n6036), .ZN(U2802) );
  NOR2_X1 U6701 ( .A1(n6064), .A2(n6049), .ZN(n6050) );
  NOR2_X1 U6702 ( .A1(n6050), .A2(n6038), .ZN(n6039) );
  OR2_X1 U6703 ( .A1(n6023), .A2(n6039), .ZN(n6434) );
  AOI21_X1 U6704 ( .B1(n6041), .B2(n6059), .A(n6040), .ZN(n6549) );
  NAND2_X1 U6705 ( .A1(n6971), .A2(n6042), .ZN(n6054) );
  AOI22_X1 U6706 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n7035), .B1(
        EBX_REG_24__SCAN_IN), .B2(n7053), .ZN(n6043) );
  OAI221_X1 U6707 ( .B1(REIP_REG_24__SCAN_IN), .B2(n6044), .C1(n6702), .C2(
        n6054), .A(n6043), .ZN(n6047) );
  INV_X1 U6708 ( .A(n6045), .ZN(n6436) );
  NOR2_X1 U6709 ( .A1(n7060), .A2(n6436), .ZN(n6046) );
  AOI211_X1 U6710 ( .C1(n6549), .C2(n7056), .A(n6047), .B(n6046), .ZN(n6048)
         );
  OAI21_X1 U6711 ( .B1(n6434), .B2(n7014), .A(n6048), .ZN(U2803) );
  AND2_X1 U6712 ( .A1(n6064), .A2(n6049), .ZN(n6051) );
  OAI22_X1 U6713 ( .A1(n6052), .A2(n7050), .B1(n7060), .B2(n6443), .ZN(n6057)
         );
  INV_X1 U6714 ( .A(n6053), .ZN(n6055) );
  INV_X1 U6715 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6700) );
  AOI21_X1 U6716 ( .B1(n6055), .B2(n6700), .A(n6054), .ZN(n6056) );
  AOI211_X1 U6717 ( .C1(EBX_REG_23__SCAN_IN), .C2(n7053), .A(n6057), .B(n6056), 
        .ZN(n6062) );
  AOI21_X1 U6718 ( .B1(n6060), .B2(n6058), .A(n4611), .ZN(n6557) );
  NAND2_X1 U6719 ( .A1(n6557), .A2(n7056), .ZN(n6061) );
  OAI211_X1 U6720 ( .C1(n6447), .C2(n7014), .A(n6062), .B(n6061), .ZN(U2804)
         );
  AOI21_X1 U6721 ( .B1(n6065), .B2(n6063), .A(n6037), .ZN(n6454) );
  INV_X1 U6722 ( .A(n6454), .ZN(n6379) );
  OAI21_X1 U6723 ( .B1(n3446), .B2(n6066), .A(n6058), .ZN(n6567) );
  INV_X1 U6724 ( .A(n6567), .ZN(n6075) );
  INV_X1 U6725 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6696) );
  NAND2_X1 U6726 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n7041) );
  NOR2_X1 U6727 ( .A1(n6696), .A2(n7041), .ZN(n6068) );
  NOR2_X1 U6728 ( .A1(n6958), .A2(n6067), .ZN(n7021) );
  NAND3_X1 U6729 ( .A1(n6068), .A2(n7042), .A3(n7049), .ZN(n7047) );
  OAI21_X1 U6730 ( .B1(n6951), .B2(n6069), .A(n6971), .ZN(n7048) );
  AOI21_X1 U6731 ( .B1(n7047), .B2(n7048), .A(n6353), .ZN(n6074) );
  INV_X1 U6732 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6129) );
  INV_X1 U6733 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6452) );
  OAI22_X1 U6734 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6070), .B1(n6452), .B2(
        n7050), .ZN(n6071) );
  AOI21_X1 U6735 ( .B1(n7017), .B2(n6450), .A(n6071), .ZN(n6072) );
  OAI21_X1 U6736 ( .B1(n7025), .B2(n6129), .A(n6072), .ZN(n6073) );
  AOI211_X1 U6737 ( .C1(n6075), .C2(n7056), .A(n6074), .B(n6073), .ZN(n6076)
         );
  OAI21_X1 U6738 ( .B1(n6379), .B2(n7014), .A(n6076), .ZN(U2805) );
  AND2_X1 U6739 ( .A1(n6140), .A2(n6077), .ZN(n6079) );
  OR2_X1 U6740 ( .A1(n6079), .A2(n6078), .ZN(n6467) );
  NAND2_X1 U6741 ( .A1(n6143), .A2(n6080), .ZN(n6081) );
  NAND2_X1 U6742 ( .A1(n6131), .A2(n6081), .ZN(n6586) );
  INV_X1 U6743 ( .A(n6586), .ZN(n6087) );
  INV_X1 U6744 ( .A(n6470), .ZN(n6082) );
  OAI22_X1 U6745 ( .A1(n6466), .A2(n7050), .B1(n7060), .B2(n6082), .ZN(n6086)
         );
  INV_X1 U6746 ( .A(n7041), .ZN(n6083) );
  AOI21_X1 U6747 ( .B1(n6083), .B2(n7042), .A(REIP_REG_20__SCAN_IN), .ZN(n6084) );
  INV_X1 U6748 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6135) );
  OAI22_X1 U6749 ( .A1(n6084), .A2(n7048), .B1(n6135), .B2(n7025), .ZN(n6085)
         );
  AOI211_X1 U6750 ( .C1(n7056), .C2(n6087), .A(n6086), .B(n6085), .ZN(n6088)
         );
  OAI21_X1 U6751 ( .B1(n6467), .B2(n7014), .A(n6088), .ZN(U2807) );
  INV_X1 U6752 ( .A(n6090), .ZN(n6091) );
  AOI21_X1 U6753 ( .B1(n6092), .B2(n6089), .A(n6091), .ZN(n6481) );
  INV_X1 U6754 ( .A(n6481), .ZN(n6384) );
  OAI21_X1 U6755 ( .B1(n6157), .B2(n6094), .A(n6093), .ZN(n6147) );
  INV_X1 U6756 ( .A(n6147), .ZN(n6925) );
  AOI21_X1 U6757 ( .B1(n7017), .B2(n6476), .A(n7034), .ZN(n6095) );
  OAI21_X1 U6758 ( .B1(n7050), .B2(n6479), .A(n6095), .ZN(n6100) );
  INV_X1 U6759 ( .A(n7042), .ZN(n6098) );
  OAI21_X1 U6760 ( .B1(n6958), .B2(n6096), .A(n6948), .ZN(n7036) );
  AOI22_X1 U6761 ( .A1(EBX_REG_18__SCAN_IN), .A2(n7053), .B1(
        REIP_REG_18__SCAN_IN), .B2(n7036), .ZN(n6097) );
  OAI21_X1 U6762 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6098), .A(n6097), .ZN(n6099) );
  AOI211_X1 U6763 ( .C1(n6925), .C2(n7056), .A(n6100), .B(n6099), .ZN(n6101)
         );
  OAI21_X1 U6764 ( .B1(n6384), .B2(n7014), .A(n6101), .ZN(U2809) );
  AOI21_X1 U6765 ( .B1(n6103), .B2(n5803), .A(n6102), .ZN(n6491) );
  INV_X1 U6766 ( .A(n6491), .ZN(n6388) );
  INV_X1 U6767 ( .A(n6155), .ZN(n6104) );
  AOI21_X1 U6768 ( .B1(n6106), .B2(n6105), .A(n6104), .ZN(n6904) );
  NAND2_X1 U6769 ( .A1(n7035), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6107)
         );
  OAI211_X1 U6770 ( .C1(n7060), .C2(n6489), .A(n6107), .B(n7023), .ZN(n6117)
         );
  INV_X1 U6771 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U6772 ( .A1(n6108), .A2(n6688), .ZN(n6109) );
  NOR2_X1 U6773 ( .A1(n6958), .A2(n6109), .ZN(n7010) );
  OAI21_X1 U6774 ( .B1(n7010), .B2(n7011), .A(REIP_REG_16__SCAN_IN), .ZN(n6114) );
  INV_X1 U6775 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6111) );
  NAND3_X1 U6776 ( .A1(n6112), .A2(n6111), .A3(n6110), .ZN(n6113) );
  OAI211_X1 U6777 ( .C1(n7025), .C2(n6115), .A(n6114), .B(n6113), .ZN(n6116)
         );
  AOI211_X1 U6778 ( .C1(n6904), .C2(n7056), .A(n6117), .B(n6116), .ZN(n6118)
         );
  OAI21_X1 U6779 ( .B1(n6388), .B2(n7014), .A(n6118), .ZN(U2811) );
  AOI22_X1 U6780 ( .A1(n6508), .A2(n6160), .B1(n6159), .B2(EBX_REG_29__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U6781 ( .B1(n6120), .B2(n6151), .A(n6119), .ZN(U2830) );
  AOI22_X1 U6782 ( .A1(n6522), .A2(n6160), .B1(EBX_REG_27__SCAN_IN), .B2(n6159), .ZN(n6121) );
  OAI21_X1 U6783 ( .B1(n6122), .B2(n6151), .A(n6121), .ZN(U2832) );
  OAI222_X1 U6784 ( .A1(n6125), .A2(n6150), .B1(n6148), .B2(n6124), .C1(n6123), 
        .C2(n6151), .ZN(U2833) );
  OAI222_X1 U6785 ( .A1(n6538), .A2(n6148), .B1(n6126), .B2(n6150), .C1(n6424), 
        .C2(n6151), .ZN(U2834) );
  AOI22_X1 U6786 ( .A1(n6549), .A2(n6160), .B1(EBX_REG_24__SCAN_IN), .B2(n6159), .ZN(n6127) );
  OAI21_X1 U6787 ( .B1(n6434), .B2(n6151), .A(n6127), .ZN(U2835) );
  AOI22_X1 U6788 ( .A1(n6557), .A2(n6160), .B1(n6159), .B2(EBX_REG_23__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U6789 ( .B1(n6447), .B2(n6151), .A(n6128), .ZN(U2836) );
  OAI222_X1 U6790 ( .A1(n6129), .A2(n6150), .B1(n6148), .B2(n6567), .C1(n6379), 
        .C2(n6151), .ZN(U2837) );
  OAI21_X1 U6791 ( .B1(n6078), .B2(n6130), .A(n6063), .ZN(n7054) );
  AOI21_X1 U6792 ( .B1(n6132), .B2(n6131), .A(n3446), .ZN(n7055) );
  INV_X1 U6793 ( .A(n7055), .ZN(n6133) );
  OAI222_X1 U6794 ( .A1(n7054), .A2(n6151), .B1(n6150), .B2(n6134), .C1(n6133), 
        .C2(n6148), .ZN(U2838) );
  OAI22_X1 U6795 ( .A1(n6586), .A2(n6148), .B1(n6135), .B2(n6150), .ZN(n6136)
         );
  INV_X1 U6796 ( .A(n6136), .ZN(n6137) );
  OAI21_X1 U6797 ( .B1(n6467), .B2(n6151), .A(n6137), .ZN(U2839) );
  NAND2_X1 U6798 ( .A1(n6090), .A2(n6138), .ZN(n6139) );
  AND2_X1 U6799 ( .A1(n6140), .A2(n6139), .ZN(n7200) );
  INV_X1 U6800 ( .A(n7200), .ZN(n6146) );
  NAND2_X1 U6801 ( .A1(n6093), .A2(n6141), .ZN(n6142) );
  AND2_X1 U6802 ( .A1(n6143), .A2(n6142), .ZN(n7037) );
  INV_X1 U6803 ( .A(n7037), .ZN(n6144) );
  OAI222_X1 U6804 ( .A1(n6146), .A2(n6151), .B1(n6150), .B2(n6145), .C1(n6148), 
        .C2(n6144), .ZN(U2840) );
  OAI222_X1 U6805 ( .A1(n6384), .A2(n6151), .B1(n6150), .B2(n6149), .C1(n6148), 
        .C2(n6147), .ZN(U2841) );
  OR2_X1 U6806 ( .A1(n6102), .A2(n6152), .ZN(n6153) );
  AND2_X1 U6807 ( .A1(n6089), .A2(n6153), .ZN(n7197) );
  INV_X1 U6808 ( .A(n7197), .ZN(n7029) );
  AND2_X1 U6809 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  NOR2_X1 U6810 ( .A1(n6157), .A2(n6156), .ZN(n7026) );
  AOI22_X1 U6811 ( .A1(n7026), .A2(n6160), .B1(n6159), .B2(EBX_REG_17__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U6812 ( .B1(n7029), .B2(n6151), .A(n6158), .ZN(U2842) );
  AOI22_X1 U6813 ( .A1(n6904), .A2(n6160), .B1(EBX_REG_16__SCAN_IN), .B2(n6159), .ZN(n6161) );
  OAI21_X1 U6814 ( .B1(n6388), .B2(n6151), .A(n6161), .ZN(U2843) );
  NAND2_X1 U6815 ( .A1(n6163), .A2(n6162), .ZN(n6165) );
  AOI22_X1 U6816 ( .A1(n7203), .A2(DATAI_31_), .B1(n7206), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n6164) );
  OAI21_X1 U6817 ( .B1(n6166), .B2(n6165), .A(n6164), .ZN(U2860) );
  NAND2_X1 U6818 ( .A1(n6395), .A2(n7204), .ZN(n6168) );
  AOI22_X1 U6819 ( .A1(n7203), .A2(DATAI_29_), .B1(n7206), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6167) );
  OAI211_X1 U6820 ( .C1(n6370), .C2(n7188), .A(n6168), .B(n6167), .ZN(U2862)
         );
  AOI22_X1 U6821 ( .A1(n7203), .A2(DATAI_28_), .B1(n7206), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U6822 ( .A1(n7207), .A2(DATAI_12_), .ZN(n6169) );
  OAI211_X1 U6823 ( .C1(n5845), .C2(n6387), .A(n6170), .B(n6169), .ZN(n6365)
         );
  INV_X1 U6824 ( .A(keyinput_63), .ZN(n6263) );
  INV_X1 U6825 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U6826 ( .A1(n6694), .A2(keyinput_63), .B1(n6696), .B2(keyinput_62), 
        .ZN(n6171) );
  OAI21_X1 U6827 ( .B1(n6696), .B2(keyinput_62), .A(n6171), .ZN(n6262) );
  AOI22_X1 U6828 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_59), .B1(n6353), 
        .B2(keyinput_60), .ZN(n6172) );
  OAI221_X1 U6829 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_59), .C1(n6353), 
        .C2(keyinput_60), .A(n6172), .ZN(n6259) );
  INV_X1 U6830 ( .A(keyinput_58), .ZN(n6257) );
  INV_X1 U6831 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6338) );
  INV_X1 U6832 ( .A(keyinput_49), .ZN(n6245) );
  INV_X1 U6833 ( .A(keyinput_48), .ZN(n6243) );
  INV_X1 U6834 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6334) );
  OAI22_X1 U6835 ( .A1(n4906), .A2(keyinput_45), .B1(W_R_N_REG_SCAN_IN), .B2(
        keyinput_46), .ZN(n6173) );
  AOI221_X1 U6836 ( .B1(n4906), .B2(keyinput_45), .C1(keyinput_46), .C2(
        W_R_N_REG_SCAN_IN), .A(n6173), .ZN(n6240) );
  INV_X1 U6837 ( .A(MORE_REG_SCAN_IN), .ZN(n7090) );
  INV_X1 U6838 ( .A(keyinput_44), .ZN(n6238) );
  INV_X1 U6839 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7131) );
  INV_X1 U6840 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6784) );
  XOR2_X1 U6841 ( .A(n6784), .B(keyinput_37), .Z(n6231) );
  INV_X1 U6842 ( .A(keyinput_36), .ZN(n6226) );
  INV_X1 U6843 ( .A(HOLD), .ZN(n6788) );
  INV_X1 U6844 ( .A(keyinput_35), .ZN(n6224) );
  INV_X1 U6845 ( .A(BS16_N), .ZN(n6629) );
  INV_X1 U6846 ( .A(keyinput_34), .ZN(n6222) );
  INV_X1 U6847 ( .A(NA_N), .ZN(n7134) );
  OAI22_X1 U6848 ( .A1(n6175), .A2(keyinput_32), .B1(DATAI_1_), .B2(
        keyinput_30), .ZN(n6174) );
  AOI221_X1 U6849 ( .B1(n6175), .B2(keyinput_32), .C1(keyinput_30), .C2(
        DATAI_1_), .A(n6174), .ZN(n6178) );
  OAI22_X1 U6850 ( .A1(n7157), .A2(keyinput_28), .B1(DATAI_0_), .B2(
        keyinput_31), .ZN(n6176) );
  AOI221_X1 U6851 ( .B1(n7157), .B2(keyinput_28), .C1(keyinput_31), .C2(
        DATAI_0_), .A(n6176), .ZN(n6177) );
  OAI211_X1 U6852 ( .C1(DATAI_2_), .C2(keyinput_29), .A(n6178), .B(n6177), 
        .ZN(n6179) );
  AOI21_X1 U6853 ( .B1(DATAI_2_), .B2(keyinput_29), .A(n6179), .ZN(n6219) );
  INV_X1 U6854 ( .A(keyinput_24), .ZN(n6213) );
  INV_X1 U6855 ( .A(keyinput_23), .ZN(n6211) );
  OAI22_X1 U6856 ( .A1(n7184), .A2(keyinput_19), .B1(DATAI_13_), .B2(
        keyinput_18), .ZN(n6180) );
  AOI221_X1 U6857 ( .B1(n7184), .B2(keyinput_19), .C1(keyinput_18), .C2(
        DATAI_13_), .A(n6180), .ZN(n6209) );
  INV_X1 U6858 ( .A(keyinput_17), .ZN(n6204) );
  OAI22_X1 U6859 ( .A1(n5001), .A2(keyinput_10), .B1(n4996), .B2(keyinput_9), 
        .ZN(n6181) );
  AOI221_X1 U6860 ( .B1(n5001), .B2(keyinput_10), .C1(keyinput_9), .C2(n4996), 
        .A(n6181), .ZN(n6202) );
  OAI22_X1 U6861 ( .A1(n4871), .A2(keyinput_13), .B1(n4881), .B2(keyinput_14), 
        .ZN(n6182) );
  AOI221_X1 U6862 ( .B1(n4871), .B2(keyinput_13), .C1(keyinput_14), .C2(n4881), 
        .A(n6182), .ZN(n6201) );
  OAI22_X1 U6863 ( .A1(DATAI_20_), .A2(keyinput_11), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n6183) );
  AOI221_X1 U6864 ( .B1(DATAI_20_), .B2(keyinput_11), .C1(keyinput_16), .C2(
        DATAI_15_), .A(n6183), .ZN(n6200) );
  INV_X1 U6865 ( .A(keyinput_7), .ZN(n6194) );
  XOR2_X1 U6866 ( .A(DATAI_29_), .B(keyinput_2), .Z(n6192) );
  AOI22_X1 U6867 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_31_), .B2(
        keyinput_0), .ZN(n6184) );
  OAI221_X1 U6868 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n6184), .ZN(n6191) );
  AOI22_X1 U6869 ( .A1(n6186), .A2(keyinput_6), .B1(keyinput_4), .B2(n6277), 
        .ZN(n6185) );
  OAI221_X1 U6870 ( .B1(n6186), .B2(keyinput_6), .C1(n6277), .C2(keyinput_4), 
        .A(n6185), .ZN(n6190) );
  AOI22_X1 U6871 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(n6188), .B2(keyinput_3), .ZN(n6187) );
  OAI221_X1 U6872 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(n6188), .C2(
        keyinput_3), .A(n6187), .ZN(n6189) );
  AOI211_X1 U6873 ( .C1(n6192), .C2(n6191), .A(n6190), .B(n6189), .ZN(n6193)
         );
  AOI221_X1 U6874 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n6284), .C2(n6194), 
        .A(n6193), .ZN(n6198) );
  OAI22_X1 U6875 ( .A1(n4876), .A2(keyinput_12), .B1(n4886), .B2(keyinput_8), 
        .ZN(n6195) );
  AOI221_X1 U6876 ( .B1(n4876), .B2(keyinput_12), .C1(keyinput_8), .C2(n4886), 
        .A(n6195), .ZN(n6196) );
  OAI21_X1 U6877 ( .B1(n5013), .B2(keyinput_15), .A(n6196), .ZN(n6197) );
  AOI211_X1 U6878 ( .C1(n5013), .C2(keyinput_15), .A(n6198), .B(n6197), .ZN(
        n6199) );
  NAND4_X1 U6879 ( .A1(n6202), .A2(n6201), .A3(n6200), .A4(n6199), .ZN(n6203)
         );
  OAI221_X1 U6880 ( .B1(DATAI_14_), .B2(n6204), .C1(n7192), .C2(keyinput_17), 
        .A(n6203), .ZN(n6208) );
  XNOR2_X1 U6881 ( .A(n7175), .B(keyinput_22), .ZN(n6207) );
  AOI22_X1 U6882 ( .A1(keyinput_20), .A2(DATAI_11_), .B1(n7178), .B2(
        keyinput_21), .ZN(n6205) );
  OAI221_X1 U6883 ( .B1(keyinput_20), .B2(DATAI_11_), .C1(n7178), .C2(
        keyinput_21), .A(n6205), .ZN(n6206) );
  AOI211_X1 U6884 ( .C1(n6209), .C2(n6208), .A(n6207), .B(n6206), .ZN(n6210)
         );
  AOI221_X1 U6885 ( .B1(DATAI_8_), .B2(n6211), .C1(n7172), .C2(keyinput_23), 
        .A(n6210), .ZN(n6212) );
  AOI221_X1 U6886 ( .B1(DATAI_7_), .B2(keyinput_24), .C1(n7169), .C2(n6213), 
        .A(n6212), .ZN(n6216) );
  AOI22_X1 U6887 ( .A1(DATAI_5_), .A2(keyinput_26), .B1(n7166), .B2(
        keyinput_25), .ZN(n6214) );
  OAI221_X1 U6888 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(n7166), .C2(
        keyinput_25), .A(n6214), .ZN(n6215) );
  AOI211_X1 U6889 ( .C1(n7160), .C2(keyinput_27), .A(n6216), .B(n6215), .ZN(
        n6217) );
  OAI21_X1 U6890 ( .B1(n7160), .B2(keyinput_27), .A(n6217), .ZN(n6218) );
  AOI22_X1 U6891 ( .A1(keyinput_33), .A2(n7134), .B1(n6219), .B2(n6218), .ZN(
        n6220) );
  OAI21_X1 U6892 ( .B1(n7134), .B2(keyinput_33), .A(n6220), .ZN(n6221) );
  OAI221_X1 U6893 ( .B1(BS16_N), .B2(keyinput_34), .C1(n6629), .C2(n6222), .A(
        n6221), .ZN(n6223) );
  OAI221_X1 U6894 ( .B1(READY_N), .B2(keyinput_35), .C1(n7143), .C2(n6224), 
        .A(n6223), .ZN(n6225) );
  OAI221_X1 U6895 ( .B1(HOLD), .B2(n6226), .C1(n6788), .C2(keyinput_36), .A(
        n6225), .ZN(n6230) );
  INV_X1 U6896 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U6897 ( .A(n6633), .B(keyinput_38), .ZN(n6229) );
  AOI22_X1 U6898 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_40), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .ZN(n6227) );
  OAI221_X1 U6899 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_40), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(keyinput_39), .A(n6227), .ZN(n6228) );
  AOI211_X1 U6900 ( .C1(n6231), .C2(n6230), .A(n6229), .B(n6228), .ZN(n6235)
         );
  INV_X1 U6901 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6233) );
  AOI22_X1 U6902 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_43), .B1(n6233), 
        .B2(keyinput_41), .ZN(n6232) );
  OAI221_X1 U6903 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_43), .C1(n6233), 
        .C2(keyinput_41), .A(n6232), .ZN(n6234) );
  AOI211_X1 U6904 ( .C1(n7131), .C2(keyinput_42), .A(n6235), .B(n6234), .ZN(
        n6236) );
  OAI21_X1 U6905 ( .B1(n7131), .B2(keyinput_42), .A(n6236), .ZN(n6237) );
  OAI221_X1 U6906 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_44), .C1(n7090), .C2(
        n6238), .A(n6237), .ZN(n6239) );
  OAI211_X1 U6907 ( .C1(BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_47), .A(n6240), .B(n6239), .ZN(n6241) );
  AOI21_X1 U6908 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_47), .A(n6241), 
        .ZN(n6242) );
  AOI221_X1 U6909 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6243), .C1(n6334), 
        .C2(keyinput_48), .A(n6242), .ZN(n6244) );
  AOI221_X1 U6910 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .C1(
        n6338), .C2(n6245), .A(n6244), .ZN(n6248) );
  AOI22_X1 U6911 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_50), .B1(n5933), .B2(keyinput_51), .ZN(n6246) );
  OAI221_X1 U6912 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_50), .C1(
        n5933), .C2(keyinput_51), .A(n6246), .ZN(n6247) );
  OAI22_X1 U6913 ( .A1(n6248), .A2(n6247), .B1(keyinput_52), .B2(n6715), .ZN(
        n6251) );
  INV_X1 U6914 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6711) );
  OAI22_X1 U6915 ( .A1(n6711), .A2(keyinput_54), .B1(REIP_REG_29__SCAN_IN), 
        .B2(keyinput_53), .ZN(n6249) );
  AOI221_X1 U6916 ( .B1(n6711), .B2(keyinput_54), .C1(keyinput_53), .C2(
        REIP_REG_29__SCAN_IN), .A(n6249), .ZN(n6250) );
  OAI221_X1 U6917 ( .B1(n6251), .B2(keyinput_52), .C1(n6251), .C2(n6715), .A(
        n6250), .ZN(n6254) );
  INV_X1 U6918 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6346) );
  AOI22_X1 U6919 ( .A1(n6346), .A2(keyinput_56), .B1(n6709), .B2(keyinput_55), 
        .ZN(n6252) );
  OAI221_X1 U6920 ( .B1(n6346), .B2(keyinput_56), .C1(n6709), .C2(keyinput_55), 
        .A(n6252), .ZN(n6253) );
  OAI22_X1 U6921 ( .A1(n6254), .A2(n6253), .B1(keyinput_57), .B2(
        REIP_REG_25__SCAN_IN), .ZN(n6255) );
  AOI21_X1 U6922 ( .B1(keyinput_57), .B2(REIP_REG_25__SCAN_IN), .A(n6255), 
        .ZN(n6256) );
  AOI221_X1 U6923 ( .B1(REIP_REG_24__SCAN_IN), .B2(n6257), .C1(n6702), .C2(
        keyinput_58), .A(n6256), .ZN(n6258) );
  OAI22_X1 U6924 ( .A1(keyinput_61), .A2(n7049), .B1(n6259), .B2(n6258), .ZN(
        n6260) );
  AOI21_X1 U6925 ( .B1(keyinput_61), .B2(n7049), .A(n6260), .ZN(n6261) );
  AOI211_X1 U6926 ( .C1(REIP_REG_19__SCAN_IN), .C2(n6263), .A(n6262), .B(n6261), .ZN(n6363) );
  INV_X1 U6927 ( .A(keyinput_126), .ZN(n6361) );
  INV_X1 U6928 ( .A(keyinput_122), .ZN(n6351) );
  INV_X1 U6929 ( .A(keyinput_113), .ZN(n6337) );
  INV_X1 U6930 ( .A(keyinput_112), .ZN(n6335) );
  OAI22_X1 U6931 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_111), .B1(
        keyinput_110), .B2(W_R_N_REG_SCAN_IN), .ZN(n6264) );
  AOI221_X1 U6932 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_111), .C1(
        W_R_N_REG_SCAN_IN), .C2(keyinput_110), .A(n6264), .ZN(n6331) );
  INV_X1 U6933 ( .A(keyinput_108), .ZN(n6329) );
  XNOR2_X1 U6934 ( .A(n6784), .B(keyinput_101), .ZN(n6323) );
  INV_X1 U6935 ( .A(keyinput_100), .ZN(n6317) );
  INV_X1 U6936 ( .A(keyinput_99), .ZN(n6315) );
  INV_X1 U6937 ( .A(keyinput_98), .ZN(n6313) );
  OAI22_X1 U6938 ( .A1(n7148), .A2(keyinput_95), .B1(DATAI_3_), .B2(
        keyinput_92), .ZN(n6265) );
  AOI221_X1 U6939 ( .B1(n7148), .B2(keyinput_95), .C1(keyinput_92), .C2(
        DATAI_3_), .A(n6265), .ZN(n6268) );
  OAI22_X1 U6940 ( .A1(n7151), .A2(keyinput_94), .B1(keyinput_93), .B2(
        DATAI_2_), .ZN(n6266) );
  AOI221_X1 U6941 ( .B1(n7151), .B2(keyinput_94), .C1(DATAI_2_), .C2(
        keyinput_93), .A(n6266), .ZN(n6267) );
  OAI211_X1 U6942 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_96), .A(n6268), 
        .B(n6267), .ZN(n6269) );
  AOI21_X1 U6943 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_96), .A(n6269), 
        .ZN(n6310) );
  INV_X1 U6944 ( .A(keyinput_88), .ZN(n6304) );
  INV_X1 U6945 ( .A(keyinput_87), .ZN(n6302) );
  OAI22_X1 U6946 ( .A1(n7184), .A2(keyinput_83), .B1(DATAI_13_), .B2(
        keyinput_82), .ZN(n6270) );
  AOI221_X1 U6947 ( .B1(n7184), .B2(keyinput_83), .C1(keyinput_82), .C2(
        DATAI_13_), .A(n6270), .ZN(n6300) );
  INV_X1 U6948 ( .A(keyinput_81), .ZN(n6295) );
  OAI22_X1 U6949 ( .A1(n4996), .A2(keyinput_73), .B1(n4876), .B2(keyinput_76), 
        .ZN(n6271) );
  AOI221_X1 U6950 ( .B1(n4996), .B2(keyinput_73), .C1(keyinput_76), .C2(n4876), 
        .A(n6271), .ZN(n6293) );
  OAI22_X1 U6951 ( .A1(n4886), .A2(keyinput_72), .B1(keyinput_74), .B2(
        DATAI_21_), .ZN(n6272) );
  AOI221_X1 U6952 ( .B1(n4886), .B2(keyinput_72), .C1(DATAI_21_), .C2(
        keyinput_74), .A(n6272), .ZN(n6292) );
  OAI22_X1 U6953 ( .A1(n5006), .A2(keyinput_75), .B1(keyinput_80), .B2(
        DATAI_15_), .ZN(n6273) );
  AOI221_X1 U6954 ( .B1(n5006), .B2(keyinput_75), .C1(DATAI_15_), .C2(
        keyinput_80), .A(n6273), .ZN(n6291) );
  INV_X1 U6955 ( .A(keyinput_71), .ZN(n6285) );
  XNOR2_X1 U6956 ( .A(DATAI_29_), .B(keyinput_66), .ZN(n6282) );
  AOI22_X1 U6957 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n6274) );
  OAI221_X1 U6958 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n6274), .ZN(n6281) );
  AOI22_X1 U6959 ( .A1(n6277), .A2(keyinput_68), .B1(n6276), .B2(keyinput_69), 
        .ZN(n6275) );
  OAI221_X1 U6960 ( .B1(n6277), .B2(keyinput_68), .C1(n6276), .C2(keyinput_69), 
        .A(n6275), .ZN(n6280) );
  AOI22_X1 U6961 ( .A1(DATAI_25_), .A2(keyinput_70), .B1(DATAI_28_), .B2(
        keyinput_67), .ZN(n6278) );
  OAI221_X1 U6962 ( .B1(DATAI_25_), .B2(keyinput_70), .C1(DATAI_28_), .C2(
        keyinput_67), .A(n6278), .ZN(n6279) );
  AOI211_X1 U6963 ( .C1(n6282), .C2(n6281), .A(n6280), .B(n6279), .ZN(n6283)
         );
  AOI221_X1 U6964 ( .B1(DATAI_24_), .B2(n6285), .C1(n6284), .C2(keyinput_71), 
        .A(n6283), .ZN(n6289) );
  OAI22_X1 U6965 ( .A1(n4871), .A2(keyinput_77), .B1(keyinput_78), .B2(
        DATAI_17_), .ZN(n6286) );
  AOI221_X1 U6966 ( .B1(n4871), .B2(keyinput_77), .C1(DATAI_17_), .C2(
        keyinput_78), .A(n6286), .ZN(n6287) );
  OAI21_X1 U6967 ( .B1(DATAI_16_), .B2(keyinput_79), .A(n6287), .ZN(n6288) );
  AOI211_X1 U6968 ( .C1(DATAI_16_), .C2(keyinput_79), .A(n6289), .B(n6288), 
        .ZN(n6290) );
  NAND4_X1 U6969 ( .A1(n6293), .A2(n6292), .A3(n6291), .A4(n6290), .ZN(n6294)
         );
  OAI221_X1 U6970 ( .B1(DATAI_14_), .B2(n6295), .C1(n7192), .C2(keyinput_81), 
        .A(n6294), .ZN(n6299) );
  XNOR2_X1 U6971 ( .A(n7175), .B(keyinput_86), .ZN(n6298) );
  AOI22_X1 U6972 ( .A1(DATAI_10_), .A2(keyinput_85), .B1(n7181), .B2(
        keyinput_84), .ZN(n6296) );
  OAI221_X1 U6973 ( .B1(DATAI_10_), .B2(keyinput_85), .C1(n7181), .C2(
        keyinput_84), .A(n6296), .ZN(n6297) );
  AOI211_X1 U6974 ( .C1(n6300), .C2(n6299), .A(n6298), .B(n6297), .ZN(n6301)
         );
  AOI221_X1 U6975 ( .B1(DATAI_8_), .B2(n6302), .C1(n7172), .C2(keyinput_87), 
        .A(n6301), .ZN(n6303) );
  AOI221_X1 U6976 ( .B1(DATAI_7_), .B2(n6304), .C1(n7169), .C2(keyinput_88), 
        .A(n6303), .ZN(n6307) );
  AOI22_X1 U6977 ( .A1(DATAI_4_), .A2(keyinput_91), .B1(n7166), .B2(
        keyinput_89), .ZN(n6305) );
  OAI221_X1 U6978 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(n7166), .C2(
        keyinput_89), .A(n6305), .ZN(n6306) );
  AOI211_X1 U6979 ( .C1(n7163), .C2(keyinput_90), .A(n6307), .B(n6306), .ZN(
        n6308) );
  OAI21_X1 U6980 ( .B1(n7163), .B2(keyinput_90), .A(n6308), .ZN(n6309) );
  AOI22_X1 U6981 ( .A1(n6310), .A2(n6309), .B1(keyinput_97), .B2(NA_N), .ZN(
        n6311) );
  OAI21_X1 U6982 ( .B1(keyinput_97), .B2(NA_N), .A(n6311), .ZN(n6312) );
  OAI221_X1 U6983 ( .B1(BS16_N), .B2(n6313), .C1(n6629), .C2(keyinput_98), .A(
        n6312), .ZN(n6314) );
  OAI221_X1 U6984 ( .B1(READY_N), .B2(n6315), .C1(n7143), .C2(keyinput_99), 
        .A(n6314), .ZN(n6316) );
  OAI221_X1 U6985 ( .B1(HOLD), .B2(n6317), .C1(n6788), .C2(keyinput_100), .A(
        n6316), .ZN(n6322) );
  XOR2_X1 U6986 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_104), .Z(n6321) );
  AOI22_X1 U6987 ( .A1(n6319), .A2(keyinput_103), .B1(keyinput_102), .B2(n6633), .ZN(n6318) );
  OAI221_X1 U6988 ( .B1(n6319), .B2(keyinput_103), .C1(n6633), .C2(
        keyinput_102), .A(n6318), .ZN(n6320) );
  AOI211_X1 U6989 ( .C1(n6323), .C2(n6322), .A(n6321), .B(n6320), .ZN(n6326)
         );
  AOI22_X1 U6990 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput_105), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_106), .ZN(n6324) );
  OAI221_X1 U6991 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput_105), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_106), .A(n6324), .ZN(n6325)
         );
  AOI211_X1 U6992 ( .C1(STATEBS16_REG_SCAN_IN), .C2(keyinput_107), .A(n6326), 
        .B(n6325), .ZN(n6327) );
  OAI21_X1 U6993 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_107), .A(n6327), 
        .ZN(n6328) );
  OAI221_X1 U6994 ( .B1(MORE_REG_SCAN_IN), .B2(n6329), .C1(n7090), .C2(
        keyinput_108), .A(n6328), .ZN(n6330) );
  OAI211_X1 U6995 ( .C1(FLUSH_REG_SCAN_IN), .C2(keyinput_109), .A(n6331), .B(
        n6330), .ZN(n6332) );
  AOI21_X1 U6996 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .A(n6332), .ZN(
        n6333) );
  AOI221_X1 U6997 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6335), .C1(n6334), 
        .C2(keyinput_112), .A(n6333), .ZN(n6336) );
  AOI221_X1 U6998 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_113), .C1(
        n6338), .C2(n6337), .A(n6336), .ZN(n6341) );
  AOI22_X1 U6999 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_114), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_115), .ZN(n6339) );
  OAI221_X1 U7000 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_114), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_115), .A(n6339), .ZN(n6340) );
  OAI22_X1 U7001 ( .A1(n6341), .A2(n6340), .B1(keyinput_116), .B2(n6715), .ZN(
        n6344) );
  OAI22_X1 U7002 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_117), .B1(
        REIP_REG_27__SCAN_IN), .B2(keyinput_119), .ZN(n6342) );
  AOI221_X1 U7003 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_117), .C1(
        keyinput_119), .C2(REIP_REG_27__SCAN_IN), .A(n6342), .ZN(n6343) );
  OAI221_X1 U7004 ( .B1(n6344), .B2(keyinput_116), .C1(n6344), .C2(n6715), .A(
        n6343), .ZN(n6348) );
  AOI22_X1 U7005 ( .A1(n6346), .A2(keyinput_120), .B1(n6711), .B2(keyinput_118), .ZN(n6345) );
  OAI221_X1 U7006 ( .B1(n6346), .B2(keyinput_120), .C1(n6711), .C2(
        keyinput_118), .A(n6345), .ZN(n6347) );
  OAI22_X1 U7007 ( .A1(keyinput_121), .A2(n6707), .B1(n6348), .B2(n6347), .ZN(
        n6349) );
  AOI21_X1 U7008 ( .B1(keyinput_121), .B2(n6707), .A(n6349), .ZN(n6350) );
  AOI221_X1 U7009 ( .B1(REIP_REG_24__SCAN_IN), .B2(n6351), .C1(n6702), .C2(
        keyinput_122), .A(n6350), .ZN(n6355) );
  AOI22_X1 U7010 ( .A1(n6353), .A2(keyinput_124), .B1(keyinput_123), .B2(n6700), .ZN(n6352) );
  OAI221_X1 U7011 ( .B1(n6353), .B2(keyinput_124), .C1(n6700), .C2(
        keyinput_123), .A(n6352), .ZN(n6354) );
  OR2_X1 U7012 ( .A1(n6355), .A2(n6354), .ZN(n6357) );
  NAND2_X1 U7013 ( .A1(n7049), .A2(keyinput_125), .ZN(n6356) );
  OAI211_X1 U7014 ( .C1(keyinput_125), .C2(n7049), .A(n6357), .B(n6356), .ZN(
        n6360) );
  OAI22_X1 U7015 ( .A1(n6696), .A2(keyinput_126), .B1(keyinput_127), .B2(
        REIP_REG_19__SCAN_IN), .ZN(n6358) );
  AOI21_X1 U7016 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput_127), .A(n6358), 
        .ZN(n6359) );
  OAI211_X1 U7017 ( .C1(REIP_REG_20__SCAN_IN), .C2(n6361), .A(n6360), .B(n6359), .ZN(n6362) );
  NAND2_X1 U7018 ( .A1(n6363), .A2(n6362), .ZN(n6364) );
  XNOR2_X1 U7019 ( .A(n6365), .B(n6364), .ZN(U2863) );
  NAND2_X1 U7020 ( .A1(n6404), .A2(n7204), .ZN(n6367) );
  AOI22_X1 U7021 ( .A1(n7203), .A2(DATAI_27_), .B1(n7206), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6366) );
  OAI211_X1 U7022 ( .C1(n6370), .C2(n7181), .A(n6367), .B(n6366), .ZN(U2864)
         );
  NAND2_X1 U7023 ( .A1(n6413), .A2(n7204), .ZN(n6369) );
  AOI22_X1 U7024 ( .A1(n7203), .A2(DATAI_26_), .B1(n7206), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6368) );
  OAI211_X1 U7025 ( .C1(n6370), .C2(n7178), .A(n6369), .B(n6368), .ZN(U2865)
         );
  AOI22_X1 U7026 ( .A1(n7203), .A2(DATAI_25_), .B1(n7206), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7027 ( .A1(n7207), .A2(DATAI_9_), .ZN(n6371) );
  OAI211_X1 U7028 ( .C1(n6424), .C2(n6387), .A(n6372), .B(n6371), .ZN(U2866)
         );
  AOI22_X1 U7029 ( .A1(n7203), .A2(DATAI_24_), .B1(n7206), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7030 ( .A1(n7207), .A2(DATAI_8_), .ZN(n6373) );
  OAI211_X1 U7031 ( .C1(n6434), .C2(n6387), .A(n6374), .B(n6373), .ZN(U2867)
         );
  AOI22_X1 U7032 ( .A1(n7203), .A2(DATAI_23_), .B1(n7206), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7033 ( .A1(n7207), .A2(DATAI_7_), .ZN(n6375) );
  OAI211_X1 U7034 ( .C1(n6447), .C2(n6387), .A(n6376), .B(n6375), .ZN(U2868)
         );
  AOI22_X1 U7035 ( .A1(n7203), .A2(DATAI_22_), .B1(n7206), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7036 ( .A1(n7207), .A2(DATAI_6_), .ZN(n6377) );
  OAI211_X1 U7037 ( .C1(n6379), .C2(n6387), .A(n6378), .B(n6377), .ZN(U2869)
         );
  AOI22_X1 U7038 ( .A1(n7203), .A2(DATAI_20_), .B1(n7206), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U7039 ( .A1(n7207), .A2(DATAI_4_), .ZN(n6380) );
  OAI211_X1 U7040 ( .C1(n6467), .C2(n6387), .A(n6381), .B(n6380), .ZN(U2871)
         );
  AOI22_X1 U7041 ( .A1(n7203), .A2(DATAI_18_), .B1(n7206), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U7042 ( .A1(n7207), .A2(DATAI_2_), .ZN(n6382) );
  OAI211_X1 U7043 ( .C1(n6384), .C2(n6387), .A(n6383), .B(n6382), .ZN(U2873)
         );
  AOI22_X1 U7044 ( .A1(n7203), .A2(DATAI_16_), .B1(n7206), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7045 ( .A1(n7207), .A2(DATAI_0_), .ZN(n6385) );
  OAI211_X1 U7046 ( .C1(n6388), .C2(n6387), .A(n6386), .B(n6385), .ZN(U2875)
         );
  NOR2_X1 U7047 ( .A1(n6894), .A2(n6713), .ZN(n6500) );
  AOI21_X1 U7048 ( .B1(n6772), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6500), 
        .ZN(n6392) );
  OAI21_X1 U7049 ( .B1(n6393), .B2(n6778), .A(n6392), .ZN(n6394) );
  AOI21_X1 U7050 ( .B1(n6395), .B2(n6773), .A(n6394), .ZN(n6396) );
  OAI21_X1 U7051 ( .B1(n6510), .B2(n7062), .A(n6396), .ZN(U2957) );
  MUX2_X1 U7052 ( .A(n6398), .B(n6397), .S(n6474), .Z(n6400) );
  XNOR2_X1 U7053 ( .A(n6400), .B(n6399), .ZN(n6525) );
  NOR2_X1 U7054 ( .A1(n6894), .A2(n6709), .ZN(n6520) );
  AOI21_X1 U7055 ( .B1(n6772), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6520), 
        .ZN(n6401) );
  OAI21_X1 U7056 ( .B1(n6402), .B2(n6778), .A(n6401), .ZN(n6403) );
  AOI21_X1 U7057 ( .B1(n6404), .B2(n6773), .A(n6403), .ZN(n6405) );
  OAI21_X1 U7058 ( .B1(n7062), .B2(n6525), .A(n6405), .ZN(U2959) );
  OAI21_X1 U7059 ( .B1(n6474), .B2(n6529), .A(n6406), .ZN(n6408) );
  XOR2_X1 U7060 ( .A(n6408), .B(n6407), .Z(n6533) );
  NAND2_X1 U7061 ( .A1(n6477), .A2(n6409), .ZN(n6410) );
  NAND2_X1 U7062 ( .A1(n6906), .A2(REIP_REG_26__SCAN_IN), .ZN(n6528) );
  OAI211_X1 U7063 ( .C1(n6753), .C2(n6411), .A(n6410), .B(n6528), .ZN(n6412)
         );
  AOI21_X1 U7064 ( .B1(n6413), .B2(n6773), .A(n6412), .ZN(n6414) );
  OAI21_X1 U7065 ( .B1(n6533), .B2(n7062), .A(n6414), .ZN(U2960) );
  OAI22_X1 U7066 ( .A1(n6753), .A2(n6415), .B1(n6894), .B2(n6707), .ZN(n6416)
         );
  AOI21_X1 U7067 ( .B1(n6477), .B2(n6417), .A(n6416), .ZN(n6423) );
  NAND2_X1 U7068 ( .A1(n6420), .A2(n6421), .ZN(n6534) );
  NAND3_X1 U7069 ( .A1(n6419), .A2(n6534), .A3(n6774), .ZN(n6422) );
  OAI211_X1 U7070 ( .C1(n6424), .C2(n6748), .A(n6423), .B(n6422), .ZN(U2961)
         );
  XNOR2_X1 U7071 ( .A(n6428), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6593)
         );
  NAND2_X1 U7072 ( .A1(n6594), .A2(n6593), .ZN(n6592) );
  INV_X1 U7073 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6425) );
  NOR2_X1 U7074 ( .A1(n6474), .A2(n6425), .ZN(n6426) );
  INV_X1 U7075 ( .A(n6562), .ZN(n6582) );
  NAND2_X1 U7076 ( .A1(n6474), .A2(n6582), .ZN(n6427) );
  NAND2_X1 U7077 ( .A1(n6429), .A2(n6427), .ZN(n6458) );
  INV_X1 U7078 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6579) );
  XNOR2_X1 U7079 ( .A(n6428), .B(n6579), .ZN(n6457) );
  NOR2_X1 U7080 ( .A1(n6458), .A2(n6457), .ZN(n6456) );
  AOI21_X1 U7081 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3519), .A(n6456), 
        .ZN(n6449) );
  NAND3_X1 U7082 ( .A1(n6463), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7083 ( .A1(n3519), .A2(n6560), .ZN(n6431) );
  INV_X1 U7084 ( .A(n6429), .ZN(n6430) );
  NAND2_X1 U7085 ( .A1(n6430), .A2(n6564), .ZN(n6440) );
  OAI22_X1 U7086 ( .A1(n6449), .A2(n6432), .B1(n6431), .B2(n6440), .ZN(n6433)
         );
  XNOR2_X1 U7087 ( .A(n6433), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6551)
         );
  INV_X1 U7088 ( .A(n6434), .ZN(n6438) );
  NOR2_X1 U7089 ( .A1(n6894), .A2(n6702), .ZN(n6548) );
  AOI21_X1 U7090 ( .B1(n6772), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6548), 
        .ZN(n6435) );
  OAI21_X1 U7091 ( .B1(n6436), .B2(n6778), .A(n6435), .ZN(n6437) );
  AOI21_X1 U7092 ( .B1(n6438), .B2(n6773), .A(n6437), .ZN(n6439) );
  OAI21_X1 U7093 ( .B1(n6551), .B2(n7062), .A(n6439), .ZN(U2962) );
  MUX2_X1 U7094 ( .A(n6441), .B(n6440), .S(n3519), .Z(n6442) );
  XNOR2_X1 U7095 ( .A(n6442), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6553)
         );
  NAND2_X1 U7096 ( .A1(n6553), .A2(n6774), .ZN(n6446) );
  NOR2_X1 U7097 ( .A1(n6894), .A2(n6700), .ZN(n6556) );
  NOR2_X1 U7098 ( .A1(n6778), .A2(n6443), .ZN(n6444) );
  AOI211_X1 U7099 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6556), 
        .B(n6444), .ZN(n6445) );
  OAI211_X1 U7100 ( .C1(n6748), .C2(n6447), .A(n6446), .B(n6445), .ZN(U2963)
         );
  XNOR2_X1 U7101 ( .A(n3519), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6448)
         );
  XNOR2_X1 U7102 ( .A(n6449), .B(n6448), .ZN(n6570) );
  NAND2_X1 U7103 ( .A1(n6477), .A2(n6450), .ZN(n6451) );
  NAND2_X1 U7104 ( .A1(n6906), .A2(REIP_REG_22__SCAN_IN), .ZN(n6566) );
  OAI211_X1 U7105 ( .C1(n6753), .C2(n6452), .A(n6451), .B(n6566), .ZN(n6453)
         );
  AOI21_X1 U7106 ( .B1(n6454), .B2(n6773), .A(n6453), .ZN(n6455) );
  OAI21_X1 U7107 ( .B1(n6570), .B2(n7062), .A(n6455), .ZN(U2964) );
  INV_X1 U7108 ( .A(n6456), .ZN(n6573) );
  NAND2_X1 U7109 ( .A1(n6458), .A2(n6457), .ZN(n6572) );
  NAND3_X1 U7110 ( .A1(n6573), .A2(n6774), .A3(n6572), .ZN(n6462) );
  NAND2_X1 U7111 ( .A1(n6906), .A2(REIP_REG_21__SCAN_IN), .ZN(n6574) );
  INV_X1 U7112 ( .A(n6574), .ZN(n6460) );
  NOR2_X1 U7113 ( .A1(n6778), .A2(n7061), .ZN(n6459) );
  AOI211_X1 U7114 ( .C1(n6772), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n6460), 
        .B(n6459), .ZN(n6461) );
  OAI211_X1 U7115 ( .C1(n6748), .C2(n7054), .A(n6462), .B(n6461), .ZN(U2965)
         );
  NAND2_X1 U7116 ( .A1(n6592), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6464) );
  MUX2_X1 U7117 ( .A(n6592), .B(n6464), .S(n6463), .Z(n6465) );
  XOR2_X1 U7118 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(n6465), .Z(n6591) );
  NAND2_X1 U7119 ( .A1(n6906), .A2(REIP_REG_20__SCAN_IN), .ZN(n6585) );
  OAI21_X1 U7120 ( .B1(n6753), .B2(n6466), .A(n6585), .ZN(n6469) );
  NOR2_X1 U7121 ( .A1(n6467), .A2(n6748), .ZN(n6468) );
  AOI211_X1 U7122 ( .C1(n6477), .C2(n6470), .A(n6469), .B(n6468), .ZN(n6471)
         );
  OAI21_X1 U7123 ( .B1(n6591), .B2(n7062), .A(n6471), .ZN(U2966) );
  NAND2_X1 U7124 ( .A1(n6474), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U7125 ( .A1(n6474), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6603)
         );
  NAND2_X1 U7126 ( .A1(n6473), .A2(n6603), .ZN(n6607) );
  OAI21_X1 U7127 ( .B1(n6472), .B2(n6605), .A(n6607), .ZN(n6475) );
  XNOR2_X1 U7128 ( .A(n6475), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6914)
         );
  NAND2_X1 U7129 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  NAND2_X1 U7130 ( .A1(n6906), .A2(REIP_REG_18__SCAN_IN), .ZN(n6915) );
  OAI211_X1 U7131 ( .C1(n6753), .C2(n6479), .A(n6478), .B(n6915), .ZN(n6480)
         );
  AOI21_X1 U7132 ( .B1(n6481), .B2(n6773), .A(n6480), .ZN(n6482) );
  OAI21_X1 U7133 ( .B1(n6914), .B2(n7062), .A(n6482), .ZN(U2968) );
  INV_X1 U7134 ( .A(n6484), .ZN(n6486) );
  NAND2_X1 U7135 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  XNOR2_X1 U7136 ( .A(n6483), .B(n6487), .ZN(n6903) );
  AOI22_X1 U7137 ( .A1(n6772), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6906), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6488) );
  OAI21_X1 U7138 ( .B1(n6489), .B2(n6778), .A(n6488), .ZN(n6490) );
  AOI21_X1 U7139 ( .B1(n6491), .B2(n6773), .A(n6490), .ZN(n6492) );
  OAI21_X1 U7140 ( .B1(n6903), .B2(n7062), .A(n6492), .ZN(U2970) );
  INV_X1 U7141 ( .A(n6518), .ZN(n6502) );
  NAND3_X1 U7142 ( .A1(n6502), .A2(n6493), .A3(n4494), .ZN(n6494) );
  OAI211_X1 U7143 ( .C1(n6506), .C2(n4494), .A(n6495), .B(n6494), .ZN(n6496)
         );
  AOI21_X1 U7144 ( .B1(n6497), .B2(n6926), .A(n6496), .ZN(n6498) );
  OAI21_X1 U7145 ( .B1(n6499), .B2(n6590), .A(n6498), .ZN(U2988) );
  INV_X1 U7146 ( .A(n6500), .ZN(n6504) );
  NAND3_X1 U7147 ( .A1(n6502), .A2(n6501), .A3(n6505), .ZN(n6503) );
  OAI211_X1 U7148 ( .C1(n6506), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6507)
         );
  AOI21_X1 U7149 ( .B1(n6926), .B2(n6508), .A(n6507), .ZN(n6509) );
  OAI21_X1 U7150 ( .B1(n6510), .B2(n6590), .A(n6509), .ZN(U2989) );
  XNOR2_X1 U7151 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U7152 ( .B1(n6518), .B2(n6512), .A(n6511), .ZN(n6515) );
  NOR2_X1 U7153 ( .A1(n6513), .A2(n6897), .ZN(n6514) );
  AOI211_X1 U7154 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n6521), .A(n6515), .B(n6514), .ZN(n6516) );
  OAI21_X1 U7155 ( .B1(n6517), .B2(n6590), .A(n6516), .ZN(U2990) );
  NOR2_X1 U7156 ( .A1(n6518), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6519)
         );
  AOI211_X1 U7157 ( .C1(n6521), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6520), .B(n6519), .ZN(n6524) );
  NAND2_X1 U7158 ( .A1(n6522), .A2(n6926), .ZN(n6523) );
  OAI211_X1 U7159 ( .C1(n6525), .C2(n6590), .A(n6524), .B(n6523), .ZN(U2991)
         );
  XNOR2_X1 U7160 ( .A(n6529), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6526)
         );
  NAND2_X1 U7161 ( .A1(n6535), .A2(n6526), .ZN(n6527) );
  OAI211_X1 U7162 ( .C1(n6544), .C2(n6529), .A(n6528), .B(n6527), .ZN(n6530)
         );
  AOI21_X1 U7163 ( .B1(n6531), .B2(n6926), .A(n6530), .ZN(n6532) );
  OAI21_X1 U7164 ( .B1(n6533), .B2(n6590), .A(n6532), .ZN(U2992) );
  NAND3_X1 U7165 ( .A1(n6419), .A2(n6534), .A3(n6920), .ZN(n6541) );
  NAND2_X1 U7166 ( .A1(n6906), .A2(REIP_REG_25__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U7167 ( .A1(n6535), .A2(n6542), .ZN(n6536) );
  OAI211_X1 U7168 ( .C1(n6538), .C2(n6897), .A(n6537), .B(n6536), .ZN(n6539)
         );
  INV_X1 U7169 ( .A(n6539), .ZN(n6540) );
  OAI211_X1 U7170 ( .C1(n6544), .C2(n6542), .A(n6541), .B(n6540), .ZN(U2993)
         );
  INV_X1 U7171 ( .A(n6543), .ZN(n6554) );
  AOI211_X1 U7172 ( .C1(n6546), .C2(n6554), .A(n6545), .B(n6544), .ZN(n6547)
         );
  AOI211_X1 U7173 ( .C1(n6926), .C2(n6549), .A(n6548), .B(n6547), .ZN(n6550)
         );
  OAI21_X1 U7174 ( .B1(n6551), .B2(n6590), .A(n6550), .ZN(U2994) );
  INV_X1 U7175 ( .A(n6552), .ZN(n6561) );
  NAND2_X1 U7176 ( .A1(n6553), .A2(n6920), .ZN(n6559) );
  NOR2_X1 U7177 ( .A1(n6554), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6555)
         );
  AOI211_X1 U7178 ( .C1(n6557), .C2(n6926), .A(n6556), .B(n6555), .ZN(n6558)
         );
  OAI211_X1 U7179 ( .C1(n6561), .C2(n6560), .A(n6559), .B(n6558), .ZN(U2995)
         );
  OAI21_X1 U7180 ( .B1(n6562), .B2(n6874), .A(n6601), .ZN(n6571) );
  NAND2_X1 U7181 ( .A1(n6595), .A2(n6562), .ZN(n6575) );
  OR3_X1 U7182 ( .A1(n6575), .A2(n6564), .A3(n6563), .ZN(n6565) );
  OAI211_X1 U7183 ( .C1(n6567), .C2(n6897), .A(n6566), .B(n6565), .ZN(n6568)
         );
  AOI21_X1 U7184 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6571), .A(n6568), 
        .ZN(n6569) );
  OAI21_X1 U7185 ( .B1(n6570), .B2(n6590), .A(n6569), .ZN(U2996) );
  INV_X1 U7186 ( .A(n6571), .ZN(n6580) );
  NAND3_X1 U7187 ( .A1(n6573), .A2(n6920), .A3(n6572), .ZN(n6578) );
  OAI21_X1 U7188 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n6575), .A(n6574), 
        .ZN(n6576) );
  AOI21_X1 U7189 ( .B1(n7055), .B2(n6926), .A(n6576), .ZN(n6577) );
  OAI211_X1 U7190 ( .C1(n6580), .C2(n6579), .A(n6578), .B(n6577), .ZN(U2997)
         );
  INV_X1 U7191 ( .A(n6601), .ZN(n6588) );
  INV_X1 U7192 ( .A(n6581), .ZN(n6583) );
  NAND3_X1 U7193 ( .A1(n6595), .A2(n6583), .A3(n6582), .ZN(n6584) );
  OAI211_X1 U7194 ( .C1(n6586), .C2(n6897), .A(n6585), .B(n6584), .ZN(n6587)
         );
  AOI21_X1 U7195 ( .B1(n6588), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6587), 
        .ZN(n6589) );
  OAI21_X1 U7196 ( .B1(n6591), .B2(n6590), .A(n6589), .ZN(U2998) );
  INV_X1 U7197 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U7198 ( .B1(n6594), .B2(n6593), .A(n6592), .ZN(n6775) );
  NAND2_X1 U7199 ( .A1(n6775), .A2(n6920), .ZN(n6599) );
  INV_X1 U7200 ( .A(n6595), .ZN(n6596) );
  OAI22_X1 U7201 ( .A1(n6894), .A2(n6694), .B1(n6596), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6597) );
  AOI21_X1 U7202 ( .B1(n7037), .B2(n6926), .A(n6597), .ZN(n6598) );
  OAI211_X1 U7203 ( .C1(n6601), .C2(n6600), .A(n6599), .B(n6598), .ZN(U2999)
         );
  INV_X1 U7204 ( .A(n6602), .ZN(n6923) );
  INV_X1 U7205 ( .A(n6603), .ZN(n6604) );
  NAND2_X1 U7206 ( .A1(n6604), .A2(n6605), .ZN(n6606) );
  MUX2_X1 U7207 ( .A(n6606), .B(n6605), .S(n6473), .Z(n6608) );
  NAND2_X1 U7208 ( .A1(n6608), .A2(n6607), .ZN(n6769) );
  NAND2_X1 U7209 ( .A1(n6769), .A2(n6920), .ZN(n6612) );
  NAND2_X1 U7210 ( .A1(n6906), .A2(REIP_REG_17__SCAN_IN), .ZN(n6609) );
  OAI21_X1 U7211 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6916), .A(n6609), 
        .ZN(n6610) );
  AOI21_X1 U7212 ( .B1(n7026), .B2(n6926), .A(n6610), .ZN(n6611) );
  OAI211_X1 U7213 ( .C1(n6923), .C2(n6917), .A(n6612), .B(n6611), .ZN(U3001)
         );
  NOR3_X1 U7214 ( .A1(n6614), .A2(n4738), .A3(n6613), .ZN(n6615) );
  AOI21_X1 U7215 ( .B1(n7071), .B2(n3468), .A(n6615), .ZN(n6616) );
  OAI21_X1 U7216 ( .B1(n6618), .B2(n6617), .A(n6616), .ZN(n7076) );
  INV_X1 U7217 ( .A(n7076), .ZN(n6626) );
  INV_X1 U7218 ( .A(n6619), .ZN(n6625) );
  AOI22_X1 U7219 ( .A1(n6623), .A2(n6622), .B1(n6621), .B2(n6620), .ZN(n6624)
         );
  OAI21_X1 U7220 ( .B1(n6626), .B2(n6625), .A(n6624), .ZN(n6628) );
  INV_X1 U7221 ( .A(n6627), .ZN(n7069) );
  MUX2_X1 U7222 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6628), .S(n7069), 
        .Z(U3460) );
  INV_X1 U7223 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6630) );
  INV_X1 U7224 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6786) );
  INV_X2 U7225 ( .A(n7139), .ZN(n6703) );
  CLKBUF_X1 U7226 ( .A(n6631), .Z(n7124) );
  INV_X1 U7227 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U7228 ( .A1(n6789), .A2(n6786), .ZN(n6780) );
  AOI21_X1 U7229 ( .B1(n6629), .B2(n6780), .A(n7124), .ZN(n7123) );
  AOI21_X1 U7230 ( .B1(n6630), .B2(n7124), .A(n7123), .ZN(U3451) );
  AND2_X1 U7231 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n7124), .ZN(U3180) );
  AND2_X1 U7232 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n7124), .ZN(U3179) );
  AND2_X1 U7233 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6631), .ZN(U3178) );
  AND2_X1 U7234 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6631), .ZN(U3177) );
  AND2_X1 U7235 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6631), .ZN(U3176) );
  AND2_X1 U7236 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6631), .ZN(U3175) );
  AND2_X1 U7237 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6631), .ZN(U3174) );
  AND2_X1 U7238 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6631), .ZN(U3173) );
  AND2_X1 U7239 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6631), .ZN(U3172) );
  AND2_X1 U7240 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6631), .ZN(U3171) );
  AND2_X1 U7241 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6631), .ZN(U3170) );
  AND2_X1 U7242 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6631), .ZN(U3169) );
  AND2_X1 U7243 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6631), .ZN(U3168) );
  AND2_X1 U7244 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6631), .ZN(U3167) );
  AND2_X1 U7245 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6631), .ZN(U3166) );
  AND2_X1 U7246 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6631), .ZN(U3165) );
  AND2_X1 U7247 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n7124), .ZN(U3164) );
  AND2_X1 U7248 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n7124), .ZN(U3163) );
  AND2_X1 U7249 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n7124), .ZN(U3162) );
  AND2_X1 U7250 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n7124), .ZN(U3161) );
  AND2_X1 U7251 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n7124), .ZN(U3160) );
  AND2_X1 U7252 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n7124), .ZN(U3159) );
  AND2_X1 U7253 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7124), .ZN(U3158) );
  AND2_X1 U7254 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7124), .ZN(U3157) );
  AND2_X1 U7255 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7124), .ZN(U3156) );
  AND2_X1 U7256 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7124), .ZN(U3155) );
  AND2_X1 U7257 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7124), .ZN(U3154) );
  AND2_X1 U7258 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7124), .ZN(U3153) );
  AND2_X1 U7259 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7124), .ZN(U3152) );
  AND2_X1 U7260 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7124), .ZN(U3151) );
  AND2_X1 U7261 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6632), .ZN(U3019)
         );
  AND2_X1 U7262 ( .A1(n6648), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U7263 ( .A1(n7129), .A2(n6786), .ZN(n6634) );
  AOI21_X1 U7264 ( .B1(n6634), .B2(n6633), .A(n7139), .ZN(U2789) );
  AOI22_X1 U7265 ( .A1(n6666), .A2(LWORD_REG_0__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6636) );
  OAI21_X1 U7266 ( .B1(n6637), .B2(n6668), .A(n6636), .ZN(U2923) );
  AOI22_X1 U7267 ( .A1(n6666), .A2(LWORD_REG_1__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6638) );
  OAI21_X1 U7268 ( .B1(n6639), .B2(n6668), .A(n6638), .ZN(U2922) );
  AOI22_X1 U7269 ( .A1(n6666), .A2(LWORD_REG_2__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6640) );
  OAI21_X1 U7270 ( .B1(n6641), .B2(n6668), .A(n6640), .ZN(U2921) );
  AOI22_X1 U7271 ( .A1(n6666), .A2(LWORD_REG_3__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6642) );
  OAI21_X1 U7272 ( .B1(n6643), .B2(n6668), .A(n6642), .ZN(U2920) );
  AOI22_X1 U7273 ( .A1(n6666), .A2(LWORD_REG_4__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6644) );
  OAI21_X1 U7274 ( .B1(n6645), .B2(n6668), .A(n6644), .ZN(U2919) );
  AOI22_X1 U7275 ( .A1(n6666), .A2(LWORD_REG_5__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6646) );
  OAI21_X1 U7276 ( .B1(n6647), .B2(n6668), .A(n6646), .ZN(U2918) );
  AOI22_X1 U7277 ( .A1(n6666), .A2(LWORD_REG_6__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6649) );
  OAI21_X1 U7278 ( .B1(n6650), .B2(n6668), .A(n6649), .ZN(U2917) );
  AOI22_X1 U7279 ( .A1(n6666), .A2(LWORD_REG_7__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6651) );
  OAI21_X1 U7280 ( .B1(n6652), .B2(n6668), .A(n6651), .ZN(U2916) );
  AOI22_X1 U7281 ( .A1(n6666), .A2(LWORD_REG_8__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6653) );
  OAI21_X1 U7282 ( .B1(n6654), .B2(n6668), .A(n6653), .ZN(U2915) );
  AOI22_X1 U7283 ( .A1(n6666), .A2(LWORD_REG_9__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U7284 ( .B1(n6656), .B2(n6668), .A(n6655), .ZN(U2914) );
  AOI22_X1 U7285 ( .A1(n6666), .A2(LWORD_REG_10__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6657) );
  OAI21_X1 U7286 ( .B1(n6658), .B2(n6668), .A(n6657), .ZN(U2913) );
  AOI22_X1 U7287 ( .A1(n6666), .A2(LWORD_REG_11__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6659) );
  OAI21_X1 U7288 ( .B1(n6660), .B2(n6668), .A(n6659), .ZN(U2912) );
  AOI22_X1 U7289 ( .A1(n6666), .A2(LWORD_REG_12__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6661) );
  OAI21_X1 U7290 ( .B1(n4003), .B2(n6668), .A(n6661), .ZN(U2911) );
  AOI22_X1 U7291 ( .A1(n6666), .A2(LWORD_REG_13__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U7292 ( .B1(n6663), .B2(n6668), .A(n6662), .ZN(U2910) );
  AOI22_X1 U7293 ( .A1(n6666), .A2(LWORD_REG_14__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U7294 ( .B1(n6665), .B2(n6668), .A(n6664), .ZN(U2909) );
  AOI22_X1 U7295 ( .A1(n6666), .A2(LWORD_REG_15__SCAN_IN), .B1(n6648), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7296 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(U2908) );
  NOR2_X2 U7297 ( .A1(n6789), .A2(n6703), .ZN(n6716) );
  NAND2_X1 U7298 ( .A1(n6789), .A2(n7139), .ZN(n6718) );
  AOI22_X1 U7299 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6703), .ZN(n6670) );
  OAI21_X1 U7300 ( .B1(n5590), .B2(n6706), .A(n6670), .ZN(U3184) );
  AOI22_X1 U7301 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6703), .ZN(n6671) );
  OAI21_X1 U7302 ( .B1(n6949), .B2(n6718), .A(n6671), .ZN(U3185) );
  AOI22_X1 U7303 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6703), .ZN(n6672) );
  OAI21_X1 U7304 ( .B1(n6949), .B2(n6706), .A(n6672), .ZN(U3186) );
  AOI22_X1 U7305 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6703), .ZN(n6673) );
  OAI21_X1 U7306 ( .B1(n6959), .B2(n6706), .A(n6673), .ZN(U3187) );
  INV_X1 U7307 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6994) );
  AOI22_X1 U7308 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6703), .ZN(n6674) );
  OAI21_X1 U7309 ( .B1(n6994), .B2(n6718), .A(n6674), .ZN(U3188) );
  AOI22_X1 U7310 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6703), .ZN(n6675) );
  OAI21_X1 U7311 ( .B1(n7006), .B2(n6718), .A(n6675), .ZN(U3189) );
  AOI22_X1 U7312 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6703), .ZN(n6676) );
  OAI21_X1 U7313 ( .B1(n5469), .B2(n6718), .A(n6676), .ZN(U3190) );
  AOI22_X1 U7314 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6703), .ZN(n6677) );
  OAI21_X1 U7315 ( .B1(n6679), .B2(n6718), .A(n6677), .ZN(U3191) );
  AOI22_X1 U7316 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6703), .ZN(n6678) );
  OAI21_X1 U7317 ( .B1(n6679), .B2(n6706), .A(n6678), .ZN(U3192) );
  INV_X1 U7318 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7319 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6703), .ZN(n6680) );
  OAI21_X1 U7320 ( .B1(n6895), .B2(n6718), .A(n6680), .ZN(U3193) );
  AOI22_X1 U7321 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6703), .ZN(n6681) );
  OAI21_X1 U7322 ( .B1(n6682), .B2(n6718), .A(n6681), .ZN(U3194) );
  AOI22_X1 U7323 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6703), .ZN(n6683) );
  OAI21_X1 U7324 ( .B1(n6685), .B2(n6718), .A(n6683), .ZN(U3195) );
  AOI22_X1 U7325 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6703), .ZN(n6684) );
  OAI21_X1 U7326 ( .B1(n6685), .B2(n6706), .A(n6684), .ZN(U3196) );
  AOI22_X1 U7327 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6703), .ZN(n6686) );
  OAI21_X1 U7328 ( .B1(n6688), .B2(n6718), .A(n6686), .ZN(U3197) );
  AOI22_X1 U7329 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6703), .ZN(n6687) );
  OAI21_X1 U7330 ( .B1(n6688), .B2(n6706), .A(n6687), .ZN(U3198) );
  AOI22_X1 U7331 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6703), .ZN(n6689) );
  OAI21_X1 U7332 ( .B1(n6691), .B2(n6718), .A(n6689), .ZN(U3199) );
  AOI22_X1 U7333 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6703), .ZN(n6690) );
  OAI21_X1 U7334 ( .B1(n6691), .B2(n6706), .A(n6690), .ZN(U3200) );
  AOI22_X1 U7335 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6703), .ZN(n6692) );
  OAI21_X1 U7336 ( .B1(n6694), .B2(n6718), .A(n6692), .ZN(U3201) );
  AOI22_X1 U7337 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6703), .ZN(n6693) );
  OAI21_X1 U7338 ( .B1(n6694), .B2(n6706), .A(n6693), .ZN(U3202) );
  AOI22_X1 U7339 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6703), .ZN(n6695) );
  OAI21_X1 U7340 ( .B1(n6696), .B2(n6706), .A(n6695), .ZN(U3203) );
  AOI22_X1 U7341 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6703), .ZN(n6697) );
  OAI21_X1 U7342 ( .B1(n7049), .B2(n6706), .A(n6697), .ZN(U3204) );
  AOI22_X1 U7343 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6703), .ZN(n6698) );
  OAI21_X1 U7344 ( .B1(n6700), .B2(n6718), .A(n6698), .ZN(U3205) );
  AOI22_X1 U7345 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6703), .ZN(n6699) );
  OAI21_X1 U7346 ( .B1(n6700), .B2(n6706), .A(n6699), .ZN(U3206) );
  AOI22_X1 U7347 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6703), .ZN(n6701) );
  OAI21_X1 U7348 ( .B1(n6702), .B2(n6706), .A(n6701), .ZN(U3207) );
  AOI22_X1 U7349 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6704), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6703), .ZN(n6705) );
  OAI21_X1 U7350 ( .B1(n6707), .B2(n6706), .A(n6705), .ZN(U3208) );
  AOI22_X1 U7351 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6703), .ZN(n6708) );
  OAI21_X1 U7352 ( .B1(n6709), .B2(n6718), .A(n6708), .ZN(U3209) );
  AOI22_X1 U7353 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6703), .ZN(n6710) );
  OAI21_X1 U7354 ( .B1(n6711), .B2(n6718), .A(n6710), .ZN(U3210) );
  AOI22_X1 U7355 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6703), .ZN(n6712) );
  OAI21_X1 U7356 ( .B1(n6713), .B2(n6718), .A(n6712), .ZN(U3211) );
  AOI22_X1 U7357 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6703), .ZN(n6714) );
  OAI21_X1 U7358 ( .B1(n6715), .B2(n6718), .A(n6714), .ZN(U3212) );
  AOI22_X1 U7359 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6716), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6703), .ZN(n6717) );
  OAI21_X1 U7360 ( .B1(n5933), .B2(n6718), .A(n6717), .ZN(U3213) );
  MUX2_X1 U7361 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6703), .Z(U3445) );
  NOR4_X1 U7362 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6722) );
  NOR4_X1 U7363 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6721) );
  NOR4_X1 U7364 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6720) );
  NOR4_X1 U7365 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6719) );
  NAND4_X1 U7366 ( .A1(n6722), .A2(n6721), .A3(n6720), .A4(n6719), .ZN(n6728)
         );
  NOR4_X1 U7367 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6726) );
  AOI211_X1 U7368 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6725) );
  NOR4_X1 U7369 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6724) );
  NOR4_X1 U7370 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6723) );
  NAND4_X1 U7371 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6727)
         );
  NOR2_X1 U7372 ( .A1(n6728), .A2(n6727), .ZN(n6738) );
  NAND2_X1 U7373 ( .A1(n6738), .A2(n5590), .ZN(n6739) );
  INV_X1 U7374 ( .A(n6738), .ZN(n6729) );
  INV_X1 U7375 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U7376 ( .A1(n6738), .A2(n6732), .ZN(n6733) );
  NOR3_X1 U7377 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(n6733), .ZN(n6736) );
  AOI21_X1 U7378 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6729), .A(n6736), .ZN(
        n6730) );
  OAI21_X1 U7379 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6739), .A(n6730), .ZN(
        U2795) );
  MUX2_X1 U7380 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6703), .Z(U3446) );
  NOR2_X1 U7381 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .ZN(n6731) );
  AOI21_X1 U7382 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6732), .A(n6731), .ZN(
        n6735) );
  OAI211_X1 U7383 ( .C1(BYTEENABLE_REG_2__SCAN_IN), .C2(n6738), .A(n6739), .B(
        n6733), .ZN(n6734) );
  OAI21_X1 U7384 ( .B1(n6735), .B2(n6739), .A(n6734), .ZN(U3468) );
  MUX2_X1 U7385 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6703), .Z(U3447) );
  OAI22_X1 U7386 ( .A1(n6739), .A2(n6736), .B1(BYTEENABLE_REG_1__SCAN_IN), 
        .B2(n6738), .ZN(n6737) );
  INV_X1 U7387 ( .A(n6737), .ZN(U2794) );
  MUX2_X1 U7388 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6703), .Z(U3448) );
  OAI22_X1 U7389 ( .A1(n6739), .A2(REIP_REG_0__SCAN_IN), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(n6738), .ZN(n6740) );
  INV_X1 U7390 ( .A(n6740), .ZN(U3469) );
  AOI22_X1 U7391 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6772), .B1(n6906), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6747) );
  NAND2_X1 U7392 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  XOR2_X1 U7393 ( .A(n6744), .B(n6743), .Z(n6841) );
  INV_X1 U7394 ( .A(n6935), .ZN(n6745) );
  AOI22_X1 U7395 ( .A1(n6841), .A2(n6774), .B1(n6773), .B2(n6745), .ZN(n6746)
         );
  OAI211_X1 U7396 ( .C1(n6778), .C2(n6940), .A(n6747), .B(n6746), .ZN(U2984)
         );
  OAI22_X1 U7397 ( .A1(n6980), .A2(n6748), .B1(n6978), .B2(n6778), .ZN(n6749)
         );
  AOI21_X1 U7398 ( .B1(n6750), .B2(n6774), .A(n6749), .ZN(n6752) );
  OAI211_X1 U7399 ( .C1(n6753), .C2(n6975), .A(n6752), .B(n6751), .ZN(U2981)
         );
  AOI22_X1 U7400 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6772), .B1(n6906), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U7401 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  XNOR2_X1 U7402 ( .A(n6754), .B(n6757), .ZN(n6835) );
  INV_X1 U7403 ( .A(n6988), .ZN(n6758) );
  AOI22_X1 U7404 ( .A1(n6835), .A2(n6774), .B1(n6773), .B2(n6758), .ZN(n6759)
         );
  OAI211_X1 U7405 ( .C1(n6778), .C2(n6987), .A(n6760), .B(n6759), .ZN(U2980)
         );
  AOI22_X1 U7406 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6772), .B1(n6906), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6768) );
  OAI21_X1 U7407 ( .B1(n6761), .B2(n6764), .A(n6763), .ZN(n6765) );
  INV_X1 U7408 ( .A(n6765), .ZN(n6863) );
  AOI22_X1 U7409 ( .A1(n6863), .A2(n6774), .B1(n6773), .B2(n6766), .ZN(n6767)
         );
  OAI211_X1 U7410 ( .C1(n6778), .C2(n6999), .A(n6768), .B(n6767), .ZN(U2979)
         );
  AOI22_X1 U7411 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6772), .B1(n6906), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U7412 ( .A1(n6769), .A2(n6774), .B1(n6773), .B2(n7197), .ZN(n6770)
         );
  OAI211_X1 U7413 ( .C1(n6778), .C2(n7033), .A(n6771), .B(n6770), .ZN(U2969)
         );
  AOI22_X1 U7414 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6772), .B1(n6906), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7415 ( .A1(n6775), .A2(n6774), .B1(n6773), .B2(n7200), .ZN(n6776)
         );
  OAI211_X1 U7416 ( .C1(n6778), .C2(n7039), .A(n6777), .B(n6776), .ZN(U2967)
         );
  NOR2_X1 U7417 ( .A1(n7139), .A2(D_C_N_REG_SCAN_IN), .ZN(n6779) );
  AOI22_X1 U7418 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7139), .B1(n6780), .B2(
        n6779), .ZN(U2791) );
  NAND2_X1 U7419 ( .A1(n6798), .A2(n6781), .ZN(n6782) );
  OAI211_X1 U7420 ( .C1(n6798), .C2(n6784), .A(n6783), .B(n6782), .ZN(U3474)
         );
  OAI22_X1 U7421 ( .A1(n6703), .A2(n6784), .B1(W_R_N_REG_SCAN_IN), .B2(n7139), 
        .ZN(n6785) );
  INV_X1 U7422 ( .A(n6785), .ZN(U3470) );
  NAND2_X1 U7423 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7132) );
  NOR2_X1 U7424 ( .A1(n6786), .A2(n7131), .ZN(n7135) );
  NOR2_X1 U7425 ( .A1(n6787), .A2(n6788), .ZN(n7126) );
  OAI22_X1 U7426 ( .A1(n7135), .A2(n7126), .B1(n6789), .B2(n6788), .ZN(n6790)
         );
  NAND3_X1 U7427 ( .A1(n6791), .A2(n7132), .A3(n6790), .ZN(U3182) );
  OAI221_X1 U7428 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n7143), .A(n7109), .ZN(n6793) );
  OAI21_X1 U7429 ( .B1(n6794), .B2(n6793), .A(n6792), .ZN(U3150) );
  OAI211_X1 U7430 ( .C1(n4415), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n7143), .ZN(n6795) );
  OAI21_X1 U7431 ( .B1(n6796), .B2(n6795), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6797) );
  NAND2_X1 U7432 ( .A1(n6797), .A2(n7117), .ZN(n6801) );
  AOI211_X1 U7433 ( .C1(n6666), .C2(n7143), .A(n6799), .B(n6798), .ZN(n6800)
         );
  MUX2_X1 U7434 ( .A(n6801), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6800), .Z(
        U3472) );
  INV_X1 U7435 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U7436 ( .A1(n6803), .A2(n6802), .ZN(n6811) );
  AOI21_X1 U7437 ( .B1(n6805), .B2(n6926), .A(n6804), .ZN(n6810) );
  INV_X1 U7438 ( .A(n6806), .ZN(n6807) );
  AOI22_X1 U7439 ( .A1(n6808), .A2(n6920), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6807), .ZN(n6809) );
  OAI211_X1 U7440 ( .C1(n6902), .C2(n6811), .A(n6810), .B(n6809), .ZN(U3004)
         );
  AOI21_X1 U7441 ( .B1(n6926), .B2(n6813), .A(n6812), .ZN(n6821) );
  AOI22_X1 U7442 ( .A1(n6815), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n6920), 
        .B2(n6814), .ZN(n6820) );
  OAI211_X1 U7443 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6818), .A(n6817), 
        .B(n6816), .ZN(n6819) );
  NAND3_X1 U7444 ( .A1(n6821), .A2(n6820), .A3(n6819), .ZN(U3017) );
  NAND2_X1 U7445 ( .A1(n6822), .A2(n6920), .ZN(n6825) );
  AOI21_X1 U7446 ( .B1(n6926), .B2(n6960), .A(n6823), .ZN(n6824) );
  OAI211_X1 U7447 ( .C1(n4445), .C2(n6826), .A(n6825), .B(n6824), .ZN(n6827)
         );
  INV_X1 U7448 ( .A(n6827), .ZN(n6830) );
  OAI211_X1 U7449 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6831), .B(n6828), .ZN(n6829) );
  NAND2_X1 U7450 ( .A1(n6830), .A2(n6829), .ZN(U3014) );
  NAND2_X1 U7451 ( .A1(n6832), .A2(n6831), .ZN(n6856) );
  INV_X1 U7452 ( .A(n6833), .ZN(n6991) );
  AOI22_X1 U7453 ( .A1(n6926), .A2(n6991), .B1(n6906), .B2(REIP_REG_6__SCAN_IN), .ZN(n6837) );
  AOI22_X1 U7454 ( .A1(n6835), .A2(n6920), .B1(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n6834), .ZN(n6836) );
  OAI211_X1 U7455 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6856), .A(n6837), 
        .B(n6836), .ZN(U3012) );
  AOI22_X1 U7456 ( .A1(n6926), .A2(n6932), .B1(n6906), .B2(REIP_REG_2__SCAN_IN), .ZN(n6846) );
  OAI221_X1 U7457 ( .B1(n6839), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6839), .C2(n6838), .A(n6853), .ZN(n6845) );
  AOI22_X1 U7458 ( .A1(n6841), .A2(n6920), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6840), .ZN(n6844) );
  NAND3_X1 U7459 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4427), .A3(n6842), 
        .ZN(n6843) );
  NAND4_X1 U7460 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(U3016)
         );
  INV_X1 U7461 ( .A(n6847), .ZN(n6849) );
  NOR2_X1 U7462 ( .A1(n6849), .A2(n6848), .ZN(n6851) );
  AOI211_X1 U7463 ( .C1(n6853), .C2(n6852), .A(n6851), .B(n6850), .ZN(n6872)
         );
  AOI21_X1 U7464 ( .B1(n6926), .B2(n6855), .A(n6854), .ZN(n6861) );
  NOR2_X1 U7465 ( .A1(n6857), .A2(n6856), .ZN(n6867) );
  AOI21_X1 U7466 ( .B1(n6862), .B2(n6866), .A(n6873), .ZN(n6858) );
  AOI22_X1 U7467 ( .A1(n6859), .A2(n6920), .B1(n6867), .B2(n6858), .ZN(n6860)
         );
  OAI211_X1 U7468 ( .C1(n6872), .C2(n6862), .A(n6861), .B(n6860), .ZN(U3010)
         );
  AOI22_X1 U7469 ( .A1(n6926), .A2(n6996), .B1(n6906), .B2(REIP_REG_7__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7470 ( .A1(n6863), .A2(n6920), .B1(n6867), .B2(n6866), .ZN(n6864)
         );
  OAI211_X1 U7471 ( .C1(n6872), .C2(n6866), .A(n6865), .B(n6864), .ZN(U3011)
         );
  NAND2_X1 U7472 ( .A1(n6873), .A2(n6867), .ZN(n6885) );
  AOI22_X1 U7473 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6869), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6868), .ZN(n6878) );
  AOI21_X1 U7474 ( .B1(n6926), .B2(n6871), .A(n6870), .ZN(n6877) );
  OAI21_X1 U7475 ( .B1(n6874), .B2(n6873), .A(n6872), .ZN(n6881) );
  AOI22_X1 U7476 ( .A1(n6875), .A2(n6920), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6881), .ZN(n6876) );
  OAI211_X1 U7477 ( .C1(n6885), .C2(n6878), .A(n6877), .B(n6876), .ZN(U3008)
         );
  AOI22_X1 U7478 ( .A1(n6926), .A2(n6879), .B1(n6906), .B2(REIP_REG_9__SCAN_IN), .ZN(n6884) );
  INV_X1 U7479 ( .A(n6880), .ZN(n6882) );
  AOI22_X1 U7480 ( .A1(n6882), .A2(n6920), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6881), .ZN(n6883) );
  OAI211_X1 U7481 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6885), .A(n6884), 
        .B(n6883), .ZN(U3009) );
  INV_X1 U7482 ( .A(n6886), .ZN(n6888) );
  AOI21_X1 U7483 ( .B1(n6888), .B2(n6926), .A(n6887), .ZN(n6893) );
  AOI21_X1 U7484 ( .B1(n5760), .B2(n4571), .A(n6902), .ZN(n6890) );
  AOI22_X1 U7485 ( .A1(n6891), .A2(n6920), .B1(n6890), .B2(n6889), .ZN(n6892)
         );
  OAI211_X1 U7486 ( .C1(n6901), .C2(n5760), .A(n6893), .B(n6892), .ZN(U3006)
         );
  OAI22_X1 U7487 ( .A1(n6897), .A2(n6896), .B1(n6895), .B2(n6894), .ZN(n6898)
         );
  AOI21_X1 U7488 ( .B1(n6899), .B2(n6920), .A(n6898), .ZN(n6900) );
  OAI221_X1 U7489 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6902), .C1(
        n4571), .C2(n6901), .A(n6900), .ZN(U3007) );
  INV_X1 U7490 ( .A(n6903), .ZN(n6905) );
  AOI22_X1 U7491 ( .A1(n6905), .A2(n6920), .B1(n6926), .B2(n6904), .ZN(n6913)
         );
  NAND2_X1 U7492 ( .A1(n6906), .A2(REIP_REG_16__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U7493 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6907), .ZN(n6911) );
  OAI211_X1 U7494 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6909), .B(n6908), .ZN(n6910) );
  NAND4_X1 U7495 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(U3002)
         );
  INV_X1 U7496 ( .A(n6914), .ZN(n6921) );
  INV_X1 U7497 ( .A(n6915), .ZN(n6919) );
  NOR3_X1 U7498 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6917), .A3(n6916), 
        .ZN(n6918) );
  AOI211_X1 U7499 ( .C1(n6921), .C2(n6920), .A(n6919), .B(n6918), .ZN(n6929)
         );
  INV_X1 U7500 ( .A(n6922), .ZN(n6924) );
  OAI21_X1 U7501 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6924), .A(n6923), 
        .ZN(n6927) );
  AOI22_X1 U7502 ( .A1(n6927), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n6926), .B2(n6925), .ZN(n6928) );
  NAND2_X1 U7503 ( .A1(n6929), .A2(n6928), .ZN(U3000) );
  NAND2_X1 U7504 ( .A1(n6930), .A2(n6948), .ZN(n6931) );
  AOI22_X1 U7505 ( .A1(n7056), .A2(n6932), .B1(REIP_REG_2__SCAN_IN), .B2(n6931), .ZN(n6939) );
  NOR2_X1 U7506 ( .A1(n6970), .A2(n4771), .ZN(n6937) );
  NOR3_X1 U7507 ( .A1(n6958), .A2(REIP_REG_2__SCAN_IN), .A3(n5590), .ZN(n6933)
         );
  AOI21_X1 U7508 ( .B1(n7035), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6933), 
        .ZN(n6934) );
  OAI21_X1 U7509 ( .B1(n6979), .B2(n6935), .A(n6934), .ZN(n6936) );
  AOI211_X1 U7510 ( .C1(EBX_REG_2__SCAN_IN), .C2(n7053), .A(n6937), .B(n6936), 
        .ZN(n6938) );
  OAI211_X1 U7511 ( .C1(n6940), .C2(n7060), .A(n6939), .B(n6938), .ZN(U2825)
         );
  OAI22_X1 U7512 ( .A1(n6942), .A2(n7050), .B1(n7060), .B2(n6941), .ZN(n6946)
         );
  OAI22_X1 U7513 ( .A1(n6944), .A2(n7025), .B1(n6943), .B2(n6979), .ZN(n6945)
         );
  AOI211_X1 U7514 ( .C1(n6947), .C2(n4732), .A(n6946), .B(n6945), .ZN(n6954)
         );
  NAND2_X1 U7515 ( .A1(n6956), .A2(n6948), .ZN(n6972) );
  OAI21_X1 U7516 ( .B1(n6951), .B2(n6950), .A(n6949), .ZN(n6952) );
  NAND3_X1 U7517 ( .A1(n6971), .A2(n6972), .A3(n6952), .ZN(n6953) );
  OAI211_X1 U7518 ( .C1(n6955), .C2(n7028), .A(n6954), .B(n6953), .ZN(U2824)
         );
  INV_X1 U7519 ( .A(n6956), .ZN(n6957) );
  NOR2_X1 U7520 ( .A1(n6958), .A2(n6957), .ZN(n6985) );
  AOI22_X1 U7521 ( .A1(n7056), .A2(n6960), .B1(n6985), .B2(n6959), .ZN(n6969)
         );
  NAND3_X1 U7522 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6971), .A3(n6972), .ZN(n6961) );
  OAI211_X1 U7523 ( .C1(n7050), .C2(n6962), .A(n7023), .B(n6961), .ZN(n6967)
         );
  INV_X1 U7524 ( .A(n6963), .ZN(n6964) );
  OAI22_X1 U7525 ( .A1(n6965), .A2(n6979), .B1(n6964), .B2(n7060), .ZN(n6966)
         );
  AOI211_X1 U7526 ( .C1(EBX_REG_4__SCAN_IN), .C2(n7053), .A(n6967), .B(n6966), 
        .ZN(n6968) );
  OAI211_X1 U7527 ( .C1(n7064), .C2(n6970), .A(n6969), .B(n6968), .ZN(U2823)
         );
  AOI21_X1 U7528 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6985), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U7529 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n6973) );
  OAI21_X1 U7530 ( .B1(n6973), .B2(n6972), .A(n6971), .ZN(n7004) );
  INV_X1 U7531 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6974) );
  OAI22_X1 U7532 ( .A1(n6975), .A2(n7050), .B1(n6974), .B2(n7025), .ZN(n6976)
         );
  AOI211_X1 U7533 ( .C1(n7056), .C2(n6977), .A(n7034), .B(n6976), .ZN(n6983)
         );
  OAI22_X1 U7534 ( .A1(n6980), .A2(n6979), .B1(n6978), .B2(n7060), .ZN(n6981)
         );
  INV_X1 U7535 ( .A(n6981), .ZN(n6982) );
  OAI211_X1 U7536 ( .C1(n6984), .C2(n7004), .A(n6983), .B(n6982), .ZN(U2822)
         );
  NAND4_X1 U7537 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n6985), .A4(n6994), .ZN(n7005) );
  OAI211_X1 U7538 ( .C1(n7050), .C2(n6986), .A(n7023), .B(n7005), .ZN(n6990)
         );
  OAI22_X1 U7539 ( .A1(n6988), .A2(n7014), .B1(n6987), .B2(n7060), .ZN(n6989)
         );
  AOI211_X1 U7540 ( .C1(EBX_REG_6__SCAN_IN), .C2(n7053), .A(n6990), .B(n6989), 
        .ZN(n6993) );
  NAND2_X1 U7541 ( .A1(n7056), .A2(n6991), .ZN(n6992) );
  OAI211_X1 U7542 ( .C1(n7004), .C2(n6994), .A(n6993), .B(n6992), .ZN(U2821)
         );
  INV_X1 U7543 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6998) );
  AOI22_X1 U7544 ( .A1(n7056), .A2(n6996), .B1(n6995), .B2(n7006), .ZN(n6997)
         );
  OAI211_X1 U7545 ( .C1(n7050), .C2(n6998), .A(n6997), .B(n7023), .ZN(n7002)
         );
  OAI22_X1 U7546 ( .A1(n7000), .A2(n7014), .B1(n6999), .B2(n7060), .ZN(n7001)
         );
  AOI211_X1 U7547 ( .C1(EBX_REG_7__SCAN_IN), .C2(n7053), .A(n7002), .B(n7001), 
        .ZN(n7003) );
  OAI221_X1 U7548 ( .B1(n7006), .B2(n7005), .C1(n7006), .C2(n7004), .A(n7003), 
        .ZN(U2820) );
  NAND2_X1 U7549 ( .A1(n7053), .A2(EBX_REG_15__SCAN_IN), .ZN(n7008) );
  AOI21_X1 U7550 ( .B1(n7035), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7034), 
        .ZN(n7007) );
  NAND2_X1 U7551 ( .A1(n7008), .A2(n7007), .ZN(n7009) );
  NOR2_X1 U7552 ( .A1(n7010), .A2(n7009), .ZN(n7013) );
  NAND2_X1 U7553 ( .A1(n7011), .A2(REIP_REG_15__SCAN_IN), .ZN(n7012) );
  OAI211_X1 U7554 ( .C1(n7015), .C2(n7014), .A(n7013), .B(n7012), .ZN(n7016)
         );
  AOI21_X1 U7555 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7019) );
  OAI21_X1 U7556 ( .B1(n7028), .B2(n7020), .A(n7019), .ZN(U2812) );
  OAI21_X1 U7557 ( .B1(REIP_REG_17__SCAN_IN), .B2(n7021), .A(n7036), .ZN(n7022) );
  OAI211_X1 U7558 ( .C1(n7025), .C2(n7024), .A(n7023), .B(n7022), .ZN(n7031)
         );
  INV_X1 U7559 ( .A(n7026), .ZN(n7027) );
  OAI22_X1 U7560 ( .A1(n7029), .A2(n7014), .B1(n7028), .B2(n7027), .ZN(n7030)
         );
  AOI211_X1 U7561 ( .C1(PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n7035), .A(n7031), 
        .B(n7030), .ZN(n7032) );
  OAI21_X1 U7562 ( .B1(n7033), .B2(n7060), .A(n7032), .ZN(U2810) );
  AOI21_X1 U7563 ( .B1(n7035), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7034), 
        .ZN(n7046) );
  AOI22_X1 U7564 ( .A1(EBX_REG_19__SCAN_IN), .A2(n7053), .B1(
        REIP_REG_19__SCAN_IN), .B2(n7036), .ZN(n7045) );
  NAND2_X1 U7565 ( .A1(n7037), .A2(n7056), .ZN(n7038) );
  OAI21_X1 U7566 ( .B1(n7060), .B2(n7039), .A(n7038), .ZN(n7040) );
  AOI21_X1 U7567 ( .B1(n7200), .B2(n7057), .A(n7040), .ZN(n7044) );
  OAI211_X1 U7568 ( .C1(REIP_REG_18__SCAN_IN), .C2(REIP_REG_19__SCAN_IN), .A(
        n7042), .B(n7041), .ZN(n7043) );
  NAND4_X1 U7569 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(U2808)
         );
  INV_X1 U7570 ( .A(n7047), .ZN(n7052) );
  OAI22_X1 U7571 ( .A1(n4180), .A2(n7050), .B1(n7049), .B2(n7048), .ZN(n7051)
         );
  AOI211_X1 U7572 ( .C1(n7053), .C2(EBX_REG_21__SCAN_IN), .A(n7052), .B(n7051), 
        .ZN(n7059) );
  INV_X1 U7573 ( .A(n7054), .ZN(n7205) );
  AOI22_X1 U7574 ( .A1(n7205), .A2(n7057), .B1(n7056), .B2(n7055), .ZN(n7058)
         );
  OAI211_X1 U7575 ( .C1(n7061), .C2(n7060), .A(n7059), .B(n7058), .ZN(U2806)
         );
  OAI21_X1 U7576 ( .B1(n7063), .B2(n4906), .A(n7062), .ZN(U2793) );
  INV_X1 U7577 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7068) );
  NOR4_X1 U7578 ( .A1(n7064), .A2(STATE2_REG_1__SCAN_IN), .A3(n3429), .A4(
        STATE2_REG_3__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U7579 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  OAI21_X1 U7580 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(U3455) );
  INV_X1 U7581 ( .A(n7082), .ZN(n7080) );
  AOI21_X1 U7582 ( .B1(n7071), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n7070), 
        .ZN(n7072) );
  NAND2_X1 U7583 ( .A1(n7073), .A2(n7072), .ZN(n7074) );
  NOR2_X1 U7584 ( .A1(n7074), .A2(n7075), .ZN(n7079) );
  AOI22_X1 U7585 ( .A1(n7077), .A2(n7076), .B1(n7075), .B2(n7074), .ZN(n7078)
         );
  AOI211_X1 U7586 ( .C1(n7080), .C2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n7079), .B(n7078), .ZN(n7081) );
  AOI21_X1 U7587 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7088) );
  NOR2_X1 U7588 ( .A1(n7085), .A2(n7084), .ZN(n7087) );
  INV_X1 U7589 ( .A(n7085), .ZN(n7086) );
  OAI22_X1 U7590 ( .A1(n7088), .A2(n7087), .B1(n7086), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7098) );
  AOI21_X1 U7591 ( .B1(n4906), .B2(n7090), .A(n7089), .ZN(n7092) );
  OR4_X1 U7592 ( .A1(n7094), .A2(n7093), .A3(n7092), .A4(n7091), .ZN(n7095) );
  AOI211_X1 U7593 ( .C1(n7098), .C2(n7097), .A(n7096), .B(n7095), .ZN(n7121)
         );
  INV_X1 U7594 ( .A(n7121), .ZN(n7100) );
  OAI22_X1 U7595 ( .A1(n7100), .A2(n7120), .B1(n7143), .B2(n7099), .ZN(n7101)
         );
  OAI21_X1 U7596 ( .B1(n7103), .B2(n7102), .A(n7101), .ZN(n7114) );
  OAI21_X1 U7597 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7143), .A(n7114), .ZN(
        n7112) );
  OAI211_X1 U7598 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n7112), .ZN(n7108) );
  OAI21_X1 U7599 ( .B1(READY_N), .B2(n7104), .A(n7120), .ZN(n7106) );
  AOI21_X1 U7600 ( .B1(n7106), .B2(n7114), .A(n7105), .ZN(n7107) );
  NAND2_X1 U7601 ( .A1(n7108), .A2(n7107), .ZN(U3149) );
  OAI221_X1 U7602 ( .B1(n7110), .B2(STATE2_REG_0__SCAN_IN), .C1(n7110), .C2(
        n7114), .A(n7109), .ZN(U3453) );
  AOI221_X1 U7603 ( .B1(n7113), .B2(STATE2_REG_0__SCAN_IN), .C1(n7112), .C2(
        STATE2_REG_0__SCAN_IN), .A(n7111), .ZN(n7119) );
  OAI211_X1 U7604 ( .C1(n7117), .C2(n7116), .A(n7115), .B(n7114), .ZN(n7118)
         );
  OAI211_X1 U7605 ( .C1(n7121), .C2(n7120), .A(n7119), .B(n7118), .ZN(U3148)
         );
  AOI21_X1 U7606 ( .B1(n7124), .B2(STATEBS16_REG_SCAN_IN), .A(n7123), .ZN(
        n7122) );
  INV_X1 U7607 ( .A(n7122), .ZN(U2792) );
  AOI21_X1 U7608 ( .B1(n7124), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7123), .ZN(
        n7125) );
  INV_X1 U7609 ( .A(n7125), .ZN(U3452) );
  AOI221_X1 U7610 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7134), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7138) );
  AOI221_X1 U7611 ( .B1(n7126), .B2(n6703), .C1(n7131), .C2(n6703), .A(n7138), 
        .ZN(n7127) );
  OAI221_X1 U7612 ( .B1(n7128), .B2(n7132), .C1(n7128), .C2(n6788), .A(n7127), 
        .ZN(U3181) );
  OAI21_X1 U7613 ( .B1(NA_N), .B2(n7143), .A(n7129), .ZN(n7130) );
  OAI211_X1 U7614 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7131), .A(HOLD), .B(n7130), 
        .ZN(n7137) );
  INV_X1 U7615 ( .A(n7132), .ZN(n7133) );
  OAI221_X1 U7616 ( .B1(STATE_REG_2__SCAN_IN), .B2(n7135), .C1(
        STATE_REG_2__SCAN_IN), .C2(n7134), .A(n7133), .ZN(n7136) );
  OAI221_X1 U7617 ( .B1(n7138), .B2(STATE_REG_0__SCAN_IN), .C1(n7138), .C2(
        n7137), .A(n7136), .ZN(U3183) );
  OAI22_X1 U7618 ( .A1(n6703), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n7139), .ZN(n7140) );
  INV_X1 U7619 ( .A(n7140), .ZN(U3473) );
  INV_X1 U7620 ( .A(n7141), .ZN(n7142) );
  OAI21_X1 U7621 ( .B1(n7144), .B2(n7143), .A(n7142), .ZN(n7190) );
  AOI22_X1 U7622 ( .A1(n7193), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n7185), .ZN(n7146) );
  OAI21_X1 U7623 ( .B1(n7196), .B2(n7148), .A(n7146), .ZN(U2924) );
  AOI22_X1 U7624 ( .A1(n7193), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n7185), .ZN(n7147) );
  OAI21_X1 U7625 ( .B1(n7196), .B2(n7148), .A(n7147), .ZN(U2939) );
  AOI22_X1 U7626 ( .A1(n7193), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n7185), .ZN(n7149) );
  OAI21_X1 U7627 ( .B1(n7196), .B2(n7151), .A(n7149), .ZN(U2925) );
  AOI22_X1 U7628 ( .A1(n7193), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n7185), .ZN(n7150) );
  OAI21_X1 U7629 ( .B1(n7196), .B2(n7151), .A(n7150), .ZN(U2940) );
  AOI22_X1 U7630 ( .A1(n7193), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n7185), .ZN(n7152) );
  OAI21_X1 U7631 ( .B1(n7196), .B2(n7154), .A(n7152), .ZN(U2926) );
  AOI22_X1 U7632 ( .A1(n7193), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n7185), .ZN(n7153) );
  OAI21_X1 U7633 ( .B1(n7196), .B2(n7154), .A(n7153), .ZN(U2941) );
  AOI22_X1 U7634 ( .A1(n7193), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n7185), .ZN(n7155) );
  OAI21_X1 U7635 ( .B1(n7196), .B2(n7157), .A(n7155), .ZN(U2927) );
  AOI22_X1 U7636 ( .A1(n7193), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n7185), .ZN(n7156) );
  OAI21_X1 U7637 ( .B1(n7196), .B2(n7157), .A(n7156), .ZN(U2942) );
  AOI22_X1 U7638 ( .A1(n7193), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n7185), .ZN(n7158) );
  OAI21_X1 U7639 ( .B1(n7196), .B2(n7160), .A(n7158), .ZN(U2928) );
  AOI22_X1 U7640 ( .A1(n7193), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n7185), .ZN(n7159) );
  OAI21_X1 U7641 ( .B1(n7196), .B2(n7160), .A(n7159), .ZN(U2943) );
  AOI22_X1 U7642 ( .A1(n7193), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n7185), .ZN(n7161) );
  OAI21_X1 U7643 ( .B1(n7196), .B2(n7163), .A(n7161), .ZN(U2929) );
  AOI22_X1 U7644 ( .A1(n7193), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n7185), .ZN(n7162) );
  OAI21_X1 U7645 ( .B1(n7196), .B2(n7163), .A(n7162), .ZN(U2944) );
  AOI22_X1 U7646 ( .A1(n7193), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n7185), .ZN(n7164) );
  OAI21_X1 U7647 ( .B1(n7196), .B2(n7166), .A(n7164), .ZN(U2930) );
  AOI22_X1 U7648 ( .A1(n7193), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n7185), .ZN(n7165) );
  OAI21_X1 U7649 ( .B1(n7196), .B2(n7166), .A(n7165), .ZN(U2945) );
  AOI22_X1 U7650 ( .A1(n7193), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n7185), .ZN(n7167) );
  OAI21_X1 U7651 ( .B1(n7196), .B2(n7169), .A(n7167), .ZN(U2931) );
  AOI22_X1 U7652 ( .A1(n7193), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n7185), .ZN(n7168) );
  OAI21_X1 U7653 ( .B1(n7196), .B2(n7169), .A(n7168), .ZN(U2946) );
  AOI22_X1 U7654 ( .A1(n7193), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n7185), .ZN(n7170) );
  OAI21_X1 U7655 ( .B1(n7196), .B2(n7172), .A(n7170), .ZN(U2932) );
  AOI22_X1 U7656 ( .A1(n7193), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n7185), .ZN(n7171) );
  OAI21_X1 U7657 ( .B1(n7196), .B2(n7172), .A(n7171), .ZN(U2947) );
  AOI22_X1 U7658 ( .A1(n7193), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n7185), .ZN(n7173) );
  OAI21_X1 U7659 ( .B1(n7196), .B2(n7175), .A(n7173), .ZN(U2933) );
  AOI22_X1 U7660 ( .A1(n7193), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n7185), .ZN(n7174) );
  OAI21_X1 U7661 ( .B1(n7196), .B2(n7175), .A(n7174), .ZN(U2948) );
  AOI22_X1 U7662 ( .A1(n7193), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n7185), .ZN(n7176) );
  OAI21_X1 U7663 ( .B1(n7196), .B2(n7178), .A(n7176), .ZN(U2934) );
  AOI22_X1 U7664 ( .A1(n7193), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n7185), .ZN(n7177) );
  OAI21_X1 U7665 ( .B1(n7196), .B2(n7178), .A(n7177), .ZN(U2949) );
  AOI22_X1 U7666 ( .A1(n7193), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n7185), .ZN(n7179) );
  OAI21_X1 U7667 ( .B1(n7196), .B2(n7181), .A(n7179), .ZN(U2935) );
  AOI22_X1 U7668 ( .A1(n7193), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n7185), .ZN(n7180) );
  OAI21_X1 U7669 ( .B1(n7196), .B2(n7181), .A(n7180), .ZN(U2950) );
  AOI22_X1 U7670 ( .A1(n7190), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n7185), .ZN(n7182) );
  OAI21_X1 U7671 ( .B1(n7196), .B2(n7184), .A(n7182), .ZN(U2936) );
  AOI22_X1 U7672 ( .A1(n7190), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n7185), .ZN(n7183) );
  OAI21_X1 U7673 ( .B1(n7196), .B2(n7184), .A(n7183), .ZN(U2951) );
  AOI22_X1 U7674 ( .A1(n7190), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n7185), .ZN(n7186) );
  OAI21_X1 U7675 ( .B1(n7196), .B2(n7188), .A(n7186), .ZN(U2937) );
  AOI22_X1 U7676 ( .A1(n7190), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n7185), .ZN(n7187) );
  OAI21_X1 U7677 ( .B1(n7196), .B2(n7188), .A(n7187), .ZN(U2952) );
  AOI22_X1 U7678 ( .A1(n7190), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n7185), .ZN(n7189) );
  OAI21_X1 U7679 ( .B1(n7196), .B2(n7192), .A(n7189), .ZN(U2938) );
  AOI22_X1 U7680 ( .A1(n7190), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n7185), .ZN(n7191) );
  OAI21_X1 U7681 ( .B1(n7196), .B2(n7192), .A(n7191), .ZN(U2953) );
  AOI22_X1 U7682 ( .A1(n7193), .A2(LWORD_REG_15__SCAN_IN), .B1(
        EAX_REG_15__SCAN_IN), .B2(n7185), .ZN(n7194) );
  OAI21_X1 U7683 ( .B1(n7196), .B2(n7195), .A(n7194), .ZN(U2954) );
  AOI22_X1 U7684 ( .A1(n7197), .A2(n7204), .B1(n7203), .B2(DATAI_17_), .ZN(
        n7199) );
  AOI22_X1 U7685 ( .A1(n7207), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7206), .ZN(n7198) );
  NAND2_X1 U7686 ( .A1(n7199), .A2(n7198), .ZN(U2874) );
  AOI22_X1 U7687 ( .A1(n7200), .A2(n7204), .B1(n7203), .B2(DATAI_19_), .ZN(
        n7202) );
  AOI22_X1 U7688 ( .A1(n7207), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n7206), .ZN(n7201) );
  NAND2_X1 U7689 ( .A1(n7202), .A2(n7201), .ZN(U2872) );
  AOI22_X1 U7690 ( .A1(n7205), .A2(n7204), .B1(n7203), .B2(DATAI_21_), .ZN(
        n7209) );
  AOI22_X1 U7691 ( .A1(n7207), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7206), .ZN(n7208) );
  NAND2_X1 U7692 ( .A1(n7209), .A2(n7208), .ZN(U2870) );
  CLKBUF_X1 U3480 ( .A(n4320), .Z(n4151) );
  AND2_X1 U3522 ( .A1(n3776), .A2(n3777), .ZN(n3432) );
  CLKBUF_X1 U3544 ( .A(n6163), .Z(n5836) );
endmodule

