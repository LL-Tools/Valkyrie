

module b20_C_SARLock_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4413, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10253;

  INV_X2 U4918 ( .A(n9452), .ZN(n9455) );
  NAND2_X1 U4919 ( .A1(n6022), .A2(n6021), .ZN(n8527) );
  INV_X1 U4920 ( .A(n5732), .ZN(n6336) );
  INV_X2 U4921 ( .A(n7783), .ZN(n7769) );
  BUF_X2 U4922 ( .A(n6340), .Z(n4419) );
  NAND2_X1 U4924 ( .A1(n6216), .A2(n6215), .ZN(n6617) );
  CLKBUF_X2 U4925 ( .A(n5203), .Z(n7423) );
  INV_X1 U4926 ( .A(n5931), .ZN(n6104) );
  CLKBUF_X1 U4927 ( .A(n5837), .Z(n4413) );
  XNOR2_X1 U4928 ( .A(n6206), .B(n6205), .ZN(n8560) );
  CLKBUF_X2 U4929 ( .A(n5840), .Z(n4416) );
  XNOR2_X1 U4930 ( .A(n5136), .B(n5135), .ZN(n5160) );
  INV_X2 U4931 ( .A(n5837), .ZN(n5869) );
  NAND2_X1 U4932 ( .A1(n8539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4979) );
  INV_X2 U4934 ( .A(n10253), .ZN(P2_U3893) );
  AND2_X1 U4936 ( .A1(n4577), .A2(n4878), .ZN(n4576) );
  AOI21_X1 U4937 ( .B1(n4576), .B2(n4574), .A(n7794), .ZN(n4573) );
  AOI22_X1 U4938 ( .A1(n10182), .A2(keyinput14), .B1(keyinput45), .B2(n10181), 
        .ZN(n10180) );
  OAI221_X1 U4939 ( .B1(n10182), .B2(keyinput14), .C1(n10181), .C2(keyinput45), 
        .A(n10180), .ZN(n10185) );
  OAI22_X1 U4940 ( .A1(n5913), .A2(n5912), .B1(n7070), .B2(n8091), .ZN(n7093)
         );
  NAND2_X1 U4941 ( .A1(n6612), .A2(n7845), .ZN(n7783) );
  INV_X1 U4942 ( .A(n5864), .ZN(n6300) );
  NAND2_X1 U4943 ( .A1(n5826), .A2(n5834), .ZN(n6240) );
  INV_X1 U4944 ( .A(n4419), .ZN(n5662) );
  INV_X1 U4945 ( .A(n5759), .ZN(n5761) );
  AND2_X1 U4946 ( .A1(n7444), .A2(n7443), .ZN(n9111) );
  NOR2_X1 U4947 ( .A1(n6945), .A2(n9446), .ZN(n6943) );
  NAND2_X1 U4948 ( .A1(n6192), .A2(n8145), .ZN(n5845) );
  OR2_X1 U4949 ( .A1(n5259), .A2(n6376), .ZN(n5191) );
  INV_X1 U4950 ( .A(n5232), .ZN(n7420) );
  NOR2_X1 U4951 ( .A1(n8981), .A2(n9146), .ZN(n8963) );
  NAND2_X1 U4952 ( .A1(n5526), .A2(n5525), .ZN(n9187) );
  INV_X1 U4953 ( .A(n9420), .ZN(n9515) );
  OAI21_X1 U4954 ( .B1(n5235), .B2(n4638), .A(n4637), .ZN(n9446) );
  OAI21_X1 U4955 ( .B1(n5523), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5052), .ZN(
        n5053) );
  OAI211_X1 U4956 ( .C1(n7621), .C2(n8128), .A(n5959), .B(n5958), .ZN(n8004)
         );
  AND3_X1 U4957 ( .A1(n5010), .A2(n5008), .A3(n5007), .ZN(n7841) );
  INV_X1 U4958 ( .A(n8158), .ZN(n8151) );
  NOR2_X1 U4959 ( .A1(n6255), .A2(n6256), .ZN(n8272) );
  NAND2_X1 U4960 ( .A1(n6033), .A2(n6032), .ZN(n8522) );
  NAND2_X1 U4961 ( .A1(n7450), .A2(n7539), .ZN(n9062) );
  AOI21_X1 U4962 ( .B1(n9507), .B2(n9141), .A(n9140), .ZN(n9142) );
  XNOR2_X1 U4963 ( .A(n4689), .B(n9221), .ZN(n5147) );
  NAND2_X1 U4964 ( .A1(n5157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  BUF_X1 U4965 ( .A(n5127), .Z(n4418) );
  INV_X1 U4966 ( .A(n9814), .ZN(n7914) );
  NAND2_X1 U4967 ( .A1(n6191), .A2(n6190), .ZN(n8085) );
  XNOR2_X1 U4968 ( .A(n5806), .B(n5805), .ZN(n8547) );
  NAND2_X2 U4969 ( .A1(n6240), .A2(n7630), .ZN(n6239) );
  AOI21_X2 U4970 ( .B1(n7951), .B2(n7952), .A(n7868), .ZN(n7871) );
  NOR2_X1 U4971 ( .A1(n7618), .A2(n5147), .ZN(n5201) );
  XNOR2_X2 U4972 ( .A(n5159), .B(n5158), .ZN(n5549) );
  NAND2_X1 U4973 ( .A1(n5809), .A2(n8547), .ZN(n5837) );
  OAI21_X4 U4975 ( .B1(n6617), .B2(n6616), .A(n6615), .ZN(n6628) );
  AOI21_X2 U4976 ( .B1(n6212), .B2(n8560), .A(n6213), .ZN(n6222) );
  XNOR2_X2 U4977 ( .A(n5133), .B(n5132), .ZN(n5759) );
  AND2_X4 U4978 ( .A1(n7618), .A2(n5147), .ZN(n5248) );
  INV_X4 U4979 ( .A(n5595), .ZN(n6352) );
  BUF_X2 U4981 ( .A(n5840), .Z(n4417) );
  NAND2_X1 U4982 ( .A1(n8543), .A2(n8547), .ZN(n5840) );
  NAND2_X1 U4983 ( .A1(n5033), .A2(n5034), .ZN(n5127) );
  NAND2_X1 U4984 ( .A1(n7464), .A2(n8922), .ZN(n7429) );
  XNOR2_X1 U4985 ( .A(n7320), .B(n7319), .ZN(n7323) );
  NAND2_X1 U4986 ( .A1(n5719), .A2(n5718), .ZN(n6292) );
  INV_X1 U4987 ( .A(n8229), .ZN(n7866) );
  NAND2_X1 U4988 ( .A1(n6913), .A2(n4451), .ZN(n4844) );
  OR2_X1 U4989 ( .A1(n8088), .A2(n9807), .ZN(n7677) );
  INV_X1 U4990 ( .A(n8004), .ZN(n9807) );
  AND3_X1 U4991 ( .A1(n5943), .A2(n5942), .A3(n5941), .ZN(n9804) );
  CLKBUF_X2 U4992 ( .A(n5287), .Z(n6342) );
  NAND4_X1 U4993 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n9759)
         );
  NAND2_X2 U4994 ( .A1(n7512), .A2(n6727), .ZN(n6725) );
  NAND2_X1 U4995 ( .A1(n4674), .A2(n4673), .ZN(n5166) );
  CLKBUF_X2 U4996 ( .A(n5201), .Z(n6416) );
  NOR2_X1 U4997 ( .A1(n4420), .A2(n9232), .ZN(n4673) );
  OAI21_X1 U4999 ( .B1(n6345), .B2(n5764), .A(n8709), .ZN(n5789) );
  NOR2_X1 U5000 ( .A1(n9132), .A2(n4554), .ZN(n4553) );
  NOR2_X1 U5001 ( .A1(n8179), .A2(n6324), .ZN(n6369) );
  INV_X1 U5002 ( .A(n6284), .ZN(n6285) );
  OAI21_X1 U5003 ( .B1(n7557), .B2(n9129), .A(n4607), .ZN(n4706) );
  OR2_X1 U5004 ( .A1(n7883), .A2(n7884), .ZN(n7885) );
  AOI21_X1 U5005 ( .B1(n4732), .B2(n4731), .A(n4733), .ZN(n7505) );
  OAI21_X2 U5006 ( .B1(n8203), .B2(n6164), .A(n6165), .ZN(n6287) );
  NAND2_X1 U5007 ( .A1(n4798), .A2(n4799), .ZN(n8978) );
  NAND2_X1 U5008 ( .A1(n4532), .A2(n4531), .ZN(n8976) );
  OAI21_X1 U5009 ( .B1(n8291), .B2(n4999), .A(n4996), .ZN(n8270) );
  XNOR2_X1 U5010 ( .A(n7323), .B(SI_29_), .ZN(n7566) );
  NAND2_X1 U5011 ( .A1(n4652), .A2(n4423), .ZN(n4651) );
  OAI21_X1 U5012 ( .B1(n8315), .B2(n7724), .A(n7719), .ZN(n8302) );
  NAND2_X1 U5013 ( .A1(n4871), .A2(n4869), .ZN(n7320) );
  XNOR2_X1 U5014 ( .A(n4611), .B(n4872), .ZN(n7849) );
  NAND2_X1 U5015 ( .A1(n8879), .A2(n8880), .ZN(n4547) );
  NAND2_X1 U5016 ( .A1(n6252), .A2(n6251), .ZN(n8315) );
  NAND2_X1 U5017 ( .A1(n6156), .A2(n6155), .ZN(n8457) );
  NAND2_X1 U5018 ( .A1(n7893), .A2(n7894), .ZN(n4834) );
  NAND2_X1 U5019 ( .A1(n5694), .A2(n5693), .ZN(n5717) );
  NOR2_X1 U5020 ( .A1(n7310), .A2(n4552), .ZN(n8873) );
  AOI21_X1 U5021 ( .B1(n4667), .B2(n4671), .A(n4665), .ZN(n4664) );
  AND2_X1 U5022 ( .A1(n4489), .A2(n4668), .ZN(n4667) );
  AND2_X1 U5023 ( .A1(n6095), .A2(n6094), .ZN(n7603) );
  NAND2_X1 U5024 ( .A1(n5573), .A2(n5572), .ZN(n9177) );
  NAND2_X1 U5025 ( .A1(n6103), .A2(n6102), .ZN(n8486) );
  NAND2_X1 U5026 ( .A1(n9397), .A2(n7374), .ZN(n7442) );
  AOI21_X1 U5027 ( .B1(n4915), .B2(n4911), .A(n4910), .ZN(n4909) );
  NAND2_X1 U5028 ( .A1(n6085), .A2(n6084), .ZN(n8498) );
  NAND2_X1 U5029 ( .A1(n7925), .A2(n7578), .ZN(n8000) );
  NAND2_X1 U5030 ( .A1(n7229), .A2(n7227), .ZN(n9396) );
  NAND2_X1 U5031 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  AOI21_X1 U5032 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7690) );
  NAND2_X1 U5033 ( .A1(n6058), .A2(n6057), .ZN(n8509) );
  OR2_X1 U5034 ( .A1(n5570), .A2(n4428), .ZN(n4893) );
  XNOR2_X1 U5035 ( .A(n5570), .B(n5569), .ZN(n7030) );
  OR2_X1 U5036 ( .A1(n5570), .A2(n5569), .ZN(n4903) );
  NAND2_X1 U5037 ( .A1(n7149), .A2(n5945), .ZN(n7253) );
  NAND2_X1 U5038 ( .A1(n4844), .A2(n4842), .ZN(n7193) );
  OR2_X1 U5039 ( .A1(n4487), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U5040 ( .A1(n5443), .A2(n5442), .ZN(n9199) );
  OAI21_X1 U5041 ( .B1(n5461), .B2(n4612), .A(n4885), .ZN(n5496) );
  AOI21_X1 U5042 ( .B1(n4928), .B2(n4677), .A(n4477), .ZN(n4675) );
  NAND2_X1 U5043 ( .A1(n4794), .A2(n7347), .ZN(n4797) );
  NOR2_X1 U5044 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  NAND2_X1 U5045 ( .A1(n5380), .A2(n5379), .ZN(n7283) );
  OR2_X1 U5046 ( .A1(n7035), .A2(n7136), .ZN(n7360) );
  OAI21_X1 U5047 ( .B1(n5373), .B2(n5078), .A(n5081), .ZN(n5392) );
  CLKBUF_X3 U5049 ( .A(n6628), .Z(n7874) );
  INV_X2 U5050 ( .A(n6464), .ZN(n6553) );
  NAND2_X1 U5051 ( .A1(n5063), .A2(n5062), .ZN(n5327) );
  INV_X2 U5052 ( .A(n5732), .ZN(n5711) );
  NAND3_X1 U5053 ( .A1(n5825), .A2(n5824), .A3(n5024), .ZN(n9774) );
  NAND4_X1 U5054 ( .A1(n5228), .A2(n5227), .A3(n5226), .A4(n5225), .ZN(n8738)
         );
  OR2_X1 U5055 ( .A1(n6722), .A2(n5549), .ZN(n6941) );
  NAND2_X1 U5056 ( .A1(n5760), .A2(n5549), .ZN(n7558) );
  NAND2_X1 U5057 ( .A1(n5046), .A2(n5045), .ZN(n5231) );
  NAND4_X1 U5058 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n6709)
         );
  NAND2_X1 U5059 ( .A1(n6203), .A2(n6204), .ZN(n6214) );
  NAND2_X1 U5060 ( .A1(n6204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  XNOR2_X1 U5061 ( .A(n6082), .B(n4854), .ZN(n8164) );
  NAND2_X1 U5062 ( .A1(n6202), .A2(n6201), .ZN(n6204) );
  OR2_X1 U5063 ( .A1(n5230), .A2(n4861), .ZN(n4860) );
  OR2_X2 U5064 ( .A1(n5804), .A2(n5814), .ZN(n5806) );
  NOR2_X1 U5065 ( .A1(n7618), .A2(n7568), .ZN(n5202) );
  NAND2_X1 U5066 ( .A1(n5161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5133) );
  CLKBUF_X1 U5067 ( .A(n6439), .Z(n4421) );
  AND2_X1 U5068 ( .A1(n5818), .A2(n5815), .ZN(n5804) );
  OAI21_X1 U5069 ( .B1(n5161), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  INV_X1 U5070 ( .A(n5744), .ZN(n4420) );
  MUX2_X1 U5071 ( .A(n5144), .B(n5143), .S(P1_IR_REG_30__SCAN_IN), .Z(n7618)
         );
  XNOR2_X1 U5072 ( .A(n5146), .B(n5123), .ZN(n5780) );
  NAND2_X1 U5073 ( .A1(n9220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5146) );
  NOR2_X1 U5074 ( .A1(n5131), .A2(n5130), .ZN(n5134) );
  NAND2_X1 U5075 ( .A1(n5125), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U5076 ( .A(n5137), .B(n4977), .ZN(n9235) );
  NAND2_X1 U5077 ( .A1(n5140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5141) );
  OAI21_X1 U5078 ( .B1(n5047), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4517), .ZN(
        n5043) );
  AND2_X1 U5079 ( .A1(n4686), .A2(n5145), .ZN(n4685) );
  OAI21_X1 U5080 ( .B1(n5465), .B2(n4475), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5137) );
  NOR2_X1 U5081 ( .A1(n5939), .A2(n4856), .ZN(n5975) );
  XNOR2_X1 U5082 ( .A(n5039), .B(SI_1_), .ZN(n5189) );
  INV_X2 U5083 ( .A(n9226), .ZN(n7569) );
  NAND2_X2 U5084 ( .A1(n4418), .A2(P2_U3151), .ZN(n8559) );
  NOR2_X1 U5085 ( .A1(n4684), .A2(n4976), .ZN(n4975) );
  OAI21_X1 U5086 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n10033), .ZN(n5034) );
  AND4_X1 U5087 ( .A1(n4591), .A2(n5908), .A3(n5891), .A4(n4590), .ZN(n4776)
         );
  AND4_X1 U5088 ( .A1(n5135), .A2(n5118), .A3(n5156), .A4(n5158), .ZN(n5119)
         );
  AND2_X1 U5089 ( .A1(n5114), .A2(n5113), .ZN(n4793) );
  INV_X1 U5090 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5156) );
  INV_X1 U5091 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5158) );
  INV_X1 U5092 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5123) );
  NOR2_X1 U5093 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5111) );
  NOR2_X1 U5094 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5112) );
  INV_X1 U5095 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10033) );
  INV_X1 U5096 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5006) );
  INV_X1 U5097 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5891) );
  NOR2_X1 U5098 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6207) );
  INV_X1 U5099 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4590) );
  NOR2_X1 U5100 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4591) );
  INV_X1 U5101 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6205) );
  INV_X4 U5102 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5103 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5795) );
  INV_X1 U5104 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U5105 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5794) );
  NOR2_X1 U5106 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5793) );
  INV_X1 U5107 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n10054) );
  INV_X1 U5108 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5974) );
  OAI22_X1 U5109 ( .A1(n6961), .A2(n5868), .B1(n5867), .B2(n9783), .ZN(n6997)
         );
  OR2_X2 U5110 ( .A1(n6128), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6139) );
  NAND2_X4 U5111 ( .A1(n5780), .A2(n6439), .ZN(n5235) );
  NAND2_X1 U5112 ( .A1(n5166), .A2(n4446), .ZN(n6340) );
  XNOR2_X1 U5113 ( .A(n5126), .B(n5121), .ZN(n6439) );
  INV_X2 U5114 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6964) );
  MUX2_X2 U5115 ( .A(n8085), .B(n8443), .S(n7783), .Z(n7772) );
  OAI22_X2 U5116 ( .A1(n8336), .A2(n6029), .B1(n8342), .B2(n8076), .ZN(n8328)
         );
  INV_X2 U5117 ( .A(n6891), .ZN(n9472) );
  OAI211_X2 U5118 ( .C1(n5235), .C2(n6446), .A(n5214), .B(n5213), .ZN(n6891)
         );
  OR2_X2 U5119 ( .A1(n7623), .A2(n7759), .ZN(n8204) );
  AND2_X2 U5120 ( .A1(n4579), .A2(n4581), .ZN(n4444) );
  AND2_X2 U5121 ( .A1(n7793), .A2(n7795), .ZN(n4581) );
  OAI21_X1 U5122 ( .B1(n7838), .B2(n8173), .A(n7837), .ZN(n5009) );
  NOR2_X2 U5123 ( .A1(n4436), .A2(n6263), .ZN(n4526) );
  AND2_X2 U5124 ( .A1(n4877), .A2(n7769), .ZN(n4436) );
  AND2_X1 U5125 ( .A1(n8861), .A2(n8718), .ZN(n4742) );
  INV_X1 U5126 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5127 ( .A1(n4793), .A2(n4792), .ZN(n4790) );
  OR2_X1 U5128 ( .A1(n8509), .A2(n7963), .ZN(n7721) );
  OR2_X1 U5129 ( .A1(n8515), .A2(n7959), .ZN(n7719) );
  NOR2_X1 U5130 ( .A1(n8894), .A2(n4968), .ZN(n4967) );
  INV_X1 U5131 ( .A(n8893), .ZN(n4968) );
  AOI21_X1 U5132 ( .B1(n8228), .B2(n6145), .A(n6144), .ZN(n8214) );
  AND2_X1 U5133 ( .A1(n4545), .A2(n4543), .ZN(n8891) );
  NAND2_X1 U5134 ( .A1(n4544), .A2(n4441), .ZN(n4543) );
  AND2_X1 U5135 ( .A1(n4975), .A2(n5122), .ZN(n4817) );
  NAND2_X1 U5136 ( .A1(n4593), .A2(n4453), .ZN(n4592) );
  NAND2_X1 U5137 ( .A1(n7666), .A2(n7818), .ZN(n4593) );
  AND2_X1 U5138 ( .A1(n8327), .A2(n7701), .ZN(n4568) );
  OAI21_X1 U5139 ( .B1(n7364), .B2(n4713), .A(n4711), .ZN(n7375) );
  NOR2_X1 U5140 ( .A1(n4714), .A2(n4716), .ZN(n4713) );
  MUX2_X1 U5141 ( .A(n7357), .B(n7356), .S(n9130), .Z(n7364) );
  AOI21_X1 U5142 ( .B1(n7744), .B2(n4585), .A(n4584), .ZN(n4583) );
  AND2_X1 U5143 ( .A1(n7743), .A2(n7742), .ZN(n4585) );
  INV_X1 U5144 ( .A(n7747), .ZN(n4584) );
  NAND2_X1 U5145 ( .A1(n7466), .A2(n7467), .ZN(n4606) );
  NOR2_X1 U5146 ( .A1(n4872), .A2(n4868), .ZN(n4867) );
  INV_X1 U5147 ( .A(n6291), .ZN(n4868) );
  NAND2_X1 U5148 ( .A1(n7759), .A2(n7755), .ZN(n5015) );
  AND2_X1 U5149 ( .A1(n7552), .A2(n7428), .ZN(n4743) );
  INV_X1 U5150 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5095) );
  AND2_X1 U5151 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  AND2_X1 U5152 ( .A1(n5791), .A2(n5003), .ZN(n5002) );
  INV_X1 U5153 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5003) );
  OR2_X1 U5154 ( .A1(n9822), .A2(n8086), .ZN(n7688) );
  NAND2_X1 U5155 ( .A1(n9760), .A2(n9774), .ZN(n7630) );
  NAND2_X1 U5156 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4588) );
  NOR2_X1 U5157 ( .A1(n5818), .A2(n4587), .ZN(n4586) );
  INV_X1 U5158 ( .A(n6210), .ZN(n4589) );
  NAND2_X1 U5159 ( .A1(n7784), .A2(n8164), .ZN(n6613) );
  AND2_X1 U5160 ( .A1(n6258), .A2(n8251), .ZN(n7806) );
  INV_X1 U5161 ( .A(n5022), .ZN(n4747) );
  AOI21_X1 U5162 ( .B1(n4992), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5163 ( .A(n7705), .ZN(n4989) );
  INV_X1 U5164 ( .A(n4993), .ZN(n4990) );
  INV_X1 U5165 ( .A(n4992), .ZN(n4991) );
  INV_X1 U5166 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U5167 ( .A1(n9048), .A2(n4520), .ZN(n8914) );
  AND2_X1 U5168 ( .A1(n9034), .A2(n7543), .ZN(n4520) );
  NOR2_X1 U5169 ( .A1(n7489), .A2(n4953), .ZN(n4952) );
  INV_X1 U5170 ( .A(n4954), .ZN(n4953) );
  NOR2_X1 U5171 ( .A1(n4950), .A2(n7489), .ZN(n4530) );
  NAND2_X1 U5172 ( .A1(n4954), .A2(n4955), .ZN(n4950) );
  AND2_X1 U5173 ( .A1(n4958), .A2(n4454), .ZN(n4956) );
  OR2_X1 U5174 ( .A1(n9264), .A2(n8730), .ZN(n4958) );
  OR2_X1 U5175 ( .A1(n5462), .A2(n4688), .ZN(n4686) );
  AND2_X1 U5176 ( .A1(n5674), .A2(n5651), .ZN(n5672) );
  NAND2_X1 U5177 ( .A1(n4864), .A2(n4862), .ZN(n5544) );
  NOR2_X1 U5178 ( .A1(n4866), .A2(n4863), .ZN(n4862) );
  INV_X1 U5179 ( .A(n5520), .ZN(n4863) );
  AOI22_X1 U5180 ( .A1(n4900), .A2(n4899), .B1(n4901), .B2(n4898), .ZN(n4897)
         );
  INV_X1 U5181 ( .A(n5568), .ZN(n4898) );
  INV_X1 U5182 ( .A(n4902), .ZN(n4899) );
  NAND3_X1 U5183 ( .A1(n5105), .A2(n5104), .A3(n4865), .ZN(n4864) );
  INV_X1 U5184 ( .A(n5521), .ZN(n4865) );
  NOR2_X1 U5185 ( .A1(n4788), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n4678) );
  INV_X1 U5186 ( .A(n4790), .ZN(n4789) );
  INV_X1 U5187 ( .A(n8085), .ZN(n7888) );
  NAND2_X1 U5188 ( .A1(n4846), .A2(n7018), .ZN(n4845) );
  AND2_X1 U5189 ( .A1(n6907), .A2(n9759), .ZN(n6908) );
  AND4_X1 U5190 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n7963)
         );
  AND4_X1 U5191 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n7959)
         );
  INV_X1 U5192 ( .A(n8547), .ZN(n4978) );
  NAND2_X1 U5193 ( .A1(n4627), .A2(n9582), .ZN(n6756) );
  NAND2_X1 U5194 ( .A1(n6760), .A2(n4621), .ZN(n9602) );
  AND2_X1 U5195 ( .A1(n4622), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U5196 ( .A1(n9623), .A2(n5946), .ZN(n9622) );
  AND2_X1 U5197 ( .A1(n6005), .A2(n6004), .ZN(n6019) );
  NOR2_X1 U5198 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6004) );
  AND2_X1 U5199 ( .A1(n7695), .A2(n7696), .ZN(n8364) );
  NAND2_X1 U5200 ( .A1(n5845), .A2(n4418), .ZN(n5865) );
  OR2_X1 U5201 ( .A1(n8451), .A2(n8062), .ZN(n8190) );
  NAND2_X1 U5202 ( .A1(n4426), .A2(n6125), .ZN(n4752) );
  NAND2_X1 U5203 ( .A1(n4753), .A2(n4426), .ZN(n4751) );
  AOI21_X1 U5204 ( .B1(n4998), .B2(n7808), .A(n4997), .ZN(n4996) );
  INV_X1 U5205 ( .A(n7740), .ZN(n4997) );
  AND2_X1 U5206 ( .A1(n7601), .A2(n8307), .ZN(n7809) );
  INV_X1 U5207 ( .A(n5845), .ZN(n6083) );
  INV_X2 U5208 ( .A(n5865), .ZN(n7774) );
  INV_X1 U5209 ( .A(n9762), .ZN(n8355) );
  NAND2_X1 U5210 ( .A1(n5021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U5211 ( .A1(n7333), .A2(n7332), .ZN(n8861) );
  NOR2_X2 U5212 ( .A1(n8981), .A2(n4641), .ZN(n8907) );
  OR2_X1 U5213 ( .A1(n9134), .A2(n4642), .ZN(n4641) );
  AOI21_X1 U5214 ( .B1(n4967), .B2(n4965), .A(n4462), .ZN(n4964) );
  INV_X1 U5215 ( .A(n4440), .ZN(n4965) );
  NAND2_X1 U5216 ( .A1(n9039), .A2(n9030), .ZN(n9024) );
  NAND2_X1 U5217 ( .A1(n4484), .A2(n4422), .ZN(n4549) );
  NAND2_X1 U5218 ( .A1(n4946), .A2(n4424), .ZN(n4945) );
  INV_X1 U5219 ( .A(n4947), .ZN(n4946) );
  AND2_X1 U5220 ( .A1(n9406), .A2(n8727), .ZN(n4552) );
  INV_X1 U5221 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U5222 ( .A1(n5235), .A2(n9237), .ZN(n4637) );
  NAND2_X1 U5223 ( .A1(n4482), .A2(n5463), .ZN(n4976) );
  BUF_X1 U5224 ( .A(n5845), .Z(n7621) );
  INV_X1 U5225 ( .A(n7876), .ZN(n4825) );
  NAND2_X1 U5226 ( .A1(n6814), .A2(n6815), .ZN(n6813) );
  XNOR2_X1 U5227 ( .A(n10218), .B(n4633), .ZN(n4632) );
  INV_X1 U5228 ( .A(n10219), .ZN(n4633) );
  INV_X1 U5229 ( .A(n5549), .ZN(n7508) );
  NAND2_X1 U5230 ( .A1(n7677), .A2(n7682), .ZN(n4525) );
  INV_X1 U5231 ( .A(n7527), .ZN(n4723) );
  NOR2_X1 U5232 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  INV_X1 U5233 ( .A(n7361), .ZN(n4726) );
  NAND2_X1 U5234 ( .A1(n7379), .A2(n7378), .ZN(n4694) );
  NAND2_X1 U5235 ( .A1(n4696), .A2(n9130), .ZN(n4695) );
  INV_X1 U5236 ( .A(n7534), .ZN(n4696) );
  OAI21_X1 U5237 ( .B1(n7371), .B2(n7370), .A(n7445), .ZN(n4691) );
  INV_X1 U5238 ( .A(n7290), .ZN(n4912) );
  NOR2_X1 U5239 ( .A1(n5474), .A2(n4917), .ZN(n4914) );
  INV_X1 U5240 ( .A(n7398), .ZN(n4700) );
  OR2_X1 U5241 ( .A1(n6612), .A2(n7784), .ZN(n6616) );
  NOR2_X1 U5242 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n5802), .ZN(n5803) );
  INV_X1 U5243 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5800) );
  NOR2_X1 U5244 ( .A1(n4929), .A2(n4474), .ZN(n4928) );
  INV_X1 U5245 ( .A(n5317), .ZN(n4929) );
  NAND2_X1 U5246 ( .A1(n8591), .A2(n4907), .ZN(n4906) );
  INV_X1 U5247 ( .A(n5584), .ZN(n4907) );
  AOI21_X1 U5248 ( .B1(n7451), .B2(n4606), .A(n7439), .ZN(n7441) );
  AOI21_X1 U5249 ( .B1(n4902), .B2(n5569), .A(n5585), .ZN(n4900) );
  AOI21_X1 U5250 ( .B1(n5569), .B2(n5568), .A(SI_20_), .ZN(n4901) );
  NOR2_X1 U5251 ( .A1(n5090), .A2(n4883), .ZN(n4882) );
  INV_X1 U5252 ( .A(n5087), .ZN(n4883) );
  OR2_X1 U5253 ( .A1(n6859), .A2(n4449), .ZN(n4522) );
  NAND2_X1 U5254 ( .A1(n8126), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4616) );
  AND2_X1 U5255 ( .A1(n5975), .A2(n5974), .ZN(n6005) );
  NAND2_X1 U5256 ( .A1(n9662), .A2(n4509), .ZN(n8113) );
  NAND2_X1 U5257 ( .A1(n8122), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4509) );
  OAI22_X1 U5258 ( .A1(n9696), .A2(n9695), .B1(n9694), .B2(n8425), .ZN(n8115)
         );
  OAI21_X1 U5259 ( .B1(n8147), .B2(n10040), .A(n9725), .ZN(n8117) );
  INV_X1 U5260 ( .A(n7667), .ZN(n5018) );
  OR2_X1 U5261 ( .A1(n7005), .A2(n5898), .ZN(n5895) );
  AOI21_X1 U5262 ( .B1(n4760), .B2(n4759), .A(n8261), .ZN(n4758) );
  INV_X1 U5263 ( .A(n4767), .ZN(n4759) );
  INV_X1 U5264 ( .A(n8272), .ZN(n4762) );
  OR2_X1 U5265 ( .A1(n8486), .A2(n7853), .ZN(n7742) );
  OR2_X1 U5266 ( .A1(n8498), .A2(n8050), .ZN(n7736) );
  INV_X1 U5267 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U5268 ( .A1(n4850), .A2(n6180), .ZN(n4849) );
  NAND2_X1 U5269 ( .A1(n4852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4850) );
  INV_X1 U5270 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5790) );
  INV_X1 U5271 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10071) );
  AOI21_X1 U5272 ( .B1(n4743), .B2(n4739), .A(n4445), .ZN(n4729) );
  OAI21_X1 U5273 ( .B1(n7414), .B2(n8868), .A(n4740), .ZN(n4739) );
  NAND2_X1 U5274 ( .A1(n4736), .A2(n4742), .ZN(n4734) );
  NAND2_X1 U5275 ( .A1(n9128), .A2(n9130), .ZN(n4737) );
  NAND2_X1 U5276 ( .A1(n4743), .A2(n4741), .ZN(n4730) );
  NOR2_X1 U5277 ( .A1(n8924), .A2(n8868), .ZN(n4741) );
  NAND2_X1 U5278 ( .A1(n8905), .A2(n8868), .ZN(n4738) );
  INV_X1 U5279 ( .A(n4742), .ZN(n4735) );
  OR2_X1 U5280 ( .A1(n9136), .A2(n8926), .ZN(n7465) );
  NAND2_X1 U5281 ( .A1(n9136), .A2(n8926), .ZN(n7464) );
  NOR2_X1 U5282 ( .A1(n4465), .A2(n4534), .ZN(n4533) );
  INV_X1 U5283 ( .A(n4964), .ZN(n4534) );
  INV_X1 U5284 ( .A(n4813), .ZN(n4812) );
  OAI21_X1 U5285 ( .B1(n4815), .B2(n7449), .A(n4814), .ZN(n4813) );
  AOI21_X1 U5286 ( .B1(n4812), .B2(n7449), .A(n4809), .ZN(n4808) );
  AND2_X1 U5287 ( .A1(n9074), .A2(n7537), .ZN(n4815) );
  NOR2_X1 U5288 ( .A1(n4941), .A2(n4938), .ZN(n4937) );
  OR2_X1 U5289 ( .A1(n6888), .A2(n9478), .ZN(n6842) );
  NAND2_X1 U5290 ( .A1(n8873), .A2(n4974), .ZN(n4972) );
  NAND2_X1 U5291 ( .A1(n7337), .A2(n8874), .ZN(n4974) );
  NAND2_X1 U5292 ( .A1(n9276), .A2(n8872), .ZN(n4973) );
  OAI21_X1 U5293 ( .B1(n7323), .B2(n7322), .A(n7321), .ZN(n7417) );
  AND2_X1 U5294 ( .A1(n6293), .A2(n5723), .ZN(n6291) );
  NOR2_X1 U5295 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4683) );
  INV_X1 U5296 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U5297 ( .A1(n5675), .A2(n5674), .ZN(n5692) );
  AND2_X1 U5298 ( .A1(n5693), .A2(n5679), .ZN(n5691) );
  NAND2_X1 U5299 ( .A1(n5544), .A2(n5543), .ZN(n5570) );
  INV_X1 U5300 ( .A(SI_17_), .ZN(n5107) );
  NAND2_X1 U5301 ( .A1(n4888), .A2(n4887), .ZN(n5103) );
  AOI21_X1 U5302 ( .B1(n4890), .B2(n5460), .A(n4433), .ZN(n4887) );
  NAND2_X1 U5303 ( .A1(n4886), .A2(n4613), .ZN(n4885) );
  NAND2_X1 U5304 ( .A1(n4614), .A2(n4613), .ZN(n4612) );
  INV_X1 U5305 ( .A(n4890), .ZN(n4886) );
  INV_X1 U5306 ( .A(SI_15_), .ZN(n5475) );
  INV_X1 U5307 ( .A(SI_14_), .ZN(n5096) );
  AND2_X1 U5308 ( .A1(n5116), .A2(n5463), .ZN(n4934) );
  INV_X1 U5309 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5116) );
  AOI21_X1 U5310 ( .B1(n4539), .B2(n4541), .A(n4537), .ZN(n4536) );
  INV_X1 U5311 ( .A(n5077), .ZN(n4537) );
  NAND2_X1 U5312 ( .A1(n5047), .A2(n6379), .ZN(n5052) );
  OAI21_X1 U5313 ( .B1(n5047), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5048), .ZN(
        n5049) );
  NAND2_X1 U5314 ( .A1(n5047), .A2(n6378), .ZN(n5048) );
  NAND2_X1 U5315 ( .A1(n4841), .A2(n7579), .ZN(n7998) );
  INV_X1 U5316 ( .A(n8000), .ZN(n4841) );
  AND2_X1 U5317 ( .A1(n4845), .A2(n4490), .ZN(n4843) );
  NAND2_X1 U5318 ( .A1(n7792), .A2(n7793), .ZN(n5011) );
  NOR2_X1 U5319 ( .A1(n7800), .A2(n7799), .ZN(n7801) );
  OAI21_X1 U5320 ( .B1(n8434), .B2(n8178), .A(n7798), .ZN(n7799) );
  INV_X1 U5321 ( .A(n7834), .ZN(n7800) );
  AND2_X1 U5322 ( .A1(n5799), .A2(n5002), .ZN(n5001) );
  NOR2_X1 U5323 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  INV_X1 U5324 ( .A(n5900), .ZN(n6303) );
  INV_X2 U5325 ( .A(n4417), .ZN(n6186) );
  OAI21_X1 U5326 ( .B1(n6794), .B2(n6660), .A(n6661), .ZN(n6791) );
  OR2_X1 U5327 ( .A1(n6664), .A2(n6747), .ZN(n4628) );
  INV_X1 U5328 ( .A(n6757), .ZN(n4625) );
  XNOR2_X1 U5329 ( .A(n6753), .B(n4510), .ZN(n9601) );
  NAND2_X1 U5330 ( .A1(n9586), .A2(n6757), .ZN(n4623) );
  AOI21_X1 U5331 ( .B1(n6743), .B2(n9600), .A(n9596), .ZN(n6745) );
  OR2_X1 U5332 ( .A1(n6854), .A2(n6853), .ZN(n4636) );
  NAND2_X1 U5333 ( .A1(n6854), .A2(n6853), .ZN(n6983) );
  OAI22_X1 U5334 ( .A1(n8133), .A2(n8132), .B1(n8131), .B2(n8130), .ZN(n9617)
         );
  OR2_X1 U5335 ( .A1(n9622), .A2(n4486), .ZN(n4619) );
  NAND2_X1 U5336 ( .A1(n4619), .A2(n4618), .ZN(n4617) );
  INV_X1 U5337 ( .A(n9639), .ZN(n4618) );
  XNOR2_X1 U5338 ( .A(n8113), .B(n9679), .ZN(n9681) );
  NAND2_X1 U5339 ( .A1(n9715), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9714) );
  XNOR2_X1 U5340 ( .A(n8117), .B(n8152), .ZN(n9742) );
  NAND2_X1 U5341 ( .A1(n9742), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9741) );
  NOR2_X1 U5342 ( .A1(n5973), .A2(n4780), .ZN(n4779) );
  INV_X1 U5343 ( .A(n5961), .ZN(n4780) );
  NAND2_X1 U5344 ( .A1(n5019), .A2(n7818), .ZN(n7092) );
  INV_X1 U5345 ( .A(n7090), .ZN(n5019) );
  NAND2_X1 U5346 ( .A1(n6302), .A2(n6301), .ZN(n6333) );
  AND2_X1 U5347 ( .A1(n6259), .A2(n7745), .ZN(n4982) );
  AND2_X1 U5348 ( .A1(n6125), .A2(n6124), .ZN(n8250) );
  NAND2_X1 U5349 ( .A1(n6113), .A2(n7853), .ZN(n6114) );
  INV_X1 U5350 ( .A(n4765), .ZN(n4764) );
  OAI22_X1 U5351 ( .A1(n8282), .A2(n4766), .B1(n8050), .B2(n7924), .ZN(n4765)
         );
  INV_X1 U5352 ( .A(n4769), .ZN(n4766) );
  AND2_X1 U5353 ( .A1(n8503), .A2(n8307), .ZN(n4769) );
  AND2_X1 U5354 ( .A1(n7736), .A2(n7740), .ZN(n8282) );
  AND2_X1 U5355 ( .A1(n6074), .A2(n6073), .ZN(n7601) );
  NAND2_X1 U5356 ( .A1(n8302), .A2(n7735), .ZN(n6254) );
  AOI21_X1 U5357 ( .B1(n4745), .B2(n7700), .A(n4470), .ZN(n4744) );
  NAND2_X1 U5358 ( .A1(n4749), .A2(n4750), .ZN(n4748) );
  INV_X2 U5359 ( .A(n8370), .ZN(n9758) );
  OR2_X1 U5360 ( .A1(n7694), .A2(n7693), .ZN(n8359) );
  AND2_X1 U5361 ( .A1(n7695), .A2(n7686), .ZN(n4993) );
  NAND2_X1 U5362 ( .A1(n4481), .A2(n7695), .ZN(n4992) );
  NAND2_X1 U5363 ( .A1(n6248), .A2(n7686), .ZN(n4994) );
  AND2_X1 U5364 ( .A1(n5977), .A2(n5976), .ZN(n9822) );
  AND3_X1 U5365 ( .A1(n5928), .A2(n5927), .A3(n5926), .ZN(n9799) );
  INV_X1 U5366 ( .A(n5802), .ZN(n5817) );
  OR2_X1 U5367 ( .A1(n6199), .A2(n5814), .ZN(n6202) );
  INV_X1 U5368 ( .A(n5005), .ZN(n5004) );
  NAND2_X1 U5369 ( .A1(n5790), .A2(n5006), .ZN(n5005) );
  XNOR2_X1 U5370 ( .A(n5846), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6662) );
  OR2_X1 U5371 ( .A1(n5821), .A2(n5814), .ZN(n5846) );
  INV_X1 U5372 ( .A(n4916), .ZN(n4915) );
  OAI21_X1 U5373 ( .B1(n7290), .B2(n7291), .A(n5459), .ZN(n4916) );
  AND2_X1 U5374 ( .A1(n4682), .A2(n8571), .ZN(n4679) );
  INV_X1 U5375 ( .A(n8675), .ZN(n4681) );
  OAI211_X1 U5376 ( .C1(n4443), .C2(n4662), .A(n5292), .B(n4660), .ZN(n6819)
         );
  AND2_X1 U5377 ( .A1(n6580), .A2(n5272), .ZN(n4661) );
  NAND2_X1 U5378 ( .A1(n6579), .A2(n6580), .ZN(n5244) );
  NAND2_X1 U5379 ( .A1(n4651), .A2(n4464), .ZN(n8664) );
  INV_X1 U5380 ( .A(n8666), .ZN(n4648) );
  NAND2_X1 U5381 ( .A1(n7278), .A2(n5413), .ZN(n4666) );
  AOI21_X1 U5382 ( .B1(n6708), .B2(n6337), .A(n5196), .ZN(n5198) );
  NAND2_X1 U5383 ( .A1(n5549), .A2(n5160), .ZN(n6721) );
  AND2_X1 U5384 ( .A1(n5760), .A2(n5761), .ZN(n7460) );
  AND2_X1 U5385 ( .A1(n7568), .A2(n7618), .ZN(n5203) );
  NOR2_X1 U5386 ( .A1(n9292), .A2(n4503), .ZN(n9312) );
  AND2_X1 U5387 ( .A1(n7460), .A2(n8750), .ZN(n8699) );
  AOI21_X1 U5388 ( .B1(n4962), .B2(n4960), .A(n4479), .ZN(n4959) );
  INV_X1 U5389 ( .A(n4962), .ZN(n4961) );
  INV_X1 U5390 ( .A(n4967), .ZN(n4966) );
  NAND2_X1 U5391 ( .A1(n4805), .A2(n4803), .ZN(n9008) );
  AND2_X1 U5392 ( .A1(n7395), .A2(n8918), .ZN(n9010) );
  OR2_X1 U5393 ( .A1(n9177), .A2(n8888), .ZN(n9034) );
  AND2_X1 U5394 ( .A1(n7543), .A2(n7470), .ZN(n9035) );
  NOR2_X1 U5395 ( .A1(n4943), .A2(n4551), .ZN(n4546) );
  NAND2_X1 U5396 ( .A1(n4424), .A2(n4422), .ZN(n4943) );
  NOR2_X1 U5397 ( .A1(n8887), .A2(n4948), .ZN(n4947) );
  INV_X1 U5398 ( .A(n8883), .ZN(n4948) );
  INV_X1 U5399 ( .A(n4815), .ZN(n4811) );
  OR2_X1 U5400 ( .A1(n9187), .A2(n8882), .ZN(n8883) );
  OR2_X1 U5401 ( .A1(n9199), .A2(n8728), .ZN(n7307) );
  NAND2_X1 U5402 ( .A1(n5420), .A2(n5419), .ZN(n7221) );
  AOI21_X1 U5403 ( .B1(n4956), .B2(n7484), .A(n7175), .ZN(n4954) );
  INV_X1 U5404 ( .A(n4956), .ZN(n4955) );
  AND2_X1 U5405 ( .A1(n7367), .A2(n7526), .ZN(n7489) );
  INV_X1 U5406 ( .A(n6919), .ZN(n4794) );
  NAND2_X1 U5407 ( .A1(n7351), .A2(n7348), .ZN(n7480) );
  NAND2_X1 U5408 ( .A1(n9472), .A2(n6943), .ZN(n6888) );
  XNOR2_X1 U5409 ( .A(n8739), .B(n9472), .ZN(n6883) );
  INV_X1 U5410 ( .A(n9101), .ZN(n9436) );
  INV_X1 U5411 ( .A(n4785), .ZN(n4783) );
  INV_X1 U5412 ( .A(n6725), .ZN(n4784) );
  NAND2_X1 U5413 ( .A1(n6725), .A2(n4785), .ZN(n6934) );
  NAND2_X1 U5414 ( .A1(n5759), .A2(n7563), .ZN(n6723) );
  NAND2_X1 U5415 ( .A1(n5653), .A2(n5652), .ZN(n9157) );
  NAND2_X1 U5416 ( .A1(n5628), .A2(n5627), .ZN(n9161) );
  NAND2_X1 U5417 ( .A1(n5590), .A2(n5589), .ZN(n9172) );
  NAND2_X1 U5418 ( .A1(n9445), .A2(n6721), .ZN(n9544) );
  NAND2_X1 U5419 ( .A1(n9415), .A2(n9509), .ZN(n9541) );
  NAND2_X1 U5420 ( .A1(n6407), .A2(n5758), .ZN(n7559) );
  AND2_X1 U5421 ( .A1(n5166), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5758) );
  OR2_X1 U5422 ( .A1(n7417), .A2(n7416), .ZN(n7419) );
  NAND2_X1 U5423 ( .A1(n4687), .A2(n4685), .ZN(n4689) );
  OR2_X1 U5424 ( .A1(n4817), .A2(n4688), .ZN(n4687) );
  XNOR2_X1 U5425 ( .A(n5138), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U5426 ( .A1(n4596), .A2(n4597), .ZN(n5645) );
  AOI21_X1 U5427 ( .B1(n4425), .B2(n4896), .A(n4598), .ZN(n4597) );
  INV_X1 U5428 ( .A(n5619), .ZN(n4598) );
  AND2_X1 U5429 ( .A1(n5646), .A2(n5626), .ZN(n5644) );
  NAND2_X1 U5430 ( .A1(n4600), .A2(n4602), .ZN(n5621) );
  NAND2_X1 U5431 ( .A1(n4601), .A2(n4895), .ZN(n4600) );
  INV_X1 U5432 ( .A(n5544), .ZN(n4601) );
  INV_X1 U5433 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5132) );
  INV_X1 U5434 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5135) );
  INV_X1 U5435 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U5436 ( .A1(n5112), .A2(n5111), .ZN(n4788) );
  NOR2_X1 U5437 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5113) );
  XNOR2_X1 U5438 ( .A(n5043), .B(SI_2_), .ZN(n5212) );
  AND2_X1 U5439 ( .A1(n6167), .A2(n6166), .ZN(n7892) );
  INV_X1 U5440 ( .A(n7891), .ZN(n4514) );
  OR2_X1 U5441 ( .A1(n7591), .A2(n8337), .ZN(n4516) );
  NAND2_X1 U5442 ( .A1(n4829), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U5443 ( .A1(n7878), .A2(n7876), .ZN(n4829) );
  OR2_X1 U5444 ( .A1(n7878), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U5445 ( .A1(n7878), .A2(n4831), .ZN(n4830) );
  INV_X1 U5446 ( .A(n7884), .ZN(n4831) );
  AND2_X1 U5447 ( .A1(n6618), .A2(n9760), .ZN(n6619) );
  INV_X1 U5448 ( .A(n8251), .ZN(n8028) );
  NAND2_X1 U5449 ( .A1(n6605), .A2(n8373), .ZN(n8064) );
  INV_X1 U5450 ( .A(n7984), .ZN(n8239) );
  INV_X1 U5451 ( .A(n7975), .ZN(n8307) );
  INV_X1 U5452 ( .A(n7959), .ZN(n8329) );
  OR2_X1 U5453 ( .A1(n4413), .A2(n5838), .ZN(n5843) );
  NAND2_X1 U5454 ( .A1(n6798), .A2(n4519), .ZN(n6815) );
  OR2_X1 U5455 ( .A1(n6641), .A2(n6642), .ZN(n4519) );
  AND2_X1 U5456 ( .A1(n8105), .A2(n9743), .ZN(n10218) );
  OR2_X1 U5457 ( .A1(n6667), .A2(n8151), .ZN(n10220) );
  AND2_X1 U5458 ( .A1(n6870), .A2(n8151), .ZN(n10223) );
  NAND2_X1 U5459 ( .A1(n8376), .A2(n6267), .ZN(n8381) );
  NAND2_X1 U5460 ( .A1(n4594), .A2(n5866), .ZN(n6965) );
  INV_X1 U5461 ( .A(n4595), .ZN(n4594) );
  OAI22_X1 U5462 ( .A1(n5864), .A2(n10034), .B1(n7621), .B2(n6747), .ZN(n4595)
         );
  OR2_X1 U5463 ( .A1(n5864), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5824) );
  OR2_X1 U5464 ( .A1(n5865), .A2(n5819), .ZN(n5825) );
  INV_X2 U5465 ( .A(n9773), .ZN(n8376) );
  AOI21_X1 U5466 ( .B1(n6198), .B2(n8355), .A(n6197), .ZN(n8447) );
  NAND2_X1 U5467 ( .A1(n8215), .A2(n8352), .ZN(n6195) );
  INV_X1 U5468 ( .A(n6333), .ZN(n8181) );
  NOR2_X1 U5469 ( .A1(n8187), .A2(n9808), .ZN(n6324) );
  INV_X1 U5470 ( .A(n7892), .ZN(n8451) );
  OR2_X1 U5471 ( .A1(n6071), .A2(n4851), .ZN(n6177) );
  NAND2_X1 U5472 ( .A1(n4855), .A2(n10054), .ZN(n4851) );
  NAND2_X1 U5473 ( .A1(n5396), .A2(n5395), .ZN(n9264) );
  INV_X1 U5474 ( .A(n7510), .ZN(n4704) );
  AND2_X1 U5475 ( .A1(n4710), .A2(n7509), .ZN(n4708) );
  INV_X1 U5476 ( .A(n7557), .ZN(n4710) );
  NAND2_X1 U5477 ( .A1(n4706), .A2(n4709), .ZN(n4705) );
  INV_X1 U5478 ( .A(n7562), .ZN(n4607) );
  INV_X1 U5479 ( .A(n8934), .ZN(n8908) );
  NAND2_X1 U5480 ( .A1(n4820), .A2(n4818), .ZN(n9132) );
  AOI21_X1 U5481 ( .B1(n8720), .B2(n8699), .A(n4819), .ZN(n4818) );
  NAND2_X1 U5482 ( .A1(n4821), .A2(n9459), .ZN(n4820) );
  NOR2_X1 U5483 ( .A1(n8928), .A2(n8929), .ZN(n4819) );
  OAI211_X1 U5484 ( .C1(n5235), .C2(n8783), .A(n5261), .B(n5260), .ZN(n9432)
         );
  OR2_X1 U5485 ( .A1(n5232), .A2(n6383), .ZN(n5261) );
  INV_X1 U5486 ( .A(n9478), .ZN(n6829) );
  OAI211_X1 U5487 ( .C1(n7669), .C2(n7783), .A(n7674), .B(n4592), .ZN(n7681)
         );
  AOI21_X1 U5488 ( .B1(n7674), .B2(n4458), .A(n4525), .ZN(n7679) );
  AOI21_X1 U5489 ( .B1(n4723), .B2(n4720), .A(n4727), .ZN(n4719) );
  OR2_X1 U5490 ( .A1(n7365), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U5491 ( .A1(n4728), .A2(n7363), .ZN(n4721) );
  AOI21_X1 U5492 ( .B1(n4725), .B2(n4431), .A(n7226), .ZN(n4717) );
  AND2_X1 U5493 ( .A1(n7717), .A2(n7718), .ZN(n4566) );
  NAND2_X1 U5494 ( .A1(n4569), .A2(n4568), .ZN(n4567) );
  INV_X1 U5495 ( .A(n4717), .ZN(n4712) );
  INV_X1 U5496 ( .A(n4719), .ZN(n4715) );
  AOI21_X1 U5497 ( .B1(n4719), .B2(n4722), .A(n4724), .ZN(n4714) );
  NAND2_X1 U5498 ( .A1(n4723), .A2(n7521), .ZN(n4722) );
  AOI21_X1 U5499 ( .B1(n4717), .B2(n4718), .A(n9130), .ZN(n4716) );
  NAND2_X1 U5500 ( .A1(n4725), .A2(n7358), .ZN(n4718) );
  INV_X1 U5501 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U5502 ( .A1(n4691), .A2(n4724), .ZN(n4690) );
  OAI21_X1 U5503 ( .B1(n7377), .B2(n4695), .A(n4694), .ZN(n4693) );
  NAND2_X1 U5504 ( .A1(n4444), .A2(n4432), .ZN(n4577) );
  INV_X1 U5505 ( .A(n4444), .ZN(n4574) );
  NOR2_X1 U5506 ( .A1(n4605), .A2(n7429), .ZN(n7451) );
  NOR2_X1 U5507 ( .A1(n4606), .A2(n7438), .ZN(n4605) );
  INV_X1 U5508 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U5509 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4587) );
  OR2_X1 U5510 ( .A1(n6409), .A2(n6233), .ZN(n6584) );
  NAND2_X1 U5511 ( .A1(n5413), .A2(n5414), .ZN(n4672) );
  INV_X1 U5512 ( .A(n4914), .ZN(n4913) );
  NAND2_X1 U5513 ( .A1(n4670), .A2(n4669), .ZN(n4668) );
  INV_X1 U5514 ( .A(n5413), .ZN(n4669) );
  INV_X1 U5515 ( .A(n4909), .ZN(n4665) );
  NOR2_X1 U5516 ( .A1(n8563), .A2(n4918), .ZN(n4910) );
  NOR2_X1 U5517 ( .A1(n4914), .A2(n4912), .ZN(n4911) );
  OR2_X1 U5518 ( .A1(n7429), .A2(n7403), .ZN(n7407) );
  NOR2_X1 U5519 ( .A1(n7429), .A2(n4698), .ZN(n4697) );
  AOI21_X1 U5520 ( .B1(n7393), .B2(n4455), .A(n4700), .ZN(n4699) );
  NAND2_X1 U5521 ( .A1(n7466), .A2(n4429), .ZN(n4698) );
  NAND2_X1 U5522 ( .A1(n7360), .A2(n7340), .ZN(n7038) );
  AOI21_X1 U5523 ( .B1(n4870), .B2(n6297), .A(n4505), .ZN(n4869) );
  NAND2_X1 U5524 ( .A1(n6292), .A2(n4867), .ZN(n4871) );
  INV_X1 U5525 ( .A(n5603), .ZN(n5604) );
  AND2_X1 U5526 ( .A1(n5568), .A2(SI_20_), .ZN(n4902) );
  INV_X1 U5527 ( .A(n5460), .ZN(n4614) );
  AND2_X1 U5528 ( .A1(n4891), .A2(n5100), .ZN(n4890) );
  NAND2_X1 U5529 ( .A1(n5101), .A2(n5475), .ZN(n4891) );
  INV_X1 U5530 ( .A(n6616), .ZN(n7835) );
  NAND2_X1 U5531 ( .A1(n4628), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5532 ( .A1(n9578), .A2(n4461), .ZN(n6753) );
  OAI21_X1 U5533 ( .B1(n8108), .B2(n6973), .A(n8107), .ZN(n8109) );
  OAI21_X1 U5534 ( .B1(n9629), .B2(n5963), .A(n9630), .ZN(n8111) );
  AOI21_X1 U5535 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8122), .A(n9671), .ZN(
        n8099) );
  INV_X1 U5536 ( .A(SI_28_), .ZN(n9965) );
  AOI21_X1 U5537 ( .B1(n5013), .B2(n7623), .A(n4471), .ZN(n5012) );
  NAND2_X1 U5538 ( .A1(n6087), .A2(n6086), .ZN(n6096) );
  INV_X1 U5539 ( .A(n6088), .ZN(n6087) );
  OR2_X1 U5540 ( .A1(n8093), .A2(n6910), .ZN(n7007) );
  OR2_X1 U5541 ( .A1(n9759), .A2(n9783), .ZN(n7646) );
  INV_X1 U5542 ( .A(n6239), .ZN(n7634) );
  INV_X1 U5543 ( .A(n6287), .ZN(n6288) );
  AND2_X1 U5544 ( .A1(n8457), .A2(n7955), .ZN(n7759) );
  INV_X1 U5545 ( .A(n7806), .ZN(n6259) );
  OR2_X1 U5546 ( .A1(n8468), .A2(n7984), .ZN(n7804) );
  NOR2_X1 U5547 ( .A1(n8282), .A2(n4768), .ZN(n4767) );
  INV_X1 U5548 ( .A(n6081), .ZN(n4768) );
  AND2_X1 U5549 ( .A1(n8492), .A2(n7920), .ZN(n6256) );
  NAND2_X1 U5550 ( .A1(n5930), .A2(n4777), .ZN(n7149) );
  INV_X1 U5551 ( .A(n7817), .ZN(n5944) );
  AND2_X1 U5552 ( .A1(n4457), .A2(n5800), .ZN(n4781) );
  NAND2_X1 U5553 ( .A1(n6207), .A2(n5801), .ZN(n5802) );
  INV_X1 U5554 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5801) );
  INV_X1 U5555 ( .A(n6875), .ZN(n4677) );
  AOI22_X1 U5556 ( .A1(n6709), .A2(n5167), .B1(n5192), .B2(n9446), .ZN(n5182)
         );
  INV_X1 U5557 ( .A(n4658), .ZN(n4656) );
  OAI21_X1 U5558 ( .B1(n8664), .B2(n4908), .A(n4905), .ZN(n5617) );
  INV_X1 U5559 ( .A(n8591), .ZN(n4908) );
  AND2_X1 U5560 ( .A1(n4906), .A2(n5602), .ZN(n4905) );
  INV_X1 U5561 ( .A(n9449), .ZN(n4609) );
  NOR2_X1 U5562 ( .A1(n9341), .A2(n4561), .ZN(n8823) );
  NOR2_X1 U5563 ( .A1(n4563), .A2(n4562), .ZN(n4561) );
  INV_X1 U5564 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n4562) );
  INV_X1 U5565 ( .A(n9346), .ZN(n4563) );
  OR2_X1 U5566 ( .A1(n8952), .A2(n8904), .ZN(n8922) );
  NAND2_X1 U5567 ( .A1(n4644), .A2(n4643), .ZN(n4642) );
  INV_X1 U5568 ( .A(n4645), .ZN(n4644) );
  AND2_X1 U5569 ( .A1(n8903), .A2(n4963), .ZN(n4962) );
  NAND2_X1 U5570 ( .A1(n8900), .A2(n8902), .ZN(n4963) );
  INV_X1 U5571 ( .A(n8902), .ZN(n4960) );
  NAND2_X1 U5572 ( .A1(n8952), .A2(n8966), .ZN(n4645) );
  OR2_X1 U5573 ( .A1(n9146), .A2(n8901), .ZN(n7467) );
  INV_X1 U5574 ( .A(n4549), .ZN(n4544) );
  NOR2_X1 U5575 ( .A1(n7337), .A2(n9406), .ZN(n4640) );
  NAND2_X1 U5576 ( .A1(n9396), .A2(n7302), .ZN(n9397) );
  NOR2_X1 U5577 ( .A1(n7033), .A2(n4796), .ZN(n4795) );
  INV_X1 U5578 ( .A(n7345), .ZN(n4796) );
  NOR2_X1 U5579 ( .A1(n9422), .A2(n7136), .ZN(n7057) );
  AND2_X1 U5580 ( .A1(n5718), .A2(n5698), .ZN(n5716) );
  INV_X1 U5581 ( .A(n5620), .ZN(n4599) );
  AND2_X1 U5582 ( .A1(n4894), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5583 ( .A1(n4895), .A2(n4604), .ZN(n4603) );
  AOI21_X1 U5584 ( .B1(n4895), .B2(n4428), .A(n4498), .ZN(n4894) );
  INV_X1 U5585 ( .A(n5543), .ZN(n4604) );
  NAND2_X1 U5586 ( .A1(n4934), .A2(n4933), .ZN(n4932) );
  NOR2_X1 U5587 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4933) );
  INV_X1 U5588 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4647) );
  AOI21_X1 U5589 ( .B1(n4882), .B2(n5391), .A(n4435), .ZN(n4881) );
  OR2_X1 U5590 ( .A1(n5344), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5377) );
  INV_X1 U5591 ( .A(n4792), .ZN(n5253) );
  NAND2_X1 U5592 ( .A1(n5047), .A2(n6373), .ZN(n4517) );
  INV_X1 U5593 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5031) );
  AND2_X1 U5594 ( .A1(n7884), .A2(n7876), .ZN(n4828) );
  AND2_X1 U5595 ( .A1(n7860), .A2(n7858), .ZN(n4847) );
  INV_X1 U5596 ( .A(n7861), .ZN(n7982) );
  NAND2_X1 U5597 ( .A1(n8024), .A2(n7858), .ZN(n7981) );
  NAND2_X1 U5598 ( .A1(n6913), .A2(n6912), .ZN(n7021) );
  INV_X1 U5599 ( .A(n7581), .ZN(n4840) );
  NAND2_X1 U5600 ( .A1(n7998), .A2(n7581), .ZN(n7940) );
  INV_X1 U5601 ( .A(n8351), .ZN(n8076) );
  NAND2_X1 U5602 ( .A1(n4620), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6793) );
  INV_X1 U5603 ( .A(n6791), .ZN(n4620) );
  NAND2_X1 U5604 ( .A1(n4524), .A2(n4523), .ZN(n6807) );
  OR2_X1 U5605 ( .A1(n6662), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U5606 ( .A1(n6662), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5607 ( .A1(n6806), .A2(n6807), .ZN(n6805) );
  NAND2_X1 U5608 ( .A1(n6793), .A2(n6661), .ZN(n6803) );
  NAND2_X1 U5609 ( .A1(n4626), .A2(n9582), .ZN(n9584) );
  INV_X1 U5610 ( .A(n4627), .ZN(n4626) );
  XNOR2_X1 U5611 ( .A(n6748), .B(n6741), .ZN(n6746) );
  XNOR2_X1 U5612 ( .A(n4522), .B(n6853), .ZN(n6977) );
  NAND2_X1 U5613 ( .A1(n6853), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5614 ( .A1(n6977), .A2(n6976), .B1(n6975), .B2(n6974), .ZN(n6978)
         );
  INV_X1 U5615 ( .A(n4522), .ZN(n6974) );
  NAND2_X1 U5616 ( .A1(n6978), .A2(n6979), .ZN(n8107) );
  INV_X1 U5617 ( .A(n5002), .ZN(n4856) );
  XNOR2_X1 U5618 ( .A(n8111), .B(n9646), .ZN(n9648) );
  NOR2_X1 U5619 ( .A1(n8097), .A2(n9654), .ZN(n9673) );
  AND2_X1 U5620 ( .A1(n8114), .A2(n9680), .ZN(n9696) );
  NAND2_X1 U5621 ( .A1(n9714), .A2(n8103), .ZN(n9731) );
  NAND2_X1 U5622 ( .A1(n9731), .A2(n9732), .ZN(n9730) );
  NAND2_X1 U5623 ( .A1(n9741), .A2(n8118), .ZN(n10204) );
  NAND2_X1 U5624 ( .A1(n9730), .A2(n4615), .ZN(n8104) );
  NAND2_X1 U5625 ( .A1(n9738), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5626 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  OR2_X1 U5627 ( .A1(n4580), .A2(n7888), .ZN(n5025) );
  NAND2_X1 U5628 ( .A1(n6138), .A2(n6137), .ZN(n6150) );
  INV_X1 U5629 ( .A(n6139), .ZN(n6138) );
  OR2_X1 U5630 ( .A1(n6117), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6128) );
  OR2_X1 U5631 ( .A1(n6096), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U5632 ( .A1(n6105), .A2(n10107), .ZN(n6117) );
  INV_X1 U5633 ( .A(n6106), .ZN(n6105) );
  NAND2_X1 U5634 ( .A1(n6060), .A2(n6059), .ZN(n6075) );
  INV_X1 U5635 ( .A(n6061), .ZN(n6060) );
  INV_X1 U5636 ( .A(n6036), .ZN(n6035) );
  OR2_X1 U5637 ( .A1(n6048), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6061) );
  INV_X1 U5638 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U5639 ( .A1(n7769), .A2(n6194), .ZN(n8370) );
  OR2_X1 U5640 ( .A1(n5980), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5995) );
  OR2_X1 U5641 ( .A1(n5964), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5980) );
  AOI21_X1 U5642 ( .B1(n7090), .B2(n5016), .A(n5017), .ZN(n7252) );
  INV_X1 U5643 ( .A(n4442), .ZN(n5016) );
  NAND2_X1 U5644 ( .A1(n7819), .A2(n7252), .ZN(n7246) );
  OR2_X1 U5645 ( .A1(n5932), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5950) );
  OR2_X1 U5646 ( .A1(n5901), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5917) );
  AND2_X1 U5647 ( .A1(n7661), .A2(n7652), .ZN(n7815) );
  CLKBUF_X1 U5648 ( .A(n6997), .Z(n7006) );
  AND2_X1 U5649 ( .A1(n7657), .A2(n7648), .ZN(n7810) );
  INV_X1 U5650 ( .A(n6241), .ZN(n9757) );
  AND3_X1 U5651 ( .A1(n5849), .A2(n5848), .A3(n5847), .ZN(n9766) );
  NAND2_X1 U5652 ( .A1(n7634), .A2(n4980), .ZN(n6896) );
  INV_X1 U5653 ( .A(n7627), .ZN(n4980) );
  AND2_X1 U5654 ( .A1(n6265), .A2(n6674), .ZN(n9765) );
  AND2_X1 U5655 ( .A1(n7796), .A2(n6325), .ZN(n9762) );
  OR2_X1 U5656 ( .A1(n7783), .A2(n6613), .ZN(n6674) );
  AND2_X1 U5657 ( .A1(n8173), .A2(n8172), .ZN(n8435) );
  AND2_X1 U5658 ( .A1(n7624), .A2(n7760), .ZN(n8213) );
  INV_X1 U5659 ( .A(n8213), .ZN(n8211) );
  AND2_X1 U5660 ( .A1(n7804), .A2(n7803), .ZN(n8227) );
  NAND2_X1 U5661 ( .A1(n8246), .A2(n8245), .ZN(n4983) );
  INV_X1 U5662 ( .A(n8250), .ZN(n8245) );
  NAND2_X1 U5663 ( .A1(n4757), .A2(n4755), .ZN(n8263) );
  AOI21_X1 U5664 ( .B1(n4758), .B2(n4761), .A(n4756), .ZN(n4755) );
  INV_X1 U5665 ( .A(n8260), .ZN(n4756) );
  INV_X1 U5666 ( .A(n6256), .ZN(n8257) );
  NAND2_X1 U5667 ( .A1(n8270), .A2(n7743), .ZN(n8258) );
  NAND2_X1 U5668 ( .A1(n8293), .A2(n4767), .ZN(n4763) );
  NOR2_X1 U5669 ( .A1(n7693), .A2(n4772), .ZN(n4771) );
  INV_X1 U5670 ( .A(n6002), .ZN(n4772) );
  AND2_X1 U5671 ( .A1(n7703), .A2(n7702), .ZN(n8346) );
  AOI21_X1 U5672 ( .B1(n4988), .B2(n4991), .A(n4986), .ZN(n4985) );
  INV_X1 U5673 ( .A(n7704), .ZN(n4986) );
  INV_X1 U5674 ( .A(n9794), .ZN(n9808) );
  INV_X1 U5675 ( .A(n6965), .ZN(n9783) );
  NOR2_X1 U5676 ( .A1(n6594), .A2(n6593), .ZN(n6607) );
  AND2_X1 U5677 ( .A1(n6585), .A2(n6330), .ZN(n6604) );
  NAND2_X1 U5678 ( .A1(n7172), .A2(n7274), .ZN(n9821) );
  AND2_X1 U5679 ( .A1(n6590), .A2(n6597), .ZN(n6410) );
  INV_X1 U5680 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5805) );
  INV_X1 U5681 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6201) );
  AOI21_X1 U5682 ( .B1(n6071), .B2(P2_IR_REG_31__SCAN_IN), .A(n4849), .ZN(
        n4848) );
  NAND2_X1 U5683 ( .A1(n4855), .A2(n4853), .ZN(n4852) );
  AND2_X1 U5684 ( .A1(n10054), .A2(n4854), .ZN(n4853) );
  INV_X1 U5685 ( .A(n5028), .ZN(n4855) );
  INV_X1 U5686 ( .A(n5655), .ZN(n5654) );
  NOR2_X1 U5687 ( .A1(n4922), .A2(n4659), .ZN(n4658) );
  INV_X1 U5688 ( .A(n8625), .ZN(n4659) );
  NAND2_X1 U5689 ( .A1(n4925), .A2(n4924), .ZN(n4922) );
  OR2_X1 U5690 ( .A1(n4927), .A2(n4926), .ZN(n4923) );
  INV_X1 U5691 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8584) );
  OR2_X1 U5692 ( .A1(n5318), .A2(n6956), .ZN(n5337) );
  NAND2_X1 U5693 ( .A1(n8624), .A2(n8625), .ZN(n8633) );
  AND2_X1 U5694 ( .A1(n5502), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5504) );
  INV_X1 U5695 ( .A(n8655), .ZN(n4920) );
  INV_X1 U5696 ( .A(n8738), .ZN(n8659) );
  OR2_X1 U5697 ( .A1(n5337), .A2(n5336), .ZN(n5358) );
  NOR2_X1 U5698 ( .A1(n5358), .A2(n9975), .ZN(n5381) );
  OR2_X1 U5699 ( .A1(n5554), .A2(n8584), .ZN(n5574) );
  NAND2_X1 U5700 ( .A1(n4650), .A2(n4495), .ZN(n4649) );
  INV_X1 U5701 ( .A(n4654), .ZN(n4650) );
  AOI21_X1 U5702 ( .B1(n4657), .B2(n4656), .A(n4655), .ZN(n4654) );
  INV_X1 U5703 ( .A(n8580), .ZN(n4655) );
  INV_X1 U5704 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8668) );
  INV_X1 U5705 ( .A(n5167), .ZN(n5732) );
  OR2_X1 U5706 ( .A1(n5397), .A2(n10006), .ZN(n5422) );
  NOR2_X1 U5707 ( .A1(n5491), .A2(n5490), .ZN(n8708) );
  NAND2_X1 U5708 ( .A1(n4483), .A2(n4730), .ZN(n4732) );
  INV_X1 U5709 ( .A(n7463), .ZN(n7504) );
  NOR2_X1 U5710 ( .A1(n7506), .A2(n7508), .ZN(n7503) );
  NAND2_X1 U5711 ( .A1(n4610), .A2(n4608), .ZN(n7557) );
  NAND2_X1 U5712 ( .A1(n7555), .A2(n7556), .ZN(n4610) );
  OR2_X1 U5713 ( .A1(n7555), .A2(n4609), .ZN(n4608) );
  AND2_X1 U5714 ( .A1(n5472), .A2(n5471), .ZN(n7309) );
  NOR2_X1 U5715 ( .A1(n6500), .A2(n4558), .ZN(n6436) );
  NOR2_X1 U5716 ( .A1(n6509), .A2(n7118), .ZN(n4558) );
  NOR2_X1 U5717 ( .A1(n6519), .A2(n4557), .ZN(n6521) );
  AND2_X1 U5718 ( .A1(n6520), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U5719 ( .A1(n6521), .A2(n6522), .ZN(n8817) );
  NOR2_X1 U5720 ( .A1(n9243), .A2(n4559), .ZN(n9294) );
  AND2_X1 U5721 ( .A1(n8819), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4559) );
  NOR2_X1 U5722 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  NAND2_X1 U5723 ( .A1(n9312), .A2(n9313), .ZN(n9311) );
  NOR2_X1 U5724 ( .A1(n9326), .A2(n4504), .ZN(n9343) );
  NOR2_X1 U5725 ( .A1(n9343), .A2(n9342), .ZN(n9341) );
  XNOR2_X1 U5726 ( .A(n8823), .B(n9359), .ZN(n9355) );
  NOR2_X1 U5727 ( .A1(n9369), .A2(n4556), .ZN(n8827) );
  AND2_X1 U5728 ( .A1(n8826), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4556) );
  NAND2_X1 U5729 ( .A1(n8827), .A2(n8828), .ZN(n8837) );
  AND2_X1 U5730 ( .A1(n8837), .A2(n8836), .ZN(n9384) );
  NAND2_X1 U5731 ( .A1(n9384), .A2(n9385), .ZN(n9382) );
  XNOR2_X1 U5732 ( .A(n8925), .B(n8905), .ZN(n4821) );
  INV_X1 U5733 ( .A(n8923), .ZN(n8939) );
  NAND2_X1 U5734 ( .A1(n8954), .A2(n8955), .ZN(n8953) );
  INV_X1 U5735 ( .A(n8903), .ZN(n8955) );
  AOI21_X1 U5736 ( .B1(n4801), .B2(n4804), .A(n4800), .ZN(n4799) );
  INV_X1 U5737 ( .A(n8919), .ZN(n4800) );
  AND2_X1 U5738 ( .A1(n7469), .A2(n7468), .ZN(n8977) );
  AOI21_X1 U5739 ( .B1(n4533), .B2(n4966), .A(n4496), .ZN(n4531) );
  NAND2_X1 U5740 ( .A1(n4807), .A2(n4521), .ZN(n9048) );
  AND2_X1 U5741 ( .A1(n4806), .A2(n4808), .ZN(n4521) );
  NAND2_X1 U5742 ( .A1(n4812), .A2(n9093), .ZN(n4806) );
  OR2_X1 U5743 ( .A1(n5527), .A2(n8687), .ZN(n5554) );
  NAND2_X1 U5744 ( .A1(n9408), .A2(n4640), .ZN(n9102) );
  NAND2_X1 U5745 ( .A1(n9408), .A2(n9545), .ZN(n9407) );
  OR2_X1 U5746 ( .A1(n5469), .A2(n8565), .ZN(n5483) );
  NOR2_X1 U5747 ( .A1(n5422), .A2(n5421), .ZN(n5444) );
  NAND2_X1 U5748 ( .A1(n4951), .A2(n4528), .ZN(n7224) );
  NOR2_X1 U5749 ( .A1(n4530), .A2(n4529), .ZN(n4528) );
  NOR2_X1 U5750 ( .A1(n7221), .A2(n8729), .ZN(n4529) );
  NAND2_X1 U5751 ( .A1(n7057), .A2(n9527), .ZN(n7081) );
  AOI21_X1 U5752 ( .B1(n4940), .B2(n7129), .A(n4472), .ZN(n4939) );
  INV_X1 U5753 ( .A(n7051), .ZN(n4940) );
  INV_X1 U5754 ( .A(n5259), .ZN(n5551) );
  INV_X1 U5755 ( .A(n5235), .ZN(n5550) );
  NAND2_X1 U5756 ( .A1(n4639), .A2(n9515), .ZN(n9422) );
  NAND2_X1 U5757 ( .A1(n7111), .A2(n7350), .ZN(n4942) );
  NAND2_X1 U5758 ( .A1(n7345), .A2(n7347), .ZN(n7479) );
  NAND3_X2 U5759 ( .A1(n5191), .A2(n5030), .A3(n5190), .ZN(n6945) );
  NAND2_X1 U5760 ( .A1(n8699), .A2(n6709), .ZN(n6546) );
  NAND2_X1 U5761 ( .A1(n7474), .A2(n6709), .ZN(n7515) );
  INV_X1 U5762 ( .A(n6709), .ZN(n6726) );
  NAND2_X1 U5763 ( .A1(n5681), .A2(n5680), .ZN(n9152) );
  INV_X1 U5764 ( .A(n9004), .ZN(n8996) );
  NAND2_X1 U5765 ( .A1(n4972), .A2(n4973), .ZN(n9108) );
  NOR2_X1 U5766 ( .A1(n9107), .A2(n4971), .ZN(n4970) );
  INV_X1 U5767 ( .A(n4973), .ZN(n4971) );
  INV_X1 U5768 ( .A(n9544), .ZN(n9507) );
  INV_X1 U5769 ( .A(n9541), .ZN(n9501) );
  NOR2_X1 U5770 ( .A1(n9124), .A2(n9123), .ZN(n9203) );
  AND2_X1 U5771 ( .A1(n4488), .A2(n5122), .ZN(n4816) );
  AOI21_X1 U5772 ( .B1(n6292), .B2(n6291), .A(n4870), .ZN(n4611) );
  INV_X1 U5773 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5124) );
  INV_X1 U5774 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U5775 ( .A(n6292), .B(n6291), .ZN(n8550) );
  XNOR2_X1 U5776 ( .A(n5717), .B(n5716), .ZN(n8554) );
  NAND2_X1 U5777 ( .A1(n4447), .A2(n5119), .ZN(n4684) );
  NAND2_X1 U5778 ( .A1(n4893), .A2(n4897), .ZN(n5605) );
  NAND2_X1 U5779 ( .A1(n4864), .A2(n5520), .ZN(n5539) );
  NAND2_X1 U5780 ( .A1(n5104), .A2(n5105), .ZN(n5522) );
  NAND2_X1 U5781 ( .A1(n4892), .A2(n5100), .ZN(n5478) );
  INV_X1 U5782 ( .A(n4934), .ZN(n4931) );
  NAND2_X1 U5783 ( .A1(n4884), .A2(n5087), .ZN(n5416) );
  OR2_X1 U5784 ( .A1(n5392), .A2(n5391), .ZN(n4884) );
  NOR2_X1 U5785 ( .A1(n4876), .A2(n4874), .ZN(n4873) );
  INV_X1 U5786 ( .A(n5066), .ZN(n4874) );
  INV_X1 U5787 ( .A(n5072), .ZN(n4541) );
  NAND2_X1 U5788 ( .A1(n5059), .A2(n5058), .ZN(n5307) );
  OR2_X1 U5789 ( .A1(n5304), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5344) );
  INV_X1 U5790 ( .A(n8215), .ZN(n7955) );
  NAND2_X1 U5791 ( .A1(n8070), .A2(n7595), .ZN(n7962) );
  NAND2_X1 U5792 ( .A1(n4844), .A2(n4845), .ZN(n7063) );
  NAND2_X1 U5793 ( .A1(n7575), .A2(n7577), .ZN(n7578) );
  INV_X1 U5794 ( .A(n8087), .ZN(n7997) );
  INV_X1 U5795 ( .A(n6678), .ZN(n6609) );
  AND4_X1 U5796 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n8050)
         );
  NAND2_X1 U5797 ( .A1(n8026), .A2(n8025), .ZN(n8024) );
  AND2_X1 U5798 ( .A1(n4843), .A2(n7065), .ZN(n4842) );
  AND2_X1 U5799 ( .A1(n4844), .A2(n4843), .ZN(n7066) );
  AND2_X1 U5800 ( .A1(n6176), .A2(n6175), .ZN(n8062) );
  NAND2_X1 U5801 ( .A1(n4834), .A2(n4832), .ZN(n8070) );
  NOR2_X1 U5802 ( .A1(n8068), .A2(n4833), .ZN(n4832) );
  INV_X1 U5803 ( .A(n4835), .ZN(n4833) );
  NAND2_X1 U5804 ( .A1(n4834), .A2(n4835), .ZN(n8069) );
  OR2_X1 U5805 ( .A1(n6784), .A2(n7275), .ZN(n8078) );
  NAND2_X1 U5806 ( .A1(n5011), .A2(n7801), .ZN(n5010) );
  INV_X1 U5807 ( .A(n8164), .ZN(n7840) );
  XNOR2_X1 U5808 ( .A(n6183), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7845) );
  INV_X1 U5809 ( .A(n8062), .ZN(n8205) );
  OAI211_X1 U5810 ( .C1(n4417), .C2(n10120), .A(n6153), .B(n6152), .ZN(n8229)
         );
  NAND4_X1 U5811 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n8251)
         );
  NAND4_X1 U5812 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n8092)
         );
  OR2_X1 U5813 ( .A1(n4416), .A2(n5807), .ZN(n5813) );
  OR2_X1 U5814 ( .A1(n5931), .A2(n5808), .ZN(n5812) );
  OAI21_X1 U5815 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6868), .A(n6867), .ZN(n6869) );
  NAND2_X1 U5816 ( .A1(n6867), .A2(n6799), .ZN(n6798) );
  NAND2_X1 U5817 ( .A1(n6868), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U5818 ( .A1(n6813), .A2(n4511), .ZN(n6645) );
  OR2_X1 U5819 ( .A1(n6644), .A2(n6662), .ZN(n4511) );
  NAND2_X1 U5820 ( .A1(n4628), .A2(n9582), .ZN(n6666) );
  NAND2_X1 U5821 ( .A1(n6760), .A2(n4622), .ZN(n9604) );
  NAND2_X1 U5822 ( .A1(n4507), .A2(n6983), .ZN(n6985) );
  NAND2_X1 U5823 ( .A1(n4636), .A2(n6983), .ZN(n6855) );
  AOI22_X1 U5824 ( .A1(n6972), .A2(n6971), .B1(n6975), .B2(n6970), .ZN(n8133)
         );
  INV_X1 U5825 ( .A(n4619), .ZN(n9640) );
  INV_X1 U5826 ( .A(n4617), .ZN(n9638) );
  AND2_X1 U5827 ( .A1(n6030), .A2(n6020), .ZN(n9694) );
  NAND2_X1 U5828 ( .A1(n6651), .A2(n6650), .ZN(n10209) );
  OAI21_X1 U5829 ( .B1(n8139), .B2(n9703), .A(n9697), .ZN(n9716) );
  AND2_X1 U5830 ( .A1(n6136), .A2(n6135), .ZN(n8231) );
  OAI21_X1 U5831 ( .B1(n7269), .B2(n6248), .A(n7686), .ZN(n8365) );
  AND2_X1 U5832 ( .A1(n4778), .A2(n4448), .ZN(n7264) );
  NAND2_X1 U5833 ( .A1(n7092), .A2(n7667), .ZN(n7144) );
  AND2_X1 U5834 ( .A1(n7784), .A2(n7840), .ZN(n9767) );
  INV_X1 U5835 ( .A(n8373), .ZN(n9768) );
  OR2_X1 U5836 ( .A1(n6275), .A2(n6593), .ZN(n8373) );
  INV_X1 U5837 ( .A(n8180), .ZN(n8378) );
  NAND2_X1 U5838 ( .A1(n8447), .A2(n9833), .ZN(n8450) );
  NAND2_X1 U5839 ( .A1(n6147), .A2(n6146), .ZN(n8462) );
  INV_X1 U5840 ( .A(n8231), .ZN(n8468) );
  NAND2_X1 U5841 ( .A1(n6127), .A2(n6126), .ZN(n8474) );
  NAND2_X1 U5842 ( .A1(n8248), .A2(n6125), .ZN(n8237) );
  NAND2_X1 U5843 ( .A1(n6116), .A2(n6115), .ZN(n8480) );
  INV_X1 U5844 ( .A(n7603), .ZN(n8492) );
  AOI21_X1 U5845 ( .B1(n8293), .B2(n6081), .A(n4769), .ZN(n8283) );
  NAND2_X1 U5846 ( .A1(n4995), .A2(n4998), .ZN(n8280) );
  NAND2_X1 U5847 ( .A1(n8291), .A2(n7807), .ZN(n4995) );
  INV_X1 U5848 ( .A(n7601), .ZN(n8503) );
  AND2_X1 U5849 ( .A1(n8309), .A2(n8308), .ZN(n8508) );
  NAND2_X1 U5850 ( .A1(n6047), .A2(n6046), .ZN(n8515) );
  AND2_X1 U5851 ( .A1(n8320), .A2(n8319), .ZN(n8514) );
  NAND2_X1 U5852 ( .A1(n4748), .A2(n4745), .ZN(n8316) );
  NAND2_X1 U5853 ( .A1(n4987), .A2(n4992), .ZN(n8360) );
  NAND2_X1 U5854 ( .A1(n7269), .A2(n4993), .ZN(n4987) );
  INV_X1 U5855 ( .A(n6410), .ZN(n6593) );
  NAND2_X1 U5856 ( .A1(n6211), .A2(n6210), .ZN(n6213) );
  MUX2_X1 U5857 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6209), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6211) );
  NAND2_X1 U5858 ( .A1(n6199), .A2(n6207), .ZN(n6208) );
  NOR2_X1 U5859 ( .A1(n4418), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8552) );
  INV_X1 U5860 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7273) );
  INV_X1 U5861 ( .A(n7845), .ZN(n7274) );
  INV_X1 U5862 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7170) );
  INV_X1 U5863 ( .A(n6612), .ZN(n7172) );
  INV_X1 U5864 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10081) );
  INV_X1 U5865 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6775) );
  INV_X1 U5866 ( .A(n8152), .ZN(n9753) );
  INV_X1 U5867 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6551) );
  INV_X1 U5868 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10152) );
  INV_X1 U5869 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10106) );
  INV_X1 U5870 ( .A(n9614), .ZN(n8128) );
  INV_X1 U5871 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6400) );
  INV_X1 U5872 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6391) );
  INV_X1 U5873 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6387) );
  AND3_X1 U5874 ( .A1(n4836), .A2(n5004), .A3(n5891), .ZN(n5907) );
  INV_X1 U5875 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6380) );
  NOR2_X1 U5876 ( .A1(n5860), .A2(n5005), .ZN(n5890) );
  XNOR2_X1 U5877 ( .A(n5877), .B(n5006), .ZN(n9591) );
  NAND2_X1 U5878 ( .A1(n5823), .A2(n5822), .ZN(n6794) );
  NAND2_X1 U5879 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5820) );
  XNOR2_X1 U5880 ( .A(n5757), .B(n5756), .ZN(n6407) );
  INV_X1 U5881 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U5882 ( .A1(n6874), .A2(n6875), .ZN(n4930) );
  OR2_X1 U5883 ( .A1(n4919), .A2(n4918), .ZN(n8562) );
  NAND2_X1 U5884 ( .A1(n4653), .A2(n4657), .ZN(n8582) );
  NAND2_X1 U5885 ( .A1(n8624), .A2(n4658), .ZN(n4653) );
  AND2_X1 U5886 ( .A1(n6351), .A2(n5775), .ZN(n8935) );
  NAND2_X1 U5887 ( .A1(n8590), .A2(n8591), .ZN(n8589) );
  NAND2_X1 U5888 ( .A1(n8664), .A2(n5584), .ZN(n8590) );
  NAND2_X1 U5889 ( .A1(n8633), .A2(n4927), .ZN(n8634) );
  NAND2_X1 U5890 ( .A1(n5244), .A2(n4443), .ZN(n8656) );
  NAND2_X1 U5891 ( .A1(n5244), .A2(n5243), .ZN(n4921) );
  NAND2_X1 U5892 ( .A1(n4651), .A2(n4649), .ZN(n8667) );
  AOI21_X1 U5893 ( .B1(n7289), .B2(n7291), .A(n7290), .ZN(n7293) );
  NOR2_X1 U5894 ( .A1(n8674), .A2(n8675), .ZN(n8673) );
  NAND2_X1 U5895 ( .A1(n5618), .A2(n4682), .ZN(n8674) );
  INV_X1 U5896 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U5897 ( .A1(n8634), .A2(n4925), .ZN(n8684) );
  OR2_X1 U5898 ( .A1(n5783), .A2(n6721), .ZN(n9255) );
  AND2_X1 U5899 ( .A1(n5765), .A2(n5763), .ZN(n8709) );
  INV_X1 U5900 ( .A(n9267), .ZN(n8713) );
  INV_X1 U5901 ( .A(n7309), .ZN(n8727) );
  AOI22_X1 U5902 ( .A1(n5248), .A2(P1_REG1_REG_1__SCAN_IN), .B1(n5202), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U5903 ( .A1(n8787), .A2(n8788), .ZN(n8786) );
  NOR2_X1 U5904 ( .A1(n6479), .A2(n6478), .ZN(n6477) );
  AND2_X1 U5905 ( .A1(n8786), .A2(n4560), .ZN(n6479) );
  NAND2_X1 U5906 ( .A1(n6450), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4560) );
  NOR2_X1 U5907 ( .A1(n6436), .A2(n6435), .ZN(n6519) );
  INV_X1 U5908 ( .A(n9368), .ZN(n9383) );
  NAND2_X1 U5909 ( .A1(n8857), .A2(n9436), .ZN(n9119) );
  INV_X1 U5910 ( .A(n9152), .ZN(n8986) );
  NAND2_X1 U5911 ( .A1(n9008), .A2(n8918), .ZN(n8991) );
  NAND2_X1 U5912 ( .A1(n4535), .A2(n4964), .ZN(n8989) );
  OR2_X1 U5913 ( .A1(n9017), .A2(n4966), .ZN(n4535) );
  NAND2_X1 U5914 ( .A1(n4969), .A2(n8893), .ZN(n9003) );
  NAND2_X1 U5915 ( .A1(n9017), .A2(n4440), .ZN(n4969) );
  AND2_X1 U5916 ( .A1(n5611), .A2(n5610), .ZN(n9030) );
  NAND2_X1 U5917 ( .A1(n4542), .A2(n4549), .ZN(n9033) );
  NAND2_X1 U5918 ( .A1(n4944), .A2(n4424), .ZN(n9046) );
  NAND2_X1 U5919 ( .A1(n8884), .A2(n4947), .ZN(n4944) );
  INV_X1 U5920 ( .A(n4810), .ZN(n9061) );
  OAI21_X1 U5921 ( .B1(n9087), .B2(n4811), .A(n7447), .ZN(n4810) );
  NAND2_X1 U5922 ( .A1(n8884), .A2(n8883), .ZN(n9060) );
  NAND2_X1 U5923 ( .A1(n4949), .A2(n4954), .ZN(n7222) );
  OR2_X1 U5924 ( .A1(n7073), .A2(n4955), .ZN(n4949) );
  AND2_X1 U5925 ( .A1(n4957), .A2(n4454), .ZN(n7173) );
  NAND2_X1 U5926 ( .A1(n7073), .A2(n7075), .ZN(n4957) );
  NAND2_X1 U5927 ( .A1(n4797), .A2(n7345), .ZN(n7034) );
  NAND2_X1 U5928 ( .A1(n9452), .A2(n6734), .ZN(n9104) );
  AND2_X1 U5929 ( .A1(n9452), .A2(n5549), .ZN(n9440) );
  OR2_X1 U5930 ( .A1(n9121), .A2(n7559), .ZN(n7121) );
  OR2_X1 U5931 ( .A1(n5259), .A2(n6373), .ZN(n5214) );
  NAND2_X1 U5932 ( .A1(n4785), .A2(n7515), .ZN(n9458) );
  AND2_X2 U5933 ( .A1(n9203), .A2(n9125), .ZN(n9575) );
  NAND2_X1 U5934 ( .A1(n9131), .A2(n9541), .ZN(n4555) );
  OR2_X1 U5935 ( .A1(n9133), .A2(n4500), .ZN(n4554) );
  AND2_X2 U5936 ( .A1(n9203), .A2(n9202), .ZN(n9553) );
  OR2_X1 U5937 ( .A1(n7559), .A2(n6396), .ZN(n9457) );
  INV_X1 U5938 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U5939 ( .A(n7331), .B(n7330), .ZN(n9227) );
  XNOR2_X1 U5940 ( .A(n5645), .B(n5644), .ZN(n7286) );
  NOR2_X1 U5941 ( .A1(n4418), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9226) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7565) );
  INV_X1 U5943 ( .A(n5760), .ZN(n7563) );
  INV_X1 U5944 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7157) );
  OR2_X1 U5945 ( .A1(n5134), .A2(n4688), .ZN(n5136) );
  INV_X1 U5946 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7032) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10070) );
  AND3_X1 U5948 ( .A1(n4793), .A2(n4792), .A3(n4791), .ZN(n5393) );
  INV_X1 U5949 ( .A(n4788), .ZN(n4791) );
  XNOR2_X1 U5950 ( .A(n4518), .B(n4450), .ZN(n6401) );
  AOI21_X1 U5951 ( .B1(n4875), .B2(n4873), .A(n4541), .ZN(n4518) );
  NAND2_X1 U5952 ( .A1(n4875), .A2(n5066), .ZN(n5343) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6390) );
  INV_X1 U5954 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6389) );
  INV_X1 U5955 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6382) );
  INV_X1 U5956 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U5957 ( .A1(n5231), .A2(n5230), .ZN(n4859) );
  XNOR2_X1 U5958 ( .A(n4564), .B(n5229), .ZN(n8772) );
  OR2_X1 U5959 ( .A1(n4792), .A2(n4688), .ZN(n4564) );
  NOR2_X1 U5960 ( .A1(n4514), .A2(n4513), .ZN(n4512) );
  NOR2_X1 U5961 ( .A1(n7892), .A2(n8081), .ZN(n4513) );
  NAND2_X1 U5962 ( .A1(n4430), .A2(n4830), .ZN(n4823) );
  INV_X1 U5963 ( .A(n10224), .ZN(n4629) );
  AOI21_X1 U5964 ( .B1(n8169), .B2(n10223), .A(n8168), .ZN(n8170) );
  INV_X1 U5965 ( .A(n6271), .ZN(n6272) );
  OAI21_X1 U5966 ( .B1(n8454), .B2(n8381), .A(n6270), .ZN(n6271) );
  NOR2_X1 U5967 ( .A1(n8181), .A2(n8383), .ZN(n6367) );
  OAI21_X1 U5968 ( .B1(n6369), .B2(n4502), .A(n4773), .ZN(P2_U3456) );
  NOR2_X1 U5969 ( .A1(n4493), .A2(n4774), .ZN(n4773) );
  NOR2_X1 U5970 ( .A1(n9833), .A2(n4502), .ZN(n4774) );
  NAND2_X1 U5971 ( .A1(n4705), .A2(n4466), .ZN(n4701) );
  NAND2_X1 U5972 ( .A1(P1_U3973), .A2(n6709), .ZN(n6405) );
  INV_X1 U5973 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6705) );
  OR2_X1 U5974 ( .A1(n9057), .A2(n8888), .ZN(n4422) );
  NAND2_X1 U5975 ( .A1(n4897), .A2(n4468), .ZN(n4896) );
  AND2_X1 U5976 ( .A1(n4657), .A2(n4495), .ZN(n4423) );
  OR2_X1 U5977 ( .A1(n9070), .A2(n8886), .ZN(n4424) );
  AND2_X1 U5978 ( .A1(n4602), .A2(n4599), .ZN(n4425) );
  OR2_X1 U5979 ( .A1(n8474), .A2(n8251), .ZN(n4426) );
  AND2_X1 U5980 ( .A1(n4763), .A2(n4760), .ZN(n4427) );
  NOR2_X1 U5981 ( .A1(n4900), .A2(n4901), .ZN(n4428) );
  AND4_X1 U5982 ( .A1(n7400), .A2(n7467), .A3(n7469), .A4(n7399), .ZN(n4429)
         );
  AND2_X1 U5983 ( .A1(n4826), .A2(n4824), .ZN(n4430) );
  AND2_X1 U5984 ( .A1(n7440), .A2(n7455), .ZN(n8905) );
  OR2_X1 U5985 ( .A1(n8457), .A2(n7955), .ZN(n7755) );
  AND2_X1 U5986 ( .A1(n5481), .A2(n5480), .ZN(n9276) );
  OR2_X1 U5987 ( .A1(n7362), .A2(n4463), .ZN(n4431) );
  AND2_X1 U5988 ( .A1(n7772), .A2(n4580), .ZN(n4432) );
  INV_X1 U5989 ( .A(n7700), .ZN(n4750) );
  INV_X1 U5990 ( .A(n8682), .ZN(n4924) );
  OR2_X1 U5991 ( .A1(n4889), .A2(SI_16_), .ZN(n4433) );
  AND2_X1 U5992 ( .A1(n4640), .A2(n9105), .ZN(n4434) );
  AND2_X1 U5993 ( .A1(n5089), .A2(SI_12_), .ZN(n4435) );
  NAND2_X1 U5994 ( .A1(n4480), .A2(n4924), .ZN(n4657) );
  OR2_X1 U5995 ( .A1(n6853), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4437) );
  AND2_X1 U5996 ( .A1(n4975), .A2(n4816), .ZN(n4438) );
  OAI21_X1 U5997 ( .B1(n7289), .B2(n7290), .A(n4915), .ZN(n4919) );
  INV_X1 U5998 ( .A(n4896), .ZN(n4895) );
  INV_X1 U5999 ( .A(n8720), .ZN(n8926) );
  INV_X1 U6000 ( .A(n7350), .ZN(n4938) );
  INV_X1 U6001 ( .A(n6293), .ZN(n4870) );
  NOR2_X1 U6002 ( .A1(n6873), .A2(n4508), .ZN(n4439) );
  NAND4_X1 U6003 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5850)
         );
  AND2_X1 U6004 ( .A1(n5208), .A2(n5209), .ZN(n4792) );
  INV_X1 U6005 ( .A(n8878), .ZN(n4548) );
  OR2_X1 U6006 ( .A1(n9030), .A2(n8892), .ZN(n4440) );
  NAND2_X2 U6007 ( .A1(n5235), .A2(n5047), .ZN(n5232) );
  OR2_X1 U6008 ( .A1(n9043), .A2(n8889), .ZN(n4441) );
  NAND2_X1 U6009 ( .A1(n7422), .A2(n7421), .ZN(n8868) );
  INV_X1 U6010 ( .A(n8868), .ZN(n9128) );
  NOR2_X1 U6011 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5821) );
  BUF_X1 U6012 ( .A(n5192), .Z(n5287) );
  NAND2_X1 U6013 ( .A1(n5731), .A2(n6340), .ZN(n5192) );
  INV_X1 U6014 ( .A(n5202), .ZN(n5595) );
  OR2_X1 U6015 ( .A1(n5018), .A2(n7670), .ZN(n4442) );
  AND2_X1 U6016 ( .A1(n4920), .A2(n5243), .ZN(n4443) );
  AND2_X1 U6017 ( .A1(n8861), .A2(n8860), .ZN(n4445) );
  AND2_X1 U6018 ( .A1(n7558), .A2(n6722), .ZN(n4446) );
  AND4_X1 U6019 ( .A1(n4683), .A2(n5117), .A3(n5153), .A4(n5132), .ZN(n4447)
         );
  INV_X1 U6020 ( .A(n8918), .ZN(n4802) );
  OR2_X1 U6021 ( .A1(n8087), .A2(n9814), .ZN(n4448) );
  NOR2_X1 U6022 ( .A1(n5518), .A2(n5519), .ZN(n4926) );
  NAND2_X1 U6023 ( .A1(n6154), .A2(n7624), .ZN(n8203) );
  AND2_X1 U6024 ( .A1(n6860), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U6025 ( .A1(n4983), .A2(n7745), .ZN(n8236) );
  AND2_X1 U6026 ( .A1(n5077), .A2(n5076), .ZN(n4450) );
  INV_X1 U6027 ( .A(n7526), .ZN(n4727) );
  AND2_X1 U6028 ( .A1(n6912), .A2(n4846), .ZN(n4451) );
  NAND2_X1 U6029 ( .A1(n5700), .A2(n5699), .ZN(n9146) );
  INV_X1 U6030 ( .A(n9146), .ZN(n8966) );
  AND2_X1 U6031 ( .A1(n4617), .A2(n4616), .ZN(n4452) );
  NAND2_X1 U6032 ( .A1(n5501), .A2(n5500), .ZN(n9192) );
  NAND2_X1 U6033 ( .A1(n7521), .A2(n7358), .ZN(n7075) );
  AND3_X1 U6034 ( .A1(n7668), .A2(n7783), .A3(n7667), .ZN(n4453) );
  NAND2_X1 U6035 ( .A1(n4836), .A2(n5790), .ZN(n5862) );
  NAND2_X1 U6036 ( .A1(n4763), .A2(n4764), .ZN(n8271) );
  AND2_X1 U6037 ( .A1(n5468), .A2(n5467), .ZN(n9545) );
  NAND2_X1 U6038 ( .A1(n5792), .A2(n5791), .ZN(n5956) );
  OR2_X1 U6039 ( .A1(n7283), .A2(n8731), .ZN(n4454) );
  AND2_X1 U6040 ( .A1(n9010), .A2(n9019), .ZN(n4455) );
  NAND2_X1 U6041 ( .A1(n4776), .A2(n5004), .ZN(n5924) );
  AND3_X1 U6042 ( .A1(n7407), .A2(n7406), .A3(n7405), .ZN(n4456) );
  INV_X1 U6043 ( .A(n8698), .ZN(n8904) );
  AND2_X1 U6044 ( .A1(n5803), .A2(n5020), .ZN(n4457) );
  NAND2_X1 U6045 ( .A1(n7676), .A2(n7675), .ZN(n4458) );
  OR2_X1 U6046 ( .A1(n7892), .A2(n8062), .ZN(n4459) );
  OR2_X1 U6047 ( .A1(n6067), .A2(n7963), .ZN(n4460) );
  INV_X1 U6048 ( .A(n4671), .ZN(n4670) );
  NAND2_X1 U6049 ( .A1(n8606), .A2(n4672), .ZN(n4671) );
  INV_X1 U6050 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U6051 ( .A1(n4762), .A2(n4764), .ZN(n4761) );
  OR2_X1 U6052 ( .A1(n6752), .A2(n6751), .ZN(n4461) );
  INV_X1 U6053 ( .A(n4804), .ZN(n4803) );
  NAND2_X1 U6054 ( .A1(n9010), .A2(n8916), .ZN(n4804) );
  AND2_X1 U6055 ( .A1(n9161), .A2(n8895), .ZN(n4462) );
  NOR2_X1 U6056 ( .A1(n7359), .A2(n7360), .ZN(n4463) );
  AND2_X1 U6057 ( .A1(n4649), .A2(n4648), .ZN(n4464) );
  NOR2_X1 U6058 ( .A1(n9000), .A2(n8896), .ZN(n4465) );
  OR2_X1 U6059 ( .A1(n7221), .A2(n7176), .ZN(n7367) );
  INV_X1 U6060 ( .A(n7472), .ZN(n4786) );
  NAND2_X1 U6061 ( .A1(n4708), .A2(n4709), .ZN(n4466) );
  AND2_X1 U6062 ( .A1(n7445), .A2(n7533), .ZN(n9107) );
  AND2_X1 U6063 ( .A1(n8656), .A2(n5272), .ZN(n4467) );
  OR2_X1 U6064 ( .A1(n5604), .A2(SI_21_), .ZN(n4468) );
  NOR2_X1 U6065 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  OR2_X1 U6066 ( .A1(n7878), .A2(n4825), .ZN(n4469) );
  INV_X1 U6067 ( .A(n4551), .ZN(n4550) );
  NOR2_X1 U6068 ( .A1(n9083), .A2(n8881), .ZN(n4551) );
  INV_X1 U6069 ( .A(n4540), .ZN(n4539) );
  OAI21_X1 U6070 ( .B1(n4873), .B2(n4541), .A(n4450), .ZN(n4540) );
  NOR2_X1 U6071 ( .A1(n6054), .A2(n7959), .ZN(n4470) );
  NOR2_X1 U6072 ( .A1(n6319), .A2(n6318), .ZN(n4471) );
  AND2_X1 U6073 ( .A1(n7052), .A2(n9515), .ZN(n4472) );
  OR2_X1 U6074 ( .A1(n5465), .A2(n4684), .ZN(n4473) );
  INV_X1 U6075 ( .A(n4581), .ZN(n7802) );
  AND2_X1 U6076 ( .A1(n6954), .A2(n6953), .ZN(n4474) );
  OR2_X1 U6077 ( .A1(n4684), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U6078 ( .A1(n7832), .A2(n7783), .ZN(n4476) );
  INV_X1 U6079 ( .A(n4999), .ZN(n4998) );
  NAND2_X1 U6080 ( .A1(n8282), .A2(n5000), .ZN(n4999) );
  INV_X1 U6081 ( .A(n4746), .ZN(n4745) );
  NAND2_X1 U6082 ( .A1(n8317), .A2(n4747), .ZN(n4746) );
  AND2_X1 U6083 ( .A1(n5335), .A2(n5334), .ZN(n4477) );
  OAI21_X1 U6084 ( .B1(n7818), .B2(n4442), .A(n7676), .ZN(n5017) );
  NAND2_X1 U6085 ( .A1(n7586), .A2(n7938), .ZN(n4478) );
  AND2_X1 U6086 ( .A1(n8952), .A2(n8698), .ZN(n4479) );
  OAI21_X1 U6087 ( .B1(n7414), .B2(n9128), .A(n4737), .ZN(n4736) );
  OAI21_X1 U6088 ( .B1(n8250), .B2(n4754), .A(n6134), .ZN(n4753) );
  NAND2_X1 U6089 ( .A1(n4923), .A2(n8680), .ZN(n4480) );
  NAND2_X1 U6090 ( .A1(n8364), .A2(n4994), .ZN(n4481) );
  AND2_X1 U6091 ( .A1(n5120), .A2(n4977), .ZN(n4482) );
  INV_X1 U6092 ( .A(n4926), .ZN(n4925) );
  INV_X1 U6093 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6094 ( .A1(n4738), .A2(n4735), .ZN(n4483) );
  NAND2_X1 U6095 ( .A1(n9047), .A2(n4945), .ZN(n4484) );
  AND2_X1 U6096 ( .A1(n7822), .A2(n4448), .ZN(n4485) );
  AND2_X1 U6097 ( .A1(n8095), .A2(n8128), .ZN(n4486) );
  NAND2_X1 U6098 ( .A1(n7412), .A2(n7411), .ZN(n9134) );
  AND2_X1 U6099 ( .A1(n4797), .A2(n4795), .ZN(n4487) );
  NOR2_X1 U6100 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4488) );
  NOR2_X1 U6101 ( .A1(n8990), .A2(n4802), .ZN(n4801) );
  NOR2_X1 U6102 ( .A1(n7587), .A2(n4840), .ZN(n4839) );
  AND2_X1 U6103 ( .A1(n4915), .A2(n4913), .ZN(n4489) );
  NAND2_X1 U6104 ( .A1(n7064), .A2(n7067), .ZN(n4490) );
  INV_X1 U6105 ( .A(n8880), .ZN(n9270) );
  AND2_X1 U6106 ( .A1(n4430), .A2(n4469), .ZN(n4491) );
  INV_X1 U6107 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4688) );
  INV_X1 U6108 ( .A(n5014), .ZN(n5013) );
  NAND2_X1 U6109 ( .A1(n6335), .A2(n6334), .ZN(n9136) );
  INV_X1 U6110 ( .A(n9136), .ZN(n4643) );
  NAND2_X1 U6111 ( .A1(n4972), .A2(n4970), .ZN(n9106) );
  AND2_X1 U6112 ( .A1(n9408), .A2(n4434), .ZN(n4492) );
  NAND2_X1 U6113 ( .A1(n4666), .A2(n4670), .ZN(n7289) );
  NAND2_X1 U6114 ( .A1(n5155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6115 ( .A1(n6003), .A2(n6002), .ZN(n8350) );
  NAND2_X1 U6116 ( .A1(n4942), .A2(n7051), .ZN(n9414) );
  NAND2_X1 U6117 ( .A1(n4770), .A2(n7692), .ZN(n8336) );
  NAND2_X1 U6118 ( .A1(n6295), .A2(n6294), .ZN(n8443) );
  INV_X1 U6119 ( .A(n8443), .ZN(n4580) );
  INV_X1 U6120 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4977) );
  INV_X1 U6121 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4854) );
  NOR2_X1 U6122 ( .A1(n5101), .A2(n5475), .ZN(n4889) );
  INV_X1 U6123 ( .A(n4889), .ZN(n4613) );
  NAND2_X1 U6124 ( .A1(n9182), .A2(n8886), .ZN(n7539) );
  INV_X1 U6125 ( .A(n7539), .ZN(n4809) );
  NOR2_X1 U6126 ( .A1(n4790), .A2(n4646), .ZN(n5439) );
  NAND2_X1 U6127 ( .A1(n4789), .A2(n4678), .ZN(n5417) );
  NOR2_X1 U6128 ( .A1(n8181), .A2(n8433), .ZN(n4493) );
  NAND2_X1 U6129 ( .A1(n7283), .A2(n7040), .ZN(n7358) );
  OR2_X1 U6130 ( .A1(n6071), .A2(n5028), .ZN(n4494) );
  INV_X1 U6131 ( .A(n8872), .ZN(n8874) );
  AND2_X1 U6132 ( .A1(n5486), .A2(n5485), .ZN(n8872) );
  NAND2_X1 U6133 ( .A1(n5567), .A2(n5566), .ZN(n4495) );
  AND2_X1 U6134 ( .A1(n9000), .A2(n8896), .ZN(n4496) );
  NOR2_X1 U6135 ( .A1(n5417), .A2(n4932), .ZN(n5497) );
  NAND2_X1 U6136 ( .A1(n4919), .A2(n4918), .ZN(n4497) );
  AND2_X1 U6137 ( .A1(n5604), .A2(SI_21_), .ZN(n4498) );
  AND2_X1 U6138 ( .A1(n5725), .A2(n5724), .ZN(n8952) );
  INV_X1 U6139 ( .A(n8952), .ZN(n9141) );
  AND2_X1 U6140 ( .A1(n9106), .A2(n8876), .ZN(n9092) );
  AND2_X1 U6141 ( .A1(n4548), .A2(n4547), .ZN(n4499) );
  AND2_X1 U6142 ( .A1(n9134), .A2(n9507), .ZN(n4500) );
  AND2_X1 U6143 ( .A1(n4748), .A2(n4747), .ZN(n4501) );
  INV_X1 U6144 ( .A(SI_20_), .ZN(n5586) );
  INV_X1 U6145 ( .A(n7129), .ZN(n4941) );
  AND2_X1 U6146 ( .A1(n5164), .A2(n4904), .ZN(n5760) );
  INV_X1 U6147 ( .A(n6297), .ZN(n4872) );
  NAND2_X1 U6148 ( .A1(n7508), .A2(n7563), .ZN(n9130) );
  INV_X2 U6149 ( .A(n9835), .ZN(n9833) );
  NOR2_X1 U6150 ( .A1(n7119), .A2(n9506), .ZN(n4639) );
  AND2_X1 U6151 ( .A1(n9835), .A2(n10113), .ZN(n4502) );
  AND2_X1 U6152 ( .A1(n9301), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U6153 ( .A1(n4930), .A2(n5317), .ZN(n6952) );
  AND2_X1 U6154 ( .A1(n8822), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U6155 ( .A1(n5962), .A2(n5961), .ZN(n7241) );
  NAND2_X1 U6156 ( .A1(n7224), .A2(n7228), .ZN(n7308) );
  NAND2_X1 U6157 ( .A1(n5930), .A2(n5929), .ZN(n7146) );
  AND2_X1 U6158 ( .A1(n6299), .A2(n9965), .ZN(n4505) );
  INV_X1 U6159 ( .A(n9851), .ZN(n9849) );
  XNOR2_X1 U6160 ( .A(n5816), .B(n5815), .ZN(n6192) );
  NOR2_X1 U6161 ( .A1(n6192), .A2(P2_U3151), .ZN(n4506) );
  NAND2_X1 U6162 ( .A1(n5761), .A2(n5160), .ZN(n6722) );
  XNOR2_X1 U6163 ( .A(n6181), .B(n6180), .ZN(n7784) );
  NAND4_X1 U6164 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n6900)
         );
  INV_X1 U6165 ( .A(n6900), .ZN(n4981) );
  AND2_X1 U6166 ( .A1(n6730), .A2(n6729), .ZN(n9399) );
  INV_X1 U6167 ( .A(n9399), .ZN(n9459) );
  INV_X1 U6168 ( .A(n8699), .ZN(n8927) );
  INV_X1 U6169 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5020) );
  AND2_X1 U6170 ( .A1(n6603), .A2(n6602), .ZN(n8067) );
  INV_X1 U6171 ( .A(n8067), .ZN(n4824) );
  OR2_X1 U6172 ( .A1(n7561), .A2(n7560), .ZN(n4709) );
  AND2_X1 U6173 ( .A1(n4636), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4507) );
  AND2_X1 U6174 ( .A1(n10209), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4508) );
  INV_X1 U6175 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5153) );
  NOR2_X1 U6176 ( .A1(n4625), .A2(n9600), .ZN(n4624) );
  INV_X1 U6177 ( .A(n9600), .ZN(n4510) );
  NAND2_X1 U6178 ( .A1(n4623), .A2(n9600), .ZN(n6760) );
  OAI21_X1 U6179 ( .B1(n5047), .B2(n5036), .A(n5035), .ZN(n5037) );
  INV_X1 U6180 ( .A(n9062), .ZN(n4814) );
  NAND2_X1 U6181 ( .A1(n4555), .A2(n4553), .ZN(n9206) );
  NAND2_X1 U6182 ( .A1(n9648), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9647) );
  INV_X1 U6183 ( .A(n5860), .ZN(n4836) );
  AOI21_X1 U6184 ( .B1(n9746), .B2(n9745), .A(n8154), .ZN(n10206) );
  NOR2_X1 U6185 ( .A1(n5005), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4775) );
  INV_X1 U6186 ( .A(n6182), .ZN(n4782) );
  NOR2_X1 U6187 ( .A1(n6220), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6199) );
  AOI21_X1 U6188 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(n9576) );
  OAI22_X2 U6189 ( .A1(n8048), .A2(n8049), .B1(n7602), .B2(n8307), .ZN(n7916)
         );
  NOR2_X2 U6190 ( .A1(n7612), .A2(n7611), .ZN(n7855) );
  NOR2_X1 U6191 ( .A1(n6781), .A2(n6782), .ZN(n6909) );
  NAND4_X2 U6192 ( .A1(n5813), .A2(n5811), .A3(n5810), .A4(n5812), .ZN(n9760)
         );
  NAND2_X1 U6193 ( .A1(n4515), .A2(n4512), .ZN(P2_U3154) );
  NAND2_X1 U6194 ( .A1(n7886), .A2(n7885), .ZN(n4515) );
  NAND2_X1 U6195 ( .A1(n7865), .A2(n7864), .ZN(n7951) );
  NAND2_X1 U6196 ( .A1(n7574), .A2(n7573), .ZN(n7575) );
  NOR2_X1 U6197 ( .A1(n6629), .A2(n6619), .ZN(n6621) );
  OAI21_X2 U6198 ( .B1(n8017), .B2(n8018), .A(n4516), .ZN(n7893) );
  NAND2_X1 U6199 ( .A1(n4776), .A2(n4775), .ZN(n5939) );
  INV_X1 U6200 ( .A(n4875), .ZN(n4538) );
  INV_X1 U6201 ( .A(n4576), .ZN(n4575) );
  INV_X1 U6202 ( .A(n5496), .ZN(n5102) );
  NAND2_X1 U6203 ( .A1(n4567), .A2(n4566), .ZN(n4565) );
  NAND2_X1 U6204 ( .A1(n7839), .A2(n8434), .ZN(n5007) );
  NAND2_X1 U6205 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U6206 ( .A1(n7680), .A2(n7681), .ZN(n7685) );
  OAI21_X1 U6207 ( .B1(n4583), .B2(n7746), .A(n7769), .ZN(n4582) );
  NOR2_X1 U6208 ( .A1(n4879), .A2(n7782), .ZN(n4527) );
  OAI21_X1 U6209 ( .B1(n4632), .B2(n10220), .A(n4631), .ZN(n4630) );
  INV_X1 U6210 ( .A(n7442), .ZN(n4787) );
  NAND2_X1 U6211 ( .A1(n4787), .A2(n4786), .ZN(n7444) );
  NOR2_X2 U6212 ( .A1(n9018), .A2(n8915), .ZN(n9022) );
  NAND3_X1 U6213 ( .A1(n4797), .A2(n4795), .A3(n7483), .ZN(n7523) );
  AOI21_X1 U6214 ( .B1(n10222), .B2(n10223), .A(n10221), .ZN(n4631) );
  XNOR2_X1 U6215 ( .A(n4630), .B(n4629), .ZN(P2_U3200) );
  NAND2_X1 U6216 ( .A1(n7685), .A2(n7684), .ZN(n7689) );
  OAI21_X2 U6217 ( .B1(n4527), .B2(n4476), .A(n4526), .ZN(n7838) );
  NAND2_X1 U6218 ( .A1(n4578), .A2(n4581), .ZN(n7779) );
  NAND2_X1 U6219 ( .A1(n4565), .A2(n8303), .ZN(n7725) );
  INV_X1 U6220 ( .A(n5009), .ZN(n5008) );
  OAI211_X1 U6221 ( .C1(n7748), .C2(n7769), .A(n8224), .B(n4582), .ZN(n7754)
         );
  NAND2_X1 U6222 ( .A1(n7690), .A2(n7769), .ZN(n4570) );
  NAND2_X1 U6223 ( .A1(n9017), .A2(n4533), .ZN(n4532) );
  OAI21_X2 U6224 ( .B1(n4538), .B2(n4540), .A(n4536), .ZN(n5373) );
  NAND3_X1 U6225 ( .A1(n4547), .A2(n4548), .A3(n4546), .ZN(n4542) );
  NAND4_X1 U6226 ( .A1(n4547), .A2(n4441), .A3(n4548), .A4(n4546), .ZN(n4545)
         );
  NAND3_X1 U6227 ( .A1(n4547), .A2(n4548), .A3(n4550), .ZN(n8884) );
  AOI21_X1 U6228 ( .B1(n7691), .B2(n7783), .A(n8366), .ZN(n4571) );
  OR2_X1 U6229 ( .A1(n7773), .A2(n4575), .ZN(n4572) );
  NAND2_X1 U6230 ( .A1(n4572), .A2(n4573), .ZN(n4877) );
  NAND2_X1 U6231 ( .A1(n7773), .A2(n7772), .ZN(n7781) );
  OR2_X1 U6232 ( .A1(n7773), .A2(n7772), .ZN(n4578) );
  OR2_X1 U6233 ( .A1(n7772), .A2(n4580), .ZN(n4579) );
  OAI21_X2 U6234 ( .B1(n4589), .B2(n4588), .A(n4586), .ZN(n8145) );
  NAND2_X1 U6235 ( .A1(n5544), .A2(n4425), .ZN(n4596) );
  NAND2_X2 U6236 ( .A1(n5094), .A2(n5093), .ZN(n5461) );
  MUX2_X1 U6237 ( .A(n8561), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6238 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8561), .S(n7621), .Z(n6678) );
  NAND2_X1 U6239 ( .A1(n9586), .A2(n4624), .ZN(n4622) );
  NAND2_X1 U6240 ( .A1(n6664), .A2(n6747), .ZN(n9582) );
  NAND2_X1 U6241 ( .A1(n4634), .A2(n4635), .ZN(n6981) );
  NAND2_X1 U6242 ( .A1(n6854), .A2(n4437), .ZN(n4634) );
  AND3_X2 U6243 ( .A1(n9408), .A2(n9270), .A3(n4434), .ZN(n9077) );
  NOR2_X1 U6244 ( .A1(n8981), .A2(n4642), .ZN(n8934) );
  OR2_X2 U6245 ( .A1(n8981), .A2(n4645), .ZN(n8947) );
  NOR2_X2 U6246 ( .A1(n9024), .A2(n9161), .ZN(n9004) );
  NOR2_X2 U6247 ( .A1(n9051), .A2(n9172), .ZN(n9039) );
  NAND4_X1 U6248 ( .A1(n5112), .A2(n5111), .A3(n4647), .A4(n5115), .ZN(n4646)
         );
  INV_X1 U6249 ( .A(n8624), .ZN(n4652) );
  NAND2_X1 U6250 ( .A1(n6579), .A2(n4661), .ZN(n4660) );
  INV_X1 U6251 ( .A(n5272), .ZN(n4662) );
  NAND2_X1 U6252 ( .A1(n7278), .A2(n4667), .ZN(n4663) );
  NAND2_X1 U6253 ( .A1(n4663), .A2(n4664), .ZN(n5489) );
  INV_X1 U6254 ( .A(n9235), .ZN(n4674) );
  NAND3_X1 U6255 ( .A1(n5294), .A2(n6820), .A3(n4928), .ZN(n4676) );
  NAND2_X1 U6256 ( .A1(n4676), .A2(n4675), .ZN(n5350) );
  NAND2_X1 U6257 ( .A1(n5294), .A2(n6820), .ZN(n6874) );
  NAND2_X1 U6258 ( .A1(n4680), .A2(n4679), .ZN(n8570) );
  OR2_X1 U6259 ( .A1(n5617), .A2(n5616), .ZN(n4682) );
  OR2_X1 U6260 ( .A1(n8572), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U6261 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  NAND2_X1 U6262 ( .A1(n4817), .A2(n5462), .ZN(n9220) );
  AOI21_X1 U6263 ( .B1(n4692), .B2(n4690), .A(n9093), .ZN(n7382) );
  OAI21_X1 U6264 ( .B1(n4699), .B2(n8990), .A(n4697), .ZN(n7408) );
  INV_X1 U6265 ( .A(n7511), .ZN(n4707) );
  NAND3_X1 U6266 ( .A1(n4703), .A2(n4702), .A3(n4701), .ZN(P1_U3242) );
  NAND3_X1 U6267 ( .A1(n5027), .A2(n7508), .A3(n4705), .ZN(n4702) );
  NAND3_X1 U6268 ( .A1(n4707), .A2(n4705), .A3(n4704), .ZN(n4703) );
  AOI22_X1 U6269 ( .A1(n4714), .A2(n4715), .B1(n4712), .B2(n4724), .ZN(n4711)
         );
  INV_X1 U6270 ( .A(n9130), .ZN(n4724) );
  INV_X1 U6271 ( .A(n7521), .ZN(n4728) );
  NAND2_X1 U6272 ( .A1(n4734), .A2(n4729), .ZN(n4733) );
  INV_X1 U6273 ( .A(n7415), .ZN(n4731) );
  NAND2_X1 U6274 ( .A1(n8868), .A2(n4724), .ZN(n4740) );
  INV_X1 U6275 ( .A(n8328), .ZN(n4749) );
  OAI21_X2 U6276 ( .B1(n4749), .B2(n4746), .A(n4744), .ZN(n8306) );
  OAI21_X2 U6277 ( .B1(n8249), .B2(n4752), .A(n4751), .ZN(n8228) );
  INV_X1 U6278 ( .A(n6125), .ZN(n4754) );
  NAND2_X1 U6279 ( .A1(n8249), .A2(n8250), .ZN(n8248) );
  NAND2_X1 U6280 ( .A1(n8293), .A2(n4758), .ZN(n4757) );
  NAND2_X1 U6281 ( .A1(n6003), .A2(n4771), .ZN(n4770) );
  AND2_X1 U6282 ( .A1(n5944), .A2(n5929), .ZN(n4777) );
  NAND2_X1 U6283 ( .A1(n5962), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U6284 ( .A1(n4778), .A2(n4485), .ZN(n7263) );
  NAND2_X1 U6285 ( .A1(n4782), .A2(n5800), .ZN(n6220) );
  NAND2_X1 U6286 ( .A1(n4782), .A2(n4781), .ZN(n5021) );
  OAI21_X1 U6287 ( .B1(n8195), .B2(n6296), .A(n5025), .ZN(n6309) );
  NOR2_X1 U6288 ( .A1(n6997), .A2(n5895), .ZN(n7103) );
  NAND2_X1 U6289 ( .A1(n8306), .A2(n8305), .ZN(n8304) );
  INV_X1 U6290 ( .A(n5939), .ZN(n5792) );
  NAND2_X1 U6291 ( .A1(n6290), .A2(n6289), .ZN(n8195) );
  NOR2_X1 U6292 ( .A1(n7103), .A2(n7102), .ZN(n5913) );
  OAI211_X1 U6293 ( .C1(n6322), .C2(n9762), .A(n6321), .B(n6320), .ZN(n8179)
         );
  NAND2_X1 U6294 ( .A1(n8304), .A2(n4460), .ZN(n8293) );
  NAND2_X1 U6295 ( .A1(n4784), .A2(n4783), .ZN(n6935) );
  NAND2_X1 U6296 ( .A1(n6726), .A2(n9446), .ZN(n4785) );
  INV_X1 U6297 ( .A(n9022), .ZN(n4805) );
  NAND2_X1 U6298 ( .A1(n9022), .A2(n4801), .ZN(n4798) );
  NOR2_X1 U6299 ( .A1(n9022), .A2(n8917), .ZN(n9009) );
  NOR2_X1 U6300 ( .A1(n9088), .A2(n9093), .ZN(n9087) );
  NAND2_X1 U6301 ( .A1(n9088), .A2(n4812), .ZN(n4807) );
  NOR2_X1 U6302 ( .A1(n9087), .A2(n7446), .ZN(n9073) );
  AOI21_X1 U6303 ( .B1(n5462), .B2(n4438), .A(n4688), .ZN(n5143) );
  AND2_X1 U6304 ( .A1(n5462), .A2(n4975), .ZN(n5139) );
  NAND2_X1 U6305 ( .A1(n7883), .A2(n4491), .ZN(n4822) );
  OAI211_X1 U6306 ( .C1(n7883), .C2(n4823), .A(n4822), .B(n7882), .ZN(P2_U3160) );
  OR2_X1 U6307 ( .A1(n7592), .A2(n8351), .ZN(n4835) );
  NAND2_X1 U6308 ( .A1(n5821), .A2(n10071), .ZN(n5860) );
  NAND2_X1 U6309 ( .A1(n8000), .A2(n4839), .ZN(n4837) );
  NAND2_X1 U6310 ( .A1(n4837), .A2(n4838), .ZN(n7590) );
  AOI21_X1 U6311 ( .B1(n4839), .B2(n8001), .A(n4478), .ZN(n4838) );
  INV_X1 U6312 ( .A(n7020), .ZN(n4846) );
  NAND2_X1 U6313 ( .A1(n8024), .A2(n4847), .ZN(n7865) );
  OAI21_X1 U6314 ( .B1(n6071), .B2(n4852), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6181) );
  INV_X1 U6315 ( .A(n4848), .ZN(n6178) );
  INV_X4 U6316 ( .A(n5127), .ZN(n5047) );
  NAND3_X1 U6317 ( .A1(n4858), .A2(n5055), .A3(n4857), .ZN(n5284) );
  NAND3_X1 U6318 ( .A1(n5257), .A2(n4860), .A3(n4861), .ZN(n4857) );
  NAND3_X1 U6319 ( .A1(n5231), .A2(n4860), .A3(n5257), .ZN(n4858) );
  NAND2_X1 U6320 ( .A1(n4859), .A2(n5051), .ZN(n5258) );
  INV_X1 U6321 ( .A(n5051), .ZN(n4861) );
  INV_X1 U6322 ( .A(n5540), .ZN(n4866) );
  NAND2_X1 U6323 ( .A1(n5327), .A2(n5326), .ZN(n4875) );
  INV_X1 U6324 ( .A(n5026), .ZN(n4876) );
  AND2_X1 U6325 ( .A1(n7832), .A2(n7793), .ZN(n4878) );
  NOR2_X1 U6326 ( .A1(n7779), .A2(n8085), .ZN(n4879) );
  NAND2_X1 U6327 ( .A1(n5392), .A2(n4882), .ZN(n4880) );
  NAND2_X1 U6328 ( .A1(n4880), .A2(n4881), .ZN(n5438) );
  OR2_X1 U6329 ( .A1(n5461), .A2(n5460), .ZN(n4892) );
  NAND2_X1 U6330 ( .A1(n5461), .A2(n4890), .ZN(n4888) );
  NAND2_X1 U6331 ( .A1(n4903), .A2(n5568), .ZN(n5587) );
  NAND2_X1 U6332 ( .A1(n4904), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6333 ( .A1(n5163), .A2(n5162), .ZN(n4904) );
  INV_X1 U6334 ( .A(n8563), .ZN(n4917) );
  INV_X1 U6335 ( .A(n5474), .ZN(n4918) );
  AOI21_X1 U6336 ( .B1(n4921), .B2(n8655), .A(n9260), .ZN(n8657) );
  AND2_X1 U6337 ( .A1(n8635), .A2(n8632), .ZN(n4927) );
  OR3_X1 U6338 ( .A1(n5417), .A2(n4931), .A3(P1_IR_REG_12__SCAN_IN), .ZN(n5465) );
  AND2_X2 U6339 ( .A1(n5439), .A2(n5116), .ZN(n5462) );
  INV_X1 U6340 ( .A(n6708), .ZN(n6710) );
  NAND3_X1 U6341 ( .A1(n4935), .A2(n5185), .A3(n5184), .ZN(n6708) );
  NAND2_X1 U6342 ( .A1(n7111), .A2(n4937), .ZN(n4936) );
  NAND2_X1 U6343 ( .A1(n4936), .A2(n4939), .ZN(n7132) );
  NAND2_X1 U6344 ( .A1(n4952), .A2(n7073), .ZN(n4951) );
  OAI21_X1 U6345 ( .B1(n8962), .B2(n4961), .A(n4959), .ZN(n8933) );
  OAI21_X1 U6346 ( .B1(n8962), .B2(n8900), .A(n8902), .ZN(n8946) );
  NAND2_X2 U6347 ( .A1(n4978), .A2(n5809), .ZN(n5900) );
  NAND3_X1 U6348 ( .A1(n4978), .A2(n5809), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n5810) );
  XNOR2_X2 U6349 ( .A(n4979), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6350 ( .A1(n4981), .A2(n6678), .ZN(n7627) );
  NAND2_X1 U6351 ( .A1(n4983), .A2(n4982), .ZN(n8225) );
  NAND2_X1 U6352 ( .A1(n7269), .A2(n4988), .ZN(n4984) );
  NAND2_X1 U6353 ( .A1(n4984), .A2(n4985), .ZN(n8345) );
  OAI21_X1 U6354 ( .B1(n8291), .B2(n7809), .A(n7807), .ZN(n8281) );
  NAND2_X1 U6355 ( .A1(n7807), .A2(n7809), .ZN(n5000) );
  NAND2_X1 U6356 ( .A1(n5792), .A2(n5001), .ZN(n6182) );
  OAI21_X1 U6357 ( .B1(n8202), .B2(n5014), .A(n5012), .ZN(n7791) );
  OAI21_X1 U6358 ( .B1(n8202), .B2(n7759), .A(n7755), .ZN(n8189) );
  NAND2_X1 U6359 ( .A1(n6315), .A2(n5015), .ZN(n5014) );
  INV_X1 U6360 ( .A(n5021), .ZN(n5818) );
  NAND2_X1 U6361 ( .A1(n4467), .A2(n5293), .ZN(n6820) );
  MUX2_X1 U6362 ( .A(n7385), .B(n7384), .S(n9130), .Z(n7387) );
  NAND2_X1 U6363 ( .A1(n7211), .A2(n5371), .ZN(n7278) );
  NAND2_X1 U6364 ( .A1(n7158), .A2(n5367), .ZN(n7211) );
  NAND2_X1 U6365 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  XNOR2_X1 U6366 ( .A(n5350), .B(n5351), .ZN(n7160) );
  NAND2_X1 U6367 ( .A1(n6019), .A2(n10055), .ZN(n6071) );
  INV_X1 U6368 ( .A(n6348), .ZN(n6345) );
  NAND3_X1 U6369 ( .A1(n8693), .A2(n8695), .A3(n8692), .ZN(n8694) );
  NAND2_X1 U6370 ( .A1(n5131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6371 ( .A1(n6777), .A2(n6778), .ZN(n6779) );
  INV_X1 U6372 ( .A(n6722), .ZN(n5142) );
  NAND2_X1 U6373 ( .A1(n5845), .A2(n5047), .ZN(n5864) );
  INV_X1 U6374 ( .A(n5139), .ZN(n5140) );
  AND2_X1 U6375 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  INV_X1 U6376 ( .A(n6213), .ZN(n6413) );
  NOR2_X1 U6377 ( .A1(n8522), .A2(n8338), .ZN(n5022) );
  NOR2_X1 U6378 ( .A1(n5504), .A2(n5503), .ZN(n5023) );
  OR2_X1 U6379 ( .A1(n5845), .A2(n6642), .ZN(n5024) );
  AND4_X1 U6380 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n7853)
         );
  AND2_X1 U6381 ( .A1(n5072), .A2(n5071), .ZN(n5026) );
  INV_X1 U6382 ( .A(n8859), .ZN(n8697) );
  INV_X1 U6383 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5036) );
  INV_X1 U6384 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5756) );
  AND2_X1 U6385 ( .A1(n7507), .A2(n7506), .ZN(n5027) );
  NAND2_X1 U6386 ( .A1(n6070), .A2(n6069), .ZN(n5028) );
  XNOR2_X1 U6387 ( .A(n7877), .B(n9766), .ZN(n6777) );
  AND2_X1 U6388 ( .A1(n8008), .A2(n8007), .ZN(n5029) );
  INV_X1 U6389 ( .A(n8717), .ZN(n5768) );
  OR2_X1 U6390 ( .A1(n5235), .A2(n6444), .ZN(n5030) );
  NAND2_X1 U6391 ( .A1(n7429), .A2(n4724), .ZN(n7406) );
  INV_X1 U6392 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5118) );
  AND2_X1 U6393 ( .A1(n8092), .A2(n7023), .ZN(n5898) );
  NOR2_X1 U6394 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  NOR2_X1 U6395 ( .A1(n5898), .A2(n5897), .ZN(n7102) );
  INV_X1 U6396 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5791) );
  INV_X1 U6397 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5115) );
  OR2_X1 U6398 ( .A1(n7572), .A2(n8090), .ZN(n7573) );
  INV_X1 U6399 ( .A(n7576), .ZN(n7577) );
  INV_X1 U6400 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10107) );
  OR2_X1 U6401 ( .A1(n5601), .A2(n5600), .ZN(n5602) );
  INV_X1 U6402 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5336) );
  AND2_X1 U6403 ( .A1(n5121), .A2(n5124), .ZN(n5122) );
  INV_X1 U6404 ( .A(SI_22_), .ZN(n5606) );
  NAND2_X1 U6405 ( .A1(n5047), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5035) );
  INV_X1 U6406 ( .A(n7198), .ZN(n7194) );
  INV_X1 U6407 ( .A(n4415), .ZN(n6778) );
  OR2_X1 U6408 ( .A1(n7960), .A2(n8329), .ZN(n7596) );
  INV_X1 U6409 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5421) );
  INV_X1 U6410 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5482) );
  INV_X1 U6411 ( .A(n8721), .ZN(n8901) );
  AOI21_X1 U6412 ( .B1(n6396), .B2(n6404), .A(n6402), .ZN(n9120) );
  NAND2_X1 U6413 ( .A1(n8737), .A2(n9484), .ZN(n7516) );
  INV_X1 U6414 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6415 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  AND2_X1 U6416 ( .A1(n6624), .A2(n6623), .ZN(n8058) );
  NAND2_X1 U6417 ( .A1(n7593), .A2(n8338), .ZN(n7595) );
  INV_X1 U6418 ( .A(n7969), .ZN(n7599) );
  INV_X1 U6419 ( .A(n8058), .ZN(n8075) );
  INV_X1 U6420 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7945) );
  INV_X1 U6421 ( .A(n8145), .ZN(n8158) );
  OR2_X1 U6422 ( .A1(n9821), .A2(n9767), .ZN(n8341) );
  NAND2_X1 U6423 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  AND2_X1 U6424 ( .A1(n7783), .A2(n6217), .ZN(n6277) );
  AND2_X1 U6425 ( .A1(n7676), .A2(n7668), .ZN(n7817) );
  AND2_X1 U6426 ( .A1(n6783), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6597) );
  INV_X1 U6427 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8565) );
  AND2_X1 U6428 ( .A1(n5739), .A2(n5740), .ZN(n5738) );
  NOR2_X1 U6429 ( .A1(n10182), .A2(n5612), .ZN(n5629) );
  AND3_X1 U6430 ( .A1(n5770), .A2(n6407), .A3(n5166), .ZN(n6718) );
  NOR2_X1 U6431 ( .A1(n5483), .A2(n5482), .ZN(n5502) );
  NOR2_X1 U6432 ( .A1(n7504), .A2(n7503), .ZN(n7509) );
  NOR2_X1 U6433 ( .A1(n5574), .A2(n8668), .ZN(n5591) );
  INV_X1 U6434 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9975) );
  INV_X1 U6435 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10006) );
  INV_X1 U6436 ( .A(n8861), .ZN(n8856) );
  INV_X1 U6437 ( .A(n9187), .ZN(n9083) );
  NAND2_X1 U6438 ( .A1(n9445), .A2(n5160), .ZN(n9101) );
  INV_X1 U6439 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5745) );
  XNOR2_X1 U6440 ( .A(n5141), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5742) );
  NAND3_X1 U6441 ( .A1(n6413), .A2(n6219), .A3(n6412), .ZN(n6590) );
  OR2_X1 U6442 ( .A1(n6608), .A2(n6623), .ZN(n8061) );
  INV_X1 U6443 ( .A(n8061), .ZN(n8073) );
  XNOR2_X1 U6444 ( .A(n6221), .B(n5020), .ZN(n6783) );
  AND3_X1 U6445 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n7984) );
  AND4_X1 U6446 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n7975)
         );
  INV_X1 U6447 ( .A(n9597), .ZN(n10207) );
  INV_X1 U6448 ( .A(n10217), .ZN(n9740) );
  INV_X1 U6449 ( .A(n8341), .ZN(n8358) );
  INV_X1 U6450 ( .A(n8381), .ZN(n8361) );
  OAI211_X1 U6451 ( .C1(n6274), .C2(n6277), .A(n6281), .B(n6237), .ZN(n6268)
         );
  OAI21_X1 U6452 ( .B1(n8454), .B2(n8422), .A(n6283), .ZN(n6284) );
  INV_X1 U6453 ( .A(n8383), .ZN(n8428) );
  AND3_X1 U6454 ( .A1(n6588), .A2(n6330), .A3(n6329), .ZN(n6281) );
  INV_X1 U6455 ( .A(n8433), .ZN(n8534) );
  NAND2_X1 U6456 ( .A1(n7257), .A2(n9808), .ZN(n9819) );
  AND2_X1 U6457 ( .A1(n9767), .A2(n7274), .ZN(n9794) );
  INV_X1 U6458 ( .A(n6214), .ZN(n6412) );
  INV_X1 U6459 ( .A(n6222), .ZN(n6409) );
  INV_X1 U6460 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5908) );
  AND2_X1 U6461 ( .A1(n5728), .A2(n5727), .ZN(n8698) );
  AND2_X1 U6462 ( .A1(n5614), .A2(n5613), .ZN(n8892) );
  OR2_X1 U6463 ( .A1(n9291), .A2(n8752), .ZN(n9368) );
  INV_X1 U6464 ( .A(n9389), .ZN(n9347) );
  XNOR2_X1 U6465 ( .A(n8864), .B(n8856), .ZN(n8857) );
  AND2_X1 U6466 ( .A1(n7467), .A2(n8921), .ZN(n8969) );
  INV_X1 U6467 ( .A(n8915), .ZN(n9019) );
  AND2_X1 U6468 ( .A1(n7448), .A2(n7447), .ZN(n9074) );
  INV_X1 U6469 ( .A(n9104), .ZN(n9431) );
  AOI21_X1 U6470 ( .B1(n6396), .B2(n5745), .A(n6398), .ZN(n9125) );
  INV_X1 U6471 ( .A(n9106), .ZN(n9196) );
  AND2_X1 U6472 ( .A1(n5743), .A2(n5742), .ZN(n6396) );
  INV_X1 U6473 ( .A(n7620), .ZN(n6686) );
  INV_X1 U6474 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6475 ( .A1(n6590), .A2(n6411), .ZN(n6647) );
  INV_X1 U6476 ( .A(n8078), .ZN(n8053) );
  INV_X1 U6477 ( .A(n7853), .ZN(n8274) );
  OR2_X1 U6478 ( .A1(P2_U3150), .A2(n6649), .ZN(n10217) );
  INV_X1 U6479 ( .A(n10209), .ZN(n9754) );
  NAND2_X1 U6480 ( .A1(n6269), .A2(n8358), .ZN(n8180) );
  AND2_X1 U6481 ( .A1(n7266), .A2(n7265), .ZN(n9825) );
  AND2_X2 U6482 ( .A1(n6268), .A2(n8373), .ZN(n9773) );
  NOR2_X1 U6483 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  NAND2_X1 U6484 ( .A1(n9851), .A2(n9819), .ZN(n8422) );
  AND3_X2 U6485 ( .A1(n6281), .A2(n6280), .A3(n6279), .ZN(n9851) );
  NAND2_X1 U6486 ( .A1(n8450), .A2(n8449), .ZN(n8453) );
  OR2_X1 U6487 ( .A1(n9835), .A2(n9827), .ZN(n8518) );
  AND3_X1 U6488 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9848) );
  AND2_X1 U6489 ( .A1(n6332), .A2(n6331), .ZN(n9835) );
  NAND2_X1 U6490 ( .A1(n6236), .A2(n6235), .ZN(n6423) );
  INV_X1 U6491 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8558) );
  INV_X1 U6492 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6951) );
  INV_X1 U6493 ( .A(n9629), .ZN(n8126) );
  AND2_X1 U6494 ( .A1(n6408), .A2(n6437), .ZN(n9305) );
  INV_X1 U6495 ( .A(n9172), .ZN(n9043) );
  INV_X1 U6496 ( .A(n9157), .ZN(n9000) );
  NAND2_X1 U6497 ( .A1(n5772), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9267) );
  AND2_X1 U6498 ( .A1(n5767), .A2(n7121), .ZN(n8717) );
  OR2_X1 U6499 ( .A1(n9291), .A2(n8750), .ZN(n9389) );
  NAND2_X1 U6500 ( .A1(n9452), .A2(n9109), .ZN(n9086) );
  INV_X1 U6501 ( .A(n9575), .ZN(n9573) );
  INV_X1 U6502 ( .A(n9553), .ZN(n9551) );
  INV_X1 U6503 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6404) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9229) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7288) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U6507 ( .A1(n6273), .A2(n6272), .ZN(P2_U3206) );
  OAI21_X1 U6508 ( .B1(n6369), .B2(n9849), .A(n6368), .ZN(P2_U3488) );
  AND2_X2 U6509 ( .A1(n6407), .A2(n6370), .ZN(P1_U3973) );
  INV_X1 U6510 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6376) );
  INV_X1 U6511 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U6512 ( .A1(n5031), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6513 ( .A1(n5032), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5033) );
  MUX2_X1 U6514 ( .A(n6376), .B(n6386), .S(n5127), .Z(n5039) );
  NAND2_X1 U6515 ( .A1(n5037), .A2(SI_0_), .ZN(n5188) );
  INV_X1 U6516 ( .A(n5188), .ZN(n5038) );
  NAND2_X1 U6517 ( .A1(n5189), .A2(n5038), .ZN(n5042) );
  INV_X1 U6518 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6519 ( .A1(n5040), .A2(SI_1_), .ZN(n5041) );
  NAND2_X1 U6520 ( .A1(n5042), .A2(n5041), .ZN(n5211) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6375) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U6523 ( .A1(n5211), .A2(n5212), .ZN(n5046) );
  INV_X1 U6524 ( .A(n5043), .ZN(n5044) );
  NAND2_X1 U6525 ( .A1(n5044), .A2(SI_2_), .ZN(n5045) );
  INV_X1 U6526 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10034) );
  INV_X1 U6527 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6378) );
  XNOR2_X1 U6528 ( .A(n5049), .B(SI_3_), .ZN(n5230) );
  INV_X1 U6529 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6530 ( .A1(n5050), .A2(SI_3_), .ZN(n5051) );
  BUF_X4 U6531 ( .A(n5047), .Z(n5523) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6384) );
  XNOR2_X1 U6533 ( .A(n5053), .B(SI_4_), .ZN(n5257) );
  INV_X1 U6534 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6535 ( .A1(n5054), .A2(SI_4_), .ZN(n5055) );
  MUX2_X1 U6536 ( .A(n6380), .B(n6382), .S(n5047), .Z(n5056) );
  XNOR2_X1 U6537 ( .A(n5056), .B(SI_5_), .ZN(n5283) );
  NAND2_X1 U6538 ( .A1(n5284), .A2(n5283), .ZN(n5059) );
  INV_X1 U6539 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6540 ( .A1(n5057), .A2(SI_5_), .ZN(n5058) );
  MUX2_X1 U6541 ( .A(n6387), .B(n6389), .S(n5047), .Z(n5060) );
  XNOR2_X1 U6542 ( .A(n5060), .B(SI_6_), .ZN(n5306) );
  NAND2_X1 U6543 ( .A1(n5307), .A2(n5306), .ZN(n5063) );
  INV_X1 U6544 ( .A(n5060), .ZN(n5061) );
  NAND2_X1 U6545 ( .A1(n5061), .A2(SI_6_), .ZN(n5062) );
  MUX2_X1 U6546 ( .A(n6391), .B(n6390), .S(n5523), .Z(n5064) );
  XNOR2_X1 U6547 ( .A(n5064), .B(SI_7_), .ZN(n5326) );
  INV_X1 U6548 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6549 ( .A1(n5065), .A2(SI_7_), .ZN(n5066) );
  INV_X1 U6550 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6394) );
  INV_X1 U6551 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5067) );
  MUX2_X1 U6552 ( .A(n6394), .B(n5067), .S(n5523), .Z(n5069) );
  INV_X1 U6553 ( .A(SI_8_), .ZN(n5068) );
  NAND2_X1 U6554 ( .A1(n5069), .A2(n5068), .ZN(n5072) );
  INV_X1 U6555 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6556 ( .A1(n5070), .A2(SI_8_), .ZN(n5071) );
  INV_X1 U6557 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6399) );
  MUX2_X1 U6558 ( .A(n6400), .B(n6399), .S(n5523), .Z(n5074) );
  INV_X1 U6559 ( .A(SI_9_), .ZN(n5073) );
  NAND2_X1 U6560 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  INV_X1 U6561 ( .A(n5074), .ZN(n5075) );
  NAND2_X1 U6562 ( .A1(n5075), .A2(SI_9_), .ZN(n5076) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6426) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6425) );
  MUX2_X1 U6565 ( .A(n6426), .B(n6425), .S(n5523), .Z(n5079) );
  XNOR2_X1 U6566 ( .A(n5079), .B(SI_10_), .ZN(n5372) );
  INV_X1 U6567 ( .A(n5372), .ZN(n5078) );
  INV_X1 U6568 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6569 ( .A1(n5080), .A2(SI_10_), .ZN(n5081) );
  INV_X1 U6570 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5082) );
  MUX2_X1 U6571 ( .A(n10106), .B(n5082), .S(n5523), .Z(n5084) );
  INV_X1 U6572 ( .A(SI_11_), .ZN(n5083) );
  NAND2_X1 U6573 ( .A1(n5084), .A2(n5083), .ZN(n5087) );
  INV_X1 U6574 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6575 ( .A1(n5085), .A2(SI_11_), .ZN(n5086) );
  NAND2_X1 U6576 ( .A1(n5087), .A2(n5086), .ZN(n5391) );
  MUX2_X1 U6577 ( .A(n10152), .B(n10070), .S(n5523), .Z(n5088) );
  XNOR2_X1 U6578 ( .A(n5088), .B(SI_12_), .ZN(n5415) );
  INV_X1 U6579 ( .A(n5415), .ZN(n5090) );
  INV_X1 U6580 ( .A(n5088), .ZN(n5089) );
  MUX2_X1 U6581 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5523), .Z(n5092) );
  XNOR2_X1 U6582 ( .A(n5092), .B(SI_13_), .ZN(n5437) );
  INV_X1 U6583 ( .A(n5437), .ZN(n5091) );
  NAND2_X1 U6584 ( .A1(n5438), .A2(n5091), .ZN(n5094) );
  NAND2_X1 U6585 ( .A1(n5092), .A2(SI_13_), .ZN(n5093) );
  MUX2_X1 U6586 ( .A(n6551), .B(n5095), .S(n5523), .Z(n5097) );
  NAND2_X1 U6587 ( .A1(n5097), .A2(n5096), .ZN(n5100) );
  INV_X1 U6588 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6589 ( .A1(n5098), .A2(SI_14_), .ZN(n5099) );
  NAND2_X1 U6590 ( .A1(n5100), .A2(n5099), .ZN(n5460) );
  MUX2_X1 U6591 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5523), .Z(n5476) );
  INV_X1 U6592 ( .A(n5476), .ZN(n5101) );
  NAND2_X1 U6593 ( .A1(n5102), .A2(SI_16_), .ZN(n5105) );
  INV_X1 U6594 ( .A(SI_16_), .ZN(n5493) );
  MUX2_X1 U6595 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5523), .Z(n5494) );
  NAND2_X1 U6596 ( .A1(n5103), .A2(n5494), .ZN(n5104) );
  MUX2_X1 U6597 ( .A(n6775), .B(n5106), .S(n5523), .Z(n5108) );
  NAND2_X1 U6598 ( .A1(n5108), .A2(n5107), .ZN(n5520) );
  INV_X1 U6599 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6600 ( .A1(n5109), .A2(SI_17_), .ZN(n5110) );
  NAND2_X1 U6601 ( .A1(n5520), .A2(n5110), .ZN(n5521) );
  XNOR2_X1 U6602 ( .A(n5522), .B(n5521), .ZN(n6685) );
  NOR2_X1 U6603 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5114) );
  NAND2_X1 U6604 ( .A1(n5139), .A2(n5124), .ZN(n5125) );
  NAND2_X1 U6605 ( .A1(n6685), .A2(n7420), .ZN(n5129) );
  NAND2_X4 U6606 ( .A1(n5235), .A2(n4418), .ZN(n5259) );
  NAND2_X1 U6607 ( .A1(n5497), .A2(n5118), .ZN(n5131) );
  XNOR2_X1 U6608 ( .A(n5154), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8813) );
  AOI22_X1 U6609 ( .A1(n5551), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5550), .B2(
        n8813), .ZN(n5128) );
  NAND2_X1 U6610 ( .A1(n5129), .A2(n5128), .ZN(n8880) );
  NAND3_X1 U6611 ( .A1(n5153), .A2(n5156), .A3(n5158), .ZN(n5130) );
  NAND2_X1 U6612 ( .A1(n5134), .A2(n5135), .ZN(n5161) );
  NAND2_X1 U6613 ( .A1(n4473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  AND2_X2 U6614 ( .A1(n5142), .A2(n5166), .ZN(n5167) );
  INV_X1 U6615 ( .A(n5143), .ZN(n5144) );
  NAND2_X1 U6616 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5145) );
  NAND2_X1 U6617 ( .A1(n6416), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5152) );
  INV_X1 U6618 ( .A(n5147), .ZN(n7568) );
  NAND2_X1 U6619 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5274) );
  INV_X1 U6620 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5273) );
  NOR2_X1 U6621 ( .A1(n5274), .A2(n5273), .ZN(n5295) );
  NAND2_X1 U6622 ( .A1(n5295), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6623 ( .A1(n5381), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6624 ( .A1(n5444), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6625 ( .A1(n5504), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5527) );
  OR2_X1 U6626 ( .A1(n5504), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5148) );
  AND2_X1 U6627 ( .A1(n5527), .A2(n5148), .ZN(n9095) );
  NAND2_X1 U6628 ( .A1(n6352), .A2(n9095), .ZN(n5151) );
  NAND2_X1 U6629 ( .A1(n7423), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6630 ( .A1(n5248), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5149) );
  NAND4_X1 U6631 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n8726)
         );
  INV_X1 U6632 ( .A(n8726), .ZN(n8877) );
  NAND2_X1 U6633 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  NAND2_X1 U6634 ( .A1(n5524), .A2(n5156), .ZN(n5157) );
  INV_X1 U6635 ( .A(n6721), .ZN(n7556) );
  OR2_X1 U6636 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  NAND2_X1 U6637 ( .A1(n7556), .A2(n7563), .ZN(n5165) );
  NAND3_X2 U6638 ( .A1(n5165), .A2(n5166), .A3(n6941), .ZN(n5731) );
  OAI22_X1 U6639 ( .A1(n9270), .A2(n5732), .B1(n8877), .B2(n5731), .ZN(n5513)
         );
  INV_X1 U6640 ( .A(n5513), .ZN(n5519) );
  NAND2_X1 U6641 ( .A1(n8880), .A2(n6342), .ZN(n5169) );
  NAND2_X1 U6642 ( .A1(n8726), .A2(n6336), .ZN(n5168) );
  NAND2_X1 U6643 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  XNOR2_X1 U6644 ( .A(n5170), .B(n4419), .ZN(n5512) );
  INV_X1 U6645 ( .A(n5512), .ZN(n5518) );
  NAND2_X1 U6646 ( .A1(n5202), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6647 ( .A1(n5201), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6648 ( .A1(n5248), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6649 ( .A1(n5203), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5171) );
  INV_X2 U6650 ( .A(n5731), .ZN(n6337) );
  NAND2_X1 U6651 ( .A1(n6709), .A2(n6337), .ZN(n5179) );
  INV_X1 U6652 ( .A(SI_0_), .ZN(n5175) );
  NOR2_X1 U6653 ( .A1(n4418), .A2(n5175), .ZN(n5177) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5176) );
  XNOR2_X1 U6655 ( .A(n5177), .B(n5176), .ZN(n9237) );
  INV_X1 U6656 ( .A(n5166), .ZN(n5180) );
  AOI22_X1 U6657 ( .A1(n9446), .A2(n5167), .B1(n5180), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6658 ( .A1(n5179), .A2(n5178), .ZN(n6530) );
  NAND2_X1 U6659 ( .A1(n5180), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U6660 ( .A1(n5182), .A2(n5181), .ZN(n6531) );
  NAND2_X1 U6661 ( .A1(n6530), .A2(n6531), .ZN(n6529) );
  NAND2_X1 U6662 ( .A1(n5182), .A2(n5662), .ZN(n5183) );
  AND2_X1 U6663 ( .A1(n6529), .A2(n5183), .ZN(n6542) );
  NAND2_X1 U6664 ( .A1(n5203), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6665 ( .A1(n5201), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6666 ( .A1(n6708), .A2(n5167), .ZN(n5194) );
  INV_X1 U6667 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6668 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5186) );
  XNOR2_X1 U6669 ( .A(n5187), .B(n5186), .ZN(n6444) );
  XNOR2_X1 U6670 ( .A(n5189), .B(n5188), .ZN(n5819) );
  INV_X1 U6671 ( .A(n5819), .ZN(n6385) );
  OR2_X1 U6672 ( .A1(n5232), .A2(n6385), .ZN(n5190) );
  NAND2_X1 U6673 ( .A1(n5192), .A2(n6945), .ZN(n5193) );
  NAND2_X1 U6674 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  XNOR2_X1 U6675 ( .A(n5195), .B(n4419), .ZN(n5197) );
  AND2_X1 U6676 ( .A1(n6945), .A2(n5167), .ZN(n5196) );
  XNOR2_X1 U6677 ( .A(n5197), .B(n5198), .ZN(n6543) );
  NAND2_X1 U6678 ( .A1(n6542), .A2(n6543), .ZN(n6541) );
  INV_X1 U6679 ( .A(n5197), .ZN(n5199) );
  NAND2_X1 U6680 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6681 ( .A1(n6541), .A2(n5200), .ZN(n6566) );
  NAND2_X1 U6682 ( .A1(n5201), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6683 ( .A1(n5202), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6684 ( .A1(n5203), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6685 ( .A1(n5248), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5204) );
  NAND4_X1 U6686 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n8739)
         );
  NAND2_X1 U6687 ( .A1(n8739), .A2(n5167), .ZN(n5216) );
  OR2_X1 U6688 ( .A1(n5208), .A2(n4688), .ZN(n5210) );
  XNOR2_X1 U6689 ( .A(n5210), .B(n5209), .ZN(n6446) );
  XNOR2_X1 U6690 ( .A(n5212), .B(n5211), .ZN(n6374) );
  OR2_X1 U6691 ( .A1(n5232), .A2(n6374), .ZN(n5213) );
  NAND2_X1 U6692 ( .A1(n6891), .A2(n5287), .ZN(n5215) );
  NAND2_X1 U6693 ( .A1(n5216), .A2(n5215), .ZN(n5217) );
  XNOR2_X1 U6694 ( .A(n5217), .B(n4419), .ZN(n5220) );
  AND2_X1 U6695 ( .A1(n6891), .A2(n5167), .ZN(n5219) );
  AOI21_X1 U6696 ( .B1(n8739), .B2(n6337), .A(n5219), .ZN(n5221) );
  XNOR2_X1 U6697 ( .A(n5220), .B(n5221), .ZN(n6567) );
  NAND2_X1 U6698 ( .A1(n6566), .A2(n6567), .ZN(n5224) );
  INV_X1 U6699 ( .A(n5220), .ZN(n5222) );
  NAND2_X1 U6700 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6701 ( .A1(n5224), .A2(n5223), .ZN(n6579) );
  INV_X1 U6702 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6703 ( .A1(n6352), .A2(n5246), .ZN(n5228) );
  NAND2_X1 U6704 ( .A1(n5201), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6705 ( .A1(n5248), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6706 ( .A1(n7423), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6707 ( .A1(n8738), .A2(n5711), .ZN(n5237) );
  INV_X1 U6708 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5229) );
  XNOR2_X1 U6709 ( .A(n5231), .B(n5230), .ZN(n6377) );
  OR2_X1 U6710 ( .A1(n5232), .A2(n6377), .ZN(n5234) );
  OR2_X1 U6711 ( .A1(n5259), .A2(n6378), .ZN(n5233) );
  OAI211_X1 U6712 ( .C1(n5235), .C2(n8772), .A(n5234), .B(n5233), .ZN(n9478)
         );
  NAND2_X1 U6713 ( .A1(n9478), .A2(n5287), .ZN(n5236) );
  NAND2_X1 U6714 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  XNOR2_X1 U6715 ( .A(n5238), .B(n4419), .ZN(n5240) );
  AND2_X1 U6716 ( .A1(n9478), .A2(n6336), .ZN(n5239) );
  AOI21_X1 U6717 ( .B1(n8738), .B2(n6337), .A(n5239), .ZN(n5241) );
  XNOR2_X1 U6718 ( .A(n5240), .B(n5241), .ZN(n6580) );
  INV_X1 U6719 ( .A(n5240), .ZN(n5242) );
  NAND2_X1 U6720 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6721 ( .A1(n5201), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5252) );
  INV_X1 U6722 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6723 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  AND2_X1 U6724 ( .A1(n5247), .A2(n5274), .ZN(n9430) );
  NAND2_X1 U6725 ( .A1(n6352), .A2(n9430), .ZN(n5251) );
  NAND2_X1 U6726 ( .A1(n7423), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6727 ( .A1(n5248), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5249) );
  NAND4_X1 U6728 ( .A1(n5252), .A2(n5251), .A3(n5250), .A4(n5249), .ZN(n8737)
         );
  NAND2_X1 U6729 ( .A1(n8737), .A2(n5711), .ZN(n5263) );
  NOR2_X1 U6730 ( .A1(n5253), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5302) );
  OR2_X1 U6731 ( .A1(n5302), .A2(n4688), .ZN(n5255) );
  INV_X1 U6732 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6733 ( .A1(n5255), .A2(n5254), .ZN(n5280) );
  OR2_X1 U6734 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U6735 ( .A1(n5280), .A2(n5256), .ZN(n8783) );
  XNOR2_X1 U6736 ( .A(n5258), .B(n5257), .ZN(n6383) );
  OR2_X1 U6737 ( .A1(n5259), .A2(n6379), .ZN(n5260) );
  NAND2_X1 U6738 ( .A1(n9432), .A2(n5287), .ZN(n5262) );
  NAND2_X1 U6739 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  XNOR2_X1 U6740 ( .A(n5264), .B(n4419), .ZN(n5267) );
  NAND2_X1 U6741 ( .A1(n8737), .A2(n6337), .ZN(n5266) );
  NAND2_X1 U6742 ( .A1(n9432), .A2(n5711), .ZN(n5265) );
  NAND2_X1 U6743 ( .A1(n5266), .A2(n5265), .ZN(n5268) );
  NAND2_X1 U6744 ( .A1(n5267), .A2(n5268), .ZN(n5272) );
  INV_X1 U6745 ( .A(n5267), .ZN(n5270) );
  INV_X1 U6746 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6747 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  NAND2_X1 U6748 ( .A1(n5272), .A2(n5271), .ZN(n8655) );
  NAND2_X1 U6749 ( .A1(n5201), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6750 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  NOR2_X1 U6751 ( .A1(n5295), .A2(n5275), .ZN(n6927) );
  NAND2_X1 U6752 ( .A1(n6352), .A2(n6927), .ZN(n5278) );
  NAND2_X1 U6753 ( .A1(n5248), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6754 ( .A1(n7423), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5276) );
  NAND4_X1 U6755 ( .A1(n5279), .A2(n5278), .A3(n5277), .A4(n5276), .ZN(n8736)
         );
  NAND2_X1 U6756 ( .A1(n8736), .A2(n6336), .ZN(n5289) );
  NAND2_X1 U6757 ( .A1(n5280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5282) );
  INV_X1 U6758 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5281) );
  XNOR2_X1 U6759 ( .A(n5282), .B(n5281), .ZN(n6476) );
  XNOR2_X1 U6760 ( .A(n5284), .B(n5283), .ZN(n6381) );
  OR2_X1 U6761 ( .A1(n5232), .A2(n6381), .ZN(n5286) );
  OR2_X1 U6762 ( .A1(n5259), .A2(n6382), .ZN(n5285) );
  OAI211_X1 U6763 ( .C1(n5235), .C2(n6476), .A(n5286), .B(n5285), .ZN(n6928)
         );
  NAND2_X1 U6764 ( .A1(n6928), .A2(n5287), .ZN(n5288) );
  NAND2_X1 U6765 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  XNOR2_X1 U6766 ( .A(n5290), .B(n4419), .ZN(n5292) );
  AND2_X1 U6767 ( .A1(n6928), .A2(n6336), .ZN(n5291) );
  AOI21_X1 U6768 ( .B1(n8736), .B2(n6337), .A(n5291), .ZN(n6821) );
  NAND2_X1 U6769 ( .A1(n6819), .A2(n6821), .ZN(n5294) );
  INV_X1 U6770 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6771 ( .A1(n5201), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6772 ( .A1(n5295), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5296) );
  AND2_X1 U6773 ( .A1(n5318), .A2(n5296), .ZN(n6845) );
  NAND2_X1 U6774 ( .A1(n6352), .A2(n6845), .ZN(n5299) );
  NAND2_X1 U6775 ( .A1(n7423), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6776 ( .A1(n5248), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5297) );
  NAND4_X1 U6777 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n8735)
         );
  NAND2_X1 U6778 ( .A1(n8735), .A2(n6336), .ZN(n5311) );
  NOR2_X1 U6779 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5301) );
  NAND2_X1 U6780 ( .A1(n5302), .A2(n5301), .ZN(n5304) );
  NAND2_X1 U6781 ( .A1(n5304), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5303) );
  MUX2_X1 U6782 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5303), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5305) );
  NAND2_X1 U6783 ( .A1(n5305), .A2(n5344), .ZN(n6489) );
  XNOR2_X1 U6784 ( .A(n5307), .B(n5306), .ZN(n6388) );
  OR2_X1 U6785 ( .A1(n5232), .A2(n6388), .ZN(n5309) );
  OR2_X1 U6786 ( .A1(n5259), .A2(n6389), .ZN(n5308) );
  OAI211_X1 U6787 ( .C1(n5235), .C2(n6489), .A(n5309), .B(n5308), .ZN(n9497)
         );
  NAND2_X1 U6788 ( .A1(n9497), .A2(n5287), .ZN(n5310) );
  NAND2_X1 U6789 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  XNOR2_X1 U6790 ( .A(n5312), .B(n4419), .ZN(n5314) );
  AND2_X1 U6791 ( .A1(n9497), .A2(n5711), .ZN(n5313) );
  AOI21_X1 U6792 ( .B1(n8735), .B2(n6337), .A(n5313), .ZN(n5315) );
  XNOR2_X1 U6793 ( .A(n5314), .B(n5315), .ZN(n6875) );
  INV_X1 U6794 ( .A(n5314), .ZN(n5316) );
  NAND2_X1 U6795 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6796 ( .A1(n6416), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6797 ( .A1(n5318), .A2(n6956), .ZN(n5319) );
  AND2_X1 U6798 ( .A1(n5337), .A2(n5319), .ZN(n7120) );
  NAND2_X1 U6799 ( .A1(n6352), .A2(n7120), .ZN(n5322) );
  NAND2_X1 U6800 ( .A1(n7423), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6801 ( .A1(n5248), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5320) );
  NAND4_X1 U6802 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n8734)
         );
  NAND2_X1 U6803 ( .A1(n8734), .A2(n5711), .ZN(n5331) );
  NAND2_X1 U6804 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5325) );
  INV_X1 U6805 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5324) );
  XNOR2_X1 U6806 ( .A(n5325), .B(n5324), .ZN(n6509) );
  XNOR2_X1 U6807 ( .A(n5327), .B(n5326), .ZN(n6392) );
  OR2_X1 U6808 ( .A1(n5232), .A2(n6392), .ZN(n5329) );
  OR2_X1 U6809 ( .A1(n5259), .A2(n6390), .ZN(n5328) );
  OAI211_X1 U6810 ( .C1(n5235), .C2(n6509), .A(n5329), .B(n5328), .ZN(n9506)
         );
  NAND2_X1 U6811 ( .A1(n9506), .A2(n6342), .ZN(n5330) );
  NAND2_X1 U6812 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  XNOR2_X1 U6813 ( .A(n5332), .B(n5662), .ZN(n6954) );
  AND2_X1 U6814 ( .A1(n9506), .A2(n5711), .ZN(n5333) );
  AOI21_X1 U6815 ( .B1(n8734), .B2(n6337), .A(n5333), .ZN(n6953) );
  INV_X1 U6816 ( .A(n6954), .ZN(n5335) );
  INV_X1 U6817 ( .A(n6953), .ZN(n5334) );
  NAND2_X1 U6818 ( .A1(n6416), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6819 ( .A1(n5337), .A2(n5336), .ZN(n5338) );
  NAND2_X1 U6820 ( .A1(n5358), .A2(n5338), .ZN(n7165) );
  INV_X1 U6821 ( .A(n7165), .ZN(n9419) );
  NAND2_X1 U6822 ( .A1(n6352), .A2(n9419), .ZN(n5341) );
  NAND2_X1 U6823 ( .A1(n7423), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6824 ( .A1(n5248), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5339) );
  NAND4_X1 U6825 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n8733)
         );
  NAND2_X1 U6826 ( .A1(n8733), .A2(n6336), .ZN(n5348) );
  XNOR2_X1 U6827 ( .A(n5343), .B(n5026), .ZN(n6395) );
  OR2_X1 U6828 ( .A1(n6395), .A2(n5232), .ZN(n5346) );
  NAND2_X1 U6829 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5353) );
  XNOR2_X1 U6830 ( .A(n5353), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U6831 ( .A1(n5551), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5550), .B2(
        n6520), .ZN(n5345) );
  NAND2_X1 U6832 ( .A1(n5346), .A2(n5345), .ZN(n9420) );
  NAND2_X1 U6833 ( .A1(n9420), .A2(n5192), .ZN(n5347) );
  NAND2_X1 U6834 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  XNOR2_X1 U6835 ( .A(n5349), .B(n5662), .ZN(n5351) );
  AOI22_X1 U6836 ( .A1(n8733), .A2(n6337), .B1(n6336), .B2(n9420), .ZN(n7159)
         );
  INV_X1 U6837 ( .A(n5350), .ZN(n5352) );
  NAND2_X1 U6838 ( .A1(n5352), .A2(n5351), .ZN(n7210) );
  OR2_X1 U6839 ( .A1(n6401), .A2(n5232), .ZN(n5357) );
  INV_X1 U6840 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6841 ( .A1(n5353), .A2(n5375), .ZN(n5354) );
  NAND2_X1 U6842 ( .A1(n5354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5355) );
  XNOR2_X1 U6843 ( .A(n5355), .B(P1_IR_REG_9__SCAN_IN), .ZN(n8818) );
  AOI22_X1 U6844 ( .A1(n5551), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5550), .B2(
        n8818), .ZN(n5356) );
  NAND2_X1 U6845 ( .A1(n5357), .A2(n5356), .ZN(n7136) );
  NAND2_X1 U6846 ( .A1(n7136), .A2(n5192), .ZN(n5365) );
  NAND2_X1 U6847 ( .A1(n6416), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5363) );
  AND2_X1 U6848 ( .A1(n5358), .A2(n9975), .ZN(n5359) );
  NOR2_X1 U6849 ( .A1(n5381), .A2(n5359), .ZN(n7218) );
  NAND2_X1 U6850 ( .A1(n6352), .A2(n7218), .ZN(n5362) );
  NAND2_X1 U6851 ( .A1(n7423), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6852 ( .A1(n5248), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5360) );
  NAND4_X1 U6853 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n8732)
         );
  NAND2_X1 U6854 ( .A1(n8732), .A2(n6336), .ZN(n5364) );
  NAND2_X1 U6855 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  XNOR2_X1 U6856 ( .A(n5366), .B(n4419), .ZN(n5368) );
  AOI22_X1 U6857 ( .A1(n7136), .A2(n5711), .B1(n8732), .B2(n6337), .ZN(n5369)
         );
  XNOR2_X1 U6858 ( .A(n5368), .B(n5369), .ZN(n7212) );
  AND2_X1 U6859 ( .A1(n7210), .A2(n7212), .ZN(n5367) );
  INV_X1 U6860 ( .A(n5368), .ZN(n5370) );
  OR2_X1 U6861 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  XNOR2_X1 U6862 ( .A(n5373), .B(n5372), .ZN(n6424) );
  NAND2_X1 U6863 ( .A1(n6424), .A2(n7420), .ZN(n5380) );
  INV_X1 U6864 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6865 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  OAI21_X1 U6866 ( .B1(n5377), .B2(n5376), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5378) );
  XNOR2_X1 U6867 ( .A(n5378), .B(P1_IR_REG_10__SCAN_IN), .ZN(n8819) );
  AOI22_X1 U6868 ( .A1(n5551), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5550), .B2(
        n8819), .ZN(n5379) );
  OR2_X1 U6869 ( .A1(n5381), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5382) );
  AND2_X1 U6870 ( .A1(n5382), .A2(n5397), .ZN(n7055) );
  NAND2_X1 U6871 ( .A1(n6352), .A2(n7055), .ZN(n5386) );
  NAND2_X1 U6872 ( .A1(n5201), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6873 ( .A1(n5248), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6874 ( .A1(n7423), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5383) );
  NAND4_X1 U6875 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n8731)
         );
  AND2_X1 U6876 ( .A1(n8731), .A2(n6337), .ZN(n5387) );
  AOI21_X1 U6877 ( .B1(n7283), .B2(n5711), .A(n5387), .ZN(n8602) );
  NAND2_X1 U6878 ( .A1(n7283), .A2(n6342), .ZN(n5389) );
  NAND2_X1 U6879 ( .A1(n8731), .A2(n5711), .ZN(n5388) );
  NAND2_X1 U6880 ( .A1(n5389), .A2(n5388), .ZN(n5390) );
  XNOR2_X1 U6881 ( .A(n5390), .B(n5662), .ZN(n8600) );
  XNOR2_X1 U6882 ( .A(n5392), .B(n5391), .ZN(n6428) );
  NAND2_X1 U6883 ( .A1(n6428), .A2(n7420), .ZN(n5396) );
  OR2_X1 U6884 ( .A1(n5393), .A2(n4688), .ZN(n5394) );
  XNOR2_X1 U6885 ( .A(n5394), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9301) );
  AOI22_X1 U6886 ( .A1(n5551), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5550), .B2(
        n9301), .ZN(n5395) );
  NAND2_X1 U6887 ( .A1(n9264), .A2(n6342), .ZN(n5404) );
  NAND2_X1 U6888 ( .A1(n6416), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6889 ( .A1(n5397), .A2(n10006), .ZN(n5398) );
  NAND2_X1 U6890 ( .A1(n5422), .A2(n5398), .ZN(n9266) );
  INV_X1 U6891 ( .A(n9266), .ZN(n7083) );
  NAND2_X1 U6892 ( .A1(n6352), .A2(n7083), .ZN(n5401) );
  NAND2_X1 U6893 ( .A1(n7423), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6894 ( .A1(n5248), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5399) );
  NAND4_X1 U6895 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n8730)
         );
  NAND2_X1 U6896 ( .A1(n8730), .A2(n5711), .ZN(n5403) );
  NAND2_X1 U6897 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  XNOR2_X1 U6898 ( .A(n5405), .B(n4419), .ZN(n5408) );
  NAND2_X1 U6899 ( .A1(n9264), .A2(n5711), .ZN(n5407) );
  NAND2_X1 U6900 ( .A1(n8730), .A2(n6337), .ZN(n5406) );
  NAND2_X1 U6901 ( .A1(n5407), .A2(n5406), .ZN(n5409) );
  NAND2_X1 U6902 ( .A1(n5408), .A2(n5409), .ZN(n8604) );
  OAI21_X1 U6903 ( .B1(n8602), .B2(n8600), .A(n8604), .ZN(n5414) );
  NAND3_X1 U6904 ( .A1(n8604), .A2(n8602), .A3(n8600), .ZN(n5412) );
  INV_X1 U6905 ( .A(n5408), .ZN(n5411) );
  INV_X1 U6906 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6907 ( .A1(n5411), .A2(n5410), .ZN(n8605) );
  AND2_X1 U6908 ( .A1(n5412), .A2(n8605), .ZN(n5413) );
  XNOR2_X1 U6909 ( .A(n5416), .B(n5415), .ZN(n6534) );
  NAND2_X1 U6910 ( .A1(n6534), .A2(n7420), .ZN(n5420) );
  NAND2_X1 U6911 ( .A1(n5417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U6912 ( .A(n5418), .B(P1_IR_REG_12__SCAN_IN), .ZN(n8821) );
  AOI22_X1 U6913 ( .A1(n5551), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5550), .B2(
        n8821), .ZN(n5419) );
  NAND2_X1 U6914 ( .A1(n7221), .A2(n6342), .ZN(n5429) );
  NAND2_X1 U6915 ( .A1(n6416), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5427) );
  AND2_X1 U6916 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  NOR2_X1 U6917 ( .A1(n5444), .A2(n5423), .ZN(n8612) );
  NAND2_X1 U6918 ( .A1(n6352), .A2(n8612), .ZN(n5426) );
  NAND2_X1 U6919 ( .A1(n7423), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6920 ( .A1(n5248), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5424) );
  NAND4_X1 U6921 ( .A1(n5427), .A2(n5426), .A3(n5425), .A4(n5424), .ZN(n8729)
         );
  NAND2_X1 U6922 ( .A1(n8729), .A2(n5711), .ZN(n5428) );
  NAND2_X1 U6923 ( .A1(n5429), .A2(n5428), .ZN(n5430) );
  XNOR2_X1 U6924 ( .A(n5430), .B(n5662), .ZN(n5432) );
  AND2_X1 U6925 ( .A1(n8729), .A2(n6337), .ZN(n5431) );
  AOI21_X1 U6926 ( .B1(n7221), .B2(n5711), .A(n5431), .ZN(n5433) );
  NAND2_X1 U6927 ( .A1(n5432), .A2(n5433), .ZN(n7291) );
  INV_X1 U6928 ( .A(n5432), .ZN(n5435) );
  INV_X1 U6929 ( .A(n5433), .ZN(n5434) );
  NAND2_X1 U6930 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  AND2_X1 U6931 ( .A1(n7291), .A2(n5436), .ZN(n8606) );
  XNOR2_X1 U6932 ( .A(n5438), .B(n5437), .ZN(n6536) );
  NAND2_X1 U6933 ( .A1(n6536), .A2(n7420), .ZN(n5443) );
  INV_X1 U6934 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6935 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X1 U6936 ( .A(n5441), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8822) );
  AOI22_X1 U6937 ( .A1(n5551), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5550), .B2(
        n8822), .ZN(n5442) );
  NAND2_X1 U6938 ( .A1(n9199), .A2(n6342), .ZN(n5451) );
  NAND2_X1 U6939 ( .A1(n6416), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5449) );
  OR2_X1 U6940 ( .A1(n5444), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5445) );
  AND2_X1 U6941 ( .A1(n5469), .A2(n5445), .ZN(n7297) );
  NAND2_X1 U6942 ( .A1(n6352), .A2(n7297), .ZN(n5448) );
  NAND2_X1 U6943 ( .A1(n5248), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6944 ( .A1(n7423), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5446) );
  NAND4_X1 U6945 ( .A1(n5449), .A2(n5448), .A3(n5447), .A4(n5446), .ZN(n8728)
         );
  NAND2_X1 U6946 ( .A1(n8728), .A2(n6336), .ZN(n5450) );
  NAND2_X1 U6947 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  XNOR2_X1 U6948 ( .A(n5452), .B(n5662), .ZN(n5454) );
  AND2_X1 U6949 ( .A1(n8728), .A2(n6337), .ZN(n5453) );
  AOI21_X1 U6950 ( .B1(n9199), .B2(n6336), .A(n5453), .ZN(n5455) );
  NAND2_X1 U6951 ( .A1(n5454), .A2(n5455), .ZN(n5459) );
  INV_X1 U6952 ( .A(n5454), .ZN(n5457) );
  INV_X1 U6953 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U6954 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U6955 ( .A1(n5459), .A2(n5458), .ZN(n7290) );
  XNOR2_X1 U6956 ( .A(n5461), .B(n5460), .ZN(n6539) );
  NAND2_X1 U6957 ( .A1(n6539), .A2(n7420), .ZN(n5468) );
  OR2_X1 U6958 ( .A1(n5462), .A2(n4688), .ZN(n5464) );
  MUX2_X1 U6959 ( .A(n5464), .B(P1_IR_REG_31__SCAN_IN), .S(n5463), .Z(n5466)
         );
  AND2_X1 U6960 ( .A1(n5466), .A2(n5465), .ZN(n9346) );
  AOI22_X1 U6961 ( .A1(n5551), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5550), .B2(
        n9346), .ZN(n5467) );
  INV_X1 U6962 ( .A(n6342), .ZN(n5729) );
  AOI22_X1 U6963 ( .A1(n6416), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7423), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6964 ( .A1(n5469), .A2(n8565), .ZN(n5470) );
  AND2_X1 U6965 ( .A1(n5483), .A2(n5470), .ZN(n9405) );
  AOI22_X1 U6966 ( .A1(n6352), .A2(n9405), .B1(n5248), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n5471) );
  OAI22_X1 U6967 ( .A1(n9545), .A2(n5729), .B1(n7309), .B2(n5732), .ZN(n5473)
         );
  XNOR2_X1 U6968 ( .A(n5473), .B(n4419), .ZN(n5474) );
  INV_X1 U6969 ( .A(n9545), .ZN(n9406) );
  AOI22_X1 U6970 ( .A1(n9406), .A2(n5711), .B1(n6337), .B2(n8727), .ZN(n8563)
         );
  XNOR2_X1 U6971 ( .A(n5476), .B(n5475), .ZN(n5477) );
  XNOR2_X1 U6972 ( .A(n5478), .B(n5477), .ZN(n6573) );
  NAND2_X1 U6973 ( .A1(n6573), .A2(n7420), .ZN(n5481) );
  NAND2_X1 U6974 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5479) );
  XNOR2_X1 U6975 ( .A(n5479), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8824) );
  AOI22_X1 U6976 ( .A1(n5551), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5550), .B2(
        n8824), .ZN(n5480) );
  AOI22_X1 U6977 ( .A1(n6416), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n5248), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n5486) );
  AND2_X1 U6978 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  NOR2_X1 U6979 ( .A1(n5502), .A2(n5484), .ZN(n8714) );
  AOI22_X1 U6980 ( .A1(n6352), .A2(n8714), .B1(n7423), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n5485) );
  OAI22_X1 U6981 ( .A1(n9276), .A2(n5729), .B1(n8872), .B2(n5732), .ZN(n5487)
         );
  XNOR2_X1 U6982 ( .A(n5487), .B(n4419), .ZN(n5488) );
  NOR2_X1 U6983 ( .A1(n5489), .A2(n5488), .ZN(n5491) );
  INV_X1 U6984 ( .A(n9276), .ZN(n7337) );
  AOI22_X1 U6985 ( .A1(n7337), .A2(n6336), .B1(n6337), .B2(n8874), .ZN(n8707)
         );
  NAND2_X1 U6986 ( .A1(n8708), .A2(n8707), .ZN(n8706) );
  INV_X1 U6987 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U6988 ( .A1(n8706), .A2(n5492), .ZN(n8624) );
  XNOR2_X1 U6989 ( .A(n5494), .B(n5493), .ZN(n5495) );
  XNOR2_X1 U6990 ( .A(n5496), .B(n5495), .ZN(n6681) );
  NAND2_X1 U6991 ( .A1(n6681), .A2(n7420), .ZN(n5501) );
  INV_X1 U6992 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6993 ( .A1(n5498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5499) );
  XNOR2_X1 U6994 ( .A(n5499), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8826) );
  AOI22_X1 U6995 ( .A1(n5551), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5550), .B2(
        n8826), .ZN(n5500) );
  INV_X1 U6996 ( .A(n9192), .ZN(n9105) );
  NAND2_X1 U6997 ( .A1(n6416), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5508) );
  NOR2_X1 U6998 ( .A1(n5502), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6999 ( .A1(n6352), .A2(n5023), .ZN(n5507) );
  NAND2_X1 U7000 ( .A1(n7423), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7001 ( .A1(n5248), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5505) );
  NAND4_X1 U7002 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n8875)
         );
  INV_X1 U7003 ( .A(n8875), .ZN(n7335) );
  OAI22_X1 U7004 ( .A1(n9105), .A2(n5732), .B1(n7335), .B2(n5731), .ZN(n5515)
         );
  NAND2_X1 U7005 ( .A1(n9192), .A2(n6342), .ZN(n5510) );
  NAND2_X1 U7006 ( .A1(n8875), .A2(n6336), .ZN(n5509) );
  NAND2_X1 U7007 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  XNOR2_X1 U7008 ( .A(n5511), .B(n4419), .ZN(n5514) );
  XOR2_X1 U7009 ( .A(n5515), .B(n5514), .Z(n8625) );
  XOR2_X1 U7010 ( .A(n5513), .B(n5512), .Z(n8635) );
  INV_X1 U7011 ( .A(n5514), .ZN(n5517) );
  INV_X1 U7012 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U7013 ( .A1(n5517), .A2(n5516), .ZN(n8632) );
  MUX2_X1 U7014 ( .A(n6951), .B(n10098), .S(n5523), .Z(n5541) );
  XNOR2_X1 U7015 ( .A(n5541), .B(SI_18_), .ZN(n5540) );
  XNOR2_X1 U7016 ( .A(n5539), .B(n5540), .ZN(n6950) );
  NAND2_X1 U7017 ( .A1(n6950), .A2(n7420), .ZN(n5526) );
  XNOR2_X1 U7018 ( .A(n5524), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8843) );
  AOI22_X1 U7019 ( .A1(n5551), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5550), .B2(
        n8843), .ZN(n5525) );
  NAND2_X1 U7020 ( .A1(n9187), .A2(n6342), .ZN(n5534) );
  NAND2_X1 U7021 ( .A1(n6416), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7022 ( .A1(n5527), .A2(n8687), .ZN(n5528) );
  AND2_X1 U7023 ( .A1(n5554), .A2(n5528), .ZN(n9080) );
  NAND2_X1 U7024 ( .A1(n6352), .A2(n9080), .ZN(n5531) );
  NAND2_X1 U7025 ( .A1(n7423), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7026 ( .A1(n5248), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5529) );
  NAND4_X1 U7027 ( .A1(n5532), .A2(n5531), .A3(n5530), .A4(n5529), .ZN(n8882)
         );
  NAND2_X1 U7028 ( .A1(n8882), .A2(n5711), .ZN(n5533) );
  NAND2_X1 U7029 ( .A1(n5534), .A2(n5533), .ZN(n5535) );
  XNOR2_X1 U7030 ( .A(n5535), .B(n5662), .ZN(n5538) );
  AND2_X1 U7031 ( .A1(n8882), .A2(n6337), .ZN(n5536) );
  AOI21_X1 U7032 ( .B1(n9187), .B2(n5711), .A(n5536), .ZN(n5537) );
  NAND2_X1 U7033 ( .A1(n5538), .A2(n5537), .ZN(n8680) );
  NOR2_X1 U7034 ( .A1(n5538), .A2(n5537), .ZN(n8682) );
  INV_X1 U7035 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7036 ( .A1(n5542), .A2(SI_18_), .ZN(n5543) );
  MUX2_X1 U7037 ( .A(n10081), .B(n7032), .S(n5523), .Z(n5546) );
  INV_X1 U7038 ( .A(SI_19_), .ZN(n5545) );
  NAND2_X1 U7039 ( .A1(n5546), .A2(n5545), .ZN(n5568) );
  INV_X1 U7040 ( .A(n5546), .ZN(n5547) );
  NAND2_X1 U7041 ( .A1(n5547), .A2(SI_19_), .ZN(n5548) );
  NAND2_X1 U7042 ( .A1(n5568), .A2(n5548), .ZN(n5569) );
  NAND2_X1 U7043 ( .A1(n7030), .A2(n7420), .ZN(n5553) );
  AOI22_X1 U7044 ( .A1(n5551), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7508), .B2(
        n5550), .ZN(n5552) );
  NAND2_X2 U7045 ( .A1(n5553), .A2(n5552), .ZN(n9182) );
  NAND2_X1 U7046 ( .A1(n9182), .A2(n6342), .ZN(n5561) );
  NAND2_X1 U7047 ( .A1(n6416), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7048 ( .A1(n5554), .A2(n8584), .ZN(n5555) );
  NAND2_X1 U7049 ( .A1(n5574), .A2(n5555), .ZN(n8583) );
  INV_X1 U7050 ( .A(n8583), .ZN(n9067) );
  NAND2_X1 U7051 ( .A1(n6352), .A2(n9067), .ZN(n5558) );
  NAND2_X1 U7052 ( .A1(n5248), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7053 ( .A1(n7423), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5556) );
  NAND4_X1 U7054 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n8885)
         );
  NAND2_X1 U7055 ( .A1(n8885), .A2(n6336), .ZN(n5560) );
  NAND2_X1 U7056 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  XNOR2_X1 U7057 ( .A(n5562), .B(n5662), .ZN(n5567) );
  INV_X1 U7058 ( .A(n5567), .ZN(n5565) );
  AND2_X1 U7059 ( .A1(n8885), .A2(n6337), .ZN(n5563) );
  AOI21_X1 U7060 ( .B1(n9182), .B2(n6336), .A(n5563), .ZN(n5566) );
  INV_X1 U7061 ( .A(n5566), .ZN(n5564) );
  NAND2_X1 U7062 ( .A1(n5565), .A2(n5564), .ZN(n8580) );
  MUX2_X1 U7063 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5523), .Z(n5585) );
  XNOR2_X1 U7064 ( .A(n5585), .B(n5586), .ZN(n5571) );
  XNOR2_X1 U7065 ( .A(n5587), .B(n5571), .ZN(n7088) );
  NAND2_X1 U7066 ( .A1(n7088), .A2(n7420), .ZN(n5573) );
  INV_X1 U7067 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7089) );
  OR2_X1 U7068 ( .A1(n5259), .A2(n7089), .ZN(n5572) );
  NAND2_X1 U7069 ( .A1(n9177), .A2(n6342), .ZN(n5579) );
  AND2_X1 U7070 ( .A1(n5574), .A2(n8668), .ZN(n5575) );
  OR2_X1 U7071 ( .A1(n5575), .A2(n5591), .ZN(n9053) );
  AOI22_X1 U7072 ( .A1(n6416), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n7423), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7073 ( .A1(n5248), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U7074 ( .C1(n9053), .C2(n5595), .A(n5577), .B(n5576), .ZN(n8725)
         );
  NAND2_X1 U7075 ( .A1(n8725), .A2(n5711), .ZN(n5578) );
  NAND2_X1 U7076 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  XNOR2_X1 U7077 ( .A(n5580), .B(n5662), .ZN(n5583) );
  AND2_X1 U7078 ( .A1(n8725), .A2(n6337), .ZN(n5581) );
  AOI21_X1 U7079 ( .B1(n9177), .B2(n5711), .A(n5581), .ZN(n5582) );
  NAND2_X1 U7080 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  OAI21_X1 U7081 ( .B1(n5583), .B2(n5582), .A(n5584), .ZN(n8666) );
  MUX2_X1 U7082 ( .A(n7170), .B(n7157), .S(n5523), .Z(n5603) );
  XNOR2_X1 U7083 ( .A(n5603), .B(SI_21_), .ZN(n5588) );
  XNOR2_X1 U7084 ( .A(n5605), .B(n5588), .ZN(n7156) );
  NAND2_X1 U7085 ( .A1(n7156), .A2(n7420), .ZN(n5590) );
  OR2_X1 U7086 ( .A1(n5259), .A2(n7157), .ZN(n5589) );
  NAND2_X1 U7087 ( .A1(n9172), .A2(n6342), .ZN(n5597) );
  OR2_X1 U7088 ( .A1(n5591), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7089 ( .A1(n5591), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7090 ( .A1(n5592), .A2(n5612), .ZN(n8593) );
  AOI22_X1 U7091 ( .A1(n6416), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5248), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7092 ( .A1(n7423), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7093 ( .C1(n8593), .C2(n5595), .A(n5594), .B(n5593), .ZN(n8724)
         );
  NAND2_X1 U7094 ( .A1(n8724), .A2(n5711), .ZN(n5596) );
  NAND2_X1 U7095 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  XNOR2_X1 U7096 ( .A(n5598), .B(n4419), .ZN(n5601) );
  AOI22_X1 U7097 ( .A1(n9172), .A2(n6336), .B1(n6337), .B2(n8724), .ZN(n5599)
         );
  XNOR2_X1 U7098 ( .A(n5601), .B(n5599), .ZN(n8591) );
  INV_X1 U7099 ( .A(n5599), .ZN(n5600) );
  MUX2_X1 U7100 ( .A(n7273), .B(n7565), .S(n5523), .Z(n5607) );
  NAND2_X1 U7101 ( .A1(n5607), .A2(n5606), .ZN(n5619) );
  INV_X1 U7102 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7103 ( .A1(n5608), .A2(SI_22_), .ZN(n5609) );
  NAND2_X1 U7104 ( .A1(n5619), .A2(n5609), .ZN(n5620) );
  XNOR2_X1 U7105 ( .A(n5621), .B(n5620), .ZN(n7272) );
  NAND2_X1 U7106 ( .A1(n7272), .A2(n7420), .ZN(n5611) );
  OR2_X1 U7107 ( .A1(n5259), .A2(n7565), .ZN(n5610) );
  AOI22_X1 U7108 ( .A1(n6416), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n7423), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5614) );
  INV_X1 U7109 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10182) );
  AOI21_X1 U7110 ( .B1(n10182), .B2(n5612), .A(n5629), .ZN(n9027) );
  AOI22_X1 U7111 ( .A1(n6352), .A2(n9027), .B1(n5248), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5613) );
  OAI22_X1 U7112 ( .A1(n9030), .A2(n5729), .B1(n8892), .B2(n5732), .ZN(n5615)
         );
  XOR2_X1 U7113 ( .A(n4419), .B(n5615), .Z(n5616) );
  OAI22_X1 U7114 ( .A1(n9030), .A2(n5732), .B1(n8892), .B2(n5731), .ZN(n8675)
         );
  INV_X1 U7115 ( .A(n5618), .ZN(n8572) );
  INV_X1 U7116 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5622) );
  MUX2_X1 U7117 ( .A(n5622), .B(n7288), .S(n5523), .Z(n5624) );
  INV_X1 U7118 ( .A(SI_23_), .ZN(n5623) );
  NAND2_X1 U7119 ( .A1(n5624), .A2(n5623), .ZN(n5646) );
  INV_X1 U7120 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7121 ( .A1(n5625), .A2(SI_23_), .ZN(n5626) );
  NAND2_X1 U7122 ( .A1(n7286), .A2(n7420), .ZN(n5628) );
  OR2_X1 U7123 ( .A1(n5259), .A2(n7288), .ZN(n5627) );
  NAND2_X1 U7124 ( .A1(n9161), .A2(n6342), .ZN(n5636) );
  NAND2_X1 U7125 ( .A1(n6416), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5634) );
  INV_X1 U7126 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8576) );
  INV_X1 U7127 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7128 ( .A1(n5629), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5655) );
  AOI21_X1 U7129 ( .B1(n8576), .B2(n5630), .A(n5654), .ZN(n9005) );
  NAND2_X1 U7130 ( .A1(n6352), .A2(n9005), .ZN(n5633) );
  NAND2_X1 U7131 ( .A1(n7423), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7132 ( .A1(n5248), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5631) );
  NAND4_X1 U7133 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n8895)
         );
  NAND2_X1 U7134 ( .A1(n8895), .A2(n6336), .ZN(n5635) );
  NAND2_X1 U7135 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  XNOR2_X1 U7136 ( .A(n5637), .B(n5662), .ZN(n5639) );
  AND2_X1 U7137 ( .A1(n8895), .A2(n6337), .ZN(n5638) );
  AOI21_X1 U7138 ( .B1(n9161), .B2(n5711), .A(n5638), .ZN(n5640) );
  NAND2_X1 U7139 ( .A1(n5639), .A2(n5640), .ZN(n8642) );
  INV_X1 U7140 ( .A(n5639), .ZN(n5642) );
  INV_X1 U7141 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7142 ( .A1(n5642), .A2(n5641), .ZN(n5643) );
  AND2_X1 U7143 ( .A1(n8642), .A2(n5643), .ZN(n8571) );
  NAND2_X1 U7144 ( .A1(n8570), .A2(n8642), .ZN(n5670) );
  NAND2_X1 U7145 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  NAND2_X1 U7146 ( .A1(n5647), .A2(n5646), .ZN(n5673) );
  INV_X1 U7147 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7570) );
  INV_X1 U7148 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7318) );
  MUX2_X1 U7149 ( .A(n7570), .B(n7318), .S(n5523), .Z(n5649) );
  INV_X1 U7150 ( .A(SI_24_), .ZN(n5648) );
  NAND2_X1 U7151 ( .A1(n5649), .A2(n5648), .ZN(n5674) );
  INV_X1 U7152 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7153 ( .A1(n5650), .A2(SI_24_), .ZN(n5651) );
  XNOR2_X1 U7154 ( .A(n5673), .B(n5672), .ZN(n7317) );
  NAND2_X1 U7155 ( .A1(n7317), .A2(n7420), .ZN(n5653) );
  OR2_X1 U7156 ( .A1(n5259), .A2(n7318), .ZN(n5652) );
  NAND2_X1 U7157 ( .A1(n9157), .A2(n6342), .ZN(n5661) );
  NAND2_X1 U7158 ( .A1(n6416), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5659) );
  INV_X1 U7159 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U7160 ( .A1(n5654), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5683) );
  INV_X1 U7161 ( .A(n5683), .ZN(n5682) );
  AOI21_X1 U7162 ( .B1(n8651), .B2(n5655), .A(n5682), .ZN(n8997) );
  NAND2_X1 U7163 ( .A1(n6352), .A2(n8997), .ZN(n5658) );
  NAND2_X1 U7164 ( .A1(n7423), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7165 ( .A1(n5248), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5656) );
  NAND4_X1 U7166 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n8722)
         );
  NAND2_X1 U7167 ( .A1(n8722), .A2(n5711), .ZN(n5660) );
  NAND2_X1 U7168 ( .A1(n5661), .A2(n5660), .ZN(n5663) );
  XNOR2_X1 U7169 ( .A(n5663), .B(n5662), .ZN(n5665) );
  AND2_X1 U7170 ( .A1(n8722), .A2(n6337), .ZN(n5664) );
  AOI21_X1 U7171 ( .B1(n9157), .B2(n6336), .A(n5664), .ZN(n5666) );
  NAND2_X1 U7172 ( .A1(n5665), .A2(n5666), .ZN(n5671) );
  INV_X1 U7173 ( .A(n5665), .ZN(n5668) );
  INV_X1 U7174 ( .A(n5666), .ZN(n5667) );
  NAND2_X1 U7175 ( .A1(n5668), .A2(n5667), .ZN(n5669) );
  AND2_X1 U7176 ( .A1(n5671), .A2(n5669), .ZN(n8643) );
  NAND2_X1 U7177 ( .A1(n5670), .A2(n8643), .ZN(n8646) );
  NAND2_X1 U7178 ( .A1(n8646), .A2(n5671), .ZN(n8615) );
  NAND2_X1 U7179 ( .A1(n5673), .A2(n5672), .ZN(n5675) );
  INV_X1 U7180 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9234) );
  MUX2_X1 U7181 ( .A(n8558), .B(n9234), .S(n5523), .Z(n5677) );
  INV_X1 U7182 ( .A(SI_25_), .ZN(n5676) );
  NAND2_X1 U7183 ( .A1(n5677), .A2(n5676), .ZN(n5693) );
  INV_X1 U7184 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7185 ( .A1(n5678), .A2(SI_25_), .ZN(n5679) );
  XNOR2_X1 U7186 ( .A(n5692), .B(n5691), .ZN(n8556) );
  NAND2_X1 U7187 ( .A1(n8556), .A2(n7420), .ZN(n5681) );
  OR2_X1 U7188 ( .A1(n5259), .A2(n9234), .ZN(n5680) );
  NAND2_X1 U7189 ( .A1(n6416), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5687) );
  INV_X1 U7190 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U7191 ( .A1(n5682), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5702) );
  INV_X1 U7192 ( .A(n5702), .ZN(n5701) );
  AOI21_X1 U7193 ( .B1(n8620), .B2(n5683), .A(n5701), .ZN(n8983) );
  NAND2_X1 U7194 ( .A1(n6352), .A2(n8983), .ZN(n5686) );
  NAND2_X1 U7195 ( .A1(n7423), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7196 ( .A1(n5248), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U7197 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n8897)
         );
  INV_X1 U7198 ( .A(n8897), .ZN(n8898) );
  OAI22_X1 U7199 ( .A1(n8986), .A2(n5732), .B1(n8898), .B2(n5731), .ZN(n5713)
         );
  NAND2_X1 U7200 ( .A1(n9152), .A2(n6342), .ZN(n5689) );
  NAND2_X1 U7201 ( .A1(n8897), .A2(n6336), .ZN(n5688) );
  NAND2_X1 U7202 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  XNOR2_X1 U7203 ( .A(n5690), .B(n4419), .ZN(n5712) );
  XOR2_X1 U7204 ( .A(n5713), .B(n5712), .Z(n8616) );
  NAND2_X1 U7205 ( .A1(n8615), .A2(n8616), .ZN(n8693) );
  NAND2_X1 U7206 ( .A1(n5692), .A2(n5691), .ZN(n5694) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8555) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U7209 ( .A(n8555), .B(n9231), .S(n5047), .Z(n5696) );
  INV_X1 U7210 ( .A(SI_26_), .ZN(n5695) );
  NAND2_X1 U7211 ( .A1(n5696), .A2(n5695), .ZN(n5718) );
  INV_X1 U7212 ( .A(n5696), .ZN(n5697) );
  NAND2_X1 U7213 ( .A1(n5697), .A2(SI_26_), .ZN(n5698) );
  NAND2_X1 U7214 ( .A1(n8554), .A2(n7420), .ZN(n5700) );
  OR2_X1 U7215 ( .A1(n5259), .A2(n9231), .ZN(n5699) );
  NAND2_X1 U7216 ( .A1(n9146), .A2(n6342), .ZN(n5708) );
  NAND2_X1 U7217 ( .A1(n6416), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5706) );
  INV_X1 U7218 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U7219 ( .A1(n5701), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5726) );
  INV_X1 U7220 ( .A(n5726), .ZN(n5773) );
  AOI21_X1 U7221 ( .B1(n8702), .B2(n5702), .A(n5773), .ZN(n8964) );
  NAND2_X1 U7222 ( .A1(n6352), .A2(n8964), .ZN(n5705) );
  NAND2_X1 U7223 ( .A1(n7423), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7224 ( .A1(n5248), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5703) );
  NAND4_X1 U7225 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n8721)
         );
  NAND2_X1 U7226 ( .A1(n8721), .A2(n5167), .ZN(n5707) );
  NAND2_X1 U7227 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  XNOR2_X1 U7228 ( .A(n5709), .B(n4419), .ZN(n5737) );
  AND2_X1 U7229 ( .A1(n8721), .A2(n6337), .ZN(n5710) );
  AOI21_X1 U7230 ( .B1(n9146), .B2(n5167), .A(n5710), .ZN(n5735) );
  XNOR2_X1 U7231 ( .A(n5737), .B(n5735), .ZN(n8695) );
  INV_X1 U7232 ( .A(n5712), .ZN(n5715) );
  INV_X1 U7233 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7234 ( .A1(n5715), .A2(n5714), .ZN(n8692) );
  NAND2_X1 U7235 ( .A1(n5717), .A2(n5716), .ZN(n5719) );
  INV_X1 U7236 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5720) );
  MUX2_X1 U7237 ( .A(n5720), .B(n9229), .S(n5047), .Z(n5721) );
  INV_X1 U7238 ( .A(SI_27_), .ZN(n10003) );
  NAND2_X1 U7239 ( .A1(n5721), .A2(n10003), .ZN(n6293) );
  INV_X1 U7240 ( .A(n5721), .ZN(n5722) );
  NAND2_X1 U7241 ( .A1(n5722), .A2(SI_27_), .ZN(n5723) );
  NAND2_X1 U7242 ( .A1(n8550), .A2(n7420), .ZN(n5725) );
  OR2_X1 U7243 ( .A1(n5259), .A2(n9229), .ZN(n5724) );
  AOI22_X1 U7244 ( .A1(n6416), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n7423), .B2(
        P1_REG0_REG_27__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U7245 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n5726), .ZN(n8950) );
  AOI22_X1 U7246 ( .A1(n6352), .A2(n8950), .B1(n5248), .B2(
        P1_REG1_REG_27__SCAN_IN), .ZN(n5727) );
  OAI22_X1 U7247 ( .A1(n8952), .A2(n5729), .B1(n8698), .B2(n5732), .ZN(n5730)
         );
  XNOR2_X1 U7248 ( .A(n5730), .B(n4419), .ZN(n5734) );
  OAI22_X1 U7249 ( .A1(n8952), .A2(n5732), .B1(n8698), .B2(n5731), .ZN(n5733)
         );
  NOR2_X1 U7250 ( .A1(n5734), .A2(n5733), .ZN(n6349) );
  AOI21_X1 U7251 ( .B1(n5734), .B2(n5733), .A(n6349), .ZN(n5739) );
  INV_X1 U7252 ( .A(n5735), .ZN(n5736) );
  NAND2_X1 U7253 ( .A1(n5737), .A2(n5736), .ZN(n5740) );
  NAND2_X1 U7254 ( .A1(n8694), .A2(n5738), .ZN(n6348) );
  AOI21_X1 U7255 ( .B1(n8694), .B2(n5740), .A(n5739), .ZN(n5764) );
  NAND2_X1 U7256 ( .A1(n9235), .A2(P1_B_REG_SCAN_IN), .ZN(n5741) );
  MUX2_X1 U7257 ( .A(n5741), .B(P1_B_REG_SCAN_IN), .S(n5744), .Z(n5743) );
  INV_X1 U7258 ( .A(n5742), .ZN(n9232) );
  AND2_X1 U7259 ( .A1(n9232), .A2(n4420), .ZN(n6398) );
  AND2_X1 U7260 ( .A1(n9232), .A2(n9235), .ZN(n6402) );
  NOR2_X1 U7261 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n5749) );
  NOR4_X1 U7262 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n5748) );
  NOR4_X1 U7263 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5747) );
  NOR4_X1 U7264 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5746) );
  NAND4_X1 U7265 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n5755)
         );
  NOR4_X1 U7266 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5753) );
  NOR4_X1 U7267 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5752) );
  NOR4_X1 U7268 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5751) );
  NOR4_X1 U7269 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5750) );
  NAND4_X1 U7270 ( .A1(n5753), .A2(n5752), .A3(n5751), .A4(n5750), .ZN(n5754)
         );
  OAI21_X1 U7271 ( .B1(n5755), .B2(n5754), .A(n6396), .ZN(n6716) );
  NAND3_X1 U7272 ( .A1(n9125), .A2(n9120), .A3(n6716), .ZN(n5769) );
  NOR2_X1 U7273 ( .A1(n5769), .A2(n7559), .ZN(n5765) );
  INV_X1 U7274 ( .A(n6723), .ZN(n9445) );
  INV_X1 U7275 ( .A(n7460), .ZN(n5762) );
  AND2_X1 U7276 ( .A1(n9544), .A2(n5762), .ZN(n5763) );
  INV_X1 U7277 ( .A(n5765), .ZN(n5783) );
  NOR2_X1 U7278 ( .A1(n6723), .A2(n5160), .ZN(n6734) );
  INV_X1 U7279 ( .A(n6734), .ZN(n5766) );
  OR2_X1 U7280 ( .A1(n5783), .A2(n5766), .ZN(n5767) );
  AND2_X1 U7281 ( .A1(n7508), .A2(n5160), .ZN(n9449) );
  NAND2_X1 U7282 ( .A1(n9445), .A2(n9449), .ZN(n9121) );
  NAND2_X1 U7283 ( .A1(n9141), .A2(n5768), .ZN(n5787) );
  OAI21_X1 U7284 ( .B1(n6734), .B2(n9544), .A(n5769), .ZN(n5771) );
  NAND2_X1 U7285 ( .A1(n7460), .A2(n6721), .ZN(n5770) );
  NAND2_X1 U7286 ( .A1(n5771), .A2(n6718), .ZN(n5772) );
  NAND2_X1 U7287 ( .A1(n6416), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5779) );
  NAND3_X1 U7288 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .A3(n5773), .ZN(n6351) );
  INV_X1 U7289 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U7290 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5773), .ZN(n5774) );
  NAND2_X1 U7291 ( .A1(n9964), .A2(n5774), .ZN(n5775) );
  NAND2_X1 U7292 ( .A1(n6352), .A2(n8935), .ZN(n5778) );
  NAND2_X1 U7293 ( .A1(n7423), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7294 ( .A1(n5248), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5776) );
  NAND4_X1 U7295 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n8720)
         );
  AND2_X2 U7296 ( .A1(n7460), .A2(n5780), .ZN(n8859) );
  NAND2_X1 U7297 ( .A1(n8720), .A2(n8859), .ZN(n5782) );
  INV_X1 U7298 ( .A(n5780), .ZN(n8750) );
  NAND2_X1 U7299 ( .A1(n8721), .A2(n8699), .ZN(n5781) );
  AND2_X1 U7300 ( .A1(n5782), .A2(n5781), .ZN(n8956) );
  INV_X1 U7301 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5784) );
  OAI22_X1 U7302 ( .A1(n8956), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5784), .ZN(n5785) );
  AOI21_X1 U7303 ( .B1(n8713), .B2(n8950), .A(n5785), .ZN(n5786) );
  AND2_X1 U7304 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  NAND2_X1 U7305 ( .A1(n5789), .A2(n5788), .ZN(P1_U3214) );
  INV_X1 U7306 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6238) );
  NOR2_X1 U7307 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5796) );
  NAND4_X1 U7308 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n5798)
         );
  INV_X2 U7309 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6180) );
  NAND4_X1 U7310 ( .A1(n10054), .A2(n6180), .A3(n5974), .A4(n6042), .ZN(n5797)
         );
  NAND2_X1 U7311 ( .A1(n5804), .A2(n5805), .ZN(n8539) );
  INV_X1 U7312 ( .A(n5809), .ZN(n8543) );
  INV_X1 U7313 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5807) );
  OR2_X2 U7314 ( .A1(n5809), .A2(n8547), .ZN(n5931) );
  INV_X1 U7315 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7316 ( .A1(n5869), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5811) );
  INV_X1 U7317 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6897) );
  INV_X1 U7318 ( .A(n9760), .ZN(n5826) );
  INV_X1 U7319 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7320 ( .A1(n6199), .A2(n5817), .ZN(n6210) );
  MUX2_X1 U7321 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5820), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5823) );
  INV_X1 U7322 ( .A(n5821), .ZN(n5822) );
  INV_X1 U7323 ( .A(n6794), .ZN(n6642) );
  INV_X1 U7324 ( .A(n9774), .ZN(n5834) );
  NAND2_X1 U7325 ( .A1(n6186), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5832) );
  INV_X1 U7326 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5827) );
  OR2_X1 U7327 ( .A1(n5837), .A2(n5827), .ZN(n5831) );
  INV_X1 U7328 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7329 ( .A1(n5931), .A2(n5828), .ZN(n5830) );
  INV_X1 U7330 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6872) );
  OR2_X1 U7331 ( .A1(n5900), .A2(n6872), .ZN(n5829) );
  NAND2_X1 U7332 ( .A1(n4418), .A2(SI_0_), .ZN(n5833) );
  XNOR2_X1 U7333 ( .A(n5833), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U7334 ( .A1(n6900), .A2(n6678), .ZN(n6898) );
  NAND2_X1 U7335 ( .A1(n6239), .A2(n6898), .ZN(n5836) );
  OR2_X1 U7336 ( .A1(n9760), .A2(n5834), .ZN(n5835) );
  NAND2_X1 U7337 ( .A1(n5836), .A2(n5835), .ZN(n9756) );
  NAND2_X1 U7338 ( .A1(n6104), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5844) );
  INV_X1 U7339 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5838) );
  INV_X1 U7340 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6638) );
  OR2_X1 U7341 ( .A1(n5900), .A2(n6638), .ZN(n5842) );
  INV_X1 U7342 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5839) );
  OR2_X1 U7343 ( .A1(n4416), .A2(n5839), .ZN(n5841) );
  OR2_X1 U7344 ( .A1(n5864), .A2(n6375), .ZN(n5849) );
  OR2_X1 U7345 ( .A1(n5865), .A2(n6374), .ZN(n5848) );
  NAND2_X1 U7346 ( .A1(n6083), .A2(n6662), .ZN(n5847) );
  OR2_X1 U7347 ( .A1(n4415), .A2(n9766), .ZN(n7638) );
  NAND2_X1 U7348 ( .A1(n4415), .A2(n9766), .ZN(n7639) );
  NAND2_X1 U7349 ( .A1(n7638), .A2(n7639), .ZN(n6241) );
  NAND2_X1 U7350 ( .A1(n9756), .A2(n6241), .ZN(n5853) );
  INV_X1 U7351 ( .A(n9766), .ZN(n5851) );
  OR2_X1 U7352 ( .A1(n4415), .A2(n5851), .ZN(n5852) );
  NAND2_X1 U7353 ( .A1(n5853), .A2(n5852), .ZN(n6961) );
  NAND2_X1 U7354 ( .A1(n6104), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5859) );
  INV_X1 U7355 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7356 ( .A1(n4413), .A2(n5854), .ZN(n5858) );
  OR2_X1 U7357 ( .A1(n5900), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5857) );
  INV_X1 U7358 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7359 ( .A1(n4416), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U7360 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7361 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5861), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5863) );
  NAND2_X1 U7362 ( .A1(n5863), .A2(n5862), .ZN(n6747) );
  OR2_X1 U7363 ( .A1(n5865), .A2(n6377), .ZN(n5866) );
  NOR2_X1 U7364 ( .A1(n9759), .A2(n6965), .ZN(n5868) );
  INV_X1 U7365 ( .A(n9759), .ZN(n5867) );
  NAND2_X1 U7366 ( .A1(n5869), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5876) );
  INV_X1 U7367 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6751) );
  OR2_X1 U7368 ( .A1(n5931), .A2(n6751), .ZN(n5875) );
  INV_X1 U7369 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7370 ( .A1(n6964), .A2(n5870), .ZN(n5883) );
  NAND2_X1 U7371 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5871) );
  AND2_X1 U7372 ( .A1(n5883), .A2(n5871), .ZN(n7001) );
  OR2_X1 U7373 ( .A1(n5900), .A2(n7001), .ZN(n5874) );
  INV_X1 U7374 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7375 ( .A1(n4416), .A2(n5872), .ZN(n5873) );
  NAND4_X1 U7376 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n8093)
         );
  NAND2_X1 U7377 ( .A1(n5862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7378 ( .A1(n5865), .A2(n6383), .ZN(n5879) );
  OR2_X1 U7379 ( .A1(n5864), .A2(n6384), .ZN(n5878) );
  OAI211_X1 U7380 ( .C1(n7621), .C2(n9591), .A(n5879), .B(n5878), .ZN(n6910)
         );
  AND2_X1 U7381 ( .A1(n8093), .A2(n6910), .ZN(n7005) );
  NAND2_X1 U7382 ( .A1(n6104), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5889) );
  INV_X1 U7383 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5880) );
  OR2_X1 U7384 ( .A1(n4413), .A2(n5880), .ZN(n5888) );
  INV_X1 U7385 ( .A(n5883), .ZN(n5882) );
  INV_X1 U7386 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7387 ( .A1(n5882), .A2(n5881), .ZN(n5901) );
  NAND2_X1 U7388 ( .A1(n5883), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5884) );
  AND2_X1 U7389 ( .A1(n5901), .A2(n5884), .ZN(n7029) );
  OR2_X1 U7390 ( .A1(n5900), .A2(n7029), .ZN(n5887) );
  INV_X1 U7391 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5885) );
  OR2_X1 U7392 ( .A1(n4417), .A2(n5885), .ZN(n5886) );
  OR2_X1 U7393 ( .A1(n5890), .A2(n5814), .ZN(n5892) );
  XNOR2_X1 U7394 ( .A(n5892), .B(n5891), .ZN(n9600) );
  OR2_X1 U7395 ( .A1(n5865), .A2(n6381), .ZN(n5894) );
  OR2_X1 U7396 ( .A1(n5864), .A2(n6380), .ZN(n5893) );
  OAI211_X1 U7397 ( .C1(n7621), .C2(n9600), .A(n5894), .B(n5893), .ZN(n7023)
         );
  OR2_X1 U7398 ( .A1(n8092), .A2(n7023), .ZN(n5896) );
  AND2_X1 U7399 ( .A1(n7007), .A2(n5896), .ZN(n5897) );
  NAND2_X1 U7400 ( .A1(n6104), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5906) );
  INV_X1 U7401 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5899) );
  OR2_X1 U7402 ( .A1(n4416), .A2(n5899), .ZN(n5905) );
  NAND2_X1 U7403 ( .A1(n5901), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5902) );
  AND2_X1 U7404 ( .A1(n5917), .A2(n5902), .ZN(n7101) );
  OR2_X1 U7405 ( .A1(n5900), .A2(n7101), .ZN(n5904) );
  INV_X1 U7406 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6758) );
  OR2_X1 U7407 ( .A1(n4413), .A2(n6758), .ZN(n5903) );
  NAND4_X1 U7408 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n8091)
         );
  OR2_X1 U7409 ( .A1(n5907), .A2(n5814), .ZN(n5909) );
  XNOR2_X1 U7410 ( .A(n5909), .B(n5908), .ZN(n6860) );
  OR2_X1 U7411 ( .A1(n5865), .A2(n6388), .ZN(n5911) );
  OR2_X1 U7412 ( .A1(n5864), .A2(n6387), .ZN(n5910) );
  OAI211_X1 U7413 ( .C1(n7621), .C2(n6860), .A(n5911), .B(n5910), .ZN(n7070)
         );
  AND2_X1 U7414 ( .A1(n8091), .A2(n7070), .ZN(n5912) );
  NAND2_X1 U7415 ( .A1(n6104), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5923) );
  INV_X1 U7416 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7417 ( .A1(n4413), .A2(n5914), .ZN(n5922) );
  INV_X1 U7418 ( .A(n5917), .ZN(n5916) );
  INV_X1 U7419 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7420 ( .A1(n5916), .A2(n5915), .ZN(n5932) );
  NAND2_X1 U7421 ( .A1(n5917), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5918) );
  AND2_X1 U7422 ( .A1(n5932), .A2(n5918), .ZN(n7199) );
  OR2_X1 U7423 ( .A1(n5900), .A2(n7199), .ZN(n5921) );
  INV_X1 U7424 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5919) );
  OR2_X1 U7425 ( .A1(n4417), .A2(n5919), .ZN(n5920) );
  NAND4_X1 U7426 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n8090)
         );
  OR2_X1 U7427 ( .A1(n5865), .A2(n6392), .ZN(n5928) );
  OR2_X1 U7428 ( .A1(n5864), .A2(n6391), .ZN(n5927) );
  NAND2_X1 U7429 ( .A1(n5924), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5925) );
  XNOR2_X1 U7430 ( .A(n5925), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U7431 ( .A1(n6083), .A2(n6975), .ZN(n5926) );
  OR2_X1 U7432 ( .A1(n8090), .A2(n9799), .ZN(n7675) );
  NAND2_X1 U7433 ( .A1(n8090), .A2(n9799), .ZN(n7667) );
  NAND2_X1 U7434 ( .A1(n7675), .A2(n7667), .ZN(n7665) );
  NAND2_X1 U7435 ( .A1(n7093), .A2(n7665), .ZN(n5930) );
  INV_X1 U7436 ( .A(n9799), .ZN(n7200) );
  OR2_X1 U7437 ( .A1(n8090), .A2(n7200), .ZN(n5929) );
  NAND2_X1 U7438 ( .A1(n5869), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5938) );
  INV_X1 U7439 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6973) );
  OR2_X1 U7440 ( .A1(n5931), .A2(n6973), .ZN(n5937) );
  NAND2_X1 U7441 ( .A1(n5932), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5933) );
  AND2_X1 U7442 ( .A1(n5950), .A2(n5933), .ZN(n7929) );
  OR2_X1 U7443 ( .A1(n5900), .A2(n7929), .ZN(n5936) );
  INV_X1 U7444 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5934) );
  OR2_X1 U7445 ( .A1(n4417), .A2(n5934), .ZN(n5935) );
  NAND4_X1 U7446 ( .A1(n5938), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n8089)
         );
  OR2_X1 U7447 ( .A1(n5865), .A2(n6395), .ZN(n5943) );
  OR2_X1 U7448 ( .A1(n5864), .A2(n6394), .ZN(n5942) );
  NAND2_X1 U7449 ( .A1(n5939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7450 ( .A(n5940), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8108) );
  NAND2_X1 U7451 ( .A1(n6083), .A2(n8108), .ZN(n5941) );
  OR2_X1 U7452 ( .A1(n8089), .A2(n9804), .ZN(n7676) );
  NAND2_X1 U7453 ( .A1(n8089), .A2(n9804), .ZN(n7668) );
  INV_X1 U7454 ( .A(n9804), .ZN(n7153) );
  NAND2_X1 U7455 ( .A1(n8089), .A2(n7153), .ZN(n5945) );
  NAND2_X1 U7456 ( .A1(n6186), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5955) );
  INV_X1 U7457 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7458 ( .A1(n4413), .A2(n5946), .ZN(n5954) );
  INV_X1 U7459 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7460 ( .A1(n5931), .A2(n5947), .ZN(n5953) );
  INV_X1 U7461 ( .A(n5950), .ZN(n5949) );
  INV_X1 U7462 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7463 ( .A1(n5949), .A2(n5948), .ZN(n5964) );
  NAND2_X1 U7464 ( .A1(n5950), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5951) );
  AND2_X1 U7465 ( .A1(n5964), .A2(n5951), .ZN(n7258) );
  OR2_X1 U7466 ( .A1(n5900), .A2(n7258), .ZN(n5952) );
  NAND4_X1 U7467 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n8088)
         );
  NAND2_X1 U7468 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  XNOR2_X1 U7469 ( .A(n5957), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9614) );
  OR2_X1 U7470 ( .A1(n5865), .A2(n6401), .ZN(n5959) );
  OR2_X1 U7471 ( .A1(n5864), .A2(n6400), .ZN(n5958) );
  OR2_X1 U7472 ( .A1(n8088), .A2(n8004), .ZN(n5960) );
  NAND2_X1 U7473 ( .A1(n7253), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7474 ( .A1(n8088), .A2(n8004), .ZN(n5961) );
  NAND2_X1 U7475 ( .A1(n6186), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5969) );
  INV_X1 U7476 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8096) );
  OR2_X1 U7477 ( .A1(n4413), .A2(n8096), .ZN(n5968) );
  INV_X1 U7478 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5963) );
  OR2_X1 U7479 ( .A1(n5931), .A2(n5963), .ZN(n5967) );
  NAND2_X1 U7480 ( .A1(n5964), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5965) );
  AND2_X1 U7481 ( .A1(n5980), .A2(n5965), .ZN(n7908) );
  OR2_X1 U7482 ( .A1(n5900), .A2(n7908), .ZN(n5966) );
  NAND4_X1 U7483 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n8087)
         );
  OR2_X1 U7484 ( .A1(n5975), .A2(n5814), .ZN(n5970) );
  XNOR2_X1 U7485 ( .A(n5970), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U7486 ( .A1(n6424), .A2(n7774), .ZN(n5972) );
  NAND2_X1 U7487 ( .A1(n6300), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n5971) );
  OAI211_X1 U7488 ( .C1(n7621), .C2(n8126), .A(n5972), .B(n5971), .ZN(n9814)
         );
  AND2_X1 U7489 ( .A1(n8087), .A2(n9814), .ZN(n5973) );
  NAND2_X1 U7490 ( .A1(n6428), .A2(n7774), .ZN(n5977) );
  OR2_X1 U7491 ( .A1(n6005), .A2(n5814), .ZN(n5988) );
  XNOR2_X1 U7492 ( .A(n5988), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9646) );
  AOI22_X1 U7493 ( .A1(n6300), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6083), .B2(
        n9646), .ZN(n5976) );
  NAND2_X1 U7494 ( .A1(n6186), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5985) );
  INV_X1 U7495 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7496 ( .A1(n4413), .A2(n5978), .ZN(n5984) );
  INV_X1 U7497 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7498 ( .A1(n5931), .A2(n5979), .ZN(n5983) );
  NAND2_X1 U7499 ( .A1(n5980), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5981) );
  AND2_X1 U7500 ( .A1(n5995), .A2(n5981), .ZN(n8037) );
  OR2_X1 U7501 ( .A1(n5900), .A2(n8037), .ZN(n5982) );
  NAND4_X1 U7502 ( .A1(n5985), .A2(n5984), .A3(n5983), .A4(n5982), .ZN(n8086)
         );
  NAND2_X1 U7503 ( .A1(n9822), .A2(n8086), .ZN(n7686) );
  NAND2_X1 U7504 ( .A1(n7688), .A2(n7686), .ZN(n7822) );
  INV_X1 U7505 ( .A(n9822), .ZN(n8044) );
  NAND2_X1 U7506 ( .A1(n8044), .A2(n8086), .ZN(n5986) );
  NAND2_X1 U7507 ( .A1(n7263), .A2(n5986), .ZN(n8367) );
  NAND2_X1 U7508 ( .A1(n6534), .A2(n7774), .ZN(n5992) );
  INV_X1 U7509 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7510 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7511 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5990) );
  XNOR2_X1 U7512 ( .A(n5990), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9661) );
  AOI22_X1 U7513 ( .A1(n6300), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6083), .B2(
        n9661), .ZN(n5991) );
  NAND2_X1 U7514 ( .A1(n5992), .A2(n5991), .ZN(n9831) );
  NAND2_X1 U7515 ( .A1(n6186), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6000) );
  INV_X1 U7516 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8375) );
  OR2_X1 U7517 ( .A1(n4413), .A2(n8375), .ZN(n5999) );
  INV_X1 U7518 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5993) );
  OR2_X1 U7519 ( .A1(n5931), .A2(n5993), .ZN(n5998) );
  INV_X1 U7520 ( .A(n5995), .ZN(n5994) );
  NAND2_X1 U7521 ( .A1(n5994), .A2(n7945), .ZN(n6013) );
  NAND2_X1 U7522 ( .A1(n5995), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5996) );
  AND2_X1 U7523 ( .A1(n6013), .A2(n5996), .ZN(n8374) );
  OR2_X1 U7524 ( .A1(n5900), .A2(n8374), .ZN(n5997) );
  NAND4_X1 U7525 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n8353)
         );
  OR2_X1 U7526 ( .A1(n9831), .A2(n8353), .ZN(n6001) );
  NAND2_X1 U7527 ( .A1(n8367), .A2(n6001), .ZN(n6003) );
  NAND2_X1 U7528 ( .A1(n9831), .A2(n8353), .ZN(n6002) );
  NAND2_X1 U7529 ( .A1(n6536), .A2(n7774), .ZN(n6008) );
  OR2_X1 U7530 ( .A1(n6019), .A2(n5814), .ZN(n6006) );
  XNOR2_X1 U7531 ( .A(n6006), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9679) );
  AOI22_X1 U7532 ( .A1(n6300), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6083), .B2(
        n9679), .ZN(n6007) );
  NAND2_X1 U7533 ( .A1(n6008), .A2(n6007), .ZN(n8533) );
  NAND2_X1 U7534 ( .A1(n6186), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6018) );
  INV_X1 U7535 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7536 ( .A1(n5931), .A2(n6009), .ZN(n6017) );
  INV_X1 U7537 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7538 ( .A1(n4413), .A2(n6010), .ZN(n6016) );
  INV_X1 U7539 ( .A(n6013), .ZN(n6012) );
  NAND2_X1 U7540 ( .A1(n6012), .A2(n6011), .ZN(n6023) );
  NAND2_X1 U7541 ( .A1(n6013), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6014) );
  AND2_X1 U7542 ( .A1(n6023), .A2(n6014), .ZN(n8349) );
  OR2_X1 U7543 ( .A1(n5900), .A2(n8349), .ZN(n6015) );
  NAND4_X1 U7544 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n8337)
         );
  AND2_X1 U7545 ( .A1(n8533), .A2(n8337), .ZN(n7693) );
  OR2_X1 U7546 ( .A1(n8533), .A2(n8337), .ZN(n7692) );
  NAND2_X1 U7547 ( .A1(n6539), .A2(n7774), .ZN(n6022) );
  NAND2_X1 U7548 ( .A1(n6071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7549 ( .A1(n6044), .A2(n6042), .ZN(n6030) );
  OR2_X1 U7550 ( .A1(n6044), .A2(n6042), .ZN(n6020) );
  AOI22_X1 U7551 ( .A1(n6300), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6083), .B2(
        n9694), .ZN(n6021) );
  NAND2_X1 U7552 ( .A1(n5869), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6028) );
  INV_X1 U7553 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8425) );
  OR2_X1 U7554 ( .A1(n5931), .A2(n8425), .ZN(n6027) );
  OR2_X2 U7555 ( .A1(n6023), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7556 ( .A1(n6023), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6024) );
  AND2_X1 U7557 ( .A1(n6036), .A2(n6024), .ZN(n8340) );
  OR2_X1 U7558 ( .A1(n5900), .A2(n8340), .ZN(n6026) );
  INV_X1 U7559 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10082) );
  OR2_X1 U7560 ( .A1(n4416), .A2(n10082), .ZN(n6025) );
  NAND4_X1 U7561 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n8351)
         );
  NOR2_X1 U7562 ( .A1(n8527), .A2(n8351), .ZN(n6029) );
  INV_X1 U7563 ( .A(n8527), .ZN(n8342) );
  NAND2_X1 U7564 ( .A1(n6573), .A2(n7774), .ZN(n6033) );
  NAND2_X1 U7565 ( .A1(n6030), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  XNOR2_X1 U7566 ( .A(n6031), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8141) );
  AOI22_X1 U7567 ( .A1(n6300), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6083), .B2(
        n8141), .ZN(n6032) );
  NAND2_X1 U7568 ( .A1(n6186), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6041) );
  INV_X1 U7569 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10085) );
  OR2_X1 U7570 ( .A1(n5931), .A2(n10085), .ZN(n6040) );
  INV_X1 U7571 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8331) );
  OR2_X1 U7572 ( .A1(n4413), .A2(n8331), .ZN(n6039) );
  INV_X1 U7573 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7574 ( .A1(n6035), .A2(n6034), .ZN(n6048) );
  NAND2_X1 U7575 ( .A1(n6036), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6037) );
  AND2_X1 U7576 ( .A1(n6048), .A2(n6037), .ZN(n8072) );
  OR2_X1 U7577 ( .A1(n5900), .A2(n8072), .ZN(n6038) );
  NAND4_X1 U7578 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n8338)
         );
  AND2_X1 U7579 ( .A1(n8522), .A2(n8338), .ZN(n7700) );
  NAND2_X1 U7580 ( .A1(n6681), .A2(n7774), .ZN(n6047) );
  NAND2_X1 U7581 ( .A1(n6042), .A2(n10016), .ZN(n6068) );
  NAND2_X1 U7582 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7583 ( .A1(n6044), .A2(n6043), .ZN(n6055) );
  INV_X1 U7584 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U7585 ( .A(n6055), .B(n6045), .ZN(n8147) );
  AOI22_X1 U7586 ( .A1(n6300), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6083), .B2(
        n8147), .ZN(n6046) );
  NAND2_X1 U7587 ( .A1(n6186), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6053) );
  INV_X1 U7588 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8321) );
  OR2_X1 U7589 ( .A1(n4413), .A2(n8321), .ZN(n6052) );
  INV_X1 U7590 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10040) );
  OR2_X1 U7591 ( .A1(n5931), .A2(n10040), .ZN(n6051) );
  NAND2_X1 U7592 ( .A1(n6048), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6049) );
  AND2_X1 U7593 ( .A1(n6061), .A2(n6049), .ZN(n8322) );
  OR2_X1 U7594 ( .A1(n5900), .A2(n8322), .ZN(n6050) );
  NAND2_X1 U7595 ( .A1(n8515), .A2(n7959), .ZN(n6253) );
  NAND2_X1 U7596 ( .A1(n7719), .A2(n6253), .ZN(n8317) );
  INV_X1 U7597 ( .A(n8515), .ZN(n6054) );
  NAND2_X1 U7598 ( .A1(n6685), .A2(n7774), .ZN(n6058) );
  OAI21_X1 U7599 ( .B1(n6055), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6056) );
  XNOR2_X1 U7600 ( .A(n6056), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8152) );
  AOI22_X1 U7601 ( .A1(n6300), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6083), .B2(
        n8152), .ZN(n6057) );
  NAND2_X1 U7602 ( .A1(n6186), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6066) );
  INV_X1 U7603 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8417) );
  OR2_X1 U7604 ( .A1(n5931), .A2(n8417), .ZN(n6065) );
  INV_X1 U7605 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8310) );
  OR2_X1 U7606 ( .A1(n5837), .A2(n8310), .ZN(n6064) );
  INV_X1 U7607 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7608 ( .A1(n6061), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6062) );
  AND2_X1 U7609 ( .A1(n6075), .A2(n6062), .ZN(n8311) );
  OR2_X1 U7610 ( .A1(n5900), .A2(n8311), .ZN(n6063) );
  NAND2_X1 U7611 ( .A1(n8509), .A2(n7963), .ZN(n7735) );
  NAND2_X1 U7612 ( .A1(n7721), .A2(n7735), .ZN(n8305) );
  INV_X1 U7613 ( .A(n8509), .ZN(n6067) );
  NAND2_X1 U7614 ( .A1(n6950), .A2(n7774), .ZN(n6074) );
  INV_X1 U7615 ( .A(n6068), .ZN(n6070) );
  NOR2_X1 U7616 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6069) );
  NAND2_X1 U7617 ( .A1(n4494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U7618 ( .A(n6072), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U7619 ( .A1(n6300), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6083), .B2(
        n10211), .ZN(n6073) );
  NAND2_X1 U7620 ( .A1(n5869), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6080) );
  INV_X1 U7621 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8414) );
  OR2_X1 U7622 ( .A1(n5931), .A2(n8414), .ZN(n6079) );
  OR2_X2 U7623 ( .A1(n6075), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7624 ( .A1(n6075), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6076) );
  AND2_X1 U7625 ( .A1(n6088), .A2(n6076), .ZN(n8297) );
  OR2_X1 U7626 ( .A1(n5900), .A2(n8297), .ZN(n6078) );
  INV_X1 U7627 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10168) );
  OR2_X1 U7628 ( .A1(n4417), .A2(n10168), .ZN(n6077) );
  NAND2_X1 U7629 ( .A1(n7601), .A2(n7975), .ZN(n6081) );
  NAND2_X1 U7630 ( .A1(n7030), .A2(n7774), .ZN(n6085) );
  NAND2_X1 U7631 ( .A1(n6177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6082) );
  AOI22_X1 U7632 ( .A1(n6300), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7840), .B2(
        n6083), .ZN(n6084) );
  NAND2_X1 U7633 ( .A1(n6186), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6093) );
  INV_X1 U7634 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8286) );
  OR2_X1 U7635 ( .A1(n5837), .A2(n8286), .ZN(n6092) );
  INV_X1 U7636 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9986) );
  OR2_X1 U7637 ( .A1(n5931), .A2(n9986), .ZN(n6091) );
  INV_X1 U7638 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7639 ( .A1(n6088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6089) );
  AND2_X1 U7640 ( .A1(n6096), .A2(n6089), .ZN(n7918) );
  OR2_X1 U7641 ( .A1(n5900), .A2(n7918), .ZN(n6090) );
  NAND2_X1 U7642 ( .A1(n8498), .A2(n8050), .ZN(n7740) );
  INV_X1 U7643 ( .A(n8498), .ZN(n7924) );
  NAND2_X1 U7644 ( .A1(n7088), .A2(n7774), .ZN(n6095) );
  NAND2_X1 U7645 ( .A1(n6300), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7646 ( .A1(n5869), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6101) );
  INV_X1 U7647 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8409) );
  OR2_X1 U7648 ( .A1(n5931), .A2(n8409), .ZN(n6100) );
  NAND2_X1 U7649 ( .A1(n6096), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6097) );
  AND2_X1 U7650 ( .A1(n6106), .A2(n6097), .ZN(n8011) );
  OR2_X1 U7651 ( .A1(n5900), .A2(n8011), .ZN(n6099) );
  INV_X1 U7652 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8491) );
  OR2_X1 U7653 ( .A1(n4416), .A2(n8491), .ZN(n6098) );
  NAND4_X1 U7654 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n8284)
         );
  AND2_X1 U7655 ( .A1(n7603), .A2(n8284), .ZN(n6255) );
  INV_X1 U7656 ( .A(n8284), .ZN(n7920) );
  NOR2_X1 U7657 ( .A1(n8492), .A2(n8284), .ZN(n8261) );
  NAND2_X1 U7658 ( .A1(n7156), .A2(n7774), .ZN(n6103) );
  NAND2_X1 U7659 ( .A1(n6300), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7660 ( .A1(n6104), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6112) );
  INV_X1 U7661 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8485) );
  OR2_X1 U7662 ( .A1(n4416), .A2(n8485), .ZN(n6111) );
  NAND2_X1 U7663 ( .A1(n6106), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6107) );
  AND2_X1 U7664 ( .A1(n6117), .A2(n6107), .ZN(n8266) );
  OR2_X1 U7665 ( .A1(n5900), .A2(n8266), .ZN(n6110) );
  INV_X1 U7666 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7667 ( .A1(n5837), .A2(n6108), .ZN(n6109) );
  NAND2_X1 U7668 ( .A1(n8486), .A2(n7853), .ZN(n7731) );
  NAND2_X1 U7669 ( .A1(n7742), .A2(n7731), .ZN(n8260) );
  INV_X1 U7670 ( .A(n8486), .ZN(n6113) );
  NAND2_X1 U7671 ( .A1(n8263), .A2(n6114), .ZN(n8249) );
  NAND2_X1 U7672 ( .A1(n7272), .A2(n7774), .ZN(n6116) );
  NAND2_X1 U7673 ( .A1(n6300), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7674 ( .A1(n6117), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7675 ( .A1(n6128), .A2(n6118), .ZN(n8247) );
  NAND2_X1 U7676 ( .A1(n6303), .A2(n8247), .ZN(n6123) );
  INV_X1 U7677 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7678 ( .A1(n4413), .A2(n6119), .ZN(n6122) );
  INV_X1 U7679 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8403) );
  OR2_X1 U7680 ( .A1(n5931), .A2(n8403), .ZN(n6121) );
  INV_X1 U7681 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8479) );
  OR2_X1 U7682 ( .A1(n4417), .A2(n8479), .ZN(n6120) );
  NAND4_X1 U7683 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n8264)
         );
  OR2_X1 U7684 ( .A1(n8480), .A2(n8264), .ZN(n6125) );
  NAND2_X1 U7685 ( .A1(n8480), .A2(n8264), .ZN(n6124) );
  NAND2_X1 U7686 ( .A1(n7286), .A2(n7774), .ZN(n6127) );
  NAND2_X1 U7687 ( .A1(n6300), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7688 ( .A1(n6128), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7689 ( .A1(n6139), .A2(n6129), .ZN(n8242) );
  NAND2_X1 U7690 ( .A1(n8242), .A2(n6303), .ZN(n6133) );
  NAND2_X1 U7691 ( .A1(n5869), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7692 ( .A1(n6104), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7693 ( .A1(n6186), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7694 ( .A1(n8474), .A2(n8251), .ZN(n6134) );
  NAND2_X1 U7695 ( .A1(n7317), .A2(n7774), .ZN(n6136) );
  NAND2_X1 U7696 ( .A1(n6300), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6135) );
  INV_X1 U7697 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7698 ( .A1(n6139), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7699 ( .A1(n6150), .A2(n6140), .ZN(n8233) );
  NAND2_X1 U7700 ( .A1(n8233), .A2(n6303), .ZN(n6143) );
  AOI22_X1 U7701 ( .A1(n5869), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n6104), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7702 ( .A1(n6186), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7703 ( .A1(n8231), .A2(n7984), .ZN(n6145) );
  NOR2_X1 U7704 ( .A1(n8231), .A2(n7984), .ZN(n6144) );
  NAND2_X1 U7705 ( .A1(n8556), .A2(n7774), .ZN(n6147) );
  NAND2_X1 U7706 ( .A1(n6300), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6146) );
  INV_X1 U7707 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10120) );
  INV_X1 U7708 ( .A(n6150), .ZN(n6149) );
  INV_X1 U7709 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7710 ( .A1(n6149), .A2(n6148), .ZN(n6157) );
  NAND2_X1 U7711 ( .A1(n6150), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7712 ( .A1(n6157), .A2(n6151), .ZN(n8217) );
  NAND2_X1 U7713 ( .A1(n8217), .A2(n6303), .ZN(n6153) );
  AOI22_X1 U7714 ( .A1(n5869), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n6104), .B2(
        P2_REG1_REG_25__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7715 ( .A1(n8462), .A2(n8229), .ZN(n7760) );
  NAND2_X1 U7716 ( .A1(n8214), .A2(n7760), .ZN(n6154) );
  OR2_X1 U7717 ( .A1(n8462), .A2(n8229), .ZN(n7624) );
  NAND2_X1 U7718 ( .A1(n8554), .A2(n7774), .ZN(n6156) );
  NAND2_X1 U7719 ( .A1(n6300), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6155) );
  OR2_X2 U7720 ( .A1(n6157), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7721 ( .A1(n6157), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7722 ( .A1(n6170), .A2(n6158), .ZN(n8208) );
  NAND2_X1 U7723 ( .A1(n8208), .A2(n6303), .ZN(n6163) );
  INV_X1 U7724 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U7725 ( .A1(n5869), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7726 ( .A1(n6104), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7727 ( .C1(n8456), .C2(n4416), .A(n6160), .B(n6159), .ZN(n6161)
         );
  INV_X1 U7728 ( .A(n6161), .ZN(n6162) );
  NAND2_X2 U7729 ( .A1(n6163), .A2(n6162), .ZN(n8215) );
  NOR2_X1 U7730 ( .A1(n8457), .A2(n8215), .ZN(n6164) );
  NAND2_X1 U7731 ( .A1(n8457), .A2(n8215), .ZN(n6165) );
  NAND2_X1 U7732 ( .A1(n8550), .A2(n7774), .ZN(n6167) );
  NAND2_X1 U7733 ( .A1(n6300), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6166) );
  INV_X1 U7734 ( .A(n6170), .ZN(n6169) );
  INV_X1 U7735 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7736 ( .A1(n6169), .A2(n6168), .ZN(n6184) );
  NAND2_X1 U7737 ( .A1(n6170), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7738 ( .A1(n6184), .A2(n6171), .ZN(n7890) );
  NAND2_X1 U7739 ( .A1(n7890), .A2(n6303), .ZN(n6176) );
  INV_X1 U7740 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U7741 ( .A1(n6104), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7742 ( .A1(n5869), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6172) );
  OAI211_X1 U7743 ( .C1(n8448), .C2(n4417), .A(n6173), .B(n6172), .ZN(n6174)
         );
  INV_X1 U7744 ( .A(n6174), .ZN(n6175) );
  NAND2_X1 U7745 ( .A1(n8451), .A2(n8062), .ZN(n8188) );
  NAND2_X1 U7746 ( .A1(n8190), .A2(n8188), .ZN(n7831) );
  XOR2_X1 U7747 ( .A(n6287), .B(n7831), .Z(n6198) );
  NAND2_X1 U7748 ( .A1(n6178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7749 ( .A(n6179), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6612) );
  INV_X1 U7750 ( .A(n7784), .ZN(n6263) );
  NAND2_X1 U7751 ( .A1(n6612), .A2(n6263), .ZN(n7796) );
  NAND2_X1 U7752 ( .A1(n6182), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7753 ( .A1(n7840), .A2(n7845), .ZN(n6325) );
  OR2_X2 U7754 ( .A1(n6184), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U7755 ( .A1(n6184), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7756 ( .A1(n8174), .A2(n6185), .ZN(n8199) );
  NAND2_X1 U7757 ( .A1(n8199), .A2(n6303), .ZN(n6191) );
  INV_X1 U7758 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U7759 ( .A1(n6186), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7760 ( .A1(n6104), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7761 ( .C1(n4413), .C2(n8198), .A(n6188), .B(n6187), .ZN(n6189)
         );
  INV_X1 U7762 ( .A(n6189), .ZN(n6190) );
  INV_X1 U7763 ( .A(n6192), .ZN(n7842) );
  NAND2_X1 U7764 ( .A1(n7842), .A2(n8158), .ZN(n6193) );
  NAND2_X1 U7765 ( .A1(n7621), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7766 ( .A1(n8085), .A2(n9758), .ZN(n6196) );
  INV_X1 U7767 ( .A(n6194), .ZN(n6623) );
  AND2_X2 U7768 ( .A1(n6623), .A2(n7769), .ZN(n8352) );
  INV_X1 U7769 ( .A(n6202), .ZN(n6200) );
  NAND2_X1 U7770 ( .A1(n6200), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U7771 ( .A(n6214), .B(P2_B_REG_SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7772 ( .A1(n6208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6209) );
  INV_X1 U7773 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U7774 ( .A1(n6222), .A2(n6415), .ZN(n6216) );
  NAND2_X1 U7775 ( .A1(n6213), .A2(n6214), .ZN(n6215) );
  INV_X1 U7776 ( .A(n6617), .ZN(n6274) );
  NAND3_X1 U7777 ( .A1(n6263), .A2(n7845), .A3(n8164), .ZN(n6217) );
  INV_X1 U7778 ( .A(n6613), .ZN(n6218) );
  OR2_X1 U7779 ( .A1(n7783), .A2(n6218), .ZN(n6588) );
  INV_X1 U7780 ( .A(n8560), .ZN(n6219) );
  NAND2_X1 U7781 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6221) );
  NOR2_X1 U7782 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n6226) );
  NOR4_X1 U7783 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6225) );
  NOR4_X1 U7784 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6224) );
  NOR4_X1 U7785 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6223) );
  NAND4_X1 U7786 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6223), .ZN(n6232)
         );
  NOR4_X1 U7787 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7788 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6229) );
  NOR4_X1 U7789 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6228) );
  NOR4_X1 U7790 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6227) );
  NAND4_X1 U7791 ( .A1(n6230), .A2(n6229), .A3(n6228), .A4(n6227), .ZN(n6231)
         );
  NOR2_X1 U7792 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  AND2_X1 U7793 ( .A1(n6410), .A2(n6584), .ZN(n6330) );
  INV_X1 U7794 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7795 ( .A1(n6222), .A2(n6234), .ZN(n6236) );
  NAND2_X1 U7796 ( .A1(n8560), .A2(n6213), .ZN(n6235) );
  OR2_X1 U7797 ( .A1(n6423), .A2(n6617), .ZN(n6329) );
  NAND2_X1 U7798 ( .A1(n6277), .A2(n6423), .ZN(n6237) );
  NAND2_X1 U7799 ( .A1(n9794), .A2(n7172), .ZN(n6275) );
  MUX2_X1 U7800 ( .A(n6238), .B(n8447), .S(n8376), .Z(n6273) );
  NAND2_X1 U7801 ( .A1(n6896), .A2(n6240), .ZN(n9755) );
  NAND2_X1 U7802 ( .A1(n9755), .A2(n9757), .ZN(n6242) );
  NAND2_X1 U7803 ( .A1(n6242), .A2(n7638), .ZN(n6963) );
  XNOR2_X1 U7804 ( .A(n9759), .B(n6965), .ZN(n7814) );
  NAND2_X1 U7805 ( .A1(n6963), .A2(n7814), .ZN(n6243) );
  NAND2_X1 U7806 ( .A1(n6243), .A2(n7646), .ZN(n6999) );
  INV_X1 U7807 ( .A(n6910), .ZN(n9787) );
  NAND2_X1 U7808 ( .A1(n8093), .A2(n9787), .ZN(n7648) );
  NAND2_X1 U7809 ( .A1(n6999), .A2(n7648), .ZN(n6244) );
  OR2_X1 U7810 ( .A1(n8093), .A2(n9787), .ZN(n7657) );
  NAND2_X1 U7811 ( .A1(n6244), .A2(n7657), .ZN(n7010) );
  INV_X1 U7812 ( .A(n7023), .ZN(n9790) );
  NAND2_X1 U7813 ( .A1(n8092), .A2(n9790), .ZN(n7647) );
  NAND2_X1 U7814 ( .A1(n7010), .A2(n7647), .ZN(n6245) );
  OR2_X1 U7815 ( .A1(n8092), .A2(n9790), .ZN(n7651) );
  NAND2_X1 U7816 ( .A1(n6245), .A2(n7651), .ZN(n7100) );
  INV_X1 U7817 ( .A(n7070), .ZN(n9795) );
  OR2_X1 U7818 ( .A1(n8091), .A2(n9795), .ZN(n7661) );
  NAND2_X1 U7819 ( .A1(n8091), .A2(n9795), .ZN(n7652) );
  NAND2_X1 U7820 ( .A1(n7100), .A2(n7815), .ZN(n6246) );
  NAND2_X1 U7821 ( .A1(n6246), .A2(n7661), .ZN(n7090) );
  INV_X1 U7822 ( .A(n7668), .ZN(n7670) );
  NAND2_X1 U7823 ( .A1(n8088), .A2(n9807), .ZN(n7247) );
  AND2_X2 U7824 ( .A1(n7677), .A2(n7247), .ZN(n7819) );
  NAND2_X1 U7825 ( .A1(n8087), .A2(n7914), .ZN(n7684) );
  AND2_X1 U7826 ( .A1(n7247), .A2(n7684), .ZN(n7678) );
  NAND2_X1 U7827 ( .A1(n7246), .A2(n7678), .ZN(n6247) );
  OR2_X1 U7828 ( .A1(n8087), .A2(n7914), .ZN(n7682) );
  NAND2_X1 U7829 ( .A1(n6247), .A2(n7682), .ZN(n7269) );
  INV_X1 U7830 ( .A(n7688), .ZN(n6248) );
  INV_X1 U7831 ( .A(n8353), .ZN(n8042) );
  OR2_X1 U7832 ( .A1(n9831), .A2(n8042), .ZN(n7695) );
  NAND2_X1 U7833 ( .A1(n9831), .A2(n8042), .ZN(n7696) );
  INV_X1 U7834 ( .A(n8337), .ZN(n8369) );
  OR2_X1 U7835 ( .A1(n8533), .A2(n8369), .ZN(n7705) );
  NAND2_X1 U7836 ( .A1(n8533), .A2(n8369), .ZN(n7704) );
  OR2_X1 U7837 ( .A1(n8527), .A2(n8076), .ZN(n7703) );
  NAND2_X1 U7838 ( .A1(n8345), .A2(n7703), .ZN(n6249) );
  NAND2_X1 U7839 ( .A1(n8527), .A2(n8076), .ZN(n7702) );
  NAND2_X1 U7840 ( .A1(n6249), .A2(n7702), .ZN(n8326) );
  INV_X1 U7841 ( .A(n8338), .ZN(n7594) );
  OR2_X1 U7842 ( .A1(n8522), .A2(n7594), .ZN(n6250) );
  NAND2_X1 U7843 ( .A1(n8326), .A2(n6250), .ZN(n6252) );
  NAND2_X1 U7844 ( .A1(n8522), .A2(n7594), .ZN(n6251) );
  INV_X1 U7845 ( .A(n6253), .ZN(n7724) );
  NAND2_X1 U7846 ( .A1(n6254), .A2(n7721), .ZN(n8291) );
  NAND2_X1 U7847 ( .A1(n8503), .A2(n7975), .ZN(n7807) );
  INV_X1 U7848 ( .A(n6255), .ZN(n7743) );
  AND2_X1 U7849 ( .A1(n7731), .A2(n8257), .ZN(n7729) );
  NAND2_X1 U7850 ( .A1(n8258), .A2(n7729), .ZN(n6257) );
  NAND2_X1 U7851 ( .A1(n6257), .A2(n7742), .ZN(n8246) );
  INV_X1 U7852 ( .A(n8264), .ZN(n7856) );
  OR2_X1 U7853 ( .A1(n8480), .A2(n7856), .ZN(n7745) );
  INV_X1 U7854 ( .A(n8474), .ZN(n6258) );
  NAND2_X1 U7855 ( .A1(n8468), .A2(n7984), .ZN(n7803) );
  NAND2_X1 U7856 ( .A1(n8474), .A2(n8028), .ZN(n8224) );
  AND2_X1 U7857 ( .A1(n7803), .A2(n8224), .ZN(n7753) );
  NAND2_X1 U7858 ( .A1(n8225), .A2(n7753), .ZN(n6260) );
  NAND2_X1 U7859 ( .A1(n6260), .A2(n7804), .ZN(n8212) );
  NOR2_X1 U7860 ( .A1(n8462), .A2(n7866), .ZN(n6262) );
  NAND2_X1 U7861 ( .A1(n8462), .A2(n7866), .ZN(n6261) );
  OAI21_X2 U7862 ( .B1(n8212), .B2(n6262), .A(n6261), .ZN(n8202) );
  XOR2_X1 U7863 ( .A(n7831), .B(n8189), .Z(n8454) );
  AOI21_X1 U7864 ( .B1(n6263), .B2(n7274), .A(n7840), .ZN(n6264) );
  AND2_X1 U7865 ( .A1(n9821), .A2(n6264), .ZN(n6265) );
  INV_X1 U7866 ( .A(n9765), .ZN(n7257) );
  AND2_X1 U7867 ( .A1(n9767), .A2(n6612), .ZN(n6894) );
  INV_X1 U7868 ( .A(n6894), .ZN(n6266) );
  NAND2_X1 U7869 ( .A1(n7257), .A2(n6266), .ZN(n6267) );
  INV_X1 U7870 ( .A(n6268), .ZN(n6269) );
  AOI22_X1 U7871 ( .A1(n8451), .A2(n8378), .B1(n9768), .B2(n7890), .ZN(n6270)
         );
  INV_X1 U7872 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7873 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7874 ( .A1(n6276), .A2(n6277), .ZN(n6280) );
  INV_X1 U7875 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U7876 ( .A1(n6278), .A2(n6423), .ZN(n6279) );
  MUX2_X1 U7877 ( .A(n6282), .B(n8447), .S(n9851), .Z(n6286) );
  INV_X1 U7878 ( .A(n9821), .ZN(n9832) );
  NAND2_X1 U7879 ( .A1(n9851), .A2(n9832), .ZN(n8383) );
  NAND2_X1 U7880 ( .A1(n8451), .A2(n8428), .ZN(n6283) );
  NAND2_X1 U7881 ( .A1(n6286), .A2(n6285), .ZN(P2_U3486) );
  NAND2_X1 U7882 ( .A1(n6288), .A2(n4459), .ZN(n6290) );
  NAND2_X1 U7883 ( .A1(n7892), .A2(n8062), .ZN(n6289) );
  MUX2_X1 U7884 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5047), .Z(n6298) );
  XNOR2_X1 U7885 ( .A(n6298), .B(n9965), .ZN(n6297) );
  NAND2_X1 U7886 ( .A1(n7849), .A2(n7774), .ZN(n6295) );
  NAND2_X1 U7887 ( .A1(n6300), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6294) );
  NOR2_X1 U7888 ( .A1(n8443), .A2(n8085), .ZN(n6296) );
  INV_X1 U7889 ( .A(n6298), .ZN(n6299) );
  INV_X1 U7890 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8545) );
  INV_X1 U7891 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7567) );
  MUX2_X1 U7892 ( .A(n8545), .B(n7567), .S(n5047), .Z(n7319) );
  NAND2_X1 U7893 ( .A1(n7566), .A2(n7774), .ZN(n6302) );
  NAND2_X1 U7894 ( .A1(n6300), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6301) );
  INV_X1 U7895 ( .A(n8174), .ZN(n6304) );
  NAND2_X1 U7896 ( .A1(n6304), .A2(n6303), .ZN(n7790) );
  INV_X1 U7897 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10113) );
  NAND2_X1 U7898 ( .A1(n6104), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7899 ( .A1(n5869), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6305) );
  OAI211_X1 U7900 ( .C1(n4416), .C2(n10113), .A(n6306), .B(n6305), .ZN(n6307)
         );
  INV_X1 U7901 ( .A(n6307), .ZN(n6308) );
  AND2_X2 U7902 ( .A1(n7790), .A2(n6308), .ZN(n8084) );
  OR2_X2 U7903 ( .A1(n6333), .A2(n8084), .ZN(n7793) );
  NAND2_X1 U7904 ( .A1(n6333), .A2(n8084), .ZN(n7795) );
  XNOR2_X1 U7905 ( .A(n6309), .B(n7802), .ZN(n6322) );
  INV_X1 U7906 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U7907 ( .A1(n5869), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7908 ( .A1(n6104), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6310) );
  OAI211_X1 U7909 ( .C1(n8440), .C2(n4417), .A(n6311), .B(n6310), .ZN(n6312)
         );
  INV_X1 U7910 ( .A(n6312), .ZN(n6313) );
  NAND2_X1 U7911 ( .A1(n7790), .A2(n6313), .ZN(n8083) );
  AND2_X1 U7912 ( .A1(n7621), .A2(P2_B_REG_SCAN_IN), .ZN(n6314) );
  NOR2_X1 U7913 ( .A1(n8370), .A2(n6314), .ZN(n8172) );
  AOI22_X1 U7914 ( .A1(n8352), .A2(n8085), .B1(n8083), .B2(n8172), .ZN(n6321)
         );
  NAND2_X1 U7915 ( .A1(n8443), .A2(n7888), .ZN(n6316) );
  AND2_X1 U7916 ( .A1(n8188), .A2(n6316), .ZN(n6315) );
  INV_X1 U7917 ( .A(n6316), .ZN(n6319) );
  OR2_X1 U7918 ( .A1(n8443), .A2(n7888), .ZN(n6317) );
  AND2_X1 U7919 ( .A1(n8190), .A2(n6317), .ZN(n6318) );
  XNOR2_X1 U7920 ( .A(n7791), .B(n7802), .ZN(n6323) );
  NAND2_X1 U7921 ( .A1(n6323), .A2(n9765), .ZN(n6320) );
  INV_X1 U7922 ( .A(n6323), .ZN(n8187) );
  INV_X1 U7923 ( .A(n6325), .ZN(n6326) );
  NAND2_X1 U7924 ( .A1(n7835), .A2(n6326), .ZN(n6328) );
  AND2_X1 U7925 ( .A1(n7783), .A2(n9821), .ZN(n6327) );
  NAND2_X1 U7926 ( .A1(n6328), .A2(n6327), .ZN(n6599) );
  NAND2_X1 U7927 ( .A1(n6599), .A2(n8341), .ZN(n6587) );
  NAND3_X1 U7928 ( .A1(n6423), .A2(n6617), .A3(n6584), .ZN(n6594) );
  NAND2_X1 U7929 ( .A1(n6587), .A2(n6607), .ZN(n6332) );
  INV_X1 U7930 ( .A(n6674), .ZN(n6606) );
  INV_X1 U7931 ( .A(n6328), .ZN(n6601) );
  INV_X1 U7932 ( .A(n6329), .ZN(n6585) );
  OAI21_X1 U7933 ( .B1(n6606), .B2(n6601), .A(n6604), .ZN(n6331) );
  OR2_X1 U7934 ( .A1(n9835), .A2(n9821), .ZN(n8433) );
  NAND2_X1 U7935 ( .A1(n7849), .A2(n7420), .ZN(n6335) );
  INV_X1 U7936 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7850) );
  OR2_X1 U7937 ( .A1(n5259), .A2(n7850), .ZN(n6334) );
  NAND2_X1 U7938 ( .A1(n9136), .A2(n5167), .ZN(n6339) );
  NAND2_X1 U7939 ( .A1(n8720), .A2(n6337), .ZN(n6338) );
  NAND2_X1 U7940 ( .A1(n6339), .A2(n6338), .ZN(n6341) );
  XNOR2_X1 U7941 ( .A(n6341), .B(n4419), .ZN(n6344) );
  AOI22_X1 U7942 ( .A1(n9136), .A2(n6342), .B1(n5167), .B2(n8720), .ZN(n6343)
         );
  XNOR2_X1 U7943 ( .A(n6344), .B(n6343), .ZN(n6350) );
  NAND3_X1 U7944 ( .A1(n6345), .A2(n6350), .A3(n8709), .ZN(n6364) );
  INV_X1 U7945 ( .A(n6349), .ZN(n6347) );
  INV_X1 U7946 ( .A(n6350), .ZN(n6346) );
  NAND4_X1 U7947 ( .A1(n6348), .A2(n6347), .A3(n6346), .A4(n8709), .ZN(n6363)
         );
  NAND3_X1 U7948 ( .A1(n6350), .A2(n8709), .A3(n6349), .ZN(n6362) );
  OR2_X1 U7949 ( .A1(n8698), .A2(n8927), .ZN(n6358) );
  NAND2_X1 U7950 ( .A1(n6416), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6356) );
  INV_X1 U7951 ( .A(n6351), .ZN(n8909) );
  NAND2_X1 U7952 ( .A1(n6352), .A2(n8909), .ZN(n6355) );
  NAND2_X1 U7953 ( .A1(n7423), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7954 ( .A1(n5248), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6353) );
  NAND4_X1 U7955 ( .A1(n6356), .A2(n6355), .A3(n6354), .A4(n6353), .ZN(n8719)
         );
  NAND2_X1 U7956 ( .A1(n8719), .A2(n8859), .ZN(n6357) );
  AND2_X1 U7957 ( .A1(n6358), .A2(n6357), .ZN(n8940) );
  OAI22_X1 U7958 ( .A1(n8940), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9964), .ZN(n6360) );
  NOR2_X1 U7959 ( .A1(n4643), .A2(n8717), .ZN(n6359) );
  AOI211_X1 U7960 ( .C1(n8713), .C2(n8935), .A(n6360), .B(n6359), .ZN(n6361)
         );
  NAND4_X1 U7961 ( .A1(n6364), .A2(n6363), .A3(n6362), .A4(n6361), .ZN(
        P1_U3220) );
  INV_X1 U7962 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6365) );
  NOR2_X1 U7963 ( .A1(n9851), .A2(n6365), .ZN(n6366) );
  INV_X4 U7964 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7965 ( .A1(n5166), .A2(P1_U3086), .ZN(n6370) );
  INV_X1 U7966 ( .A(n6783), .ZN(n6411) );
  NAND2_X1 U7967 ( .A1(n7783), .A2(n6590), .ZN(n6371) );
  NAND2_X1 U7968 ( .A1(n6371), .A2(n6783), .ZN(n6652) );
  NAND2_X1 U7969 ( .A1(n6652), .A2(n7621), .ZN(n6372) );
  NAND2_X1 U7970 ( .A1(n6372), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X2 U7971 ( .A1(n4418), .A2(P1_U3086), .ZN(n7620) );
  OAI222_X1 U7972 ( .A1(n7620), .A2(n6373), .B1(n7569), .B2(n6374), .C1(
        P1_U3086), .C2(n6446), .ZN(P1_U3353) );
  INV_X2 U7973 ( .A(n8552), .ZN(n8557) );
  OAI222_X1 U7974 ( .A1(n8557), .A2(n10034), .B1(n8559), .B2(n6377), .C1(n6747), .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U7975 ( .A(n6662), .ZN(n6809) );
  OAI222_X1 U7976 ( .A1(n8557), .A2(n6375), .B1(n8559), .B2(n6374), .C1(n6809), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  OAI222_X1 U7977 ( .A1(n7620), .A2(n6376), .B1(n6444), .B2(P1_U3086), .C1(
        n7569), .C2(n6385), .ZN(P1_U3354) );
  OAI222_X1 U7978 ( .A1(n7620), .A2(n6378), .B1(n7569), .B2(n6377), .C1(
        P1_U3086), .C2(n8772), .ZN(P1_U3352) );
  OAI222_X1 U7979 ( .A1(n7620), .A2(n6379), .B1(n7569), .B2(n6383), .C1(
        P1_U3086), .C2(n8783), .ZN(P1_U3351) );
  OAI222_X1 U7980 ( .A1(n9600), .A2(P2_U3151), .B1(n8559), .B2(n6381), .C1(
        n6380), .C2(n8557), .ZN(P2_U3290) );
  OAI222_X1 U7981 ( .A1(n7620), .A2(n6382), .B1(n7569), .B2(n6381), .C1(
        P1_U3086), .C2(n6476), .ZN(P1_U3350) );
  OAI222_X1 U7982 ( .A1(n8557), .A2(n6384), .B1(n8559), .B2(n6383), .C1(n9591), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  OAI222_X1 U7983 ( .A1(n6794), .A2(P2_U3151), .B1(n8557), .B2(n6386), .C1(
        n8559), .C2(n6385), .ZN(P2_U3294) );
  OAI222_X1 U7984 ( .A1(n6860), .A2(P2_U3151), .B1(n8559), .B2(n6388), .C1(
        n6387), .C2(n8557), .ZN(P2_U3289) );
  OAI222_X1 U7985 ( .A1(n7620), .A2(n6389), .B1(n7569), .B2(n6388), .C1(
        P1_U3086), .C2(n6489), .ZN(P1_U3349) );
  OAI222_X1 U7986 ( .A1(n7620), .A2(n6390), .B1(n7569), .B2(n6392), .C1(
        P1_U3086), .C2(n6509), .ZN(P1_U3348) );
  INV_X1 U7987 ( .A(n6975), .ZN(n6853) );
  OAI222_X1 U7988 ( .A1(n6853), .A2(P2_U3151), .B1(n8559), .B2(n6392), .C1(
        n6391), .C2(n8557), .ZN(P2_U3288) );
  AOI22_X1 U7989 ( .A1(n6520), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6686), .ZN(n6393) );
  OAI21_X1 U7990 ( .B1(n6395), .B2(n7569), .A(n6393), .ZN(P1_U3347) );
  INV_X1 U7991 ( .A(n8108), .ZN(n8130) );
  OAI222_X1 U7992 ( .A1(n8130), .A2(P2_U3151), .B1(n8559), .B2(n6395), .C1(
        n6394), .C2(n8557), .ZN(P2_U3287) );
  NAND2_X1 U7993 ( .A1(n9457), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U7994 ( .B1(n9457), .B2(n6398), .A(n6397), .ZN(P1_U3439) );
  INV_X1 U7995 ( .A(n8818), .ZN(n6524) );
  OAI222_X1 U7996 ( .A1(n7569), .A2(n6401), .B1(n6524), .B2(P1_U3086), .C1(
        n6399), .C2(n7620), .ZN(P1_U3346) );
  OAI222_X1 U7997 ( .A1(P2_U3151), .A2(n8128), .B1(n8559), .B2(n6401), .C1(
        n6400), .C2(n8557), .ZN(P2_U3286) );
  INV_X1 U7998 ( .A(n9457), .ZN(n9456) );
  OR2_X1 U7999 ( .A1(n9457), .A2(n6402), .ZN(n6403) );
  OAI21_X1 U8000 ( .B1(n9456), .B2(n6404), .A(n6403), .ZN(P1_U3440) );
  OAI21_X1 U8001 ( .B1(P1_U3973), .B2(n5036), .A(n6405), .ZN(P1_U3554) );
  NAND2_X1 U8002 ( .A1(n6407), .A2(n7460), .ZN(n6406) );
  AND2_X1 U8003 ( .A1(n6406), .A2(n5235), .ZN(n6438) );
  INV_X1 U8004 ( .A(n6438), .ZN(n6408) );
  OR2_X1 U8005 ( .A1(n6407), .A2(P1_U3086), .ZN(n7562) );
  NAND2_X1 U8006 ( .A1(n7562), .A2(n7559), .ZN(n6437) );
  NOR2_X1 U8007 ( .A1(n9305), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8008 ( .A1(n6410), .A2(n6409), .ZN(n6464) );
  NOR4_X1 U8009 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(P2_U3151), .ZN(n6414) );
  AOI21_X1 U8010 ( .B1(n6464), .B2(n6415), .A(n6414), .ZN(P2_U3376) );
  INV_X1 U8011 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8012 ( .A1(n6416), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8013 ( .A1(n5248), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8014 ( .A1(n7423), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6417) );
  AND3_X1 U8015 ( .A1(n6419), .A2(n6418), .A3(n6417), .ZN(n8860) );
  INV_X1 U8016 ( .A(n8860), .ZN(n7427) );
  NAND2_X1 U8017 ( .A1(n7427), .A2(P1_U3973), .ZN(n6420) );
  OAI21_X1 U8018 ( .B1(P1_U3973), .B2(n6421), .A(n6420), .ZN(P1_U3585) );
  NAND2_X1 U8019 ( .A1(n6593), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U8020 ( .B1(n6593), .B2(n6423), .A(n6422), .ZN(P2_U3377) );
  INV_X1 U8021 ( .A(n6424), .ZN(n6427) );
  INV_X1 U8022 ( .A(n8819), .ZN(n9249) );
  OAI222_X1 U8023 ( .A1(n7569), .A2(n6427), .B1(n9249), .B2(P1_U3086), .C1(
        n6425), .C2(n7620), .ZN(P1_U3345) );
  OAI222_X1 U8024 ( .A1(P2_U3151), .A2(n8126), .B1(n8559), .B2(n6427), .C1(
        n6426), .C2(n8557), .ZN(P2_U3285) );
  INV_X1 U8025 ( .A(n6428), .ZN(n6463) );
  AOI22_X1 U8026 ( .A1(n9301), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6686), .ZN(n6429) );
  OAI21_X1 U8027 ( .B1(n6463), .B2(n7569), .A(n6429), .ZN(P1_U3344) );
  INV_X1 U8028 ( .A(n6489), .ZN(n6434) );
  INV_X1 U8029 ( .A(n6476), .ZN(n6431) );
  INV_X1 U8030 ( .A(n8783), .ZN(n6450) );
  INV_X1 U8031 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6733) );
  INV_X1 U8032 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9976) );
  INV_X1 U8033 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6430) );
  XNOR2_X1 U8034 ( .A(n6444), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8741) );
  AND2_X1 U8035 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8754) );
  NAND2_X1 U8036 ( .A1(n8741), .A2(n8754), .ZN(n8740) );
  OAI21_X1 U8037 ( .B1(n6444), .B2(n6430), .A(n8740), .ZN(n8765) );
  XNOR2_X1 U8038 ( .A(n6446), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U8039 ( .A1(n8765), .A2(n8766), .ZN(n8764) );
  OAI21_X1 U8040 ( .B1(n9976), .B2(n6446), .A(n8764), .ZN(n8778) );
  MUX2_X1 U8041 ( .A(n6733), .B(P1_REG2_REG_3__SCAN_IN), .S(n8772), .Z(n8779)
         );
  NAND2_X1 U8042 ( .A1(n8778), .A2(n8779), .ZN(n8777) );
  OAI21_X1 U8043 ( .B1(n6733), .B2(n8772), .A(n8777), .ZN(n8787) );
  INV_X1 U8044 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10117) );
  MUX2_X1 U8045 ( .A(n10117), .B(P1_REG2_REG_4__SCAN_IN), .S(n8783), .Z(n8788)
         );
  XOR2_X1 U8046 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6476), .Z(n6478) );
  AOI21_X1 U8047 ( .B1(n6431), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6477), .ZN(
        n6492) );
  INV_X1 U8048 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6432) );
  MUX2_X1 U8049 ( .A(n6432), .B(P1_REG2_REG_6__SCAN_IN), .S(n6489), .Z(n6433)
         );
  INV_X1 U8050 ( .A(n6433), .ZN(n6491) );
  NOR2_X1 U8051 ( .A1(n6492), .A2(n6491), .ZN(n6490) );
  AOI21_X1 U8052 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6434), .A(n6490), .ZN(
        n6502) );
  INV_X1 U8053 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7118) );
  MUX2_X1 U8054 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7118), .S(n6509), .Z(n6501)
         );
  NOR2_X1 U8055 ( .A1(n6502), .A2(n6501), .ZN(n6500) );
  XNOR2_X1 U8056 ( .A(n6520), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6435) );
  INV_X1 U8057 ( .A(n6435), .ZN(n6441) );
  INV_X1 U8058 ( .A(n6436), .ZN(n6440) );
  NAND2_X1 U8059 ( .A1(n6438), .A2(n6437), .ZN(n9291) );
  OR2_X1 U8060 ( .A1(n5780), .A2(n4421), .ZN(n8752) );
  OAI21_X1 U8061 ( .B1(n6441), .B2(n6440), .A(n9383), .ZN(n6462) );
  INV_X1 U8062 ( .A(n9305), .ZN(n9393) );
  INV_X1 U8063 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8064 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7163) );
  OAI21_X1 U8065 ( .B1(n9393), .B2(n6442), .A(n7163), .ZN(n6443) );
  AOI21_X1 U8066 ( .B1(n6520), .B2(n9347), .A(n6443), .ZN(n6461) );
  INV_X1 U8067 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9566) );
  MUX2_X1 U8068 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9566), .S(n6520), .Z(n6459)
         );
  INV_X1 U8069 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10181) );
  MUX2_X1 U8070 ( .A(n10181), .B(P1_REG1_REG_1__SCAN_IN), .S(n6444), .Z(n8745)
         );
  AND2_X1 U8071 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8744) );
  NAND2_X1 U8072 ( .A1(n8745), .A2(n8744), .ZN(n8743) );
  INV_X1 U8073 ( .A(n6444), .ZN(n8742) );
  NAND2_X1 U8074 ( .A1(n8742), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U8075 ( .A1(n8743), .A2(n6445), .ZN(n8762) );
  XNOR2_X1 U8076 ( .A(n6446), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U8077 ( .A1(n8762), .A2(n8763), .ZN(n8761) );
  INV_X1 U8078 ( .A(n6446), .ZN(n8760) );
  NAND2_X1 U8079 ( .A1(n8760), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8080 ( .A1(n8761), .A2(n6447), .ZN(n8775) );
  XNOR2_X1 U8081 ( .A(n8772), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U8082 ( .A1(n8775), .A2(n8776), .ZN(n8774) );
  INV_X1 U8083 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8084 ( .A1(n8772), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U8085 ( .A1(n8774), .A2(n6449), .ZN(n8790) );
  INV_X1 U8086 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9560) );
  MUX2_X1 U8087 ( .A(n9560), .B(P1_REG1_REG_4__SCAN_IN), .S(n8783), .Z(n8791)
         );
  NAND2_X1 U8088 ( .A1(n8790), .A2(n8791), .ZN(n8789) );
  NAND2_X1 U8089 ( .A1(n6450), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U8090 ( .A1(n8789), .A2(n6451), .ZN(n6481) );
  XNOR2_X1 U8091 ( .A(n6476), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8092 ( .A1(n6481), .A2(n6482), .ZN(n6480) );
  INV_X1 U8093 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6452) );
  OR2_X1 U8094 ( .A1(n6476), .A2(n6452), .ZN(n6453) );
  NAND2_X1 U8095 ( .A1(n6480), .A2(n6453), .ZN(n6494) );
  INV_X1 U8096 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U8097 ( .A(n9563), .B(P1_REG1_REG_6__SCAN_IN), .S(n6489), .Z(n6495)
         );
  NAND2_X1 U8098 ( .A1(n6494), .A2(n6495), .ZN(n6493) );
  OR2_X1 U8099 ( .A1(n6489), .A2(n9563), .ZN(n6454) );
  NAND2_X1 U8100 ( .A1(n6493), .A2(n6454), .ZN(n6504) );
  XNOR2_X1 U8101 ( .A(n6509), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U8102 ( .A1(n6504), .A2(n6505), .ZN(n6503) );
  INV_X1 U8103 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6455) );
  OR2_X1 U8104 ( .A1(n6509), .A2(n6455), .ZN(n6456) );
  NAND2_X1 U8105 ( .A1(n6503), .A2(n6456), .ZN(n6458) );
  INV_X1 U8106 ( .A(n4421), .ZN(n6457) );
  NOR2_X2 U8107 ( .A1(n9291), .A2(n6457), .ZN(n9379) );
  NAND2_X1 U8108 ( .A1(n6458), .A2(n6459), .ZN(n6514) );
  OAI211_X1 U8109 ( .C1(n6459), .C2(n6458), .A(n9379), .B(n6514), .ZN(n6460)
         );
  OAI211_X1 U8110 ( .C1(n6519), .C2(n6462), .A(n6461), .B(n6460), .ZN(P1_U3251) );
  INV_X1 U8111 ( .A(n9646), .ZN(n8124) );
  OAI222_X1 U8112 ( .A1(n8124), .A2(P2_U3151), .B1(n8559), .B2(n6463), .C1(
        n10106), .C2(n8557), .ZN(P2_U3284) );
  INV_X1 U8113 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U8114 ( .A1(n6553), .A2(n6465), .ZN(P2_U3246) );
  INV_X1 U8115 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10032) );
  NOR2_X1 U8116 ( .A1(n6553), .A2(n10032), .ZN(P2_U3255) );
  INV_X1 U8117 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U8118 ( .A1(n6553), .A2(n6466), .ZN(P2_U3250) );
  INV_X1 U8119 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6467) );
  NOR2_X1 U8120 ( .A1(n6553), .A2(n6467), .ZN(P2_U3251) );
  INV_X1 U8121 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U8122 ( .A1(n6553), .A2(n6468), .ZN(P2_U3256) );
  INV_X1 U8123 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U8124 ( .A1(n6553), .A2(n6469), .ZN(P2_U3247) );
  INV_X1 U8125 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U8126 ( .A1(n6553), .A2(n6470), .ZN(P2_U3253) );
  INV_X1 U8127 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U8128 ( .A1(n6553), .A2(n10183), .ZN(P2_U3252) );
  INV_X1 U8129 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6471) );
  NOR2_X1 U8130 ( .A1(n6553), .A2(n6471), .ZN(P2_U3249) );
  INV_X1 U8131 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U8132 ( .A1(n6553), .A2(n6472), .ZN(P2_U3248) );
  INV_X1 U8133 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U8134 ( .A1(n6553), .A2(n6473), .ZN(P2_U3254) );
  INV_X1 U8135 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9962) );
  NOR2_X1 U8136 ( .A1(n6553), .A2(n9962), .ZN(P2_U3257) );
  NAND2_X1 U8137 ( .A1(n9305), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U8138 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n6474) );
  OAI211_X1 U8139 ( .C1(n9389), .C2(n6476), .A(n6475), .B(n6474), .ZN(n6486)
         );
  AOI211_X1 U8140 ( .C1(n6479), .C2(n6478), .A(n6477), .B(n9368), .ZN(n6485)
         );
  OAI211_X1 U8141 ( .C1(n6482), .C2(n6481), .A(n9379), .B(n6480), .ZN(n6483)
         );
  INV_X1 U8142 ( .A(n6483), .ZN(n6484) );
  OR3_X1 U8143 ( .A1(n6486), .A2(n6485), .A3(n6484), .ZN(P1_U3248) );
  NAND2_X1 U8144 ( .A1(n9305), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8145 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6487) );
  OAI211_X1 U8146 ( .C1(n9389), .C2(n6489), .A(n6488), .B(n6487), .ZN(n6499)
         );
  AOI211_X1 U8147 ( .C1(n6492), .C2(n6491), .A(n6490), .B(n9368), .ZN(n6498)
         );
  OAI211_X1 U8148 ( .C1(n6495), .C2(n6494), .A(n9379), .B(n6493), .ZN(n6496)
         );
  INV_X1 U8149 ( .A(n6496), .ZN(n6497) );
  OR3_X1 U8150 ( .A1(n6499), .A2(n6498), .A3(n6497), .ZN(P1_U3249) );
  AOI211_X1 U8151 ( .C1(n6502), .C2(n6501), .A(n9368), .B(n6500), .ZN(n6512)
         );
  OAI211_X1 U8152 ( .C1(n6505), .C2(n6504), .A(n9379), .B(n6503), .ZN(n6506)
         );
  INV_X1 U8153 ( .A(n6506), .ZN(n6511) );
  NAND2_X1 U8154 ( .A1(n9305), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8155 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6507) );
  OAI211_X1 U8156 ( .C1(n9389), .C2(n6509), .A(n6508), .B(n6507), .ZN(n6510)
         );
  OR3_X1 U8157 ( .A1(n6512), .A2(n6511), .A3(n6510), .ZN(P1_U3250) );
  INV_X1 U8158 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U8159 ( .A(n10031), .B(P1_REG1_REG_9__SCAN_IN), .S(n8818), .Z(n6517)
         );
  NAND2_X1 U8160 ( .A1(n6520), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8161 ( .A1(n6514), .A2(n6513), .ZN(n6516) );
  OR2_X1 U8162 ( .A1(n6516), .A2(n6517), .ZN(n8802) );
  INV_X1 U8163 ( .A(n8802), .ZN(n6515) );
  AOI21_X1 U8164 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6528) );
  INV_X1 U8165 ( .A(n9379), .ZN(n9295) );
  NOR2_X1 U8166 ( .A1(n8818), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6518) );
  AOI21_X1 U8167 ( .B1(n8818), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6518), .ZN(
        n6522) );
  OAI21_X1 U8168 ( .B1(n6522), .B2(n6521), .A(n8817), .ZN(n6523) );
  NAND2_X1 U8169 ( .A1(n6523), .A2(n9383), .ZN(n6527) );
  NOR2_X1 U8170 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9975), .ZN(n7217) );
  NOR2_X1 U8171 ( .A1(n9389), .A2(n6524), .ZN(n6525) );
  AOI211_X1 U8172 ( .C1(n9305), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7217), .B(
        n6525), .ZN(n6526) );
  OAI211_X1 U8173 ( .C1(n6528), .C2(n9295), .A(n6527), .B(n6526), .ZN(P1_U3252) );
  OAI21_X1 U8174 ( .B1(n6531), .B2(n6530), .A(n6529), .ZN(n8751) );
  INV_X1 U8175 ( .A(n8709), .ZN(n9260) );
  NAND2_X1 U8176 ( .A1(n9267), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8177 ( .A1(n6708), .A2(n8859), .ZN(n9461) );
  INV_X1 U8178 ( .A(n9446), .ZN(n7474) );
  OAI22_X1 U8179 ( .A1(n9255), .A2(n9461), .B1(n8717), .B2(n7474), .ZN(n6532)
         );
  AOI21_X1 U8180 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6569), .A(n6532), .ZN(
        n6533) );
  OAI21_X1 U8181 ( .B1(n8751), .B2(n9260), .A(n6533), .ZN(P1_U3232) );
  INV_X1 U8182 ( .A(n6534), .ZN(n6535) );
  INV_X1 U8183 ( .A(n8821), .ZN(n9317) );
  OAI222_X1 U8184 ( .A1(n7569), .A2(n6535), .B1(n9317), .B2(P1_U3086), .C1(
        n10070), .C2(n7620), .ZN(P1_U3343) );
  INV_X1 U8185 ( .A(n9661), .ZN(n8122) );
  OAI222_X1 U8186 ( .A1(P2_U3151), .A2(n8122), .B1(n8559), .B2(n6535), .C1(
        n10152), .C2(n8557), .ZN(P2_U3283) );
  INV_X1 U8187 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9945) );
  INV_X1 U8188 ( .A(n6536), .ZN(n6538) );
  INV_X1 U8189 ( .A(n8822), .ZN(n9332) );
  OAI222_X1 U8190 ( .A1(n7620), .A2(n9945), .B1(n7569), .B2(n6538), .C1(
        P1_U3086), .C2(n9332), .ZN(P1_U3342) );
  INV_X1 U8191 ( .A(n9679), .ZN(n8120) );
  INV_X1 U8192 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6537) );
  OAI222_X1 U8193 ( .A1(n8120), .A2(P2_U3151), .B1(n8559), .B2(n6538), .C1(
        n6537), .C2(n8557), .ZN(P2_U3282) );
  INV_X1 U8194 ( .A(n6539), .ZN(n6552) );
  AOI22_X1 U8195 ( .A1(n9346), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6686), .ZN(n6540) );
  OAI21_X1 U8196 ( .B1(n6552), .B2(n7569), .A(n6540), .ZN(P1_U3341) );
  INV_X1 U8197 ( .A(n6569), .ZN(n6550) );
  INV_X1 U8198 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6549) );
  OAI21_X1 U8199 ( .B1(n6543), .B2(n6542), .A(n6541), .ZN(n6544) );
  NAND2_X1 U8200 ( .A1(n6544), .A2(n8709), .ZN(n6548) );
  NAND2_X1 U8201 ( .A1(n8739), .A2(n8859), .ZN(n6545) );
  NAND2_X1 U8202 ( .A1(n6546), .A2(n6545), .ZN(n6936) );
  INV_X1 U8203 ( .A(n9255), .ZN(n8660) );
  AOI22_X1 U8204 ( .A1(n6945), .A2(n5768), .B1(n6936), .B2(n8660), .ZN(n6547)
         );
  OAI211_X1 U8205 ( .C1(n6550), .C2(n6549), .A(n6548), .B(n6547), .ZN(P1_U3222) );
  INV_X1 U8206 ( .A(n9694), .ZN(n9703) );
  OAI222_X1 U8207 ( .A1(n9703), .A2(P2_U3151), .B1(n8559), .B2(n6552), .C1(
        n6551), .C2(n8557), .ZN(P2_U3281) );
  INV_X1 U8208 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U8209 ( .A1(n6553), .A2(n10149), .ZN(P2_U3261) );
  INV_X1 U8210 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n6554) );
  NOR2_X1 U8211 ( .A1(n6553), .A2(n6554), .ZN(P2_U3245) );
  INV_X1 U8212 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6555) );
  NOR2_X1 U8213 ( .A1(n6553), .A2(n6555), .ZN(P2_U3258) );
  INV_X1 U8214 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6556) );
  NOR2_X1 U8215 ( .A1(n6553), .A2(n6556), .ZN(P2_U3263) );
  INV_X1 U8216 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6557) );
  NOR2_X1 U8217 ( .A1(n6553), .A2(n6557), .ZN(P2_U3262) );
  INV_X1 U8218 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6558) );
  NOR2_X1 U8219 ( .A1(n6553), .A2(n6558), .ZN(P2_U3235) );
  INV_X1 U8220 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6559) );
  NOR2_X1 U8221 ( .A1(n6553), .A2(n6559), .ZN(P2_U3260) );
  INV_X1 U8222 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U8223 ( .A1(n6553), .A2(n10161), .ZN(P2_U3259) );
  INV_X1 U8224 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6560) );
  NOR2_X1 U8225 ( .A1(n6553), .A2(n6560), .ZN(P2_U3240) );
  INV_X1 U8226 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U8227 ( .A1(n6553), .A2(n10092), .ZN(P2_U3241) );
  INV_X1 U8228 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U8229 ( .A1(n6553), .A2(n6561), .ZN(P2_U3237) );
  INV_X1 U8230 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6562) );
  NOR2_X1 U8231 ( .A1(n6553), .A2(n6562), .ZN(P2_U3234) );
  INV_X1 U8232 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U8233 ( .A1(n6553), .A2(n6563), .ZN(P2_U3236) );
  INV_X1 U8234 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10177) );
  NOR2_X1 U8235 ( .A1(n6553), .A2(n10177), .ZN(P2_U3242) );
  INV_X1 U8236 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6564) );
  NOR2_X1 U8237 ( .A1(n6553), .A2(n6564), .ZN(P2_U3244) );
  INV_X1 U8238 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U8239 ( .A1(n6553), .A2(n9990), .ZN(P2_U3243) );
  INV_X1 U8240 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U8241 ( .A1(n6553), .A2(n10014), .ZN(P2_U3239) );
  INV_X1 U8242 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6565) );
  NOR2_X1 U8243 ( .A1(n6553), .A2(n6565), .ZN(P2_U3238) );
  XOR2_X1 U8244 ( .A(n6566), .B(n6567), .Z(n6571) );
  AOI22_X1 U8245 ( .A1(n8699), .A2(n6708), .B1(n8738), .B2(n8859), .ZN(n6885)
         );
  OAI22_X1 U8246 ( .A1(n6885), .A2(n9255), .B1(n9472), .B2(n8717), .ZN(n6568)
         );
  AOI21_X1 U8247 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6569), .A(n6568), .ZN(
        n6570) );
  OAI21_X1 U8248 ( .B1(n6571), .B2(n9260), .A(n6570), .ZN(P1_U3237) );
  NAND2_X1 U8249 ( .A1(n6900), .A2(P2_U3893), .ZN(n6572) );
  OAI21_X1 U8250 ( .B1(P2_U3893), .B2(n5176), .A(n6572), .ZN(P2_U3491) );
  INV_X1 U8251 ( .A(n6573), .ZN(n6575) );
  INV_X1 U8252 ( .A(n8824), .ZN(n9359) );
  INV_X1 U8253 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10171) );
  OAI222_X1 U8254 ( .A1(n7569), .A2(n6575), .B1(n9359), .B2(P1_U3086), .C1(
        n10171), .C2(n7620), .ZN(P1_U3340) );
  INV_X1 U8255 ( .A(n8141), .ZN(n9723) );
  INV_X1 U8256 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6574) );
  OAI222_X1 U8257 ( .A1(P2_U3151), .A2(n9723), .B1(n8559), .B2(n6575), .C1(
        n6574), .C2(n8557), .ZN(P2_U3280) );
  INV_X1 U8258 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U8259 ( .A1(n6900), .A2(n6609), .ZN(n7633) );
  NAND2_X1 U8260 ( .A1(n7627), .A2(n7633), .ZN(n7811) );
  OAI21_X1 U8261 ( .B1(n8355), .B2(n9819), .A(n7811), .ZN(n6576) );
  NAND2_X1 U8262 ( .A1(n9760), .A2(n9758), .ZN(n6675) );
  OAI211_X1 U8263 ( .C1(n9821), .C2(n6609), .A(n6576), .B(n6675), .ZN(n8432)
         );
  NAND2_X1 U8264 ( .A1(n8432), .A2(n9833), .ZN(n6577) );
  OAI21_X1 U8265 ( .B1(n6578), .B2(n9833), .A(n6577), .ZN(P2_U3390) );
  XOR2_X1 U8266 ( .A(n6579), .B(n6580), .Z(n6583) );
  INV_X1 U8267 ( .A(n8737), .ZN(n6832) );
  INV_X1 U8268 ( .A(n8739), .ZN(n6713) );
  OAI22_X1 U8269 ( .A1(n6832), .A2(n8697), .B1(n6713), .B2(n8927), .ZN(n6731)
         );
  AOI22_X1 U8270 ( .A1(n6731), .A2(n8660), .B1(n9478), .B2(n5768), .ZN(n6582)
         );
  MUX2_X1 U8271 ( .A(n9267), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6581) );
  OAI211_X1 U8272 ( .C1(n6583), .C2(n9260), .A(n6582), .B(n6581), .ZN(P1_U3218) );
  NAND2_X1 U8273 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  NAND2_X1 U8274 ( .A1(n6587), .A2(n6586), .ZN(n6591) );
  NAND2_X1 U8275 ( .A1(n6601), .A2(n6594), .ZN(n6589) );
  NAND4_X1 U8276 ( .A1(n6591), .A2(n6590), .A3(n6589), .A4(n6588), .ZN(n6592)
         );
  NAND2_X1 U8277 ( .A1(n6592), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6596) );
  NOR2_X1 U8278 ( .A1(n6674), .A2(n6593), .ZN(n7843) );
  NAND2_X1 U8279 ( .A1(n7843), .A2(n6594), .ZN(n6595) );
  NAND2_X1 U8280 ( .A1(n6596), .A2(n6595), .ZN(n6784) );
  INV_X1 U8281 ( .A(n6597), .ZN(n6598) );
  NOR2_X1 U8282 ( .A1(n6784), .A2(n6598), .ZN(n6639) );
  INV_X1 U8283 ( .A(n6599), .ZN(n6600) );
  NAND2_X1 U8284 ( .A1(n6600), .A2(n6604), .ZN(n6603) );
  NAND2_X1 U8285 ( .A1(n6607), .A2(n6601), .ZN(n6602) );
  NAND2_X1 U8286 ( .A1(n6604), .A2(n9832), .ZN(n6605) );
  INV_X1 U8287 ( .A(n8064), .ZN(n8081) );
  AND2_X1 U8288 ( .A1(n6607), .A2(n6606), .ZN(n6624) );
  INV_X1 U8289 ( .A(n6624), .ZN(n6608) );
  OAI22_X1 U8290 ( .A1(n8081), .A2(n6609), .B1(n5826), .B2(n8061), .ZN(n6610)
         );
  AOI21_X1 U8291 ( .B1(n7811), .B2(n4824), .A(n6610), .ZN(n6611) );
  OAI21_X1 U8292 ( .B1(n6639), .B2(n6872), .A(n6611), .ZN(P2_U3172) );
  NAND2_X1 U8293 ( .A1(n6612), .A2(n7784), .ZN(n6614) );
  XNOR2_X1 U8294 ( .A(n6628), .B(n9774), .ZN(n6618) );
  NOR2_X1 U8295 ( .A1(n6618), .A2(n9760), .ZN(n6629) );
  OAI21_X1 U8296 ( .B1(n6678), .B2(n7874), .A(n7627), .ZN(n6620) );
  NAND2_X1 U8297 ( .A1(n6621), .A2(n6620), .ZN(n6631) );
  OAI21_X1 U8298 ( .B1(n6621), .B2(n6620), .A(n6631), .ZN(n6622) );
  NAND2_X1 U8299 ( .A1(n6622), .A2(n4824), .ZN(n6627) );
  OAI22_X1 U8300 ( .A1(n8075), .A2(n4981), .B1(n8081), .B2(n9774), .ZN(n6625)
         );
  AOI21_X1 U8301 ( .B1(n8073), .B2(n4415), .A(n6625), .ZN(n6626) );
  OAI211_X1 U8302 ( .C1(n6639), .C2(n6897), .A(n6627), .B(n6626), .ZN(P2_U3162) );
  INV_X4 U8303 ( .A(n6628), .ZN(n7877) );
  XNOR2_X1 U8304 ( .A(n6777), .B(n4415), .ZN(n6633) );
  INV_X1 U8305 ( .A(n6629), .ZN(n6630) );
  NAND2_X1 U8306 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  NAND2_X1 U8307 ( .A1(n6632), .A2(n6633), .ZN(n6780) );
  OAI21_X1 U8308 ( .B1(n6633), .B2(n6632), .A(n6780), .ZN(n6634) );
  NAND2_X1 U8309 ( .A1(n6634), .A2(n4824), .ZN(n6637) );
  OAI22_X1 U8310 ( .A1(n8075), .A2(n5826), .B1(n9766), .B2(n8081), .ZN(n6635)
         );
  AOI21_X1 U8311 ( .B1(n8073), .B2(n9759), .A(n6635), .ZN(n6636) );
  OAI211_X1 U8312 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(P2_U3177) );
  MUX2_X1 U8313 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8151), .Z(n6738) );
  XNOR2_X1 U8314 ( .A(n6738), .B(n6747), .ZN(n6646) );
  MUX2_X1 U8315 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8145), .Z(n6643) );
  INV_X1 U8316 ( .A(n6643), .ZN(n6644) );
  MUX2_X1 U8317 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8145), .Z(n6640) );
  INV_X1 U8318 ( .A(n6640), .ZN(n6641) );
  XNOR2_X1 U8319 ( .A(n6640), .B(n6642), .ZN(n6799) );
  MUX2_X1 U8320 ( .A(n5827), .B(n5828), .S(n8145), .Z(n6868) );
  XNOR2_X1 U8321 ( .A(n6643), .B(n6662), .ZN(n6814) );
  NOR2_X1 U8322 ( .A1(n6645), .A2(n6646), .ZN(n6739) );
  AOI21_X1 U8323 ( .B1(n6646), .B2(n6645), .A(n6739), .ZN(n6673) );
  NAND2_X1 U8324 ( .A1(P2_U3893), .A2(n6192), .ZN(n9597) );
  INV_X1 U8325 ( .A(n6647), .ZN(n6649) );
  NOR2_X1 U8326 ( .A1(n8151), .A2(P2_U3151), .ZN(n8551) );
  AND2_X1 U8327 ( .A1(n6192), .A2(n8551), .ZN(n6648) );
  NAND2_X1 U8328 ( .A1(n6652), .A2(n6648), .ZN(n6651) );
  NAND2_X1 U8329 ( .A1(n4506), .A2(n6649), .ZN(n6650) );
  OAI22_X1 U8330 ( .A1(n9754), .A2(n6747), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6964), .ZN(n6671) );
  AND2_X1 U8331 ( .A1(n6652), .A2(n4506), .ZN(n6870) );
  INV_X1 U8332 ( .A(n10223), .ZN(n9607) );
  INV_X1 U8333 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U8334 ( .A1(n5821), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U8335 ( .A1(n6794), .A2(n6657), .ZN(n6656) );
  NAND2_X1 U8336 ( .A1(n4590), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6654) );
  OR2_X1 U8337 ( .A1(n6654), .A2(n5821), .ZN(n6655) );
  NAND2_X1 U8338 ( .A1(n6656), .A2(n6655), .ZN(n6789) );
  NAND2_X1 U8339 ( .A1(n6789), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U8340 ( .A1(n6658), .A2(n6657), .ZN(n6806) );
  NAND2_X1 U8341 ( .A1(n6809), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8342 ( .A1(n6805), .A2(n6659), .ZN(n6748) );
  INV_X1 U8343 ( .A(n6747), .ZN(n6741) );
  XOR2_X1 U8344 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6746), .Z(n6669) );
  AND2_X1 U8345 ( .A1(n4590), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8346 ( .A1(n5821), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6661) );
  INV_X1 U8347 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6790) );
  XNOR2_X1 U8348 ( .A(n6662), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8349 ( .A1(n6803), .A2(n6804), .ZN(n6802) );
  NAND2_X1 U8350 ( .A1(n6809), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8351 ( .A1(n6802), .A2(n6663), .ZN(n6664) );
  INV_X1 U8352 ( .A(n9584), .ZN(n6665) );
  AOI21_X1 U8353 ( .B1(n5854), .B2(n6666), .A(n6665), .ZN(n6668) );
  INV_X1 U8354 ( .A(n6870), .ZN(n6667) );
  OAI22_X1 U8355 ( .A1(n9607), .A2(n6669), .B1(n6668), .B2(n10220), .ZN(n6670)
         );
  AOI211_X1 U8356 ( .C1(n9740), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6671), .B(
        n6670), .ZN(n6672) );
  OAI21_X1 U8357 ( .B1(n6673), .B2(n9597), .A(n6672), .ZN(P2_U3185) );
  NAND3_X1 U8358 ( .A1(n7811), .A2(n6674), .A3(n9821), .ZN(n6676) );
  OAI211_X1 U8359 ( .C1(n6872), .C2(n8373), .A(n6676), .B(n6675), .ZN(n6677)
         );
  NAND2_X1 U8360 ( .A1(n6677), .A2(n8376), .ZN(n6680) );
  AOI22_X1 U8361 ( .A1(n8378), .A2(n6678), .B1(P2_REG2_REG_0__SCAN_IN), .B2(
        n9773), .ZN(n6679) );
  NAND2_X1 U8362 ( .A1(n6680), .A2(n6679), .ZN(P2_U3233) );
  INV_X1 U8363 ( .A(n6681), .ZN(n6683) );
  INV_X1 U8364 ( .A(n8826), .ZN(n9367) );
  INV_X1 U8365 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6682) );
  OAI222_X1 U8366 ( .A1(n7569), .A2(n6683), .B1(n9367), .B2(P1_U3086), .C1(
        n6682), .C2(n7620), .ZN(P1_U3339) );
  INV_X1 U8367 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6684) );
  INV_X1 U8368 ( .A(n8147), .ZN(n9738) );
  OAI222_X1 U8369 ( .A1(n8557), .A2(n6684), .B1(P2_U3151), .B2(n9738), .C1(
        n6683), .C2(n8559), .ZN(P2_U3279) );
  INV_X1 U8370 ( .A(n6685), .ZN(n6776) );
  AOI22_X1 U8371 ( .A1(n8813), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6686), .ZN(n6687) );
  OAI21_X1 U8372 ( .B1(n6776), .B2(n7569), .A(n6687), .ZN(P1_U3338) );
  INV_X1 U8373 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U8374 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6688) );
  AOI21_X1 U8375 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6688), .ZN(n9866) );
  NOR2_X1 U8376 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6689) );
  AOI21_X1 U8377 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6689), .ZN(n9869) );
  NOR2_X1 U8378 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n6690) );
  AOI21_X1 U8379 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n6690), .ZN(n9872) );
  NOR2_X1 U8380 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6691) );
  AOI21_X1 U8381 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6691), .ZN(n9875) );
  NOR2_X1 U8382 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6692) );
  AOI21_X1 U8383 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6692), .ZN(n9878) );
  NOR2_X1 U8384 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n6693) );
  AOI21_X1 U8385 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n6693), .ZN(n9881) );
  NOR2_X1 U8386 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6694) );
  AOI21_X1 U8387 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6694), .ZN(n9884) );
  NOR2_X1 U8388 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6695) );
  AOI21_X1 U8389 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6695), .ZN(n9887) );
  NOR2_X1 U8390 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .ZN(n6696) );
  AOI21_X1 U8391 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n6696), .ZN(n10233) );
  NOR2_X1 U8392 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .ZN(n6697) );
  AOI21_X1 U8393 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n6697), .ZN(n10239) );
  NOR2_X1 U8394 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .ZN(n6698) );
  AOI21_X1 U8395 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n6698), .ZN(n10236) );
  NOR2_X1 U8396 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6699) );
  AOI21_X1 U8397 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6699), .ZN(n10227) );
  NOR2_X1 U8398 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n6700) );
  AOI21_X1 U8399 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n6700), .ZN(n10230) );
  INV_X1 U8400 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9859) );
  INV_X1 U8401 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9858) );
  NOR2_X1 U8402 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  NOR2_X1 U8403 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9857), .ZN(n9853) );
  INV_X1 U8404 ( .A(n9853), .ZN(n9854) );
  INV_X1 U8405 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9856) );
  NAND3_X1 U8406 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U8407 ( .A1(n9856), .A2(n9855), .ZN(n9852) );
  NAND2_X1 U8408 ( .A1(n9854), .A2(n9852), .ZN(n10242) );
  NAND2_X1 U8409 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6701) );
  OAI21_X1 U8410 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6701), .ZN(n10241) );
  NOR2_X1 U8411 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  AOI21_X1 U8412 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10240), .ZN(n10245) );
  NAND2_X1 U8413 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6702) );
  OAI21_X1 U8414 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6702), .ZN(n10244) );
  NOR2_X1 U8415 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  AOI21_X1 U8416 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10243), .ZN(n10248) );
  NOR2_X1 U8417 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6703) );
  AOI21_X1 U8418 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n6703), .ZN(n10247) );
  NAND2_X1 U8419 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  OAI21_X1 U8420 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10246), .ZN(n10229) );
  NAND2_X1 U8421 ( .A1(n10230), .A2(n10229), .ZN(n10228) );
  OAI21_X1 U8422 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10228), .ZN(n10226) );
  NAND2_X1 U8423 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  OAI21_X1 U8424 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10225), .ZN(n10235) );
  NAND2_X1 U8425 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  OAI21_X1 U8426 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10234), .ZN(n10238) );
  NAND2_X1 U8427 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  OAI21_X1 U8428 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10237), .ZN(n10232) );
  NAND2_X1 U8429 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  OAI21_X1 U8430 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10231), .ZN(n9886) );
  NAND2_X1 U8431 ( .A1(n9887), .A2(n9886), .ZN(n9885) );
  OAI21_X1 U8432 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9885), .ZN(n9883) );
  NAND2_X1 U8433 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U8434 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9882), .ZN(n9880) );
  NAND2_X1 U8435 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  OAI21_X1 U8436 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9879), .ZN(n9877) );
  NAND2_X1 U8437 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  OAI21_X1 U8438 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9876), .ZN(n9874) );
  NAND2_X1 U8439 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  OAI21_X1 U8440 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9873), .ZN(n9871) );
  NAND2_X1 U8441 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  OAI21_X1 U8442 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9870), .ZN(n9868) );
  NAND2_X1 U8443 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  OAI21_X1 U8444 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9867), .ZN(n9865) );
  NAND2_X1 U8445 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  OAI21_X1 U8446 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9864), .ZN(n9862) );
  NOR2_X1 U8447 ( .A1(n9861), .A2(n9862), .ZN(n6704) );
  NAND2_X1 U8448 ( .A1(n9861), .A2(n9862), .ZN(n9860) );
  OAI21_X1 U8449 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6704), .A(n9860), .ZN(
        n6707) );
  XNOR2_X1 U8450 ( .A(n6705), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6706) );
  XNOR2_X1 U8451 ( .A(n6707), .B(n6706), .ZN(ADD_1068_U4) );
  NAND2_X1 U8452 ( .A1(n8659), .A2(n9478), .ZN(n6837) );
  NAND2_X1 U8453 ( .A1(n8738), .A2(n6829), .ZN(n7513) );
  NAND2_X1 U8454 ( .A1(n6837), .A2(n7513), .ZN(n7473) );
  INV_X1 U8455 ( .A(n6945), .ZN(n9464) );
  NAND2_X1 U8456 ( .A1(n6708), .A2(n9464), .ZN(n7512) );
  NAND2_X1 U8457 ( .A1(n6710), .A2(n6945), .ZN(n6727) );
  NAND2_X1 U8458 ( .A1(n6709), .A2(n9446), .ZN(n6938) );
  NAND2_X1 U8459 ( .A1(n6725), .A2(n6938), .ZN(n6712) );
  NAND2_X1 U8460 ( .A1(n6710), .A2(n9464), .ZN(n6711) );
  NAND2_X1 U8461 ( .A1(n6712), .A2(n6711), .ZN(n6882) );
  NAND2_X1 U8462 ( .A1(n6882), .A2(n6883), .ZN(n6715) );
  NAND2_X1 U8463 ( .A1(n6713), .A2(n9472), .ZN(n6714) );
  NAND2_X1 U8464 ( .A1(n6715), .A2(n6714), .ZN(n6828) );
  XOR2_X1 U8465 ( .A(n7473), .B(n6828), .Z(n9481) );
  AND2_X1 U8466 ( .A1(n6716), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8467 ( .A1(n6718), .A2(n6717), .ZN(n9124) );
  INV_X1 U8468 ( .A(n9125), .ZN(n9202) );
  NAND2_X1 U8469 ( .A1(n9202), .A2(n9120), .ZN(n6719) );
  OR2_X1 U8470 ( .A1(n9124), .A2(n6719), .ZN(n6720) );
  AND2_X1 U8471 ( .A1(n7558), .A2(n6721), .ZN(n6724) );
  OAI21_X1 U8472 ( .B1(n6722), .B2(n7558), .A(n6723), .ZN(n9444) );
  OR2_X1 U8473 ( .A1(n6724), .A2(n9444), .ZN(n9415) );
  NAND2_X1 U8474 ( .A1(n9415), .A2(n6941), .ZN(n9109) );
  NAND2_X1 U8475 ( .A1(n6935), .A2(n6727), .ZN(n6884) );
  NOR2_X1 U8476 ( .A1(n8739), .A2(n9472), .ZN(n6728) );
  NAND2_X1 U8477 ( .A1(n8739), .A2(n9472), .ZN(n7514) );
  OAI21_X1 U8478 ( .B1(n6884), .B2(n6728), .A(n7514), .ZN(n6838) );
  XNOR2_X1 U8479 ( .A(n7473), .B(n6838), .ZN(n6732) );
  NAND2_X1 U8480 ( .A1(n5760), .A2(n7508), .ZN(n6730) );
  OR2_X1 U8481 ( .A1(n5759), .A2(n5160), .ZN(n6729) );
  AOI21_X1 U8482 ( .B1(n6732), .B2(n9459), .A(n6731), .ZN(n9480) );
  MUX2_X1 U8483 ( .A(n6733), .B(n9480), .S(n9452), .Z(n6737) );
  INV_X1 U8484 ( .A(n6842), .ZN(n9438) );
  AOI211_X1 U8485 ( .C1(n9478), .C2(n6888), .A(n9101), .B(n9438), .ZN(n9477)
         );
  OAI22_X1 U8486 ( .A1(n9104), .A2(n6829), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n7121), .ZN(n6735) );
  AOI21_X1 U8487 ( .B1(n9477), .B2(n9440), .A(n6735), .ZN(n6736) );
  OAI211_X1 U8488 ( .C1(n9481), .C2(n9086), .A(n6737), .B(n6736), .ZN(P1_U3290) );
  MUX2_X1 U8489 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8151), .Z(n6743) );
  INV_X1 U8490 ( .A(n6738), .ZN(n6740) );
  MUX2_X1 U8491 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8151), .Z(n6742) );
  INV_X1 U8492 ( .A(n9591), .ZN(n6752) );
  XNOR2_X1 U8493 ( .A(n6742), .B(n6752), .ZN(n9577) );
  AOI22_X1 U8494 ( .A1(n9576), .A2(n9577), .B1(n6742), .B2(n9591), .ZN(n9598)
         );
  XNOR2_X1 U8495 ( .A(n6743), .B(n9600), .ZN(n9599) );
  NOR2_X1 U8496 ( .A1(n9598), .A2(n9599), .ZN(n9596) );
  MUX2_X1 U8497 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8151), .Z(n6850) );
  XOR2_X1 U8498 ( .A(n6860), .B(n6850), .Z(n6744) );
  NAND2_X1 U8499 ( .A1(n6745), .A2(n6744), .ZN(n6849) );
  OAI21_X1 U8500 ( .B1(n6745), .B2(n6744), .A(n6849), .ZN(n6773) );
  INV_X1 U8501 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9842) );
  MUX2_X1 U8502 ( .A(n9842), .B(P2_REG1_REG_6__SCAN_IN), .S(n6860), .Z(n6755)
         );
  NAND2_X1 U8503 ( .A1(n6746), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U8504 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND2_X1 U8505 ( .A1(n6750), .A2(n6749), .ZN(n9579) );
  MUX2_X1 U8506 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6751), .S(n9591), .Z(n9580)
         );
  NAND2_X1 U8507 ( .A1(n9579), .A2(n9580), .ZN(n9578) );
  AOI22_X1 U8508 ( .A1(n9601), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n9600), .B2(
        n6753), .ZN(n6754) );
  NOR2_X1 U8509 ( .A1(n6754), .A2(n6755), .ZN(n6859) );
  AOI21_X1 U8510 ( .B1(n6755), .B2(n6754), .A(n6859), .ZN(n6766) );
  INV_X1 U8511 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U8512 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7000), .S(n9591), .Z(n9581)
         );
  NAND2_X1 U8513 ( .A1(n6756), .A2(n9581), .ZN(n9586) );
  NAND2_X1 U8514 ( .A1(n9591), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6757) );
  INV_X1 U8515 ( .A(n6760), .ZN(n6759) );
  XNOR2_X1 U8516 ( .A(n6860), .B(n6758), .ZN(n6761) );
  NOR2_X1 U8517 ( .A1(n6759), .A2(n6761), .ZN(n6764) );
  NAND2_X1 U8518 ( .A1(n9602), .A2(n6760), .ZN(n6762) );
  NAND2_X1 U8519 ( .A1(n6762), .A2(n6761), .ZN(n6852) );
  INV_X1 U8520 ( .A(n6852), .ZN(n6763) );
  AOI21_X1 U8521 ( .B1(n6764), .B2(n9602), .A(n6763), .ZN(n6765) );
  OAI22_X1 U8522 ( .A1(n9607), .A2(n6766), .B1(n6765), .B2(n10220), .ZN(n6772)
         );
  INV_X1 U8523 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6770) );
  INV_X1 U8524 ( .A(n6860), .ZN(n6768) );
  INV_X1 U8525 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6767) );
  NOR2_X1 U8526 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6767), .ZN(n7069) );
  AOI21_X1 U8527 ( .B1(n10209), .B2(n6768), .A(n7069), .ZN(n6769) );
  OAI21_X1 U8528 ( .B1(n10217), .B2(n6770), .A(n6769), .ZN(n6771) );
  AOI211_X1 U8529 ( .C1(n6773), .C2(n10207), .A(n6772), .B(n6771), .ZN(n6774)
         );
  INV_X1 U8530 ( .A(n6774), .ZN(P2_U3188) );
  OAI222_X1 U8531 ( .A1(n9753), .A2(P2_U3151), .B1(n8559), .B2(n6776), .C1(
        n6775), .C2(n8557), .ZN(P2_U3278) );
  XNOR2_X1 U8532 ( .A(n7877), .B(n6965), .ZN(n6907) );
  XNOR2_X1 U8533 ( .A(n6907), .B(n9759), .ZN(n6782) );
  NAND2_X1 U8534 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  AOI211_X1 U8535 ( .C1(n6782), .C2(n6781), .A(n8067), .B(n6909), .ZN(n6788)
         );
  INV_X1 U8536 ( .A(n8093), .ZN(n7025) );
  OR2_X1 U8537 ( .A1(n6783), .A2(P2_U3151), .ZN(n7847) );
  INV_X1 U8538 ( .A(n7847), .ZN(n7275) );
  MUX2_X1 U8539 ( .A(n8053), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6786) );
  AOI22_X1 U8540 ( .A1(n8058), .A2(n4415), .B1(n6965), .B2(n8064), .ZN(n6785)
         );
  OAI211_X1 U8541 ( .C1(n7025), .C2(n8061), .A(n6786), .B(n6785), .ZN(n6787)
         );
  OR2_X1 U8542 ( .A1(n6788), .A2(n6787), .ZN(P2_U3158) );
  XNOR2_X1 U8543 ( .A(n6789), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8544 ( .A1(n6791), .A2(n6790), .ZN(n6792) );
  AOI21_X1 U8545 ( .B1(n6793), .B2(n6792), .A(n10220), .ZN(n6796) );
  OAI22_X1 U8546 ( .A1(n9754), .A2(n6794), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6897), .ZN(n6795) );
  AOI211_X1 U8547 ( .C1(n10223), .C2(n6797), .A(n6796), .B(n6795), .ZN(n6801)
         );
  OAI211_X1 U8548 ( .C1(n6799), .C2(n6867), .A(n6798), .B(n10207), .ZN(n6800)
         );
  OAI211_X1 U8549 ( .C1(n9856), .C2(n10217), .A(n6801), .B(n6800), .ZN(
        P2_U3183) );
  INV_X1 U8550 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6818) );
  INV_X1 U8551 ( .A(n10220), .ZN(n9749) );
  OAI21_X1 U8552 ( .B1(n6804), .B2(n6803), .A(n6802), .ZN(n6812) );
  OAI21_X1 U8553 ( .B1(n6807), .B2(n6806), .A(n6805), .ZN(n6808) );
  AND2_X1 U8554 ( .A1(n10223), .A2(n6808), .ZN(n6811) );
  OAI22_X1 U8555 ( .A1(n9754), .A2(n6809), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6638), .ZN(n6810) );
  AOI211_X1 U8556 ( .C1(n9749), .C2(n6812), .A(n6811), .B(n6810), .ZN(n6817)
         );
  OAI211_X1 U8557 ( .C1(n6815), .C2(n6814), .A(n6813), .B(n10207), .ZN(n6816)
         );
  OAI211_X1 U8558 ( .C1(n10217), .C2(n6818), .A(n6817), .B(n6816), .ZN(
        P2_U3184) );
  NAND2_X1 U8559 ( .A1(n6820), .A2(n6819), .ZN(n6822) );
  XNOR2_X1 U8560 ( .A(n6822), .B(n6821), .ZN(n6827) );
  NAND2_X1 U8561 ( .A1(n8737), .A2(n8699), .ZN(n6824) );
  NAND2_X1 U8562 ( .A1(n8735), .A2(n8859), .ZN(n6823) );
  NAND2_X1 U8563 ( .A1(n6824), .A2(n6823), .ZN(n6921) );
  AOI22_X1 U8564 ( .A1(n6921), .A2(n8660), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6826) );
  AOI22_X1 U8565 ( .A1(n5768), .A2(n6928), .B1(n6927), .B2(n8713), .ZN(n6825)
         );
  OAI211_X1 U8566 ( .C1(n6827), .C2(n9260), .A(n6826), .B(n6825), .ZN(P1_U3227) );
  NAND2_X1 U8567 ( .A1(n6828), .A2(n7473), .ZN(n6831) );
  NAND2_X1 U8568 ( .A1(n8659), .A2(n6829), .ZN(n6830) );
  NAND2_X1 U8569 ( .A1(n6831), .A2(n6830), .ZN(n9433) );
  NAND2_X1 U8570 ( .A1(n6832), .A2(n9432), .ZN(n7344) );
  INV_X1 U8571 ( .A(n9432), .ZN(n9484) );
  NAND2_X1 U8572 ( .A1(n7344), .A2(n7516), .ZN(n9434) );
  NAND2_X1 U8573 ( .A1(n9433), .A2(n9434), .ZN(n6834) );
  NAND2_X1 U8574 ( .A1(n6832), .A2(n9484), .ZN(n6833) );
  NAND2_X1 U8575 ( .A1(n6834), .A2(n6833), .ZN(n6924) );
  INV_X1 U8576 ( .A(n8736), .ZN(n8658) );
  NAND2_X1 U8577 ( .A1(n8658), .A2(n6928), .ZN(n7345) );
  INV_X1 U8578 ( .A(n6928), .ZN(n9492) );
  NAND2_X1 U8579 ( .A1(n8736), .A2(n9492), .ZN(n7347) );
  NAND2_X1 U8580 ( .A1(n6924), .A2(n7479), .ZN(n6836) );
  NAND2_X1 U8581 ( .A1(n8658), .A2(n9492), .ZN(n6835) );
  NAND2_X1 U8582 ( .A1(n6836), .A2(n6835), .ZN(n7045) );
  INV_X1 U8583 ( .A(n8735), .ZN(n7047) );
  NAND2_X1 U8584 ( .A1(n7047), .A2(n9497), .ZN(n7351) );
  INV_X1 U8585 ( .A(n9497), .ZN(n7046) );
  NAND2_X1 U8586 ( .A1(n8735), .A2(n7046), .ZN(n7348) );
  XOR2_X1 U8587 ( .A(n7045), .B(n7480), .Z(n9500) );
  NAND2_X1 U8588 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  NAND2_X1 U8589 ( .A1(n6839), .A2(n7513), .ZN(n9427) );
  NAND2_X1 U8590 ( .A1(n9427), .A2(n7344), .ZN(n6840) );
  NAND2_X1 U8591 ( .A1(n6840), .A2(n7516), .ZN(n6919) );
  INV_X1 U8592 ( .A(n7347), .ZN(n7517) );
  XOR2_X1 U8593 ( .A(n7480), .B(n7034), .Z(n6841) );
  INV_X1 U8594 ( .A(n8734), .ZN(n7050) );
  OAI22_X1 U8595 ( .A1(n8658), .A2(n8927), .B1(n7050), .B2(n8697), .ZN(n6876)
         );
  AOI21_X1 U8596 ( .B1(n6841), .B2(n9459), .A(n6876), .ZN(n9499) );
  MUX2_X1 U8597 ( .A(n6432), .B(n9499), .S(n9452), .Z(n6848) );
  NOR2_X2 U8598 ( .A1(n6842), .A2(n9432), .ZN(n9435) );
  AND2_X1 U8599 ( .A1(n9435), .A2(n9492), .ZN(n6925) );
  INV_X1 U8600 ( .A(n6925), .ZN(n6844) );
  NAND2_X1 U8601 ( .A1(n6925), .A2(n7046), .ZN(n7119) );
  INV_X1 U8602 ( .A(n7119), .ZN(n6843) );
  AOI211_X1 U8603 ( .C1(n9497), .C2(n6844), .A(n9101), .B(n6843), .ZN(n9496)
         );
  INV_X1 U8604 ( .A(n6845), .ZN(n6878) );
  OAI22_X1 U8605 ( .A1(n9104), .A2(n7046), .B1(n7121), .B2(n6878), .ZN(n6846)
         );
  AOI21_X1 U8606 ( .B1(n9496), .B2(n9440), .A(n6846), .ZN(n6847) );
  OAI211_X1 U8607 ( .C1(n9500), .C2(n9086), .A(n6848), .B(n6847), .ZN(P1_U3287) );
  MUX2_X1 U8608 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8151), .Z(n6969) );
  XNOR2_X1 U8609 ( .A(n6969), .B(n6975), .ZN(n6971) );
  OAI21_X1 U8610 ( .B1(n6850), .B2(n6860), .A(n6849), .ZN(n6972) );
  XOR2_X1 U8611 ( .A(n6971), .B(n6972), .Z(n6866) );
  NAND2_X1 U8612 ( .A1(n6860), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U8613 ( .A1(n6852), .A2(n6851), .ZN(n6854) );
  NAND2_X1 U8614 ( .A1(n6855), .A2(n5914), .ZN(n6856) );
  NAND2_X1 U8615 ( .A1(n6985), .A2(n6856), .ZN(n6864) );
  INV_X1 U8616 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6858) );
  AND2_X1 U8617 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7201) );
  AOI21_X1 U8618 ( .B1(n10209), .B2(n6975), .A(n7201), .ZN(n6857) );
  OAI21_X1 U8619 ( .B1(n10217), .B2(n6858), .A(n6857), .ZN(n6863) );
  XNOR2_X1 U8620 ( .A(n6977), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n6861) );
  NOR2_X1 U8621 ( .A1(n6861), .A2(n9607), .ZN(n6862) );
  AOI211_X1 U8622 ( .C1(n9749), .C2(n6864), .A(n6863), .B(n6862), .ZN(n6865)
         );
  OAI21_X1 U8623 ( .B1(n6866), .B2(n9597), .A(n6865), .ZN(P2_U3189) );
  OAI21_X1 U8624 ( .B1(n6870), .B2(n10207), .A(n6869), .ZN(n6871) );
  OAI21_X1 U8625 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6872), .A(n6871), .ZN(n6873) );
  OAI21_X1 U8626 ( .B1(n10217), .B2(n9858), .A(n4439), .ZN(P2_U3182) );
  XOR2_X1 U8627 ( .A(n6874), .B(n6875), .Z(n6881) );
  AOI22_X1 U8628 ( .A1(n6876), .A2(n8660), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6877) );
  OAI21_X1 U8629 ( .B1(n6878), .B2(n9267), .A(n6877), .ZN(n6879) );
  AOI21_X1 U8630 ( .B1(n9497), .B2(n5768), .A(n6879), .ZN(n6880) );
  OAI21_X1 U8631 ( .B1(n6881), .B2(n9260), .A(n6880), .ZN(P1_U3239) );
  INV_X1 U8632 ( .A(n6883), .ZN(n7475) );
  XNOR2_X1 U8633 ( .A(n6882), .B(n7475), .ZN(n9470) );
  XNOR2_X1 U8634 ( .A(n6884), .B(n6883), .ZN(n6886) );
  OAI21_X1 U8635 ( .B1(n6886), .B2(n9399), .A(n6885), .ZN(n9473) );
  NAND2_X1 U8636 ( .A1(n9473), .A2(n9452), .ZN(n6893) );
  INV_X1 U8637 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6887) );
  OAI22_X1 U8638 ( .A1(n9452), .A2(n9976), .B1(n6887), .B2(n7121), .ZN(n6890)
         );
  INV_X1 U8639 ( .A(n9440), .ZN(n8871) );
  OAI211_X1 U8640 ( .C1(n6943), .C2(n9472), .A(n6888), .B(n9436), .ZN(n9471)
         );
  NOR2_X1 U8641 ( .A1(n8871), .A2(n9471), .ZN(n6889) );
  AOI211_X1 U8642 ( .C1(n9431), .C2(n6891), .A(n6890), .B(n6889), .ZN(n6892)
         );
  OAI211_X1 U8643 ( .C1(n9470), .C2(n9086), .A(n6893), .B(n6892), .ZN(P1_U3291) );
  NAND2_X1 U8644 ( .A1(n8376), .A2(n6894), .ZN(n8186) );
  INV_X1 U8645 ( .A(n8186), .ZN(n9770) );
  NAND2_X1 U8646 ( .A1(n6239), .A2(n7627), .ZN(n6895) );
  NAND2_X1 U8647 ( .A1(n6896), .A2(n6895), .ZN(n9777) );
  OAI22_X1 U8648 ( .A1(n8180), .A2(n9774), .B1(n6897), .B2(n8373), .ZN(n6905)
         );
  INV_X1 U8649 ( .A(n6898), .ZN(n6899) );
  XNOR2_X1 U8650 ( .A(n6239), .B(n6899), .ZN(n6903) );
  NAND2_X1 U8651 ( .A1(n9777), .A2(n9765), .ZN(n6902) );
  INV_X1 U8652 ( .A(n8352), .ZN(n8372) );
  AOI22_X1 U8653 ( .A1(n8352), .A2(n6900), .B1(n4415), .B2(n9758), .ZN(n6901)
         );
  OAI211_X1 U8654 ( .C1(n9762), .C2(n6903), .A(n6902), .B(n6901), .ZN(n9775)
         );
  MUX2_X1 U8655 ( .A(n9775), .B(P2_REG2_REG_1__SCAN_IN), .S(n9773), .Z(n6904)
         );
  AOI211_X1 U8656 ( .C1(n9770), .C2(n9777), .A(n6905), .B(n6904), .ZN(n6906)
         );
  INV_X1 U8657 ( .A(n6906), .ZN(P2_U3232) );
  NOR2_X2 U8658 ( .A1(n6909), .A2(n6908), .ZN(n6913) );
  XNOR2_X1 U8659 ( .A(n7877), .B(n6910), .ZN(n6911) );
  NOR2_X1 U8660 ( .A1(n6911), .A2(n8093), .ZN(n7018) );
  AOI21_X1 U8661 ( .B1(n6911), .B2(n8093), .A(n7018), .ZN(n6912) );
  OAI21_X1 U8662 ( .B1(n6913), .B2(n6912), .A(n7021), .ZN(n6914) );
  NAND2_X1 U8663 ( .A1(n6914), .A2(n4824), .ZN(n6918) );
  NAND2_X1 U8664 ( .A1(n8058), .A2(n9759), .ZN(n6915) );
  NAND2_X1 U8665 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9589) );
  OAI211_X1 U8666 ( .C1(n9787), .C2(n8081), .A(n6915), .B(n9589), .ZN(n6916)
         );
  AOI21_X1 U8667 ( .B1(n8073), .B2(n8092), .A(n6916), .ZN(n6917) );
  OAI211_X1 U8668 ( .C1(n7001), .C2(n8053), .A(n6918), .B(n6917), .ZN(P2_U3170) );
  XNOR2_X1 U8669 ( .A(n6919), .B(n7479), .ZN(n6920) );
  NAND2_X1 U8670 ( .A1(n6920), .A2(n9459), .ZN(n6923) );
  INV_X1 U8671 ( .A(n6921), .ZN(n6922) );
  NAND2_X1 U8672 ( .A1(n6923), .A2(n6922), .ZN(n9495) );
  INV_X1 U8673 ( .A(n9495), .ZN(n6933) );
  XNOR2_X1 U8674 ( .A(n6924), .B(n7479), .ZN(n9490) );
  INV_X1 U8675 ( .A(n9086), .ZN(n9441) );
  OAI21_X1 U8676 ( .B1(n9435), .B2(n9492), .A(n9436), .ZN(n6926) );
  OR2_X1 U8677 ( .A1(n6926), .A2(n6925), .ZN(n9491) );
  INV_X2 U8678 ( .A(n7121), .ZN(n9447) );
  AOI22_X1 U8679 ( .A1(n9455), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6927), .B2(
        n9447), .ZN(n6930) );
  NAND2_X1 U8680 ( .A1(n9431), .A2(n6928), .ZN(n6929) );
  OAI211_X1 U8681 ( .C1(n9491), .C2(n8871), .A(n6930), .B(n6929), .ZN(n6931)
         );
  AOI21_X1 U8682 ( .B1(n9490), .B2(n9441), .A(n6931), .ZN(n6932) );
  OAI21_X1 U8683 ( .B1(n6933), .B2(n9455), .A(n6932), .ZN(P1_U3288) );
  NAND2_X1 U8684 ( .A1(n6935), .A2(n6934), .ZN(n6937) );
  AOI21_X1 U8685 ( .B1(n6937), .B2(n9459), .A(n6936), .ZN(n6940) );
  XNOR2_X1 U8686 ( .A(n6725), .B(n6938), .ZN(n9466) );
  INV_X1 U8687 ( .A(n9415), .ZN(n9513) );
  NAND2_X1 U8688 ( .A1(n9466), .A2(n9513), .ZN(n6939) );
  AND2_X1 U8689 ( .A1(n6940), .A2(n6939), .ZN(n9468) );
  NOR2_X1 U8690 ( .A1(n9455), .A2(n6941), .ZN(n9424) );
  NAND2_X1 U8691 ( .A1(n6945), .A2(n9446), .ZN(n6942) );
  NAND2_X1 U8692 ( .A1(n6942), .A2(n9436), .ZN(n6944) );
  OR2_X1 U8693 ( .A1(n6944), .A2(n6943), .ZN(n9463) );
  AOI22_X1 U8694 ( .A1(n9455), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9447), .ZN(n6947) );
  NAND2_X1 U8695 ( .A1(n9431), .A2(n6945), .ZN(n6946) );
  OAI211_X1 U8696 ( .C1(n8871), .C2(n9463), .A(n6947), .B(n6946), .ZN(n6948)
         );
  AOI21_X1 U8697 ( .B1(n9466), .B2(n9424), .A(n6948), .ZN(n6949) );
  OAI21_X1 U8698 ( .B1(n9468), .B2(n9455), .A(n6949), .ZN(P1_U3292) );
  INV_X1 U8699 ( .A(n6950), .ZN(n6996) );
  INV_X1 U8700 ( .A(n10211), .ZN(n8155) );
  OAI222_X1 U8701 ( .A1(n8557), .A2(n6951), .B1(n8559), .B2(n6996), .C1(
        P2_U3151), .C2(n8155), .ZN(P2_U3277) );
  XNOR2_X1 U8702 ( .A(n6954), .B(n6953), .ZN(n6955) );
  XNOR2_X1 U8703 ( .A(n6952), .B(n6955), .ZN(n6960) );
  INV_X1 U8704 ( .A(n9506), .ZN(n7123) );
  NOR2_X1 U8705 ( .A1(n8717), .A2(n7123), .ZN(n6958) );
  AOI22_X1 U8706 ( .A1(n8699), .A2(n8735), .B1(n8733), .B2(n8859), .ZN(n7115)
         );
  OAI22_X1 U8707 ( .A1(n7115), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6956), .ZN(n6957) );
  AOI211_X1 U8708 ( .C1(n8713), .C2(n7120), .A(n6958), .B(n6957), .ZN(n6959)
         );
  OAI21_X1 U8709 ( .B1(n6960), .B2(n9260), .A(n6959), .ZN(P1_U3213) );
  XOR2_X1 U8710 ( .A(n6961), .B(n7814), .Z(n6962) );
  AOI222_X1 U8711 ( .A1(n8355), .A2(n6962), .B1(n4415), .B2(n8352), .C1(n8093), 
        .C2(n9758), .ZN(n9782) );
  XNOR2_X1 U8712 ( .A(n6963), .B(n7814), .ZN(n9785) );
  AOI22_X1 U8713 ( .A1(n8378), .A2(n6965), .B1(n9768), .B2(n6964), .ZN(n6966)
         );
  OAI21_X1 U8714 ( .B1(n5854), .B2(n8376), .A(n6966), .ZN(n6967) );
  AOI21_X1 U8715 ( .B1(n9785), .B2(n8361), .A(n6967), .ZN(n6968) );
  OAI21_X1 U8716 ( .B1(n9782), .B2(n9773), .A(n6968), .ZN(P2_U3230) );
  MUX2_X1 U8717 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8151), .Z(n8131) );
  XOR2_X1 U8718 ( .A(n8108), .B(n8131), .Z(n8132) );
  INV_X1 U8719 ( .A(n6969), .ZN(n6970) );
  XOR2_X1 U8720 ( .A(n8132), .B(n8133), .Z(n6995) );
  MUX2_X1 U8721 ( .A(n6973), .B(P2_REG1_REG_8__SCAN_IN), .S(n8108), .Z(n6979)
         );
  INV_X1 U8722 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6976) );
  OAI21_X1 U8723 ( .B1(n6979), .B2(n6978), .A(n8107), .ZN(n6993) );
  INV_X1 U8724 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8725 ( .A(n6980), .B(P2_REG2_REG_8__SCAN_IN), .S(n8108), .Z(n6982)
         );
  NAND2_X1 U8726 ( .A1(n6981), .A2(n6982), .ZN(n8094) );
  INV_X1 U8727 ( .A(n6982), .ZN(n6984) );
  NAND3_X1 U8728 ( .A1(n6985), .A2(n6984), .A3(n6983), .ZN(n6986) );
  AND2_X1 U8729 ( .A1(n8094), .A2(n6986), .ZN(n6987) );
  NOR2_X1 U8730 ( .A1(n10220), .A2(n6987), .ZN(n6992) );
  INV_X1 U8731 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6990) );
  INV_X1 U8732 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6988) );
  NOR2_X1 U8733 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6988), .ZN(n7930) );
  AOI21_X1 U8734 ( .B1(n10209), .B2(n8108), .A(n7930), .ZN(n6989) );
  OAI21_X1 U8735 ( .B1(n10217), .B2(n6990), .A(n6989), .ZN(n6991) );
  AOI211_X1 U8736 ( .C1(n6993), .C2(n10223), .A(n6992), .B(n6991), .ZN(n6994)
         );
  OAI21_X1 U8737 ( .B1(n6995), .B2(n9597), .A(n6994), .ZN(P2_U3190) );
  INV_X1 U8738 ( .A(n8843), .ZN(n9388) );
  OAI222_X1 U8739 ( .A1(n7620), .A2(n10098), .B1(n9388), .B2(P1_U3086), .C1(
        n7569), .C2(n6996), .ZN(P1_U3337) );
  XNOR2_X1 U8740 ( .A(n7006), .B(n7810), .ZN(n6998) );
  AOI222_X1 U8741 ( .A1(n8355), .A2(n6998), .B1(n8092), .B2(n9758), .C1(n9759), 
        .C2(n8352), .ZN(n9786) );
  XNOR2_X1 U8742 ( .A(n6999), .B(n7810), .ZN(n9789) );
  NOR2_X1 U8743 ( .A1(n8376), .A2(n7000), .ZN(n7003) );
  OAI22_X1 U8744 ( .A1(n8180), .A2(n9787), .B1(n7001), .B2(n8373), .ZN(n7002)
         );
  AOI211_X1 U8745 ( .C1(n9789), .C2(n8361), .A(n7003), .B(n7002), .ZN(n7004)
         );
  OAI21_X1 U8746 ( .B1(n9786), .B2(n9773), .A(n7004), .ZN(P2_U3229) );
  OR2_X1 U8747 ( .A1(n7006), .A2(n7005), .ZN(n7008) );
  NAND2_X1 U8748 ( .A1(n7008), .A2(n7007), .ZN(n7009) );
  XNOR2_X1 U8749 ( .A(n7023), .B(n8092), .ZN(n7813) );
  XNOR2_X1 U8750 ( .A(n7009), .B(n7813), .ZN(n7013) );
  XNOR2_X1 U8751 ( .A(n7010), .B(n7813), .ZN(n9793) );
  NAND2_X1 U8752 ( .A1(n9793), .A2(n9765), .ZN(n7012) );
  AOI22_X1 U8753 ( .A1(n8352), .A2(n8093), .B1(n8091), .B2(n9758), .ZN(n7011)
         );
  OAI211_X1 U8754 ( .C1(n9762), .C2(n7013), .A(n7012), .B(n7011), .ZN(n9791)
         );
  INV_X1 U8755 ( .A(n9791), .ZN(n7017) );
  NOR2_X1 U8756 ( .A1(n8376), .A2(n5880), .ZN(n7015) );
  OAI22_X1 U8757 ( .A1(n8180), .A2(n9790), .B1(n7029), .B2(n8373), .ZN(n7014)
         );
  AOI211_X1 U8758 ( .C1(n9793), .C2(n9770), .A(n7015), .B(n7014), .ZN(n7016)
         );
  OAI21_X1 U8759 ( .B1(n7017), .B2(n9773), .A(n7016), .ZN(P2_U3228) );
  INV_X1 U8760 ( .A(n7018), .ZN(n7019) );
  XNOR2_X1 U8761 ( .A(n7877), .B(n7023), .ZN(n7062) );
  XNOR2_X1 U8762 ( .A(n7062), .B(n8092), .ZN(n7020) );
  AND3_X1 U8763 ( .A1(n7021), .A2(n7020), .A3(n7019), .ZN(n7022) );
  OAI21_X1 U8764 ( .B1(n7063), .B2(n7022), .A(n4824), .ZN(n7028) );
  AND2_X1 U8765 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9610) );
  AOI21_X1 U8766 ( .B1(n8064), .B2(n7023), .A(n9610), .ZN(n7024) );
  OAI21_X1 U8767 ( .B1(n8075), .B2(n7025), .A(n7024), .ZN(n7026) );
  AOI21_X1 U8768 ( .B1(n8073), .B2(n8091), .A(n7026), .ZN(n7027) );
  OAI211_X1 U8769 ( .C1(n7029), .C2(n8053), .A(n7028), .B(n7027), .ZN(P2_U3167) );
  INV_X1 U8770 ( .A(n7030), .ZN(n7031) );
  OAI222_X1 U8771 ( .A1(P2_U3151), .A2(n8164), .B1(n8559), .B2(n7031), .C1(
        n10081), .C2(n8557), .ZN(P2_U3276) );
  OAI222_X1 U8772 ( .A1(n7620), .A2(n7032), .B1(n7569), .B2(n7031), .C1(
        P1_U3086), .C2(n5549), .ZN(P1_U3336) );
  INV_X1 U8773 ( .A(n7351), .ZN(n7033) );
  INV_X1 U8774 ( .A(n8732), .ZN(n7035) );
  NAND2_X1 U8775 ( .A1(n8733), .A2(n9515), .ZN(n7340) );
  INV_X1 U8776 ( .A(n7038), .ZN(n7353) );
  INV_X1 U8777 ( .A(n8733), .ZN(n7052) );
  NAND2_X1 U8778 ( .A1(n7052), .A2(n9420), .ZN(n7342) );
  NAND2_X1 U8779 ( .A1(n7050), .A2(n9506), .ZN(n7127) );
  NAND2_X1 U8780 ( .A1(n7342), .A2(n7127), .ZN(n7354) );
  NAND2_X1 U8781 ( .A1(n7035), .A2(n7136), .ZN(n7363) );
  INV_X1 U8782 ( .A(n7363), .ZN(n7036) );
  AOI21_X1 U8783 ( .B1(n7353), .B2(n7354), .A(n7036), .ZN(n7483) );
  NAND2_X1 U8784 ( .A1(n8734), .A2(n7123), .ZN(n7339) );
  INV_X1 U8785 ( .A(n7339), .ZN(n7037) );
  NOR2_X1 U8786 ( .A1(n7038), .A2(n7037), .ZN(n7482) );
  NAND2_X1 U8787 ( .A1(n7482), .A2(n7348), .ZN(n7039) );
  NAND2_X1 U8788 ( .A1(n7483), .A2(n7039), .ZN(n7520) );
  NAND2_X1 U8789 ( .A1(n7523), .A2(n7520), .ZN(n7041) );
  INV_X1 U8790 ( .A(n8731), .ZN(n7040) );
  OR2_X1 U8791 ( .A1(n7283), .A2(n7040), .ZN(n7521) );
  XNOR2_X1 U8792 ( .A(n7041), .B(n7075), .ZN(n7044) );
  NAND2_X1 U8793 ( .A1(n8730), .A2(n8859), .ZN(n7043) );
  NAND2_X1 U8794 ( .A1(n8732), .A2(n8699), .ZN(n7042) );
  NAND2_X1 U8795 ( .A1(n7043), .A2(n7042), .ZN(n7279) );
  AOI21_X1 U8796 ( .B1(n7044), .B2(n9459), .A(n7279), .ZN(n9526) );
  NAND2_X1 U8797 ( .A1(n7045), .A2(n7480), .ZN(n7049) );
  NAND2_X1 U8798 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  NAND2_X1 U8799 ( .A1(n7049), .A2(n7048), .ZN(n7111) );
  NAND2_X1 U8800 ( .A1(n7127), .A2(n7339), .ZN(n7350) );
  NAND2_X1 U8801 ( .A1(n7050), .A2(n7123), .ZN(n7051) );
  NAND2_X1 U8802 ( .A1(n7342), .A2(n7340), .ZN(n7129) );
  NAND2_X1 U8803 ( .A1(n7360), .A2(n7363), .ZN(n7133) );
  NAND2_X1 U8804 ( .A1(n7132), .A2(n7133), .ZN(n7054) );
  OR2_X1 U8805 ( .A1(n8732), .A2(n7136), .ZN(n7053) );
  NAND2_X1 U8806 ( .A1(n7054), .A2(n7053), .ZN(n7073) );
  XNOR2_X1 U8807 ( .A(n7073), .B(n7075), .ZN(n9529) );
  NAND2_X1 U8808 ( .A1(n9529), .A2(n9441), .ZN(n7061) );
  INV_X1 U8809 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7056) );
  INV_X1 U8810 ( .A(n7055), .ZN(n7281) );
  OAI22_X1 U8811 ( .A1(n9452), .A2(n7056), .B1(n7281), .B2(n7121), .ZN(n7059)
         );
  INV_X1 U8812 ( .A(n7283), .ZN(n9527) );
  OAI211_X1 U8813 ( .C1(n7057), .C2(n9527), .A(n7081), .B(n9436), .ZN(n9525)
         );
  NOR2_X1 U8814 ( .A1(n9525), .A2(n8871), .ZN(n7058) );
  AOI211_X1 U8815 ( .C1(n9431), .C2(n7283), .A(n7059), .B(n7058), .ZN(n7060)
         );
  OAI211_X1 U8816 ( .C1(n9526), .C2(n9455), .A(n7061), .B(n7060), .ZN(P1_U3283) );
  INV_X1 U8817 ( .A(n8092), .ZN(n7067) );
  INV_X1 U8818 ( .A(n7062), .ZN(n7064) );
  XNOR2_X1 U8819 ( .A(n7874), .B(n7070), .ZN(n7191) );
  XNOR2_X1 U8820 ( .A(n7191), .B(n8091), .ZN(n7065) );
  OAI211_X1 U8821 ( .C1(n7066), .C2(n7065), .A(n7193), .B(n4824), .ZN(n7072)
         );
  INV_X1 U8822 ( .A(n8090), .ZN(n7147) );
  OAI22_X1 U8823 ( .A1(n8075), .A2(n7067), .B1(n7147), .B2(n8061), .ZN(n7068)
         );
  AOI211_X1 U8824 ( .C1(n7070), .C2(n8064), .A(n7069), .B(n7068), .ZN(n7071)
         );
  OAI211_X1 U8825 ( .C1(n7101), .C2(n8053), .A(n7072), .B(n7071), .ZN(P2_U3179) );
  INV_X1 U8826 ( .A(n8730), .ZN(n7174) );
  OR2_X1 U8827 ( .A1(n9264), .A2(n7174), .ZN(n7366) );
  NAND2_X1 U8828 ( .A1(n9264), .A2(n7174), .ZN(n7361) );
  NAND2_X1 U8829 ( .A1(n7366), .A2(n7361), .ZN(n7486) );
  INV_X1 U8830 ( .A(n7486), .ZN(n7074) );
  XNOR2_X1 U8831 ( .A(n7173), .B(n7074), .ZN(n9534) );
  INV_X1 U8832 ( .A(n7075), .ZN(n7484) );
  NAND3_X1 U8833 ( .A1(n7523), .A2(n7484), .A3(n7520), .ZN(n7177) );
  NAND2_X1 U8834 ( .A1(n7177), .A2(n7358), .ZN(n7076) );
  XNOR2_X1 U8835 ( .A(n7076), .B(n7486), .ZN(n7079) );
  NAND2_X1 U8836 ( .A1(n8729), .A2(n8859), .ZN(n7078) );
  NAND2_X1 U8837 ( .A1(n8731), .A2(n8699), .ZN(n7077) );
  AND2_X1 U8838 ( .A1(n7078), .A2(n7077), .ZN(n9256) );
  OAI21_X1 U8839 ( .B1(n7079), .B2(n9399), .A(n9256), .ZN(n7080) );
  AOI21_X1 U8840 ( .B1(n9534), .B2(n9513), .A(n7080), .ZN(n9536) );
  AOI21_X1 U8841 ( .B1(n7081), .B2(n9264), .A(n9101), .ZN(n7082) );
  OR2_X2 U8842 ( .A1(n7081), .A2(n9264), .ZN(n7183) );
  NAND2_X1 U8843 ( .A1(n7082), .A2(n7183), .ZN(n9531) );
  AOI22_X1 U8844 ( .A1(n9455), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7083), .B2(
        n9447), .ZN(n7085) );
  NAND2_X1 U8845 ( .A1(n9264), .A2(n9431), .ZN(n7084) );
  OAI211_X1 U8846 ( .C1(n9531), .C2(n8871), .A(n7085), .B(n7084), .ZN(n7086)
         );
  AOI21_X1 U8847 ( .B1(n9534), .B2(n9424), .A(n7086), .ZN(n7087) );
  OAI21_X1 U8848 ( .B1(n9536), .B2(n9455), .A(n7087), .ZN(P1_U3282) );
  INV_X1 U8849 ( .A(n7088), .ZN(n7143) );
  OAI222_X1 U8850 ( .A1(n7569), .A2(n7143), .B1(n5160), .B2(P1_U3086), .C1(
        n7089), .C2(n7620), .ZN(P1_U3335) );
  NAND2_X1 U8851 ( .A1(n7090), .A2(n7665), .ZN(n7091) );
  NAND2_X1 U8852 ( .A1(n7092), .A2(n7091), .ZN(n9800) );
  XNOR2_X1 U8853 ( .A(n7093), .B(n7665), .ZN(n7094) );
  NAND2_X1 U8854 ( .A1(n7094), .A2(n8355), .ZN(n7096) );
  AOI22_X1 U8855 ( .A1(n8352), .A2(n8091), .B1(n8089), .B2(n9758), .ZN(n7095)
         );
  OAI211_X1 U8856 ( .C1(n9800), .C2(n7257), .A(n7096), .B(n7095), .ZN(n9802)
         );
  NAND2_X1 U8857 ( .A1(n9802), .A2(n8376), .ZN(n7099) );
  OAI22_X1 U8858 ( .A1(n8376), .A2(n5914), .B1(n7199), .B2(n8373), .ZN(n7097)
         );
  AOI21_X1 U8859 ( .B1(n8378), .B2(n7200), .A(n7097), .ZN(n7098) );
  OAI211_X1 U8860 ( .C1(n9800), .C2(n8186), .A(n7099), .B(n7098), .ZN(P2_U3226) );
  XNOR2_X1 U8861 ( .A(n7100), .B(n7815), .ZN(n9798) );
  OAI22_X1 U8862 ( .A1(n8180), .A2(n9795), .B1(n7101), .B2(n8373), .ZN(n7109)
         );
  XNOR2_X1 U8863 ( .A(n7104), .B(n7815), .ZN(n7105) );
  NAND2_X1 U8864 ( .A1(n7105), .A2(n8355), .ZN(n7107) );
  AOI22_X1 U8865 ( .A1(n8352), .A2(n8092), .B1(n8090), .B2(n9758), .ZN(n7106)
         );
  NAND2_X1 U8866 ( .A1(n7107), .A2(n7106), .ZN(n9796) );
  MUX2_X1 U8867 ( .A(n9796), .B(P2_REG2_REG_6__SCAN_IN), .S(n9773), .Z(n7108)
         );
  AOI211_X1 U8868 ( .C1(n8361), .C2(n9798), .A(n7109), .B(n7108), .ZN(n7110)
         );
  INV_X1 U8869 ( .A(n7110), .ZN(P2_U3227) );
  XNOR2_X1 U8870 ( .A(n7111), .B(n4938), .ZN(n9510) );
  INV_X1 U8871 ( .A(n7348), .ZN(n7112) );
  INV_X1 U8872 ( .A(n7114), .ZN(n7341) );
  NAND2_X1 U8873 ( .A1(n7341), .A2(n4938), .ZN(n7128) );
  INV_X1 U8874 ( .A(n7128), .ZN(n7113) );
  AOI21_X1 U8875 ( .B1(n7350), .B2(n7114), .A(n7113), .ZN(n7116) );
  OAI21_X1 U8876 ( .B1(n7116), .B2(n9399), .A(n7115), .ZN(n9504) );
  INV_X1 U8877 ( .A(n9504), .ZN(n7117) );
  MUX2_X1 U8878 ( .A(n7118), .B(n7117), .S(n9452), .Z(n7126) );
  AOI211_X1 U8879 ( .C1(n9506), .C2(n7119), .A(n9101), .B(n4639), .ZN(n9505)
         );
  INV_X1 U8880 ( .A(n7120), .ZN(n7122) );
  OAI22_X1 U8881 ( .A1(n9104), .A2(n7123), .B1(n7122), .B2(n7121), .ZN(n7124)
         );
  AOI21_X1 U8882 ( .B1(n9505), .B2(n9440), .A(n7124), .ZN(n7125) );
  OAI211_X1 U8883 ( .C1(n9510), .C2(n9086), .A(n7126), .B(n7125), .ZN(P1_U3286) );
  NAND2_X1 U8884 ( .A1(n7128), .A2(n7127), .ZN(n9413) );
  NAND2_X1 U8885 ( .A1(n9413), .A2(n4941), .ZN(n9412) );
  NAND2_X1 U8886 ( .A1(n9412), .A2(n7342), .ZN(n7130) );
  XNOR2_X1 U8887 ( .A(n7130), .B(n7133), .ZN(n7131) );
  NAND2_X1 U8888 ( .A1(n8733), .A2(n8699), .ZN(n7214) );
  OAI21_X1 U8889 ( .B1(n7131), .B2(n9399), .A(n7214), .ZN(n9522) );
  INV_X1 U8890 ( .A(n9522), .ZN(n7141) );
  XNOR2_X1 U8891 ( .A(n7132), .B(n7133), .ZN(n9524) );
  INV_X1 U8892 ( .A(n7136), .ZN(n9521) );
  XNOR2_X1 U8893 ( .A(n9422), .B(n9521), .ZN(n7135) );
  NAND2_X1 U8894 ( .A1(n8731), .A2(n8859), .ZN(n7215) );
  INV_X1 U8895 ( .A(n7215), .ZN(n7134) );
  AOI21_X1 U8896 ( .B1(n7135), .B2(n9436), .A(n7134), .ZN(n9520) );
  AOI22_X1 U8897 ( .A1(n9455), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7218), .B2(
        n9447), .ZN(n7138) );
  NAND2_X1 U8898 ( .A1(n9431), .A2(n7136), .ZN(n7137) );
  OAI211_X1 U8899 ( .C1(n9520), .C2(n8871), .A(n7138), .B(n7137), .ZN(n7139)
         );
  AOI21_X1 U8900 ( .B1(n9524), .B2(n9441), .A(n7139), .ZN(n7140) );
  OAI21_X1 U8901 ( .B1(n7141), .B2(n9455), .A(n7140), .ZN(P1_U3284) );
  INV_X1 U8902 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7142) );
  OAI222_X1 U8903 ( .A1(n7784), .A2(P2_U3151), .B1(n8559), .B2(n7143), .C1(
        n7142), .C2(n8557), .ZN(P2_U3275) );
  XOR2_X1 U8904 ( .A(n7817), .B(n7144), .Z(n9806) );
  INV_X1 U8905 ( .A(n9806), .ZN(n7155) );
  NAND2_X1 U8906 ( .A1(n9773), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7145) );
  OAI21_X1 U8907 ( .B1(n7929), .B2(n8373), .A(n7145), .ZN(n7152) );
  AOI21_X1 U8908 ( .B1(n7146), .B2(n7817), .A(n9762), .ZN(n7150) );
  INV_X1 U8909 ( .A(n8088), .ZN(n7933) );
  OAI22_X1 U8910 ( .A1(n7147), .A2(n8372), .B1(n7933), .B2(n8370), .ZN(n7148)
         );
  AOI21_X1 U8911 ( .B1(n7150), .B2(n7149), .A(n7148), .ZN(n9803) );
  NOR2_X1 U8912 ( .A1(n9803), .A2(n9773), .ZN(n7151) );
  AOI211_X1 U8913 ( .C1(n8378), .C2(n7153), .A(n7152), .B(n7151), .ZN(n7154)
         );
  OAI21_X1 U8914 ( .B1(n7155), .B2(n8381), .A(n7154), .ZN(P2_U3225) );
  INV_X1 U8915 ( .A(n7156), .ZN(n7171) );
  OAI222_X1 U8916 ( .A1(n7569), .A2(n7171), .B1(n5759), .B2(P1_U3086), .C1(
        n7157), .C2(n7620), .ZN(P1_U3334) );
  OAI21_X1 U8917 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7168) );
  NOR2_X1 U8918 ( .A1(n8717), .A2(n9515), .ZN(n7167) );
  NAND2_X1 U8919 ( .A1(n8734), .A2(n8699), .ZN(n7162) );
  NAND2_X1 U8920 ( .A1(n8732), .A2(n8859), .ZN(n7161) );
  NAND2_X1 U8921 ( .A1(n7162), .A2(n7161), .ZN(n9417) );
  NAND2_X1 U8922 ( .A1(n9417), .A2(n8660), .ZN(n7164) );
  OAI211_X1 U8923 ( .C1(n9267), .C2(n7165), .A(n7164), .B(n7163), .ZN(n7166)
         );
  AOI211_X1 U8924 ( .C1(n7168), .C2(n8709), .A(n7167), .B(n7166), .ZN(n7169)
         );
  INV_X1 U8925 ( .A(n7169), .ZN(P1_U3221) );
  OAI222_X1 U8926 ( .A1(n7172), .A2(P2_U3151), .B1(n8559), .B2(n7171), .C1(
        n7170), .C2(n8557), .ZN(P2_U3274) );
  INV_X1 U8927 ( .A(n9264), .ZN(n9532) );
  NOR2_X1 U8928 ( .A1(n9532), .A2(n7174), .ZN(n7175) );
  INV_X1 U8929 ( .A(n8729), .ZN(n7176) );
  NAND2_X1 U8930 ( .A1(n7221), .A2(n7176), .ZN(n7526) );
  XNOR2_X1 U8931 ( .A(n7222), .B(n7489), .ZN(n9542) );
  INV_X1 U8932 ( .A(n9542), .ZN(n7189) );
  AND2_X1 U8933 ( .A1(n7361), .A2(n7358), .ZN(n7524) );
  NAND2_X1 U8934 ( .A1(n7177), .A2(n7524), .ZN(n7178) );
  NAND2_X1 U8935 ( .A1(n7178), .A2(n7366), .ZN(n7179) );
  NAND2_X1 U8936 ( .A1(n7179), .A2(n7489), .ZN(n7229) );
  OAI211_X1 U8937 ( .C1(n7489), .C2(n7179), .A(n7229), .B(n9459), .ZN(n7182)
         );
  NAND2_X1 U8938 ( .A1(n8728), .A2(n8859), .ZN(n7181) );
  NAND2_X1 U8939 ( .A1(n8730), .A2(n8699), .ZN(n7180) );
  AND2_X1 U8940 ( .A1(n7181), .A2(n7180), .ZN(n8610) );
  NAND2_X1 U8941 ( .A1(n7182), .A2(n8610), .ZN(n9540) );
  INV_X1 U8942 ( .A(n7221), .ZN(n9538) );
  INV_X1 U8943 ( .A(n7183), .ZN(n7184) );
  NOR2_X2 U8944 ( .A1(n7183), .A2(n7221), .ZN(n7235) );
  INV_X1 U8945 ( .A(n7235), .ZN(n7236) );
  OAI211_X1 U8946 ( .C1(n9538), .C2(n7184), .A(n7236), .B(n9436), .ZN(n9537)
         );
  AOI22_X1 U8947 ( .A1(n9455), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8612), .B2(
        n9447), .ZN(n7186) );
  NAND2_X1 U8948 ( .A1(n7221), .A2(n9431), .ZN(n7185) );
  OAI211_X1 U8949 ( .C1(n9537), .C2(n8871), .A(n7186), .B(n7185), .ZN(n7187)
         );
  AOI21_X1 U8950 ( .B1(n9540), .B2(n9452), .A(n7187), .ZN(n7188) );
  OAI21_X1 U8951 ( .B1(n7189), .B2(n9086), .A(n7188), .ZN(P1_U3281) );
  XNOR2_X1 U8952 ( .A(n9799), .B(n7874), .ZN(n7572) );
  XNOR2_X1 U8953 ( .A(n7572), .B(n8090), .ZN(n7198) );
  INV_X1 U8954 ( .A(n8091), .ZN(n7190) );
  NAND2_X1 U8955 ( .A1(n7193), .A2(n7192), .ZN(n7197) );
  INV_X1 U8956 ( .A(n7197), .ZN(n7195) );
  NAND2_X1 U8957 ( .A1(n7195), .A2(n7194), .ZN(n7574) );
  INV_X1 U8958 ( .A(n7574), .ZN(n7196) );
  AOI21_X1 U8959 ( .B1(n7198), .B2(n7197), .A(n7196), .ZN(n7209) );
  INV_X1 U8960 ( .A(n7199), .ZN(n7207) );
  NAND2_X1 U8961 ( .A1(n8073), .A2(n8089), .ZN(n7205) );
  NAND2_X1 U8962 ( .A1(n8058), .A2(n8091), .ZN(n7204) );
  NAND2_X1 U8963 ( .A1(n8064), .A2(n7200), .ZN(n7203) );
  INV_X1 U8964 ( .A(n7201), .ZN(n7202) );
  NAND4_X1 U8965 ( .A1(n7205), .A2(n7204), .A3(n7203), .A4(n7202), .ZN(n7206)
         );
  AOI21_X1 U8966 ( .B1(n7207), .B2(n8078), .A(n7206), .ZN(n7208) );
  OAI21_X1 U8967 ( .B1(n7209), .B2(n8067), .A(n7208), .ZN(P2_U3153) );
  AND2_X1 U8968 ( .A1(n7210), .A2(n7158), .ZN(n7213) );
  OAI211_X1 U8969 ( .C1(n7213), .C2(n7212), .A(n8709), .B(n7211), .ZN(n7220)
         );
  AOI21_X1 U8970 ( .B1(n7215), .B2(n7214), .A(n9255), .ZN(n7216) );
  AOI211_X1 U8971 ( .C1(n8713), .C2(n7218), .A(n7217), .B(n7216), .ZN(n7219)
         );
  OAI211_X1 U8972 ( .C1(n9521), .C2(n8717), .A(n7220), .B(n7219), .ZN(P1_U3231) );
  INV_X1 U8973 ( .A(n8728), .ZN(n7223) );
  OR2_X1 U8974 ( .A1(n9199), .A2(n7223), .ZN(n7368) );
  NAND2_X1 U8975 ( .A1(n9199), .A2(n7223), .ZN(n9395) );
  NAND2_X1 U8976 ( .A1(n7368), .A2(n9395), .ZN(n7228) );
  OAI21_X1 U8977 ( .B1(n7224), .B2(n7228), .A(n7308), .ZN(n7225) );
  INV_X1 U8978 ( .A(n7225), .ZN(n9201) );
  INV_X1 U8979 ( .A(n7367), .ZN(n7226) );
  NOR2_X1 U8980 ( .A1(n7228), .A2(n7226), .ZN(n7227) );
  INV_X1 U8981 ( .A(n9396), .ZN(n7231) );
  INV_X1 U8982 ( .A(n7228), .ZN(n7490) );
  AOI21_X1 U8983 ( .B1(n7229), .B2(n7367), .A(n7490), .ZN(n7230) );
  OAI21_X1 U8984 ( .B1(n7231), .B2(n7230), .A(n9459), .ZN(n7234) );
  OR2_X1 U8985 ( .A1(n7309), .A2(n8697), .ZN(n7233) );
  NAND2_X1 U8986 ( .A1(n8729), .A2(n8699), .ZN(n7232) );
  AND2_X1 U8987 ( .A1(n7233), .A2(n7232), .ZN(n7294) );
  NAND2_X1 U8988 ( .A1(n7234), .A2(n7294), .ZN(n9197) );
  INV_X1 U8989 ( .A(n9199), .ZN(n7300) );
  AND2_X2 U8990 ( .A1(n7235), .A2(n7300), .ZN(n9408) );
  AOI211_X1 U8991 ( .C1(n9199), .C2(n7236), .A(n9101), .B(n9408), .ZN(n9198)
         );
  NAND2_X1 U8992 ( .A1(n9198), .A2(n9440), .ZN(n7238) );
  AOI22_X1 U8993 ( .A1(n9455), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7297), .B2(
        n9447), .ZN(n7237) );
  OAI211_X1 U8994 ( .C1(n7300), .C2(n9104), .A(n7238), .B(n7237), .ZN(n7239)
         );
  AOI21_X1 U8995 ( .B1(n9452), .B2(n9197), .A(n7239), .ZN(n7240) );
  OAI21_X1 U8996 ( .B1(n9201), .B2(n9086), .A(n7240), .ZN(P1_U3280) );
  NAND2_X1 U8997 ( .A1(n7682), .A2(n7684), .ZN(n7821) );
  INV_X1 U8998 ( .A(n7821), .ZN(n7242) );
  XNOR2_X1 U8999 ( .A(n7241), .B(n7242), .ZN(n7243) );
  NAND2_X1 U9000 ( .A1(n7243), .A2(n8355), .ZN(n7245) );
  AOI22_X1 U9001 ( .A1(n8352), .A2(n8088), .B1(n8086), .B2(n9758), .ZN(n7244)
         );
  AND2_X1 U9002 ( .A1(n7245), .A2(n7244), .ZN(n9817) );
  NAND2_X1 U9003 ( .A1(n7246), .A2(n7247), .ZN(n7248) );
  XNOR2_X1 U9004 ( .A(n7248), .B(n7821), .ZN(n9813) );
  NOR2_X1 U9005 ( .A1(n8180), .A2(n7914), .ZN(n7250) );
  OAI22_X1 U9006 ( .A1(n8376), .A2(n8096), .B1(n7908), .B2(n8373), .ZN(n7249)
         );
  AOI211_X1 U9007 ( .C1(n9813), .C2(n8361), .A(n7250), .B(n7249), .ZN(n7251)
         );
  OAI21_X1 U9008 ( .B1(n9817), .B2(n9773), .A(n7251), .ZN(P2_U3223) );
  OAI21_X1 U9009 ( .B1(n7252), .B2(n7819), .A(n7246), .ZN(n9809) );
  AOI22_X1 U9010 ( .A1(n8352), .A2(n8089), .B1(n8087), .B2(n9758), .ZN(n7256)
         );
  XNOR2_X1 U9011 ( .A(n7253), .B(n7819), .ZN(n7254) );
  NAND2_X1 U9012 ( .A1(n7254), .A2(n8355), .ZN(n7255) );
  OAI211_X1 U9013 ( .C1(n9809), .C2(n7257), .A(n7256), .B(n7255), .ZN(n9811)
         );
  INV_X1 U9014 ( .A(n7258), .ZN(n7993) );
  AOI22_X1 U9015 ( .A1(n9773), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9768), .B2(
        n7993), .ZN(n7260) );
  OR2_X1 U9016 ( .A1(n8180), .A2(n9807), .ZN(n7259) );
  OAI211_X1 U9017 ( .C1(n9809), .C2(n8186), .A(n7260), .B(n7259), .ZN(n7261)
         );
  AOI21_X1 U9018 ( .B1(n9811), .B2(n8376), .A(n7261), .ZN(n7262) );
  INV_X1 U9019 ( .A(n7262), .ZN(P2_U3224) );
  OAI211_X1 U9020 ( .C1(n7264), .C2(n7822), .A(n7263), .B(n8355), .ZN(n7266)
         );
  AOI22_X1 U9021 ( .A1(n8352), .A2(n8087), .B1(n8353), .B2(n9758), .ZN(n7265)
         );
  OAI22_X1 U9022 ( .A1(n8376), .A2(n5978), .B1(n8037), .B2(n8373), .ZN(n7267)
         );
  AOI21_X1 U9023 ( .B1(n8378), .B2(n8044), .A(n7267), .ZN(n7271) );
  INV_X1 U9024 ( .A(n7822), .ZN(n7268) );
  XNOR2_X1 U9025 ( .A(n7269), .B(n7268), .ZN(n9820) );
  NAND2_X1 U9026 ( .A1(n9820), .A2(n8361), .ZN(n7270) );
  OAI211_X1 U9027 ( .C1(n9825), .C2(n9773), .A(n7271), .B(n7270), .ZN(P2_U3222) );
  INV_X1 U9028 ( .A(n7272), .ZN(n7564) );
  OAI222_X1 U9029 ( .A1(P2_U3151), .A2(n7274), .B1(n8559), .B2(n7564), .C1(
        n7273), .C2(n8557), .ZN(P2_U3273) );
  INV_X1 U9030 ( .A(n7286), .ZN(n7277) );
  AOI21_X1 U9031 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8552), .A(n7275), .ZN(
        n7276) );
  OAI21_X1 U9032 ( .B1(n7277), .B2(n8559), .A(n7276), .ZN(P2_U3272) );
  XOR2_X1 U9033 ( .A(n7278), .B(n8600), .Z(n8603) );
  XNOR2_X1 U9034 ( .A(n8603), .B(n8602), .ZN(n7285) );
  NAND2_X1 U9035 ( .A1(n7279), .A2(n8660), .ZN(n7280) );
  NAND2_X1 U9036 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9251) );
  OAI211_X1 U9037 ( .C1(n9267), .C2(n7281), .A(n7280), .B(n9251), .ZN(n7282)
         );
  AOI21_X1 U9038 ( .B1(n7283), .B2(n5768), .A(n7282), .ZN(n7284) );
  OAI21_X1 U9039 ( .B1(n7285), .B2(n9260), .A(n7284), .ZN(P1_U3217) );
  NAND2_X1 U9040 ( .A1(n7286), .A2(n9226), .ZN(n7287) );
  OAI211_X1 U9041 ( .C1(n7288), .C2(n7620), .A(n7287), .B(n7562), .ZN(P1_U3332) );
  AND3_X1 U9042 ( .A1(n7289), .A2(n7291), .A3(n7290), .ZN(n7292) );
  OAI21_X1 U9043 ( .B1(n7293), .B2(n7292), .A(n8709), .ZN(n7299) );
  NAND2_X1 U9044 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9334) );
  INV_X1 U9045 ( .A(n9334), .ZN(n7296) );
  NOR2_X1 U9046 ( .A1(n7294), .A2(n9255), .ZN(n7295) );
  AOI211_X1 U9047 ( .C1(n8713), .C2(n7297), .A(n7296), .B(n7295), .ZN(n7298)
         );
  OAI211_X1 U9048 ( .C1(n7300), .C2(n8717), .A(n7299), .B(n7298), .ZN(P1_U3234) );
  OR2_X1 U9049 ( .A1(n9545), .A2(n8727), .ZN(n7372) );
  NAND2_X1 U9050 ( .A1(n9545), .A2(n8727), .ZN(n7374) );
  NAND2_X1 U9051 ( .A1(n7372), .A2(n7374), .ZN(n9401) );
  INV_X1 U9052 ( .A(n9395), .ZN(n7301) );
  NOR2_X1 U9053 ( .A1(n9401), .A2(n7301), .ZN(n7302) );
  OR2_X1 U9054 ( .A1(n9276), .A2(n8874), .ZN(n7443) );
  NAND2_X1 U9055 ( .A1(n9276), .A2(n8874), .ZN(n7376) );
  NAND2_X1 U9056 ( .A1(n7443), .A2(n7376), .ZN(n7472) );
  XNOR2_X1 U9057 ( .A(n7442), .B(n7472), .ZN(n7306) );
  OR2_X1 U9058 ( .A1(n7309), .A2(n8927), .ZN(n7304) );
  NAND2_X1 U9059 ( .A1(n8875), .A2(n8859), .ZN(n7303) );
  AND2_X1 U9060 ( .A1(n7304), .A2(n7303), .ZN(n8711) );
  INV_X1 U9061 ( .A(n8711), .ZN(n7305) );
  AOI21_X1 U9062 ( .B1(n7306), .B2(n9459), .A(n7305), .ZN(n9275) );
  NAND2_X1 U9063 ( .A1(n7308), .A2(n7307), .ZN(n9394) );
  AOI21_X1 U9064 ( .B1(n7309), .B2(n9545), .A(n9394), .ZN(n7310) );
  XNOR2_X1 U9065 ( .A(n8873), .B(n7472), .ZN(n9278) );
  NAND2_X1 U9066 ( .A1(n9278), .A2(n9441), .ZN(n7316) );
  INV_X1 U9067 ( .A(n9407), .ZN(n7311) );
  OAI211_X1 U9068 ( .C1(n7311), .C2(n9276), .A(n9436), .B(n9102), .ZN(n9274)
         );
  INV_X1 U9069 ( .A(n9274), .ZN(n7314) );
  AOI22_X1 U9070 ( .A1(n9455), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8714), .B2(
        n9447), .ZN(n7312) );
  OAI21_X1 U9071 ( .B1(n9276), .B2(n9104), .A(n7312), .ZN(n7313) );
  AOI21_X1 U9072 ( .B1(n7314), .B2(n9440), .A(n7313), .ZN(n7315) );
  OAI211_X1 U9073 ( .C1(n9455), .C2(n9275), .A(n7316), .B(n7315), .ZN(P1_U3278) );
  INV_X1 U9074 ( .A(n7317), .ZN(n7571) );
  OAI222_X1 U9075 ( .A1(n7569), .A2(n7571), .B1(n4420), .B2(P1_U3086), .C1(
        n7318), .C2(n7620), .ZN(P1_U3331) );
  INV_X1 U9076 ( .A(SI_29_), .ZN(n7322) );
  OR2_X1 U9077 ( .A1(n7320), .A2(n7319), .ZN(n7321) );
  INV_X1 U9078 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7619) );
  INV_X1 U9079 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10086) );
  MUX2_X1 U9080 ( .A(n7619), .B(n10086), .S(n4418), .Z(n7325) );
  INV_X1 U9081 ( .A(SI_30_), .ZN(n7324) );
  NAND2_X1 U9082 ( .A1(n7325), .A2(n7324), .ZN(n7328) );
  INV_X1 U9083 ( .A(n7325), .ZN(n7326) );
  NAND2_X1 U9084 ( .A1(n7326), .A2(SI_30_), .ZN(n7327) );
  NAND2_X1 U9085 ( .A1(n7328), .A2(n7327), .ZN(n7416) );
  NAND2_X1 U9086 ( .A1(n7419), .A2(n7328), .ZN(n7331) );
  INV_X1 U9087 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9223) );
  MUX2_X1 U9088 ( .A(n9223), .B(n6421), .S(n4418), .Z(n7329) );
  XNOR2_X1 U9089 ( .A(n7329), .B(SI_31_), .ZN(n7330) );
  NAND2_X1 U9090 ( .A1(n9227), .A2(n7420), .ZN(n7333) );
  OR2_X1 U9091 ( .A1(n5259), .A2(n9223), .ZN(n7332) );
  OR2_X1 U9092 ( .A1(n9192), .A2(n7335), .ZN(n7445) );
  INV_X1 U9093 ( .A(n7443), .ZN(n7334) );
  NAND2_X1 U9094 ( .A1(n7445), .A2(n7334), .ZN(n7336) );
  NAND2_X1 U9095 ( .A1(n9192), .A2(n7335), .ZN(n7533) );
  OAI211_X1 U9096 ( .C1(n7337), .C2(n9130), .A(n7336), .B(n7533), .ZN(n7379)
         );
  INV_X1 U9097 ( .A(n7533), .ZN(n7338) );
  OAI21_X1 U9098 ( .B1(n7338), .B2(n8872), .A(n4724), .ZN(n7378) );
  OAI211_X1 U9099 ( .C1(n7341), .C2(n7350), .A(n7340), .B(n7339), .ZN(n7343)
         );
  NAND3_X1 U9100 ( .A1(n7343), .A2(n7363), .A3(n7342), .ZN(n7357) );
  INV_X1 U9101 ( .A(n7516), .ZN(n7346) );
  OAI211_X1 U9102 ( .C1(n9427), .C2(n7346), .A(n7345), .B(n7344), .ZN(n7349)
         );
  NAND3_X1 U9103 ( .A1(n7349), .A2(n7348), .A3(n7347), .ZN(n7352) );
  AOI21_X1 U9104 ( .B1(n7352), .B2(n7351), .A(n7350), .ZN(n7355) );
  OAI21_X1 U9105 ( .B1(n7355), .B2(n7354), .A(n7353), .ZN(n7356) );
  INV_X1 U9106 ( .A(n7358), .ZN(n7359) );
  NAND2_X1 U9107 ( .A1(n7366), .A2(n7521), .ZN(n7362) );
  INV_X1 U9108 ( .A(n7524), .ZN(n7365) );
  NAND2_X1 U9109 ( .A1(n7367), .A2(n7366), .ZN(n7527) );
  AND2_X1 U9110 ( .A1(n7374), .A2(n7368), .ZN(n7531) );
  INV_X1 U9111 ( .A(n7531), .ZN(n7369) );
  AOI21_X1 U9112 ( .B1(n7375), .B2(n9395), .A(n7369), .ZN(n7371) );
  AND2_X1 U9113 ( .A1(n7443), .A2(n7372), .ZN(n7529) );
  NAND2_X1 U9114 ( .A1(n7533), .A2(n7529), .ZN(n7370) );
  NAND2_X1 U9115 ( .A1(n7372), .A2(n9395), .ZN(n7373) );
  AOI22_X1 U9116 ( .A1(n7375), .A2(n7531), .B1(n7374), .B2(n7373), .ZN(n7377)
         );
  NAND2_X1 U9117 ( .A1(n7445), .A2(n7376), .ZN(n7534) );
  OR2_X1 U9118 ( .A1(n8880), .A2(n8877), .ZN(n7537) );
  NAND2_X1 U9119 ( .A1(n8880), .A2(n8877), .ZN(n7381) );
  NAND2_X1 U9120 ( .A1(n7537), .A2(n7381), .ZN(n9093) );
  INV_X1 U9121 ( .A(n8882), .ZN(n8881) );
  OR2_X1 U9122 ( .A1(n9187), .A2(n8881), .ZN(n7448) );
  INV_X1 U9123 ( .A(n7448), .ZN(n7494) );
  INV_X1 U9124 ( .A(n7537), .ZN(n7446) );
  NOR3_X1 U9125 ( .A1(n7382), .A2(n7494), .A3(n7446), .ZN(n7380) );
  INV_X1 U9126 ( .A(n8885), .ZN(n8886) );
  NAND2_X1 U9127 ( .A1(n9187), .A2(n8881), .ZN(n7447) );
  INV_X1 U9128 ( .A(n7447), .ZN(n7449) );
  NOR3_X1 U9129 ( .A1(n7380), .A2(n4809), .A3(n7449), .ZN(n7385) );
  NAND2_X1 U9130 ( .A1(n7447), .A2(n7381), .ZN(n7536) );
  NOR2_X1 U9131 ( .A1(n7382), .A2(n7536), .ZN(n7383) );
  OR2_X1 U9132 ( .A1(n9182), .A2(n8886), .ZN(n7450) );
  NAND2_X1 U9133 ( .A1(n7450), .A2(n7448), .ZN(n7540) );
  INV_X1 U9134 ( .A(n8725), .ZN(n8888) );
  NAND2_X1 U9135 ( .A1(n9177), .A2(n8888), .ZN(n7471) );
  OAI211_X1 U9136 ( .C1(n7383), .C2(n7540), .A(n7471), .B(n7539), .ZN(n7384)
         );
  AOI21_X1 U9137 ( .B1(n9034), .B2(n7450), .A(n9130), .ZN(n7386) );
  NOR2_X1 U9138 ( .A1(n7387), .A2(n7386), .ZN(n7391) );
  INV_X1 U9139 ( .A(n8724), .ZN(n8889) );
  NAND2_X1 U9140 ( .A1(n9172), .A2(n8889), .ZN(n7470) );
  NAND2_X1 U9141 ( .A1(n7470), .A2(n7471), .ZN(n7433) );
  OR2_X1 U9142 ( .A1(n9172), .A2(n8889), .ZN(n7543) );
  NAND2_X1 U9143 ( .A1(n7543), .A2(n9034), .ZN(n7388) );
  MUX2_X1 U9144 ( .A(n7433), .B(n7388), .S(n9130), .Z(n7390) );
  MUX2_X1 U9145 ( .A(n7470), .B(n7543), .S(n4724), .Z(n7389) );
  OAI21_X1 U9146 ( .B1(n7391), .B2(n7390), .A(n7389), .ZN(n7393) );
  INV_X1 U9147 ( .A(n8892), .ZN(n8723) );
  OR2_X1 U9148 ( .A1(n9030), .A2(n8723), .ZN(n7434) );
  NAND2_X1 U9149 ( .A1(n9030), .A2(n8723), .ZN(n8916) );
  NAND2_X1 U9150 ( .A1(n7434), .A2(n8916), .ZN(n8915) );
  INV_X1 U9151 ( .A(n8895), .ZN(n7392) );
  OR2_X1 U9152 ( .A1(n9161), .A2(n7392), .ZN(n7395) );
  NAND2_X1 U9153 ( .A1(n9161), .A2(n7392), .ZN(n8918) );
  NAND2_X1 U9154 ( .A1(n7395), .A2(n8916), .ZN(n7394) );
  NAND2_X1 U9155 ( .A1(n7394), .A2(n8918), .ZN(n7430) );
  INV_X1 U9156 ( .A(n7434), .ZN(n7396) );
  OAI21_X1 U9157 ( .B1(n4802), .B2(n7396), .A(n7395), .ZN(n7397) );
  MUX2_X1 U9158 ( .A(n7430), .B(n7397), .S(n9130), .Z(n7398) );
  INV_X1 U9159 ( .A(n8722), .ZN(n8896) );
  OR2_X1 U9160 ( .A1(n9157), .A2(n8896), .ZN(n8919) );
  NAND2_X1 U9161 ( .A1(n9157), .A2(n8896), .ZN(n7435) );
  NAND2_X1 U9162 ( .A1(n8919), .A2(n7435), .ZN(n8990) );
  NAND2_X1 U9163 ( .A1(n8952), .A2(n8904), .ZN(n7466) );
  NAND2_X1 U9164 ( .A1(n9146), .A2(n8901), .ZN(n8921) );
  NAND2_X1 U9165 ( .A1(n9152), .A2(n8898), .ZN(n7468) );
  AND2_X1 U9166 ( .A1(n8921), .A2(n7468), .ZN(n7400) );
  OR2_X1 U9167 ( .A1(n9152), .A2(n8898), .ZN(n7469) );
  MUX2_X1 U9168 ( .A(n8919), .B(n7435), .S(n9130), .Z(n7399) );
  INV_X1 U9169 ( .A(n7467), .ZN(n7402) );
  INV_X1 U9170 ( .A(n7469), .ZN(n8920) );
  INV_X1 U9171 ( .A(n7400), .ZN(n7404) );
  NAND2_X1 U9172 ( .A1(n7404), .A2(n7467), .ZN(n7401) );
  OAI211_X1 U9173 ( .C1(n7402), .C2(n8920), .A(n7401), .B(n9130), .ZN(n7403)
         );
  NAND4_X1 U9174 ( .A1(n7466), .A2(n4724), .A3(n7467), .A4(n7404), .ZN(n7405)
         );
  NAND2_X1 U9175 ( .A1(n7408), .A2(n4456), .ZN(n7410) );
  OAI21_X1 U9176 ( .B1(n7429), .B2(n7466), .A(n7465), .ZN(n7409) );
  AOI22_X1 U9177 ( .A1(n7410), .A2(n7465), .B1(n9130), .B2(n7409), .ZN(n7415)
         );
  NAND2_X1 U9178 ( .A1(n7566), .A2(n7420), .ZN(n7412) );
  OR2_X1 U9179 ( .A1(n5259), .A2(n7567), .ZN(n7411) );
  INV_X1 U9180 ( .A(n8719), .ZN(n7413) );
  OR2_X1 U9181 ( .A1(n9134), .A2(n7413), .ZN(n7440) );
  NAND2_X1 U9182 ( .A1(n9134), .A2(n7413), .ZN(n7455) );
  INV_X1 U9183 ( .A(n8905), .ZN(n8924) );
  MUX2_X1 U9184 ( .A(n7455), .B(n7440), .S(n9130), .Z(n7414) );
  NAND2_X1 U9185 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  NAND2_X1 U9186 ( .A1(n7419), .A2(n7418), .ZN(n7775) );
  NAND2_X1 U9187 ( .A1(n7775), .A2(n7420), .ZN(n7422) );
  OR2_X1 U9188 ( .A1(n5259), .A2(n7619), .ZN(n7421) );
  OR2_X1 U9189 ( .A1(n8861), .A2(n8860), .ZN(n7552) );
  NAND2_X1 U9190 ( .A1(n6416), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9191 ( .A1(n5248), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7425) );
  NAND2_X1 U9192 ( .A1(n7423), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7424) );
  AND3_X1 U9193 ( .A1(n7426), .A2(n7425), .A3(n7424), .ZN(n8928) );
  INV_X1 U9194 ( .A(n8928), .ZN(n8718) );
  NAND2_X1 U9195 ( .A1(n8718), .A2(n7427), .ZN(n7428) );
  AOI21_X1 U9196 ( .B1(n4724), .B2(n4445), .A(n7505), .ZN(n7511) );
  OAI211_X1 U9197 ( .C1(n7552), .C2(n5549), .A(n5761), .B(n7563), .ZN(n7510)
         );
  INV_X1 U9198 ( .A(n7428), .ZN(n7459) );
  INV_X1 U9199 ( .A(n7430), .ZN(n7431) );
  NAND2_X1 U9200 ( .A1(n7431), .A2(n7435), .ZN(n7432) );
  AND3_X1 U9201 ( .A1(n7469), .A2(n8919), .A3(n7432), .ZN(n7544) );
  NAND2_X1 U9202 ( .A1(n7433), .A2(n7543), .ZN(n8913) );
  NAND4_X1 U9203 ( .A1(n7435), .A2(n8918), .A3(n7434), .A4(n8913), .ZN(n7437)
         );
  INV_X1 U9204 ( .A(n7468), .ZN(n7436) );
  AOI21_X1 U9205 ( .B1(n7544), .B2(n7437), .A(n7436), .ZN(n7438) );
  INV_X1 U9206 ( .A(n7465), .ZN(n7439) );
  AND2_X1 U9207 ( .A1(n7441), .A2(n7440), .ZN(n7545) );
  INV_X1 U9208 ( .A(n9107), .ZN(n9110) );
  OAI21_X1 U9209 ( .B1(n9111), .B2(n9110), .A(n7533), .ZN(n9088) );
  INV_X1 U9210 ( .A(n7544), .ZN(n7454) );
  INV_X1 U9211 ( .A(n7451), .ZN(n7453) );
  INV_X1 U9212 ( .A(n8921), .ZN(n7452) );
  NOR2_X1 U9213 ( .A1(n7453), .A2(n7452), .ZN(n7548) );
  OAI21_X1 U9214 ( .B1(n8914), .B2(n7454), .A(n7548), .ZN(n7457) );
  AND2_X1 U9215 ( .A1(n8868), .A2(n8928), .ZN(n7501) );
  INV_X1 U9216 ( .A(n7501), .ZN(n7456) );
  NAND2_X1 U9217 ( .A1(n7456), .A2(n7455), .ZN(n7549) );
  AOI21_X1 U9218 ( .B1(n7545), .B2(n7457), .A(n7549), .ZN(n7458) );
  AOI211_X1 U9219 ( .C1(n9128), .C2(n7459), .A(n4445), .B(n7458), .ZN(n7462)
         );
  OAI21_X1 U9220 ( .B1(n9128), .B2(n8861), .A(n7552), .ZN(n7461) );
  OAI211_X1 U9221 ( .C1(n7462), .C2(n7461), .A(n7460), .B(n5549), .ZN(n7463)
         );
  AOI21_X1 U9222 ( .B1(n9128), .B2(n8718), .A(n4445), .ZN(n7551) );
  NAND2_X1 U9223 ( .A1(n7465), .A2(n7464), .ZN(n8923) );
  NAND2_X1 U9224 ( .A1(n8922), .A2(n7466), .ZN(n8903) );
  INV_X1 U9225 ( .A(n9010), .ZN(n7498) );
  NAND2_X1 U9226 ( .A1(n9034), .A2(n7471), .ZN(n9047) );
  INV_X1 U9227 ( .A(n9047), .ZN(n7496) );
  NOR2_X1 U9228 ( .A1(n7473), .A2(n6725), .ZN(n7478) );
  INV_X1 U9229 ( .A(n9434), .ZN(n7477) );
  NOR2_X1 U9230 ( .A1(n9458), .A2(n5761), .ZN(n7476) );
  NAND4_X1 U9231 ( .A1(n7478), .A2(n7477), .A3(n7476), .A4(n7475), .ZN(n7481)
         );
  NOR3_X1 U9232 ( .A1(n7481), .A2(n7480), .A3(n7479), .ZN(n7485) );
  NAND4_X1 U9233 ( .A1(n7485), .A2(n7484), .A3(n7483), .A4(n7482), .ZN(n7487)
         );
  NOR2_X1 U9234 ( .A1(n7487), .A2(n7486), .ZN(n7488) );
  NAND3_X1 U9235 ( .A1(n7490), .A2(n7489), .A3(n7488), .ZN(n7491) );
  NOR2_X1 U9236 ( .A1(n9401), .A2(n7491), .ZN(n7492) );
  NAND4_X1 U9237 ( .A1(n7537), .A2(n9107), .A3(n4786), .A4(n7492), .ZN(n7493)
         );
  NOR4_X1 U9238 ( .A1(n9062), .A2(n7494), .A3(n7536), .A4(n7493), .ZN(n7495)
         );
  NAND3_X1 U9239 ( .A1(n9035), .A2(n7496), .A3(n7495), .ZN(n7497) );
  NOR4_X1 U9240 ( .A1(n7498), .A2(n8990), .A3(n8915), .A4(n7497), .ZN(n7499)
         );
  NAND4_X1 U9241 ( .A1(n8955), .A2(n8969), .A3(n8977), .A4(n7499), .ZN(n7500)
         );
  NOR4_X1 U9242 ( .A1(n8924), .A2(n7501), .A3(n8923), .A4(n7500), .ZN(n7502)
         );
  NAND3_X1 U9243 ( .A1(n7552), .A2(n7551), .A3(n7502), .ZN(n7506) );
  OAI21_X1 U9244 ( .B1(n7505), .B2(n7563), .A(n5761), .ZN(n7507) );
  INV_X1 U9245 ( .A(n5160), .ZN(n9129) );
  NAND3_X1 U9246 ( .A1(n7513), .A2(n7512), .A3(n5761), .ZN(n7519) );
  NAND3_X1 U9247 ( .A1(n7516), .A2(n7515), .A3(n7514), .ZN(n7518) );
  NOR3_X1 U9248 ( .A1(n7519), .A2(n7518), .A3(n7517), .ZN(n7522) );
  OAI211_X1 U9249 ( .C1(n7523), .C2(n7522), .A(n7521), .B(n7520), .ZN(n7525)
         );
  AND2_X1 U9250 ( .A1(n7525), .A2(n7524), .ZN(n7528) );
  OAI211_X1 U9251 ( .C1(n7528), .C2(n7527), .A(n9395), .B(n7526), .ZN(n7532)
         );
  INV_X1 U9252 ( .A(n7529), .ZN(n7530) );
  AOI21_X1 U9253 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7535) );
  OAI21_X1 U9254 ( .B1(n7535), .B2(n7534), .A(n7533), .ZN(n7538) );
  AOI21_X1 U9255 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7541) );
  OAI21_X1 U9256 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7542) );
  NAND4_X1 U9257 ( .A1(n7544), .A2(n7543), .A3(n9034), .A4(n7542), .ZN(n7547)
         );
  INV_X1 U9258 ( .A(n7545), .ZN(n7546) );
  AOI21_X1 U9259 ( .B1(n7548), .B2(n7547), .A(n7546), .ZN(n7550) );
  NOR2_X1 U9260 ( .A1(n7550), .A2(n7549), .ZN(n7554) );
  INV_X1 U9261 ( .A(n7551), .ZN(n7553) );
  OAI21_X1 U9262 ( .B1(n7554), .B2(n7553), .A(n7552), .ZN(n7555) );
  NOR4_X1 U9263 ( .A1(n7559), .A2(n6722), .A3(n8752), .A4(n7558), .ZN(n7561)
         );
  OAI21_X1 U9264 ( .B1(n7562), .B2(n5760), .A(P1_B_REG_SCAN_IN), .ZN(n7560) );
  OAI222_X1 U9265 ( .A1(n7620), .A2(n7565), .B1(n7569), .B2(n7564), .C1(
        P1_U3086), .C2(n7563), .ZN(P1_U3333) );
  INV_X1 U9266 ( .A(n7566), .ZN(n8546) );
  OAI222_X1 U9267 ( .A1(n7569), .A2(n8546), .B1(P1_U3086), .B2(n7568), .C1(
        n7567), .C2(n7620), .ZN(P1_U3326) );
  OAI222_X1 U9268 ( .A1(n6214), .A2(P2_U3151), .B1(n8559), .B2(n7571), .C1(
        n7570), .C2(n8557), .ZN(P2_U3271) );
  XNOR2_X1 U9269 ( .A(n8486), .B(n7877), .ZN(n7851) );
  XNOR2_X1 U9270 ( .A(n7851), .B(n7853), .ZN(n7854) );
  XNOR2_X1 U9271 ( .A(n8527), .B(n7877), .ZN(n7592) );
  XNOR2_X1 U9272 ( .A(n9804), .B(n7874), .ZN(n7576) );
  XNOR2_X1 U9273 ( .A(n7575), .B(n7576), .ZN(n7926) );
  INV_X1 U9274 ( .A(n8089), .ZN(n7927) );
  XNOR2_X1 U9275 ( .A(n8004), .B(n7877), .ZN(n7580) );
  XNOR2_X1 U9276 ( .A(n7580), .B(n8088), .ZN(n8001) );
  INV_X1 U9277 ( .A(n8001), .ZN(n7579) );
  NAND2_X1 U9278 ( .A1(n7580), .A2(n8088), .ZN(n7581) );
  XNOR2_X1 U9279 ( .A(n9814), .B(n7874), .ZN(n7905) );
  XNOR2_X1 U9280 ( .A(n7822), .B(n7877), .ZN(n8034) );
  OAI21_X1 U9281 ( .B1(n7997), .B2(n7905), .A(n8034), .ZN(n7587) );
  XNOR2_X1 U9282 ( .A(n9831), .B(n7874), .ZN(n7588) );
  NAND2_X1 U9283 ( .A1(n7588), .A2(n8042), .ZN(n7938) );
  NAND3_X1 U9284 ( .A1(n7997), .A2(n9814), .A3(n7874), .ZN(n7582) );
  OAI21_X1 U9285 ( .B1(n7874), .B2(n8086), .A(n7582), .ZN(n7585) );
  NAND3_X1 U9286 ( .A1(n7997), .A2(n7914), .A3(n7877), .ZN(n7583) );
  OAI211_X1 U9287 ( .C1(n7877), .C2(n8086), .A(n7822), .B(n7583), .ZN(n7584)
         );
  OAI21_X1 U9288 ( .B1(n7822), .B2(n7585), .A(n7584), .ZN(n7586) );
  INV_X1 U9289 ( .A(n7588), .ZN(n7589) );
  NAND2_X1 U9290 ( .A1(n7589), .A2(n8353), .ZN(n7939) );
  NAND2_X1 U9291 ( .A1(n7590), .A2(n7939), .ZN(n8017) );
  XNOR2_X1 U9292 ( .A(n8533), .B(n7877), .ZN(n7591) );
  XNOR2_X1 U9293 ( .A(n7591), .B(n8337), .ZN(n8018) );
  XNOR2_X1 U9294 ( .A(n7592), .B(n8076), .ZN(n7894) );
  XNOR2_X1 U9295 ( .A(n8522), .B(n7877), .ZN(n7593) );
  XNOR2_X1 U9296 ( .A(n7593), .B(n8338), .ZN(n8068) );
  XNOR2_X1 U9297 ( .A(n8515), .B(n7877), .ZN(n7960) );
  NAND2_X1 U9298 ( .A1(n7962), .A2(n7596), .ZN(n7972) );
  NAND2_X1 U9299 ( .A1(n7960), .A2(n8329), .ZN(n7971) );
  XNOR2_X1 U9300 ( .A(n8509), .B(n7874), .ZN(n7598) );
  INV_X1 U9301 ( .A(n7598), .ZN(n7597) );
  INV_X1 U9302 ( .A(n7963), .ZN(n8318) );
  NAND2_X1 U9303 ( .A1(n7597), .A2(n8318), .ZN(n7970) );
  AND2_X1 U9304 ( .A1(n7971), .A2(n7970), .ZN(n7600) );
  NAND2_X1 U9305 ( .A1(n7598), .A2(n7963), .ZN(n7969) );
  AOI21_X2 U9306 ( .B1(n7972), .B2(n7600), .A(n7599), .ZN(n8048) );
  XNOR2_X1 U9307 ( .A(n7601), .B(n7874), .ZN(n7602) );
  XNOR2_X1 U9308 ( .A(n7602), .B(n8307), .ZN(n8049) );
  XNOR2_X1 U9309 ( .A(n8498), .B(n7874), .ZN(n7607) );
  XNOR2_X1 U9310 ( .A(n7607), .B(n8050), .ZN(n7915) );
  XNOR2_X1 U9311 ( .A(n7603), .B(n7874), .ZN(n7606) );
  INV_X1 U9312 ( .A(n7606), .ZN(n7604) );
  AND2_X1 U9313 ( .A1(n7604), .A2(n7920), .ZN(n7610) );
  OR2_X1 U9314 ( .A1(n7915), .A2(n7610), .ZN(n7605) );
  NOR2_X2 U9315 ( .A1(n7916), .A2(n7605), .ZN(n7612) );
  XNOR2_X1 U9316 ( .A(n7606), .B(n8284), .ZN(n8010) );
  INV_X1 U9317 ( .A(n8010), .ZN(n7609) );
  INV_X1 U9318 ( .A(n7607), .ZN(n7608) );
  INV_X1 U9319 ( .A(n8050), .ZN(n8294) );
  NAND2_X1 U9320 ( .A1(n7608), .A2(n8294), .ZN(n8006) );
  AND2_X1 U9321 ( .A1(n7609), .A2(n8006), .ZN(n8007) );
  NOR2_X1 U9322 ( .A1(n7610), .A2(n8007), .ZN(n7611) );
  XOR2_X1 U9323 ( .A(n7855), .B(n7854), .Z(n7617) );
  OAI22_X1 U9324 ( .A1(n7856), .A2(n8061), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10107), .ZN(n7613) );
  AOI21_X1 U9325 ( .B1(n8058), .B2(n8284), .A(n7613), .ZN(n7614) );
  OAI21_X1 U9326 ( .B1(n8053), .B2(n8266), .A(n7614), .ZN(n7615) );
  AOI21_X1 U9327 ( .B1(n8486), .B2(n8064), .A(n7615), .ZN(n7616) );
  OAI21_X1 U9328 ( .B1(n7617), .B2(n8067), .A(n7616), .ZN(P2_U3163) );
  INV_X1 U9329 ( .A(n7775), .ZN(n8544) );
  OAI222_X1 U9330 ( .A1(n7620), .A2(n7619), .B1(n7569), .B2(n8544), .C1(
        P1_U3086), .C2(n7618), .ZN(P1_U3325) );
  MUX2_X1 U9331 ( .A(n9227), .B(P1_DATAO_REG_31__SCAN_IN), .S(n5523), .Z(n7622) );
  NAND2_X1 U9332 ( .A1(n7622), .A2(n7621), .ZN(n8384) );
  INV_X1 U9333 ( .A(n8384), .ZN(n8434) );
  INV_X1 U9334 ( .A(n7755), .ZN(n7623) );
  INV_X1 U9335 ( .A(n8462), .ZN(n8219) );
  MUX2_X1 U9336 ( .A(n7866), .B(n8219), .S(n7783), .Z(n7750) );
  NAND2_X1 U9337 ( .A1(n7750), .A2(n8213), .ZN(n7625) );
  OAI22_X1 U9338 ( .A1(n8204), .A2(n7625), .B1(n7769), .B2(n7755), .ZN(n7626)
         );
  NOR2_X1 U9339 ( .A1(n7626), .A2(n7831), .ZN(n7768) );
  NAND2_X1 U9340 ( .A1(n7633), .A2(n6612), .ZN(n7628) );
  NAND2_X1 U9341 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  NAND2_X1 U9342 ( .A1(n7629), .A2(n7783), .ZN(n7635) );
  INV_X1 U9343 ( .A(n7630), .ZN(n7631) );
  OAI21_X1 U9344 ( .B1(n7635), .B2(n7631), .A(n6240), .ZN(n7632) );
  MUX2_X1 U9345 ( .A(n7632), .B(n6240), .S(n7769), .Z(n7637) );
  NAND3_X1 U9346 ( .A1(n7635), .A2(n7634), .A3(n7633), .ZN(n7636) );
  NAND3_X1 U9347 ( .A1(n7637), .A2(n9757), .A3(n7636), .ZN(n7644) );
  NAND2_X1 U9348 ( .A1(n7638), .A2(n7646), .ZN(n7641) );
  NAND2_X1 U9349 ( .A1(n9759), .A2(n9783), .ZN(n7655) );
  NAND2_X1 U9350 ( .A1(n7655), .A2(n7639), .ZN(n7640) );
  MUX2_X1 U9351 ( .A(n7641), .B(n7640), .S(n7769), .Z(n7642) );
  INV_X1 U9352 ( .A(n7642), .ZN(n7643) );
  NAND2_X1 U9353 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  NAND2_X1 U9354 ( .A1(n7645), .A2(n7810), .ZN(n7660) );
  INV_X1 U9355 ( .A(n7646), .ZN(n7650) );
  NAND2_X1 U9356 ( .A1(n7652), .A2(n7647), .ZN(n7662) );
  INV_X1 U9357 ( .A(n7662), .ZN(n7649) );
  OAI211_X1 U9358 ( .C1(n7660), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7654)
         );
  NAND2_X1 U9359 ( .A1(n7661), .A2(n7651), .ZN(n7656) );
  NAND2_X1 U9360 ( .A1(n7656), .A2(n7652), .ZN(n7653) );
  AOI21_X1 U9361 ( .B1(n7654), .B2(n7653), .A(n7665), .ZN(n7669) );
  INV_X1 U9362 ( .A(n7655), .ZN(n7659) );
  INV_X1 U9363 ( .A(n7656), .ZN(n7658) );
  OAI211_X1 U9364 ( .C1(n7660), .C2(n7659), .A(n7658), .B(n7657), .ZN(n7664)
         );
  NAND2_X1 U9365 ( .A1(n7662), .A2(n7661), .ZN(n7663) );
  NAND2_X1 U9366 ( .A1(n7664), .A2(n7663), .ZN(n7666) );
  INV_X1 U9367 ( .A(n7665), .ZN(n7818) );
  INV_X1 U9368 ( .A(n7676), .ZN(n7671) );
  MUX2_X1 U9369 ( .A(n7671), .B(n7670), .S(n7769), .Z(n7673) );
  INV_X1 U9370 ( .A(n7819), .ZN(n7672) );
  MUX2_X1 U9371 ( .A(n7679), .B(n7678), .S(n7783), .Z(n7680) );
  NAND3_X1 U9372 ( .A1(n7685), .A2(n7682), .A3(n7688), .ZN(n7683) );
  NAND2_X1 U9373 ( .A1(n7683), .A2(n7686), .ZN(n7691) );
  INV_X1 U9374 ( .A(n7686), .ZN(n7687) );
  INV_X1 U9375 ( .A(n8364), .ZN(n8366) );
  INV_X1 U9376 ( .A(n7692), .ZN(n7694) );
  NOR2_X1 U9377 ( .A1(n8351), .A2(n7769), .ZN(n7706) );
  NAND2_X1 U9378 ( .A1(n8527), .A2(n7706), .ZN(n7699) );
  NAND2_X1 U9379 ( .A1(n8351), .A2(n7769), .ZN(n7708) );
  OR2_X1 U9380 ( .A1(n8527), .A2(n7708), .ZN(n7698) );
  MUX2_X1 U9381 ( .A(n7696), .B(n7695), .S(n7769), .Z(n7697) );
  AND4_X1 U9382 ( .A1(n8359), .A2(n7699), .A3(n7698), .A4(n7697), .ZN(n7701)
         );
  OR2_X2 U9383 ( .A1(n5022), .A2(n7700), .ZN(n8327) );
  INV_X1 U9384 ( .A(n8317), .ZN(n7718) );
  MUX2_X1 U9385 ( .A(n7705), .B(n7704), .S(n7769), .Z(n7712) );
  INV_X1 U9386 ( .A(n7706), .ZN(n7707) );
  NAND2_X1 U9387 ( .A1(n8527), .A2(n7707), .ZN(n7711) );
  INV_X1 U9388 ( .A(n7708), .ZN(n7709) );
  OR2_X1 U9389 ( .A1(n8527), .A2(n7709), .ZN(n7710) );
  AOI22_X1 U9390 ( .A1(n8346), .A2(n7712), .B1(n7711), .B2(n7710), .ZN(n7716)
         );
  OAI21_X1 U9391 ( .B1(n8338), .B2(n7783), .A(n8522), .ZN(n7715) );
  AND2_X1 U9392 ( .A1(n8338), .A2(n7783), .ZN(n7713) );
  OR2_X1 U9393 ( .A1(n8522), .A2(n7713), .ZN(n7714) );
  AOI22_X1 U9394 ( .A1(n8327), .A2(n7716), .B1(n7715), .B2(n7714), .ZN(n7717)
         );
  INV_X1 U9395 ( .A(n8305), .ZN(n8303) );
  INV_X1 U9396 ( .A(n7719), .ZN(n7720) );
  NOR2_X1 U9397 ( .A1(n7725), .A2(n7720), .ZN(n7727) );
  INV_X1 U9398 ( .A(n7721), .ZN(n7722) );
  NOR2_X1 U9399 ( .A1(n7809), .A2(n7722), .ZN(n7723) );
  OAI21_X1 U9400 ( .B1(n7725), .B2(n7724), .A(n7723), .ZN(n7726) );
  MUX2_X1 U9401 ( .A(n7727), .B(n7726), .S(n7783), .Z(n7739) );
  NAND3_X1 U9402 ( .A1(n7739), .A2(n7740), .A3(n7807), .ZN(n7728) );
  NAND3_X1 U9403 ( .A1(n7728), .A2(n7743), .A3(n7736), .ZN(n7730) );
  NAND2_X1 U9404 ( .A1(n7730), .A2(n7729), .ZN(n7734) );
  MUX2_X1 U9405 ( .A(n7731), .B(n7742), .S(n7783), .Z(n7732) );
  INV_X1 U9406 ( .A(n7732), .ZN(n7733) );
  NOR2_X1 U9407 ( .A1(n8250), .A2(n7733), .ZN(n7747) );
  AOI22_X1 U9408 ( .A1(n7734), .A2(n7747), .B1(n7856), .B2(n8480), .ZN(n7748)
         );
  NAND2_X1 U9409 ( .A1(n7807), .A2(n7735), .ZN(n7738) );
  INV_X1 U9410 ( .A(n7809), .ZN(n7737) );
  OAI211_X1 U9411 ( .C1(n7739), .C2(n7738), .A(n7737), .B(n7736), .ZN(n7741)
         );
  NAND3_X1 U9412 ( .A1(n7741), .A2(n8257), .A3(n7740), .ZN(n7744) );
  NAND2_X1 U9413 ( .A1(n6259), .A2(n7745), .ZN(n7746) );
  NAND2_X1 U9414 ( .A1(n7754), .A2(n6259), .ZN(n7752) );
  NAND2_X1 U9415 ( .A1(n7803), .A2(n7783), .ZN(n7749) );
  NOR2_X1 U9416 ( .A1(n7759), .A2(n7749), .ZN(n7751) );
  INV_X1 U9417 ( .A(n7750), .ZN(n7761) );
  NAND2_X1 U9418 ( .A1(n7761), .A2(n7760), .ZN(n7756) );
  NAND3_X1 U9419 ( .A1(n7752), .A2(n7751), .A3(n7756), .ZN(n7767) );
  NAND2_X1 U9420 ( .A1(n7754), .A2(n7753), .ZN(n7758) );
  AND4_X1 U9421 ( .A1(n7756), .A2(n7769), .A3(n7755), .A4(n7804), .ZN(n7757)
         );
  NAND2_X1 U9422 ( .A1(n7758), .A2(n7757), .ZN(n7766) );
  XNOR2_X1 U9423 ( .A(n7759), .B(n7769), .ZN(n7764) );
  NAND2_X1 U9424 ( .A1(n7804), .A2(n7783), .ZN(n7763) );
  NAND3_X1 U9425 ( .A1(n7761), .A2(n7783), .A3(n7760), .ZN(n7762) );
  NAND3_X1 U9426 ( .A1(n7764), .A2(n7763), .A3(n7762), .ZN(n7765) );
  NAND4_X1 U9427 ( .A1(n7768), .A2(n7767), .A3(n7766), .A4(n7765), .ZN(n7771)
         );
  MUX2_X1 U9428 ( .A(n8188), .B(n8190), .S(n7769), .Z(n7770) );
  NAND2_X1 U9429 ( .A1(n7771), .A2(n7770), .ZN(n7773) );
  NAND2_X1 U9430 ( .A1(n7775), .A2(n7774), .ZN(n7777) );
  OR2_X1 U9431 ( .A1(n5864), .A2(n10086), .ZN(n7776) );
  NAND2_X1 U9432 ( .A1(n7777), .A2(n7776), .ZN(n8437) );
  INV_X1 U9433 ( .A(n8083), .ZN(n7778) );
  OR2_X1 U9434 ( .A1(n8437), .A2(n7778), .ZN(n7832) );
  AND2_X1 U9435 ( .A1(n8437), .A2(n7778), .ZN(n7794) );
  INV_X1 U9436 ( .A(n7794), .ZN(n7780) );
  OAI211_X1 U9437 ( .C1(n7802), .C2(n7781), .A(n7795), .B(n7780), .ZN(n7782)
         );
  INV_X1 U9438 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9439 ( .A1(n5869), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7786) );
  INV_X1 U9440 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9955) );
  OR2_X1 U9441 ( .A1(n5931), .A2(n9955), .ZN(n7785) );
  OAI211_X1 U9442 ( .C1(n7787), .C2(n4416), .A(n7786), .B(n7785), .ZN(n7788)
         );
  INV_X1 U9443 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U9444 ( .A1(n7790), .A2(n7789), .ZN(n8173) );
  NAND3_X1 U9445 ( .A1(n7838), .A2(n7832), .A3(n8173), .ZN(n7839) );
  INV_X1 U9446 ( .A(n7791), .ZN(n7792) );
  AOI21_X1 U9447 ( .B1(n8384), .B2(n8173), .A(n7794), .ZN(n7834) );
  INV_X1 U9448 ( .A(n8437), .ZN(n8178) );
  INV_X1 U9449 ( .A(n7795), .ZN(n7797) );
  XNOR2_X1 U9450 ( .A(n8443), .B(n7888), .ZN(n8194) );
  INV_X1 U9451 ( .A(n8224), .ZN(n7805) );
  NOR2_X1 U9452 ( .A1(n7806), .A2(n7805), .ZN(n8238) );
  INV_X1 U9453 ( .A(n7807), .ZN(n7808) );
  NOR2_X1 U9454 ( .A1(n7809), .A2(n7808), .ZN(n8292) );
  INV_X1 U9455 ( .A(n7810), .ZN(n7812) );
  NOR4_X1 U9456 ( .A1(n6241), .A2(n7812), .A3(n7811), .A4(n6239), .ZN(n7816)
         );
  AND4_X1 U9457 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n7820)
         );
  NAND4_X1 U9458 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n7823)
         );
  NOR3_X1 U9459 ( .A1(n7823), .A2(n7822), .A3(n7821), .ZN(n7824) );
  NAND4_X1 U9460 ( .A1(n7824), .A2(n8364), .A3(n8346), .A4(n8359), .ZN(n7826)
         );
  INV_X1 U9461 ( .A(n8327), .ZN(n7825) );
  NOR4_X1 U9462 ( .A1(n8305), .A2(n7826), .A3(n8317), .A4(n7825), .ZN(n7827)
         );
  NAND4_X1 U9463 ( .A1(n8272), .A2(n8282), .A3(n8292), .A4(n7827), .ZN(n7828)
         );
  NOR3_X1 U9464 ( .A1(n8250), .A2(n8260), .A3(n7828), .ZN(n7829) );
  NAND4_X1 U9465 ( .A1(n8211), .A2(n8227), .A3(n8238), .A4(n7829), .ZN(n7830)
         );
  NOR4_X1 U9466 ( .A1(n8194), .A2(n8204), .A3(n7831), .A4(n7830), .ZN(n7833)
         );
  NAND4_X1 U9467 ( .A1(n7834), .A2(n4581), .A3(n7833), .A4(n7832), .ZN(n7836)
         );
  NAND2_X1 U9468 ( .A1(n7836), .A2(n7835), .ZN(n7837) );
  XNOR2_X1 U9469 ( .A(n7841), .B(n7840), .ZN(n7848) );
  NAND3_X1 U9470 ( .A1(n7843), .A2(n7842), .A3(n8151), .ZN(n7844) );
  OAI211_X1 U9471 ( .C1(n7845), .C2(n7847), .A(n7844), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7846) );
  OAI21_X1 U9472 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(P2_U3296) );
  INV_X1 U9473 ( .A(n7849), .ZN(n8549) );
  OAI222_X1 U9474 ( .A1(n7569), .A2(n8549), .B1(n5780), .B2(P1_U3086), .C1(
        n7850), .C2(n7620), .ZN(P1_U3327) );
  INV_X1 U9475 ( .A(n7851), .ZN(n7852) );
  AOI22_X1 U9476 ( .A1(n7855), .A2(n7854), .B1(n7853), .B2(n7852), .ZN(n8026)
         );
  XNOR2_X1 U9477 ( .A(n8480), .B(n7877), .ZN(n7857) );
  XNOR2_X1 U9478 ( .A(n7857), .B(n7856), .ZN(n8025) );
  NAND2_X1 U9479 ( .A1(n7857), .A2(n8264), .ZN(n7858) );
  XNOR2_X1 U9480 ( .A(n8231), .B(n7877), .ZN(n7985) );
  XNOR2_X1 U9481 ( .A(n8474), .B(n7874), .ZN(n7861) );
  OAI22_X1 U9482 ( .A1(n7985), .A2(n7984), .B1(n8028), .B2(n7861), .ZN(n7859)
         );
  INV_X1 U9483 ( .A(n7859), .ZN(n7860) );
  OAI21_X1 U9484 ( .B1(n7982), .B2(n8251), .A(n8239), .ZN(n7863) );
  NOR3_X1 U9485 ( .A1(n7982), .A2(n8239), .A3(n8251), .ZN(n7862) );
  AOI21_X1 U9486 ( .B1(n7985), .B2(n7863), .A(n7862), .ZN(n7864) );
  XNOR2_X1 U9487 ( .A(n8462), .B(n7877), .ZN(n7867) );
  XNOR2_X1 U9488 ( .A(n7867), .B(n7866), .ZN(n7952) );
  NOR2_X1 U9489 ( .A1(n7867), .A2(n8229), .ZN(n7868) );
  XNOR2_X1 U9490 ( .A(n8457), .B(n7874), .ZN(n7869) );
  XNOR2_X1 U9491 ( .A(n7871), .B(n7869), .ZN(n8057) );
  NAND2_X1 U9492 ( .A1(n8057), .A2(n7955), .ZN(n7873) );
  INV_X1 U9493 ( .A(n7869), .ZN(n7870) );
  OR2_X1 U9494 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  NAND2_X1 U9495 ( .A1(n7873), .A2(n7872), .ZN(n7883) );
  XNOR2_X1 U9496 ( .A(n7892), .B(n7874), .ZN(n7875) );
  NAND2_X1 U9497 ( .A1(n7875), .A2(n8205), .ZN(n7876) );
  OAI21_X1 U9498 ( .B1(n7875), .B2(n8205), .A(n7876), .ZN(n7884) );
  XNOR2_X1 U9499 ( .A(n8194), .B(n7877), .ZN(n7878) );
  AOI22_X1 U9500 ( .A1(n8205), .A2(n8058), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7880) );
  NAND2_X1 U9501 ( .A1(n8199), .A2(n8078), .ZN(n7879) );
  OAI211_X1 U9502 ( .C1(n8084), .C2(n8061), .A(n7880), .B(n7879), .ZN(n7881)
         );
  AOI21_X1 U9503 ( .B1(n8443), .B2(n8064), .A(n7881), .ZN(n7882) );
  AOI21_X1 U9504 ( .B1(n7883), .B2(n7884), .A(n8067), .ZN(n7886) );
  AOI22_X1 U9505 ( .A1(n8215), .A2(n8058), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7887) );
  OAI21_X1 U9506 ( .B1(n7888), .B2(n8061), .A(n7887), .ZN(n7889) );
  AOI21_X1 U9507 ( .B1(n7890), .B2(n8078), .A(n7889), .ZN(n7891) );
  XOR2_X1 U9508 ( .A(n7893), .B(n7894), .Z(n7899) );
  AOI22_X1 U9509 ( .A1(n8073), .A2(n8338), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7896) );
  NAND2_X1 U9510 ( .A1(n8058), .A2(n8337), .ZN(n7895) );
  OAI211_X1 U9511 ( .C1(n8053), .C2(n8340), .A(n7896), .B(n7895), .ZN(n7897)
         );
  AOI21_X1 U9512 ( .B1(n8527), .B2(n8064), .A(n7897), .ZN(n7898) );
  OAI21_X1 U9513 ( .B1(n7899), .B2(n8067), .A(n7898), .ZN(P2_U3155) );
  XNOR2_X1 U9514 ( .A(n7981), .B(n7982), .ZN(n7983) );
  XNOR2_X1 U9515 ( .A(n7983), .B(n8028), .ZN(n7904) );
  NAND2_X1 U9516 ( .A1(n8078), .A2(n8242), .ZN(n7901) );
  AOI22_X1 U9517 ( .A1(n8058), .A2(n8264), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7900) );
  OAI211_X1 U9518 ( .C1(n7984), .C2(n8061), .A(n7901), .B(n7900), .ZN(n7902)
         );
  AOI21_X1 U9519 ( .B1(n8474), .B2(n8064), .A(n7902), .ZN(n7903) );
  OAI21_X1 U9520 ( .B1(n7904), .B2(n8067), .A(n7903), .ZN(P2_U3156) );
  XNOR2_X1 U9521 ( .A(n7940), .B(n7997), .ZN(n7906) );
  NAND2_X1 U9522 ( .A1(n7906), .A2(n7905), .ZN(n8036) );
  OAI21_X1 U9523 ( .B1(n7906), .B2(n7905), .A(n8036), .ZN(n7907) );
  NAND2_X1 U9524 ( .A1(n7907), .A2(n4824), .ZN(n7913) );
  INV_X1 U9525 ( .A(n7908), .ZN(n7911) );
  INV_X1 U9526 ( .A(n8086), .ZN(n8371) );
  NAND2_X1 U9527 ( .A1(n8058), .A2(n8088), .ZN(n7909) );
  INV_X1 U9528 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10160) );
  OR2_X1 U9529 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10160), .ZN(n9643) );
  OAI211_X1 U9530 ( .C1(n8371), .C2(n8061), .A(n7909), .B(n9643), .ZN(n7910)
         );
  AOI21_X1 U9531 ( .B1(n7911), .B2(n8078), .A(n7910), .ZN(n7912) );
  OAI211_X1 U9532 ( .C1(n7914), .C2(n8081), .A(n7913), .B(n7912), .ZN(P2_U3157) );
  AOI21_X1 U9533 ( .B1(n7916), .B2(n7915), .A(n8067), .ZN(n7917) );
  OR2_X1 U9534 ( .A1(n7916), .A2(n7915), .ZN(n8008) );
  NAND2_X1 U9535 ( .A1(n7917), .A2(n8008), .ZN(n7923) );
  INV_X1 U9536 ( .A(n7918), .ZN(n8287) );
  NAND2_X1 U9537 ( .A1(n8307), .A2(n8058), .ZN(n7919) );
  NAND2_X1 U9538 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U9539 ( .C1(n7920), .C2(n8061), .A(n7919), .B(n8163), .ZN(n7921)
         );
  AOI21_X1 U9540 ( .B1(n8287), .B2(n8078), .A(n7921), .ZN(n7922) );
  OAI211_X1 U9541 ( .C1(n7924), .C2(n8081), .A(n7923), .B(n7922), .ZN(P2_U3159) );
  OAI21_X1 U9542 ( .B1(n7927), .B2(n7926), .A(n7925), .ZN(n7928) );
  NAND2_X1 U9543 ( .A1(n7928), .A2(n4824), .ZN(n7937) );
  INV_X1 U9544 ( .A(n7929), .ZN(n7935) );
  NAND2_X1 U9545 ( .A1(n8058), .A2(n8090), .ZN(n7932) );
  INV_X1 U9546 ( .A(n7930), .ZN(n7931) );
  OAI211_X1 U9547 ( .C1(n7933), .C2(n8061), .A(n7932), .B(n7931), .ZN(n7934)
         );
  AOI21_X1 U9548 ( .B1(n7935), .B2(n8078), .A(n7934), .ZN(n7936) );
  OAI211_X1 U9549 ( .C1(n9804), .C2(n8081), .A(n7937), .B(n7936), .ZN(P2_U3161) );
  NAND2_X1 U9550 ( .A1(n7939), .A2(n7938), .ZN(n7943) );
  INV_X1 U9551 ( .A(n7940), .ZN(n7941) );
  NAND2_X1 U9552 ( .A1(n7941), .A2(n7997), .ZN(n8035) );
  NAND3_X1 U9553 ( .A1(n8036), .A2(n8034), .A3(n8035), .ZN(n8033) );
  OAI21_X1 U9554 ( .B1(n8371), .B2(n8034), .A(n8033), .ZN(n7942) );
  XOR2_X1 U9555 ( .A(n7943), .B(n7942), .Z(n7950) );
  INV_X1 U9556 ( .A(n8374), .ZN(n7944) );
  NAND2_X1 U9557 ( .A1(n8078), .A2(n7944), .ZN(n7947) );
  NOR2_X1 U9558 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7945), .ZN(n9670) );
  AOI21_X1 U9559 ( .B1(n8058), .B2(n8086), .A(n9670), .ZN(n7946) );
  OAI211_X1 U9560 ( .C1(n8369), .C2(n8061), .A(n7947), .B(n7946), .ZN(n7948)
         );
  AOI21_X1 U9561 ( .B1(n9831), .B2(n8064), .A(n7948), .ZN(n7949) );
  OAI21_X1 U9562 ( .B1(n7950), .B2(n8067), .A(n7949), .ZN(P2_U3164) );
  XOR2_X1 U9563 ( .A(n7952), .B(n7951), .Z(n7958) );
  AOI22_X1 U9564 ( .A1(n8239), .A2(n8058), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7954) );
  NAND2_X1 U9565 ( .A1(n8078), .A2(n8217), .ZN(n7953) );
  OAI211_X1 U9566 ( .C1(n7955), .C2(n8061), .A(n7954), .B(n7953), .ZN(n7956)
         );
  AOI21_X1 U9567 ( .B1(n8462), .B2(n8064), .A(n7956), .ZN(n7957) );
  OAI21_X1 U9568 ( .B1(n7958), .B2(n8067), .A(n7957), .ZN(P2_U3165) );
  XNOR2_X1 U9569 ( .A(n7960), .B(n7959), .ZN(n7961) );
  XNOR2_X1 U9570 ( .A(n7962), .B(n7961), .ZN(n7968) );
  AND2_X1 U9571 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9724) );
  NOR2_X1 U9572 ( .A1(n7963), .A2(n8061), .ZN(n7964) );
  AOI211_X1 U9573 ( .C1(n8058), .C2(n8338), .A(n9724), .B(n7964), .ZN(n7965)
         );
  OAI21_X1 U9574 ( .B1(n8322), .B2(n8053), .A(n7965), .ZN(n7966) );
  AOI21_X1 U9575 ( .B1(n8515), .B2(n8064), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9576 ( .B1(n7968), .B2(n8067), .A(n7967), .ZN(P2_U3166) );
  NAND2_X1 U9577 ( .A1(n7970), .A2(n7969), .ZN(n7974) );
  NAND2_X1 U9578 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  XOR2_X1 U9579 ( .A(n7974), .B(n7973), .Z(n7980) );
  AND2_X1 U9580 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9739) );
  NOR2_X1 U9581 ( .A1(n7975), .A2(n8061), .ZN(n7976) );
  AOI211_X1 U9582 ( .C1(n8058), .C2(n8329), .A(n9739), .B(n7976), .ZN(n7977)
         );
  OAI21_X1 U9583 ( .B1(n8311), .B2(n8053), .A(n7977), .ZN(n7978) );
  AOI21_X1 U9584 ( .B1(n8509), .B2(n8064), .A(n7978), .ZN(n7979) );
  OAI21_X1 U9585 ( .B1(n7980), .B2(n8067), .A(n7979), .ZN(P2_U3168) );
  OAI22_X1 U9586 ( .A1(n7983), .A2(n8251), .B1(n7982), .B2(n7981), .ZN(n7987)
         );
  XNOR2_X1 U9587 ( .A(n7985), .B(n7984), .ZN(n7986) );
  XNOR2_X1 U9588 ( .A(n7987), .B(n7986), .ZN(n7992) );
  AOI22_X1 U9589 ( .A1(n8229), .A2(n8073), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7989) );
  NAND2_X1 U9590 ( .A1(n8078), .A2(n8233), .ZN(n7988) );
  OAI211_X1 U9591 ( .C1(n8028), .C2(n8075), .A(n7989), .B(n7988), .ZN(n7990)
         );
  AOI21_X1 U9592 ( .B1(n8468), .B2(n8064), .A(n7990), .ZN(n7991) );
  OAI21_X1 U9593 ( .B1(n7992), .B2(n8067), .A(n7991), .ZN(P2_U3169) );
  NAND2_X1 U9594 ( .A1(n8078), .A2(n7993), .ZN(n7996) );
  NAND2_X1 U9595 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9626) );
  INV_X1 U9596 ( .A(n9626), .ZN(n7994) );
  AOI21_X1 U9597 ( .B1(n8058), .B2(n8089), .A(n7994), .ZN(n7995) );
  OAI211_X1 U9598 ( .C1(n7997), .C2(n8061), .A(n7996), .B(n7995), .ZN(n8003)
         );
  INV_X1 U9599 ( .A(n7998), .ZN(n7999) );
  AOI211_X1 U9600 ( .C1(n8001), .C2(n8000), .A(n8067), .B(n7999), .ZN(n8002)
         );
  AOI211_X1 U9601 ( .C1(n8004), .C2(n8064), .A(n8003), .B(n8002), .ZN(n8005)
         );
  INV_X1 U9602 ( .A(n8005), .ZN(P2_U3171) );
  NAND2_X1 U9603 ( .A1(n8008), .A2(n8006), .ZN(n8009) );
  AOI21_X1 U9604 ( .B1(n8010), .B2(n8009), .A(n5029), .ZN(n8016) );
  INV_X1 U9605 ( .A(n8011), .ZN(n8277) );
  NAND2_X1 U9606 ( .A1(n8078), .A2(n8277), .ZN(n8013) );
  AOI22_X1 U9607 ( .A1(n8274), .A2(n8073), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8012) );
  OAI211_X1 U9608 ( .C1(n8050), .C2(n8075), .A(n8013), .B(n8012), .ZN(n8014)
         );
  AOI21_X1 U9609 ( .B1(n8492), .B2(n8064), .A(n8014), .ZN(n8015) );
  OAI21_X1 U9610 ( .B1(n8016), .B2(n8067), .A(n8015), .ZN(P2_U3173) );
  XOR2_X1 U9611 ( .A(n8017), .B(n8018), .Z(n8023) );
  AOI22_X1 U9612 ( .A1(n8058), .A2(n8353), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8020) );
  NAND2_X1 U9613 ( .A1(n8073), .A2(n8351), .ZN(n8019) );
  OAI211_X1 U9614 ( .C1(n8053), .C2(n8349), .A(n8020), .B(n8019), .ZN(n8021)
         );
  AOI21_X1 U9615 ( .B1(n8533), .B2(n8064), .A(n8021), .ZN(n8022) );
  OAI21_X1 U9616 ( .B1(n8023), .B2(n8067), .A(n8022), .ZN(P2_U3174) );
  INV_X1 U9617 ( .A(n8480), .ZN(n8032) );
  OAI211_X1 U9618 ( .C1(n8026), .C2(n8025), .A(n8024), .B(n4824), .ZN(n8031)
         );
  AOI22_X1 U9619 ( .A1(n8274), .A2(n8058), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8027) );
  OAI21_X1 U9620 ( .B1(n8028), .B2(n8061), .A(n8027), .ZN(n8029) );
  AOI21_X1 U9621 ( .B1(n8247), .B2(n8078), .A(n8029), .ZN(n8030) );
  OAI211_X1 U9622 ( .C1(n8032), .C2(n8081), .A(n8031), .B(n8030), .ZN(P2_U3175) );
  NAND2_X1 U9623 ( .A1(n8033), .A2(n4824), .ZN(n8047) );
  AOI21_X1 U9624 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8046) );
  INV_X1 U9625 ( .A(n8037), .ZN(n8038) );
  NAND2_X1 U9626 ( .A1(n8078), .A2(n8038), .ZN(n8041) );
  NAND2_X1 U9627 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9658) );
  INV_X1 U9628 ( .A(n9658), .ZN(n8039) );
  AOI21_X1 U9629 ( .B1(n8058), .B2(n8087), .A(n8039), .ZN(n8040) );
  OAI211_X1 U9630 ( .C1(n8042), .C2(n8061), .A(n8041), .B(n8040), .ZN(n8043)
         );
  AOI21_X1 U9631 ( .B1(n8044), .B2(n8064), .A(n8043), .ZN(n8045) );
  OAI21_X1 U9632 ( .B1(n8047), .B2(n8046), .A(n8045), .ZN(P2_U3176) );
  XOR2_X1 U9633 ( .A(n8049), .B(n8048), .Z(n8056) );
  INV_X1 U9634 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10100) );
  OAI22_X1 U9635 ( .A1(n8050), .A2(n8061), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10100), .ZN(n8051) );
  AOI21_X1 U9636 ( .B1(n8058), .B2(n8318), .A(n8051), .ZN(n8052) );
  OAI21_X1 U9637 ( .B1(n8053), .B2(n8297), .A(n8052), .ZN(n8054) );
  AOI21_X1 U9638 ( .B1(n8503), .B2(n8064), .A(n8054), .ZN(n8055) );
  OAI21_X1 U9639 ( .B1(n8056), .B2(n8067), .A(n8055), .ZN(P2_U3178) );
  XNOR2_X1 U9640 ( .A(n8057), .B(n8215), .ZN(n8066) );
  AOI22_X1 U9641 ( .A1(n8229), .A2(n8058), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8060) );
  NAND2_X1 U9642 ( .A1(n8078), .A2(n8208), .ZN(n8059) );
  OAI211_X1 U9643 ( .C1(n8062), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8063)
         );
  AOI21_X1 U9644 ( .B1(n8457), .B2(n8064), .A(n8063), .ZN(n8065) );
  OAI21_X1 U9645 ( .B1(n8066), .B2(n8067), .A(n8065), .ZN(P2_U3180) );
  INV_X1 U9646 ( .A(n8522), .ZN(n8082) );
  AOI21_X1 U9647 ( .B1(n8069), .B2(n8068), .A(n8067), .ZN(n8071) );
  NAND2_X1 U9648 ( .A1(n8071), .A2(n8070), .ZN(n8080) );
  INV_X1 U9649 ( .A(n8072), .ZN(n8332) );
  AND2_X1 U9650 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9711) );
  AOI21_X1 U9651 ( .B1(n8329), .B2(n8073), .A(n9711), .ZN(n8074) );
  OAI21_X1 U9652 ( .B1(n8076), .B2(n8075), .A(n8074), .ZN(n8077) );
  AOI21_X1 U9653 ( .B1(n8332), .B2(n8078), .A(n8077), .ZN(n8079) );
  OAI211_X1 U9654 ( .C1(n8082), .C2(n8081), .A(n8080), .B(n8079), .ZN(P2_U3181) );
  MUX2_X1 U9655 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8173), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9656 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8083), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U9657 ( .A(n8084), .ZN(n8196) );
  MUX2_X1 U9658 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8196), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9659 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8085), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9660 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8205), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9661 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8215), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9662 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8229), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9663 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8239), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9664 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8251), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9665 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8264), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9666 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8274), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9667 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8284), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9668 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8294), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9669 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8307), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9670 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8318), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8329), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9672 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8338), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9673 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8351), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9674 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8337), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9675 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8353), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9676 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8086), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9677 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8087), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9678 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8088), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9679 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8089), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9680 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8090), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9681 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8091), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9682 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8092), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9683 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8093), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9684 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9759), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9685 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n4415), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9686 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9760), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9687 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8286), .S(n8164), .Z(n8159)
         );
  AOI22_X1 U9688 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9738), .B1(n8147), .B2(
        n8321), .ZN(n9732) );
  OAI21_X1 U9689 ( .B1(n8108), .B2(n6980), .A(n8094), .ZN(n8095) );
  XNOR2_X1 U9690 ( .A(n8095), .B(n8128), .ZN(n9623) );
  MUX2_X1 U9691 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8096), .S(n9629), .Z(n9639)
         );
  NOR2_X1 U9692 ( .A1(n9646), .A2(n4452), .ZN(n8097) );
  XNOR2_X1 U9693 ( .A(n9646), .B(n4452), .ZN(n9655) );
  NOR2_X1 U9694 ( .A1(n5978), .A2(n9655), .ZN(n9654) );
  MUX2_X1 U9695 ( .A(n8375), .B(P2_REG2_REG_12__SCAN_IN), .S(n9661), .Z(n8098)
         );
  INV_X1 U9696 ( .A(n8098), .ZN(n9672) );
  NOR2_X1 U9697 ( .A1(n9673), .A2(n9672), .ZN(n9671) );
  NOR2_X1 U9698 ( .A1(n9679), .A2(n8099), .ZN(n8100) );
  XNOR2_X1 U9699 ( .A(n9679), .B(n8099), .ZN(n9688) );
  NOR2_X1 U9700 ( .A1(n6010), .A2(n9688), .ZN(n9687) );
  NOR2_X1 U9701 ( .A1(n8100), .A2(n9687), .ZN(n9704) );
  INV_X1 U9702 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8101) );
  AND2_X1 U9703 ( .A1(n9694), .A2(n8101), .ZN(n9702) );
  OAI22_X1 U9704 ( .A1(n9704), .A2(n9702), .B1(n9694), .B2(n8101), .ZN(n8102)
         );
  NAND2_X1 U9705 ( .A1(n9723), .A2(n8102), .ZN(n8103) );
  XNOR2_X1 U9706 ( .A(n8102), .B(n8141), .ZN(n9715) );
  NAND2_X1 U9707 ( .A1(n9753), .A2(n8104), .ZN(n8105) );
  XNOR2_X1 U9708 ( .A(n8104), .B(n8152), .ZN(n9744) );
  NAND2_X1 U9709 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n9744), .ZN(n9743) );
  INV_X1 U9710 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8296) );
  XNOR2_X1 U9711 ( .A(n10211), .B(n8296), .ZN(n10219) );
  OAI22_X1 U9712 ( .A1(n10218), .A2(n10219), .B1(n10211), .B2(n8296), .ZN(
        n8106) );
  XOR2_X1 U9713 ( .A(n8159), .B(n8106), .Z(n8171) );
  XNOR2_X1 U9714 ( .A(n8147), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9726) );
  AOI22_X1 U9715 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8122), .B1(n9661), .B2(
        n5993), .ZN(n9664) );
  AOI22_X1 U9716 ( .A1(n9629), .A2(n5963), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n8126), .ZN(n9632) );
  NAND2_X1 U9717 ( .A1(n8109), .A2(n8128), .ZN(n8110) );
  XNOR2_X1 U9718 ( .A(n8109), .B(n9614), .ZN(n9619) );
  NAND2_X1 U9719 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n9619), .ZN(n9618) );
  NAND2_X1 U9720 ( .A1(n8110), .A2(n9618), .ZN(n9631) );
  NAND2_X1 U9721 ( .A1(n9632), .A2(n9631), .ZN(n9630) );
  NAND2_X1 U9722 ( .A1(n8124), .A2(n8111), .ZN(n8112) );
  NAND2_X1 U9723 ( .A1(n8112), .A2(n9647), .ZN(n9663) );
  NAND2_X1 U9724 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  NAND2_X1 U9725 ( .A1(n8120), .A2(n8113), .ZN(n8114) );
  NAND2_X1 U9726 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9681), .ZN(n9680) );
  XNOR2_X1 U9727 ( .A(n9694), .B(n8425), .ZN(n9695) );
  NAND2_X1 U9728 ( .A1(n9723), .A2(n8115), .ZN(n8116) );
  XNOR2_X1 U9729 ( .A(n8115), .B(n8141), .ZN(n9713) );
  NAND2_X1 U9730 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9713), .ZN(n9712) );
  NAND2_X1 U9731 ( .A1(n8116), .A2(n9712), .ZN(n9727) );
  NAND2_X1 U9732 ( .A1(n9726), .A2(n9727), .ZN(n9725) );
  NAND2_X1 U9733 ( .A1(n9753), .A2(n8117), .ZN(n8118) );
  XNOR2_X1 U9734 ( .A(n10211), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n10203) );
  OAI21_X1 U9735 ( .B1(n10211), .B2(n8414), .A(n10202), .ZN(n8119) );
  XNOR2_X1 U9736 ( .A(n8164), .B(n9986), .ZN(n8160) );
  XNOR2_X1 U9737 ( .A(n8119), .B(n8160), .ZN(n8169) );
  MUX2_X1 U9738 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8151), .Z(n8156) );
  INV_X1 U9739 ( .A(n8156), .ZN(n10205) );
  MUX2_X1 U9740 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8151), .Z(n8140) );
  XNOR2_X1 U9741 ( .A(n8140), .B(n8141), .ZN(n9717) );
  MUX2_X1 U9742 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8151), .Z(n8139) );
  XNOR2_X1 U9743 ( .A(n8139), .B(n9694), .ZN(n9699) );
  MUX2_X1 U9744 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8145), .Z(n8121) );
  OR2_X1 U9745 ( .A1(n8121), .A2(n8120), .ZN(n8138) );
  XNOR2_X1 U9746 ( .A(n8121), .B(n9679), .ZN(n9684) );
  MUX2_X1 U9747 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8145), .Z(n8123) );
  OR2_X1 U9748 ( .A1(n8123), .A2(n8122), .ZN(n8137) );
  XNOR2_X1 U9749 ( .A(n8123), .B(n9661), .ZN(n9667) );
  MUX2_X1 U9750 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8151), .Z(n8125) );
  OR2_X1 U9751 ( .A1(n8125), .A2(n8124), .ZN(n8136) );
  XNOR2_X1 U9752 ( .A(n8125), .B(n9646), .ZN(n9651) );
  MUX2_X1 U9753 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8151), .Z(n8127) );
  OR2_X1 U9754 ( .A1(n8127), .A2(n8126), .ZN(n8135) );
  XNOR2_X1 U9755 ( .A(n8127), .B(n9629), .ZN(n9635) );
  MUX2_X1 U9756 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8151), .Z(n8129) );
  OR2_X1 U9757 ( .A1(n8129), .A2(n8128), .ZN(n8134) );
  XNOR2_X1 U9758 ( .A(n8129), .B(n9614), .ZN(n9616) );
  NAND2_X1 U9759 ( .A1(n9616), .A2(n9617), .ZN(n9615) );
  NAND2_X1 U9760 ( .A1(n8134), .A2(n9615), .ZN(n9634) );
  NAND2_X1 U9761 ( .A1(n9635), .A2(n9634), .ZN(n9633) );
  NAND2_X1 U9762 ( .A1(n8135), .A2(n9633), .ZN(n9650) );
  NAND2_X1 U9763 ( .A1(n9651), .A2(n9650), .ZN(n9649) );
  NAND2_X1 U9764 ( .A1(n8136), .A2(n9649), .ZN(n9666) );
  NAND2_X1 U9765 ( .A1(n9667), .A2(n9666), .ZN(n9665) );
  NAND2_X1 U9766 ( .A1(n8137), .A2(n9665), .ZN(n9683) );
  NAND2_X1 U9767 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  NAND2_X1 U9768 ( .A1(n8138), .A2(n9682), .ZN(n9698) );
  NAND2_X1 U9769 ( .A1(n9699), .A2(n9698), .ZN(n9697) );
  NAND2_X1 U9770 ( .A1(n9717), .A2(n9716), .ZN(n8144) );
  INV_X1 U9771 ( .A(n8140), .ZN(n8142) );
  NAND2_X1 U9772 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  NAND2_X1 U9773 ( .A1(n8144), .A2(n8143), .ZN(n9729) );
  MUX2_X1 U9774 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8151), .Z(n8146) );
  XNOR2_X1 U9775 ( .A(n8146), .B(n8147), .ZN(n9728) );
  NAND2_X1 U9776 ( .A1(n9729), .A2(n9728), .ZN(n8150) );
  INV_X1 U9777 ( .A(n8146), .ZN(n8148) );
  NAND2_X1 U9778 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U9779 ( .A1(n8150), .A2(n8149), .ZN(n9746) );
  MUX2_X1 U9780 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8151), .Z(n8153) );
  XNOR2_X1 U9781 ( .A(n8153), .B(n8152), .ZN(n9745) );
  NOR2_X1 U9782 ( .A1(n8153), .A2(n9753), .ZN(n8154) );
  OAI21_X1 U9783 ( .B1(n8156), .B2(n8155), .A(n10206), .ZN(n8157) );
  OAI21_X1 U9784 ( .B1(n10211), .B2(n10205), .A(n8157), .ZN(n8162) );
  MUX2_X1 U9785 ( .A(n8160), .B(n8159), .S(n8158), .Z(n8161) );
  XNOR2_X1 U9786 ( .A(n8162), .B(n8161), .ZN(n8167) );
  OAI21_X1 U9787 ( .B1(n9754), .B2(n8164), .A(n8163), .ZN(n8165) );
  AOI21_X1 U9788 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n9740), .A(n8165), .ZN(
        n8166) );
  OAI21_X1 U9789 ( .B1(n8167), .B2(n9597), .A(n8166), .ZN(n8168) );
  OAI21_X1 U9790 ( .B1(n8171), .B2(n10220), .A(n8170), .ZN(P2_U3201) );
  NOR2_X1 U9791 ( .A1(n8174), .A2(n8373), .ZN(n8183) );
  AOI21_X1 U9792 ( .B1(n8435), .B2(n8376), .A(n8183), .ZN(n8177) );
  NAND2_X1 U9793 ( .A1(n9773), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8175) );
  OAI211_X1 U9794 ( .C1(n8384), .C2(n8180), .A(n8177), .B(n8175), .ZN(P2_U3202) );
  NAND2_X1 U9795 ( .A1(n9773), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8176) );
  OAI211_X1 U9796 ( .C1(n8178), .C2(n8180), .A(n8177), .B(n8176), .ZN(P2_U3203) );
  NAND2_X1 U9797 ( .A1(n8179), .A2(n8376), .ZN(n8185) );
  NOR2_X1 U9798 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  AOI211_X1 U9799 ( .C1(n9773), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8183), .B(
        n8182), .ZN(n8184) );
  OAI211_X1 U9800 ( .C1(n8187), .C2(n8186), .A(n8185), .B(n8184), .ZN(P2_U3204) );
  NAND2_X1 U9801 ( .A1(n8189), .A2(n8188), .ZN(n8191) );
  NAND2_X1 U9802 ( .A1(n8191), .A2(n8190), .ZN(n8193) );
  INV_X1 U9803 ( .A(n8194), .ZN(n8192) );
  XNOR2_X1 U9804 ( .A(n8193), .B(n8192), .ZN(n8446) );
  XNOR2_X1 U9805 ( .A(n8195), .B(n8194), .ZN(n8197) );
  AOI222_X2 U9806 ( .A1(n8355), .A2(n8197), .B1(n8196), .B2(n9758), .C1(n8205), 
        .C2(n8352), .ZN(n8441) );
  MUX2_X1 U9807 ( .A(n8198), .B(n8441), .S(n8376), .Z(n8201) );
  AOI22_X1 U9808 ( .A1(n8443), .A2(n8378), .B1(n9768), .B2(n8199), .ZN(n8200)
         );
  OAI211_X1 U9809 ( .C1(n8446), .C2(n8381), .A(n8201), .B(n8200), .ZN(P2_U3205) );
  XNOR2_X1 U9810 ( .A(n8202), .B(n8204), .ZN(n8460) );
  INV_X1 U9811 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8207) );
  XNOR2_X1 U9812 ( .A(n8203), .B(n8204), .ZN(n8206) );
  AOI222_X1 U9813 ( .A1(n8355), .A2(n8206), .B1(n8229), .B2(n8352), .C1(n8205), 
        .C2(n9758), .ZN(n8455) );
  MUX2_X1 U9814 ( .A(n8207), .B(n8455), .S(n8376), .Z(n8210) );
  AOI22_X1 U9815 ( .A1(n8457), .A2(n8378), .B1(n9768), .B2(n8208), .ZN(n8209)
         );
  OAI211_X1 U9816 ( .C1(n8460), .C2(n8381), .A(n8210), .B(n8209), .ZN(P2_U3207) );
  XNOR2_X1 U9817 ( .A(n8212), .B(n8211), .ZN(n8465) );
  XNOR2_X1 U9818 ( .A(n8214), .B(n8213), .ZN(n8216) );
  AOI222_X1 U9819 ( .A1(n8355), .A2(n8216), .B1(n8239), .B2(n8352), .C1(n8215), 
        .C2(n9758), .ZN(n8461) );
  INV_X1 U9820 ( .A(n8461), .ZN(n8221) );
  INV_X1 U9821 ( .A(n8217), .ZN(n8218) );
  OAI22_X1 U9822 ( .A1(n8219), .A2(n8341), .B1(n8218), .B2(n8373), .ZN(n8220)
         );
  OAI21_X1 U9823 ( .B1(n8221), .B2(n8220), .A(n8376), .ZN(n8223) );
  NAND2_X1 U9824 ( .A1(n9773), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8222) );
  OAI211_X1 U9825 ( .C1(n8465), .C2(n8381), .A(n8223), .B(n8222), .ZN(P2_U3208) );
  NAND2_X1 U9826 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  XOR2_X1 U9827 ( .A(n8227), .B(n8226), .Z(n8471) );
  XNOR2_X1 U9828 ( .A(n8228), .B(n8227), .ZN(n8230) );
  AOI222_X1 U9829 ( .A1(n8355), .A2(n8230), .B1(n8251), .B2(n8352), .C1(n8229), 
        .C2(n9758), .ZN(n8466) );
  OAI21_X1 U9830 ( .B1(n8231), .B2(n8341), .A(n8466), .ZN(n8232) );
  NAND2_X1 U9831 ( .A1(n8232), .A2(n8376), .ZN(n8235) );
  AOI22_X1 U9832 ( .A1(n9773), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9768), .B2(
        n8233), .ZN(n8234) );
  OAI211_X1 U9833 ( .C1(n8471), .C2(n8381), .A(n8235), .B(n8234), .ZN(P2_U3209) );
  XNOR2_X1 U9834 ( .A(n8236), .B(n8238), .ZN(n8477) );
  INV_X1 U9835 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8241) );
  XOR2_X1 U9836 ( .A(n8238), .B(n8237), .Z(n8240) );
  AOI222_X1 U9837 ( .A1(n8355), .A2(n8240), .B1(n8239), .B2(n9758), .C1(n8264), 
        .C2(n8352), .ZN(n8472) );
  MUX2_X1 U9838 ( .A(n8241), .B(n8472), .S(n8376), .Z(n8244) );
  AOI22_X1 U9839 ( .A1(n8474), .A2(n8378), .B1(n9768), .B2(n8242), .ZN(n8243)
         );
  OAI211_X1 U9840 ( .C1(n8477), .C2(n8381), .A(n8244), .B(n8243), .ZN(P2_U3210) );
  XNOR2_X1 U9841 ( .A(n8246), .B(n8245), .ZN(n8483) );
  INV_X1 U9842 ( .A(n8247), .ZN(n8253) );
  OAI21_X1 U9843 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8252) );
  AOI222_X1 U9844 ( .A1(n8355), .A2(n8252), .B1(n8251), .B2(n9758), .C1(n8274), 
        .C2(n8352), .ZN(n8478) );
  OAI21_X1 U9845 ( .B1(n8253), .B2(n8373), .A(n8478), .ZN(n8254) );
  NAND2_X1 U9846 ( .A1(n8254), .A2(n8376), .ZN(n8256) );
  AOI22_X1 U9847 ( .A1(n8480), .A2(n8378), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n9773), .ZN(n8255) );
  OAI211_X1 U9848 ( .C1(n8483), .C2(n8381), .A(n8256), .B(n8255), .ZN(P2_U3211) );
  NAND2_X1 U9849 ( .A1(n8258), .A2(n8257), .ZN(n8259) );
  XNOR2_X1 U9850 ( .A(n8259), .B(n8260), .ZN(n8489) );
  OR3_X1 U9851 ( .A1(n4427), .A2(n8261), .A3(n8260), .ZN(n8262) );
  NAND2_X1 U9852 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  AOI222_X1 U9853 ( .A1(n8355), .A2(n8265), .B1(n8284), .B2(n8352), .C1(n8264), 
        .C2(n9758), .ZN(n8484) );
  OAI21_X1 U9854 ( .B1(n8266), .B2(n8373), .A(n8484), .ZN(n8267) );
  NAND2_X1 U9855 ( .A1(n8267), .A2(n8376), .ZN(n8269) );
  AOI22_X1 U9856 ( .A1(n8486), .A2(n8378), .B1(P2_REG2_REG_21__SCAN_IN), .B2(
        n9773), .ZN(n8268) );
  OAI211_X1 U9857 ( .C1(n8489), .C2(n8381), .A(n8269), .B(n8268), .ZN(P2_U3212) );
  XOR2_X1 U9858 ( .A(n8272), .B(n8270), .Z(n8495) );
  INV_X1 U9859 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8276) );
  AOI21_X1 U9860 ( .B1(n8272), .B2(n8271), .A(n4427), .ZN(n8273) );
  INV_X1 U9861 ( .A(n8273), .ZN(n8275) );
  AOI222_X1 U9862 ( .A1(n8355), .A2(n8275), .B1(n8274), .B2(n9758), .C1(n8294), 
        .C2(n8352), .ZN(n8490) );
  MUX2_X1 U9863 ( .A(n8276), .B(n8490), .S(n8376), .Z(n8279) );
  AOI22_X1 U9864 ( .A1(n8492), .A2(n8378), .B1(n9768), .B2(n8277), .ZN(n8278)
         );
  OAI211_X1 U9865 ( .C1(n8495), .C2(n8381), .A(n8279), .B(n8278), .ZN(P2_U3213) );
  OAI21_X1 U9866 ( .B1(n8281), .B2(n8282), .A(n8280), .ZN(n8499) );
  INV_X1 U9867 ( .A(n8499), .ZN(n8290) );
  XOR2_X1 U9868 ( .A(n8283), .B(n8282), .Z(n8285) );
  AOI222_X1 U9869 ( .A1(n8355), .A2(n8285), .B1(n8284), .B2(n9758), .C1(n8307), 
        .C2(n8352), .ZN(n8496) );
  MUX2_X1 U9870 ( .A(n8286), .B(n8496), .S(n8376), .Z(n8289) );
  AOI22_X1 U9871 ( .A1(n8498), .A2(n8378), .B1(n9768), .B2(n8287), .ZN(n8288)
         );
  OAI211_X1 U9872 ( .C1(n8290), .C2(n8381), .A(n8289), .B(n8288), .ZN(P2_U3214) );
  XOR2_X1 U9873 ( .A(n8291), .B(n8292), .Z(n8504) );
  INV_X1 U9874 ( .A(n8504), .ZN(n8301) );
  XNOR2_X1 U9875 ( .A(n8293), .B(n8292), .ZN(n8295) );
  AOI222_X1 U9876 ( .A1(n8355), .A2(n8295), .B1(n8318), .B2(n8352), .C1(n8294), 
        .C2(n9758), .ZN(n8502) );
  MUX2_X1 U9877 ( .A(n8296), .B(n8502), .S(n8376), .Z(n8300) );
  INV_X1 U9878 ( .A(n8297), .ZN(n8298) );
  AOI22_X1 U9879 ( .A1(n8503), .A2(n8378), .B1(n9768), .B2(n8298), .ZN(n8299)
         );
  OAI211_X1 U9880 ( .C1(n8301), .C2(n8381), .A(n8300), .B(n8299), .ZN(P2_U3215) );
  XNOR2_X1 U9881 ( .A(n8302), .B(n8303), .ZN(n8512) );
  OAI211_X1 U9882 ( .C1(n8306), .C2(n8305), .A(n8304), .B(n8355), .ZN(n8309)
         );
  AOI22_X1 U9883 ( .A1(n9758), .A2(n8307), .B1(n8329), .B2(n8352), .ZN(n8308)
         );
  MUX2_X1 U9884 ( .A(n8508), .B(n8310), .S(n9773), .Z(n8314) );
  INV_X1 U9885 ( .A(n8311), .ZN(n8312) );
  AOI22_X1 U9886 ( .A1(n8509), .A2(n8378), .B1(n9768), .B2(n8312), .ZN(n8313)
         );
  OAI211_X1 U9887 ( .C1(n8512), .C2(n8381), .A(n8314), .B(n8313), .ZN(P2_U3216) );
  XNOR2_X1 U9888 ( .A(n8315), .B(n8317), .ZN(n8519) );
  OAI211_X1 U9889 ( .C1(n4501), .C2(n8317), .A(n8316), .B(n8355), .ZN(n8320)
         );
  AOI22_X1 U9890 ( .A1(n8318), .A2(n9758), .B1(n8352), .B2(n8338), .ZN(n8319)
         );
  MUX2_X1 U9891 ( .A(n8514), .B(n8321), .S(n9773), .Z(n8325) );
  INV_X1 U9892 ( .A(n8322), .ZN(n8323) );
  AOI22_X1 U9893 ( .A1(n8515), .A2(n8378), .B1(n9768), .B2(n8323), .ZN(n8324)
         );
  OAI211_X1 U9894 ( .C1(n8519), .C2(n8381), .A(n8325), .B(n8324), .ZN(P2_U3217) );
  XNOR2_X1 U9895 ( .A(n8326), .B(n8327), .ZN(n8523) );
  INV_X1 U9896 ( .A(n8523), .ZN(n8335) );
  XNOR2_X1 U9897 ( .A(n8328), .B(n8327), .ZN(n8330) );
  AOI222_X1 U9898 ( .A1(n8355), .A2(n8330), .B1(n8329), .B2(n9758), .C1(n8351), 
        .C2(n8352), .ZN(n8520) );
  MUX2_X1 U9899 ( .A(n8331), .B(n8520), .S(n8376), .Z(n8334) );
  AOI22_X1 U9900 ( .A1(n8522), .A2(n8378), .B1(n9768), .B2(n8332), .ZN(n8333)
         );
  OAI211_X1 U9901 ( .C1(n8335), .C2(n8381), .A(n8334), .B(n8333), .ZN(P2_U3218) );
  XOR2_X1 U9902 ( .A(n8336), .B(n8346), .Z(n8339) );
  AOI222_X1 U9903 ( .A1(n8355), .A2(n8339), .B1(n8338), .B2(n9758), .C1(n8337), 
        .C2(n8352), .ZN(n8526) );
  INV_X1 U9904 ( .A(n8526), .ZN(n8344) );
  OAI22_X1 U9905 ( .A1(n8342), .A2(n8341), .B1(n8340), .B2(n8373), .ZN(n8343)
         );
  OAI21_X1 U9906 ( .B1(n8344), .B2(n8343), .A(n8376), .ZN(n8348) );
  XNOR2_X1 U9907 ( .A(n8345), .B(n8346), .ZN(n8528) );
  AOI22_X1 U9908 ( .A1(n8528), .A2(n8361), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9773), .ZN(n8347) );
  NAND2_X1 U9909 ( .A1(n8348), .A2(n8347), .ZN(P2_U3219) );
  NOR2_X1 U9910 ( .A1(n8373), .A2(n8349), .ZN(n8357) );
  XNOR2_X1 U9911 ( .A(n8350), .B(n8359), .ZN(n8354) );
  AOI222_X1 U9912 ( .A1(n8355), .A2(n8354), .B1(n8353), .B2(n8352), .C1(n8351), 
        .C2(n9758), .ZN(n8531) );
  INV_X1 U9913 ( .A(n8531), .ZN(n8356) );
  AOI211_X1 U9914 ( .C1(n8358), .C2(n8533), .A(n8357), .B(n8356), .ZN(n8363)
         );
  XNOR2_X1 U9915 ( .A(n8360), .B(n8359), .ZN(n8536) );
  AOI22_X1 U9916 ( .A1(n8536), .A2(n8361), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9773), .ZN(n8362) );
  OAI21_X1 U9917 ( .B1(n8363), .B2(n9773), .A(n8362), .ZN(P2_U3220) );
  XNOR2_X1 U9918 ( .A(n8365), .B(n8364), .ZN(n9828) );
  XNOR2_X1 U9919 ( .A(n8367), .B(n8366), .ZN(n8368) );
  OAI222_X1 U9920 ( .A1(n8372), .A2(n8371), .B1(n8370), .B2(n8369), .C1(n8368), 
        .C2(n9762), .ZN(n9829) );
  NAND2_X1 U9921 ( .A1(n9829), .A2(n8376), .ZN(n8380) );
  OAI22_X1 U9922 ( .A1(n8376), .A2(n8375), .B1(n8374), .B2(n8373), .ZN(n8377)
         );
  AOI21_X1 U9923 ( .B1(n8378), .B2(n9831), .A(n8377), .ZN(n8379) );
  OAI211_X1 U9924 ( .C1(n9828), .C2(n8381), .A(n8380), .B(n8379), .ZN(P2_U3221) );
  NAND2_X1 U9925 ( .A1(n9849), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U9926 ( .A1(n8435), .A2(n9851), .ZN(n8385) );
  OAI211_X1 U9927 ( .C1(n8384), .C2(n8383), .A(n8382), .B(n8385), .ZN(P2_U3490) );
  INV_X1 U9928 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U9929 ( .A1(n8437), .A2(n8428), .ZN(n8386) );
  OAI211_X1 U9930 ( .C1(n9851), .C2(n8387), .A(n8386), .B(n8385), .ZN(P2_U3489) );
  INV_X1 U9931 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8388) );
  MUX2_X1 U9932 ( .A(n8388), .B(n8441), .S(n9851), .Z(n8390) );
  NAND2_X1 U9933 ( .A1(n8443), .A2(n8428), .ZN(n8389) );
  OAI211_X1 U9934 ( .C1(n8446), .C2(n8422), .A(n8390), .B(n8389), .ZN(P2_U3487) );
  INV_X1 U9935 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8391) );
  MUX2_X1 U9936 ( .A(n8391), .B(n8455), .S(n9851), .Z(n8393) );
  NAND2_X1 U9937 ( .A1(n8457), .A2(n8428), .ZN(n8392) );
  OAI211_X1 U9938 ( .C1(n8422), .C2(n8460), .A(n8393), .B(n8392), .ZN(P2_U3485) );
  INV_X1 U9939 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8394) );
  MUX2_X1 U9940 ( .A(n8394), .B(n8461), .S(n9851), .Z(n8396) );
  NAND2_X1 U9941 ( .A1(n8462), .A2(n8428), .ZN(n8395) );
  OAI211_X1 U9942 ( .C1(n8422), .C2(n8465), .A(n8396), .B(n8395), .ZN(P2_U3484) );
  INV_X1 U9943 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8397) );
  MUX2_X1 U9944 ( .A(n8397), .B(n8466), .S(n9851), .Z(n8399) );
  NAND2_X1 U9945 ( .A1(n8468), .A2(n8428), .ZN(n8398) );
  OAI211_X1 U9946 ( .C1(n8422), .C2(n8471), .A(n8399), .B(n8398), .ZN(P2_U3483) );
  INV_X1 U9947 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8400) );
  MUX2_X1 U9948 ( .A(n8400), .B(n8472), .S(n9851), .Z(n8402) );
  NAND2_X1 U9949 ( .A1(n8474), .A2(n8428), .ZN(n8401) );
  OAI211_X1 U9950 ( .C1(n8477), .C2(n8422), .A(n8402), .B(n8401), .ZN(P2_U3482) );
  MUX2_X1 U9951 ( .A(n8403), .B(n8478), .S(n9851), .Z(n8405) );
  NAND2_X1 U9952 ( .A1(n8480), .A2(n8428), .ZN(n8404) );
  OAI211_X1 U9953 ( .C1(n8422), .C2(n8483), .A(n8405), .B(n8404), .ZN(P2_U3481) );
  INV_X1 U9954 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8406) );
  MUX2_X1 U9955 ( .A(n8406), .B(n8484), .S(n9851), .Z(n8408) );
  NAND2_X1 U9956 ( .A1(n8486), .A2(n8428), .ZN(n8407) );
  OAI211_X1 U9957 ( .C1(n8422), .C2(n8489), .A(n8408), .B(n8407), .ZN(P2_U3480) );
  MUX2_X1 U9958 ( .A(n8409), .B(n8490), .S(n9851), .Z(n8411) );
  NAND2_X1 U9959 ( .A1(n8492), .A2(n8428), .ZN(n8410) );
  OAI211_X1 U9960 ( .C1(n8422), .C2(n8495), .A(n8411), .B(n8410), .ZN(P2_U3479) );
  MUX2_X1 U9961 ( .A(n9986), .B(n8496), .S(n9851), .Z(n8413) );
  INV_X1 U9962 ( .A(n8422), .ZN(n8429) );
  AOI22_X1 U9963 ( .A1(n8499), .A2(n8429), .B1(n8428), .B2(n8498), .ZN(n8412)
         );
  NAND2_X1 U9964 ( .A1(n8413), .A2(n8412), .ZN(P2_U3478) );
  MUX2_X1 U9965 ( .A(n8414), .B(n8502), .S(n9851), .Z(n8416) );
  AOI22_X1 U9966 ( .A1(n8504), .A2(n8429), .B1(n8428), .B2(n8503), .ZN(n8415)
         );
  NAND2_X1 U9967 ( .A1(n8416), .A2(n8415), .ZN(P2_U3477) );
  MUX2_X1 U9968 ( .A(n8508), .B(n8417), .S(n9849), .Z(n8419) );
  NAND2_X1 U9969 ( .A1(n8509), .A2(n8428), .ZN(n8418) );
  OAI211_X1 U9970 ( .C1(n8512), .C2(n8422), .A(n8419), .B(n8418), .ZN(P2_U3476) );
  MUX2_X1 U9971 ( .A(n10040), .B(n8514), .S(n9851), .Z(n8421) );
  NAND2_X1 U9972 ( .A1(n8515), .A2(n8428), .ZN(n8420) );
  OAI211_X1 U9973 ( .C1(n8422), .C2(n8519), .A(n8421), .B(n8420), .ZN(P2_U3475) );
  MUX2_X1 U9974 ( .A(n10085), .B(n8520), .S(n9851), .Z(n8424) );
  AOI22_X1 U9975 ( .A1(n8523), .A2(n8429), .B1(n8428), .B2(n8522), .ZN(n8423)
         );
  NAND2_X1 U9976 ( .A1(n8424), .A2(n8423), .ZN(P2_U3474) );
  MUX2_X1 U9977 ( .A(n8425), .B(n8526), .S(n9851), .Z(n8427) );
  AOI22_X1 U9978 ( .A1(n8528), .A2(n8429), .B1(n8428), .B2(n8527), .ZN(n8426)
         );
  NAND2_X1 U9979 ( .A1(n8427), .A2(n8426), .ZN(P2_U3473) );
  MUX2_X1 U9980 ( .A(n6009), .B(n8531), .S(n9851), .Z(n8431) );
  AOI22_X1 U9981 ( .A1(n8536), .A2(n8429), .B1(n8428), .B2(n8533), .ZN(n8430)
         );
  NAND2_X1 U9982 ( .A1(n8431), .A2(n8430), .ZN(P2_U3472) );
  MUX2_X1 U9983 ( .A(n8432), .B(P2_REG1_REG_0__SCAN_IN), .S(n9849), .Z(
        P2_U3459) );
  NAND2_X1 U9984 ( .A1(n8434), .A2(n8534), .ZN(n8436) );
  NAND2_X1 U9985 ( .A1(n8435), .A2(n9833), .ZN(n8438) );
  OAI211_X1 U9986 ( .C1(n7787), .C2(n9833), .A(n8436), .B(n8438), .ZN(P2_U3458) );
  NAND2_X1 U9987 ( .A1(n8437), .A2(n8534), .ZN(n8439) );
  OAI211_X1 U9988 ( .C1(n9833), .C2(n8440), .A(n8439), .B(n8438), .ZN(P2_U3457) );
  INV_X1 U9989 ( .A(n9819), .ZN(n9827) );
  INV_X1 U9990 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8442) );
  MUX2_X1 U9991 ( .A(n8442), .B(n8441), .S(n9833), .Z(n8445) );
  NAND2_X1 U9992 ( .A1(n8443), .A2(n8534), .ZN(n8444) );
  OAI211_X1 U9993 ( .C1(n8446), .C2(n8518), .A(n8445), .B(n8444), .ZN(P2_U3455) );
  NAND2_X1 U9994 ( .A1(n9835), .A2(n8448), .ZN(n8449) );
  NAND2_X1 U9995 ( .A1(n8451), .A2(n8534), .ZN(n8452) );
  OAI211_X1 U9996 ( .C1(n8454), .C2(n8518), .A(n8453), .B(n8452), .ZN(P2_U3454) );
  MUX2_X1 U9997 ( .A(n8456), .B(n8455), .S(n9833), .Z(n8459) );
  NAND2_X1 U9998 ( .A1(n8457), .A2(n8534), .ZN(n8458) );
  OAI211_X1 U9999 ( .C1(n8460), .C2(n8518), .A(n8459), .B(n8458), .ZN(P2_U3453) );
  MUX2_X1 U10000 ( .A(n10120), .B(n8461), .S(n9833), .Z(n8464) );
  NAND2_X1 U10001 ( .A1(n8462), .A2(n8534), .ZN(n8463) );
  OAI211_X1 U10002 ( .C1(n8465), .C2(n8518), .A(n8464), .B(n8463), .ZN(
        P2_U3452) );
  INV_X1 U10003 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8467) );
  MUX2_X1 U10004 ( .A(n8467), .B(n8466), .S(n9833), .Z(n8470) );
  NAND2_X1 U10005 ( .A1(n8468), .A2(n8534), .ZN(n8469) );
  OAI211_X1 U10006 ( .C1(n8471), .C2(n8518), .A(n8470), .B(n8469), .ZN(
        P2_U3451) );
  INV_X1 U10007 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8473) );
  MUX2_X1 U10008 ( .A(n8473), .B(n8472), .S(n9833), .Z(n8476) );
  NAND2_X1 U10009 ( .A1(n8474), .A2(n8534), .ZN(n8475) );
  OAI211_X1 U10010 ( .C1(n8477), .C2(n8518), .A(n8476), .B(n8475), .ZN(
        P2_U3450) );
  MUX2_X1 U10011 ( .A(n8479), .B(n8478), .S(n9833), .Z(n8482) );
  NAND2_X1 U10012 ( .A1(n8480), .A2(n8534), .ZN(n8481) );
  OAI211_X1 U10013 ( .C1(n8483), .C2(n8518), .A(n8482), .B(n8481), .ZN(
        P2_U3449) );
  MUX2_X1 U10014 ( .A(n8485), .B(n8484), .S(n9833), .Z(n8488) );
  NAND2_X1 U10015 ( .A1(n8486), .A2(n8534), .ZN(n8487) );
  OAI211_X1 U10016 ( .C1(n8489), .C2(n8518), .A(n8488), .B(n8487), .ZN(
        P2_U3448) );
  MUX2_X1 U10017 ( .A(n8491), .B(n8490), .S(n9833), .Z(n8494) );
  NAND2_X1 U10018 ( .A1(n8492), .A2(n8534), .ZN(n8493) );
  OAI211_X1 U10019 ( .C1(n8495), .C2(n8518), .A(n8494), .B(n8493), .ZN(
        P2_U3447) );
  INV_X1 U10020 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U10021 ( .A(n8497), .B(n8496), .S(n9833), .Z(n8501) );
  INV_X1 U10022 ( .A(n8518), .ZN(n8535) );
  AOI22_X1 U10023 ( .A1(n8499), .A2(n8535), .B1(n8534), .B2(n8498), .ZN(n8500)
         );
  NAND2_X1 U10024 ( .A1(n8501), .A2(n8500), .ZN(P2_U3446) );
  MUX2_X1 U10025 ( .A(n10168), .B(n8502), .S(n9833), .Z(n8506) );
  AOI22_X1 U10026 ( .A1(n8504), .A2(n8535), .B1(n8534), .B2(n8503), .ZN(n8505)
         );
  NAND2_X1 U10027 ( .A1(n8506), .A2(n8505), .ZN(P2_U3444) );
  INV_X1 U10028 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8507) );
  MUX2_X1 U10029 ( .A(n8508), .B(n8507), .S(n9835), .Z(n8511) );
  NAND2_X1 U10030 ( .A1(n8509), .A2(n8534), .ZN(n8510) );
  OAI211_X1 U10031 ( .C1(n8512), .C2(n8518), .A(n8511), .B(n8510), .ZN(
        P2_U3441) );
  INV_X1 U10032 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8513) );
  MUX2_X1 U10033 ( .A(n8514), .B(n8513), .S(n9835), .Z(n8517) );
  NAND2_X1 U10034 ( .A1(n8515), .A2(n8534), .ZN(n8516) );
  OAI211_X1 U10035 ( .C1(n8519), .C2(n8518), .A(n8517), .B(n8516), .ZN(
        P2_U3438) );
  INV_X1 U10036 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8521) );
  MUX2_X1 U10037 ( .A(n8521), .B(n8520), .S(n9833), .Z(n8525) );
  AOI22_X1 U10038 ( .A1(n8523), .A2(n8535), .B1(n8534), .B2(n8522), .ZN(n8524)
         );
  NAND2_X1 U10039 ( .A1(n8525), .A2(n8524), .ZN(P2_U3435) );
  MUX2_X1 U10040 ( .A(n10082), .B(n8526), .S(n9833), .Z(n8530) );
  AOI22_X1 U10041 ( .A1(n8528), .A2(n8535), .B1(n8534), .B2(n8527), .ZN(n8529)
         );
  NAND2_X1 U10042 ( .A1(n8530), .A2(n8529), .ZN(P2_U3432) );
  INV_X1 U10043 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10044 ( .A(n8532), .B(n8531), .S(n9833), .Z(n8538) );
  AOI22_X1 U10045 ( .A1(n8536), .A2(n8535), .B1(n8534), .B2(n8533), .ZN(n8537)
         );
  NAND2_X1 U10046 ( .A1(n8538), .A2(n8537), .ZN(P2_U3429) );
  INV_X1 U10047 ( .A(n9227), .ZN(n8542) );
  NOR4_X1 U10048 ( .A1(n8539), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5814), .ZN(n8540) );
  AOI21_X1 U10049 ( .B1(n8552), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8540), .ZN(
        n8541) );
  OAI21_X1 U10050 ( .B1(n8542), .B2(n8559), .A(n8541), .ZN(P2_U3264) );
  OAI222_X1 U10051 ( .A1(n8543), .A2(P2_U3151), .B1(n8559), .B2(n8544), .C1(
        n10086), .C2(n8557), .ZN(P2_U3265) );
  OAI222_X1 U10052 ( .A1(P2_U3151), .A2(n8547), .B1(n8559), .B2(n8546), .C1(
        n8545), .C2(n8557), .ZN(P2_U3266) );
  AOI21_X1 U10053 ( .B1(n8552), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n4506), .ZN(
        n8548) );
  OAI21_X1 U10054 ( .B1(n8549), .B2(n8559), .A(n8548), .ZN(P2_U3267) );
  INV_X1 U10055 ( .A(n8550), .ZN(n9230) );
  AOI21_X1 U10056 ( .B1(n8552), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8551), .ZN(
        n8553) );
  OAI21_X1 U10057 ( .B1(n9230), .B2(n8559), .A(n8553), .ZN(P2_U3268) );
  INV_X1 U10058 ( .A(n8554), .ZN(n9233) );
  OAI222_X1 U10059 ( .A1(n6213), .A2(P2_U3151), .B1(n8559), .B2(n9233), .C1(
        n8555), .C2(n8557), .ZN(P2_U3269) );
  INV_X1 U10060 ( .A(n8556), .ZN(n9236) );
  OAI222_X1 U10061 ( .A1(n8560), .A2(P2_U3151), .B1(n8559), .B2(n9236), .C1(
        n8558), .C2(n8557), .ZN(P2_U3270) );
  NAND2_X1 U10062 ( .A1(n4497), .A2(n8562), .ZN(n8564) );
  XNOR2_X1 U10063 ( .A(n8564), .B(n8563), .ZN(n8569) );
  AOI22_X1 U10064 ( .A1(n8874), .A2(n8859), .B1(n8699), .B2(n8728), .ZN(n9402)
         );
  OAI22_X1 U10065 ( .A1(n9402), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8565), .ZN(n8567) );
  NOR2_X1 U10066 ( .A1(n9545), .A2(n8717), .ZN(n8566) );
  AOI211_X1 U10067 ( .C1(n8713), .C2(n9405), .A(n8567), .B(n8566), .ZN(n8568)
         );
  OAI21_X1 U10068 ( .B1(n8569), .B2(n9260), .A(n8568), .ZN(P1_U3215) );
  INV_X1 U10069 ( .A(n9161), .ZN(n9007) );
  INV_X1 U10070 ( .A(n8570), .ZN(n8645) );
  NOR3_X1 U10071 ( .A1(n8673), .A2(n8572), .A3(n8571), .ZN(n8573) );
  OAI21_X1 U10072 ( .B1(n8645), .B2(n8573), .A(n8709), .ZN(n8579) );
  OR2_X1 U10073 ( .A1(n8892), .A2(n8927), .ZN(n8575) );
  NAND2_X1 U10074 ( .A1(n8722), .A2(n8859), .ZN(n8574) );
  AND2_X1 U10075 ( .A1(n8575), .A2(n8574), .ZN(n9011) );
  OAI22_X1 U10076 ( .A1(n9011), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8576), .ZN(n8577) );
  AOI21_X1 U10077 ( .B1(n9005), .B2(n8713), .A(n8577), .ZN(n8578) );
  OAI211_X1 U10078 ( .C1(n9007), .C2(n8717), .A(n8579), .B(n8578), .ZN(
        P1_U3216) );
  NAND2_X1 U10079 ( .A1(n4495), .A2(n8580), .ZN(n8581) );
  XNOR2_X1 U10080 ( .A(n8582), .B(n8581), .ZN(n8588) );
  NOR2_X1 U10081 ( .A1(n9267), .A2(n8583), .ZN(n8586) );
  AOI22_X1 U10082 ( .A1(n8725), .A2(n8859), .B1(n8699), .B2(n8882), .ZN(n9063)
         );
  OAI22_X1 U10083 ( .A1(n9063), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8584), .ZN(n8585) );
  AOI211_X1 U10084 ( .C1(n9182), .C2(n5768), .A(n8586), .B(n8585), .ZN(n8587)
         );
  OAI21_X1 U10085 ( .B1(n8588), .B2(n9260), .A(n8587), .ZN(P1_U3219) );
  OAI21_X1 U10086 ( .B1(n8591), .B2(n8590), .A(n8589), .ZN(n8592) );
  NAND2_X1 U10087 ( .A1(n8592), .A2(n8709), .ZN(n8599) );
  INV_X1 U10088 ( .A(n8593), .ZN(n9040) );
  OR2_X1 U10089 ( .A1(n8892), .A2(n8697), .ZN(n8595) );
  NAND2_X1 U10090 ( .A1(n8725), .A2(n8699), .ZN(n8594) );
  AND2_X1 U10091 ( .A1(n8595), .A2(n8594), .ZN(n9037) );
  INV_X1 U10092 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8596) );
  OAI22_X1 U10093 ( .A1(n9037), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8596), .ZN(n8597) );
  AOI21_X1 U10094 ( .B1(n9040), .B2(n8713), .A(n8597), .ZN(n8598) );
  OAI211_X1 U10095 ( .C1(n9043), .C2(n8717), .A(n8599), .B(n8598), .ZN(
        P1_U3223) );
  INV_X1 U10096 ( .A(n7278), .ZN(n8601) );
  OAI22_X1 U10097 ( .A1(n8603), .A2(n8602), .B1(n8601), .B2(n8600), .ZN(n9259)
         );
  NAND2_X1 U10098 ( .A1(n8604), .A2(n8605), .ZN(n9258) );
  NOR2_X1 U10099 ( .A1(n9259), .A2(n9258), .ZN(n9257) );
  INV_X1 U10100 ( .A(n8605), .ZN(n8607) );
  NOR3_X1 U10101 ( .A1(n9257), .A2(n8607), .A3(n8606), .ZN(n8609) );
  INV_X1 U10102 ( .A(n7289), .ZN(n8608) );
  OAI21_X1 U10103 ( .B1(n8609), .B2(n8608), .A(n8709), .ZN(n8614) );
  NAND2_X1 U10104 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9319) );
  OAI21_X1 U10105 ( .B1(n8610), .B2(n9255), .A(n9319), .ZN(n8611) );
  AOI21_X1 U10106 ( .B1(n8612), .B2(n8713), .A(n8611), .ZN(n8613) );
  OAI211_X1 U10107 ( .C1(n9538), .C2(n8717), .A(n8614), .B(n8613), .ZN(
        P1_U3224) );
  OAI21_X1 U10108 ( .B1(n8616), .B2(n8615), .A(n8693), .ZN(n8617) );
  NAND2_X1 U10109 ( .A1(n8617), .A2(n8709), .ZN(n8623) );
  NAND2_X1 U10110 ( .A1(n8722), .A2(n8699), .ZN(n8619) );
  NAND2_X1 U10111 ( .A1(n8721), .A2(n8859), .ZN(n8618) );
  AND2_X1 U10112 ( .A1(n8619), .A2(n8618), .ZN(n8979) );
  OAI22_X1 U10113 ( .A1(n8979), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8620), .ZN(n8621) );
  AOI21_X1 U10114 ( .B1(n8983), .B2(n8713), .A(n8621), .ZN(n8622) );
  OAI211_X1 U10115 ( .C1(n8986), .C2(n8717), .A(n8623), .B(n8622), .ZN(
        P1_U3225) );
  OAI21_X1 U10116 ( .B1(n8625), .B2(n8624), .A(n8633), .ZN(n8626) );
  NAND2_X1 U10117 ( .A1(n8626), .A2(n8709), .ZN(n8631) );
  OR2_X1 U10118 ( .A1(n8872), .A2(n8927), .ZN(n8628) );
  NAND2_X1 U10119 ( .A1(n8726), .A2(n8859), .ZN(n8627) );
  AND2_X1 U10120 ( .A1(n8628), .A2(n8627), .ZN(n9112) );
  NAND2_X1 U10121 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9375) );
  OAI21_X1 U10122 ( .B1(n9112), .B2(n9255), .A(n9375), .ZN(n8629) );
  AOI21_X1 U10123 ( .B1(n5023), .B2(n8713), .A(n8629), .ZN(n8630) );
  OAI211_X1 U10124 ( .C1(n9105), .C2(n8717), .A(n8631), .B(n8630), .ZN(
        P1_U3226) );
  AND2_X1 U10125 ( .A1(n8633), .A2(n8632), .ZN(n8636) );
  OAI211_X1 U10126 ( .C1(n8636), .C2(n8635), .A(n8709), .B(n8634), .ZN(n8641)
         );
  NAND2_X1 U10127 ( .A1(n8882), .A2(n8859), .ZN(n8638) );
  NAND2_X1 U10128 ( .A1(n8875), .A2(n8699), .ZN(n8637) );
  AND2_X1 U10129 ( .A1(n8638), .A2(n8637), .ZN(n9089) );
  NAND2_X1 U10130 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8831) );
  OAI21_X1 U10131 ( .B1(n9089), .B2(n9255), .A(n8831), .ZN(n8639) );
  AOI21_X1 U10132 ( .B1(n9095), .B2(n8713), .A(n8639), .ZN(n8640) );
  OAI211_X1 U10133 ( .C1(n9270), .C2(n8717), .A(n8641), .B(n8640), .ZN(
        P1_U3228) );
  INV_X1 U10134 ( .A(n8642), .ZN(n8644) );
  NOR3_X1 U10135 ( .A1(n8645), .A2(n8644), .A3(n8643), .ZN(n8648) );
  INV_X1 U10136 ( .A(n8646), .ZN(n8647) );
  OAI21_X1 U10137 ( .B1(n8648), .B2(n8647), .A(n8709), .ZN(n8654) );
  NAND2_X1 U10138 ( .A1(n8895), .A2(n8699), .ZN(n8650) );
  NAND2_X1 U10139 ( .A1(n8897), .A2(n8859), .ZN(n8649) );
  AND2_X1 U10140 ( .A1(n8650), .A2(n8649), .ZN(n8992) );
  OAI22_X1 U10141 ( .A1(n8992), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8651), .ZN(n8652) );
  AOI21_X1 U10142 ( .B1(n8997), .B2(n8713), .A(n8652), .ZN(n8653) );
  OAI211_X1 U10143 ( .C1(n9000), .C2(n8717), .A(n8654), .B(n8653), .ZN(
        P1_U3229) );
  NAND2_X1 U10144 ( .A1(n8657), .A2(n8656), .ZN(n8663) );
  OAI22_X1 U10145 ( .A1(n8659), .A2(n8927), .B1(n8658), .B2(n8697), .ZN(n9428)
         );
  AOI22_X1 U10146 ( .A1(n9428), .A2(n8660), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n8662) );
  AOI22_X1 U10147 ( .A1(n5768), .A2(n9432), .B1(n8713), .B2(n9430), .ZN(n8661)
         );
  NAND3_X1 U10148 ( .A1(n8663), .A2(n8662), .A3(n8661), .ZN(P1_U3230) );
  INV_X1 U10149 ( .A(n8664), .ZN(n8665) );
  AOI21_X1 U10150 ( .B1(n8667), .B2(n8666), .A(n8665), .ZN(n8672) );
  NOR2_X1 U10151 ( .A1(n9267), .A2(n9053), .ZN(n8670) );
  AOI22_X1 U10152 ( .A1(n8724), .A2(n8859), .B1(n8699), .B2(n8885), .ZN(n9049)
         );
  OAI22_X1 U10153 ( .A1(n9049), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8668), .ZN(n8669) );
  AOI211_X1 U10154 ( .C1(n9177), .C2(n5768), .A(n8670), .B(n8669), .ZN(n8671)
         );
  OAI21_X1 U10155 ( .B1(n8672), .B2(n9260), .A(n8671), .ZN(P1_U3233) );
  AOI21_X1 U10156 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8679) );
  AOI22_X1 U10157 ( .A1(n8724), .A2(n8699), .B1(n8859), .B2(n8895), .ZN(n9021)
         );
  OAI22_X1 U10158 ( .A1(n9021), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10182), .ZN(n8677) );
  NOR2_X1 U10159 ( .A1(n9030), .A2(n8717), .ZN(n8676) );
  AOI211_X1 U10160 ( .C1(n8713), .C2(n9027), .A(n8677), .B(n8676), .ZN(n8678)
         );
  OAI21_X1 U10161 ( .B1(n8679), .B2(n9260), .A(n8678), .ZN(P1_U3235) );
  INV_X1 U10162 ( .A(n8680), .ZN(n8681) );
  NOR2_X1 U10163 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  XNOR2_X1 U10164 ( .A(n8684), .B(n8683), .ZN(n8691) );
  NAND2_X1 U10165 ( .A1(n8885), .A2(n8859), .ZN(n8686) );
  NAND2_X1 U10166 ( .A1(n8726), .A2(n8699), .ZN(n8685) );
  AND2_X1 U10167 ( .A1(n8686), .A2(n8685), .ZN(n9075) );
  OAI22_X1 U10168 ( .A1(n9075), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8687), .ZN(n8689) );
  NOR2_X1 U10169 ( .A1(n9083), .A2(n8717), .ZN(n8688) );
  AOI211_X1 U10170 ( .C1(n8713), .C2(n9080), .A(n8689), .B(n8688), .ZN(n8690)
         );
  OAI21_X1 U10171 ( .B1(n8691), .B2(n9260), .A(n8690), .ZN(P1_U3238) );
  AND2_X1 U10172 ( .A1(n8693), .A2(n8692), .ZN(n8696) );
  OAI211_X1 U10173 ( .C1(n8696), .C2(n8695), .A(n8709), .B(n8694), .ZN(n8705)
         );
  OR2_X1 U10174 ( .A1(n8698), .A2(n8697), .ZN(n8701) );
  NAND2_X1 U10175 ( .A1(n8897), .A2(n8699), .ZN(n8700) );
  AND2_X1 U10176 ( .A1(n8701), .A2(n8700), .ZN(n8970) );
  OAI22_X1 U10177 ( .A1(n8970), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8702), .ZN(n8703) );
  AOI21_X1 U10178 ( .B1(n8964), .B2(n8713), .A(n8703), .ZN(n8704) );
  OAI211_X1 U10179 ( .C1(n8966), .C2(n8717), .A(n8705), .B(n8704), .ZN(
        P1_U3240) );
  OAI21_X1 U10180 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8710) );
  NAND2_X1 U10181 ( .A1(n8710), .A2(n8709), .ZN(n8716) );
  NAND2_X1 U10182 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9361) );
  OAI21_X1 U10183 ( .B1(n8711), .B2(n9255), .A(n9361), .ZN(n8712) );
  AOI21_X1 U10184 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8715) );
  OAI211_X1 U10185 ( .C1(n9276), .C2(n8717), .A(n8716), .B(n8715), .ZN(
        P1_U3241) );
  MUX2_X1 U10186 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8718), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10187 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8719), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8720), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10189 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n8904), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10190 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8721), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8897), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8722), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8895), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n8723), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n8724), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10196 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n8725), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10197 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n8885), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8882), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10199 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n8726), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8875), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8874), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10202 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8727), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10203 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8728), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10204 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8729), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10205 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8730), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10206 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8731), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10207 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8732), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10208 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8733), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10209 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8734), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10210 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8735), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10211 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8736), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10212 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8737), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10213 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8738), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10214 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8739), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10215 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6708), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10216 ( .C1(n8741), .C2(n8754), .A(n9383), .B(n8740), .ZN(n8749)
         );
  AOI22_X1 U10217 ( .A1(n9305), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8748) );
  NAND2_X1 U10218 ( .A1(n9347), .A2(n8742), .ZN(n8747) );
  OAI211_X1 U10219 ( .C1(n8745), .C2(n8744), .A(n9379), .B(n8743), .ZN(n8746)
         );
  NAND4_X1 U10220 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(
        P1_U3244) );
  NAND3_X1 U10221 ( .A1(n8751), .A2(n8750), .A3(n4421), .ZN(n8757) );
  INV_X1 U10222 ( .A(n8752), .ZN(n8755) );
  NOR2_X1 U10223 ( .A1(n4421), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8753) );
  NOR2_X1 U10224 ( .A1(n5780), .A2(n8753), .ZN(n9284) );
  NOR2_X1 U10225 ( .A1(n9284), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9283) );
  AOI21_X1 U10226 ( .B1(n8755), .B2(n8754), .A(n9283), .ZN(n8756) );
  NAND3_X1 U10227 ( .A1(n8757), .A2(P1_U3973), .A3(n8756), .ZN(n8795) );
  INV_X1 U10228 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8758) );
  OAI22_X1 U10229 ( .A1(n9393), .A2(n8758), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6887), .ZN(n8759) );
  AOI21_X1 U10230 ( .B1(n8760), .B2(n9347), .A(n8759), .ZN(n8769) );
  OAI211_X1 U10231 ( .C1(n8763), .C2(n8762), .A(n9379), .B(n8761), .ZN(n8768)
         );
  OAI211_X1 U10232 ( .C1(n8766), .C2(n8765), .A(n9383), .B(n8764), .ZN(n8767)
         );
  NAND4_X1 U10233 ( .A1(n8795), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(
        P1_U3245) );
  NAND2_X1 U10234 ( .A1(n9305), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U10235 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n8770) );
  OAI211_X1 U10236 ( .C1(n9389), .C2(n8772), .A(n8771), .B(n8770), .ZN(n8773)
         );
  INV_X1 U10237 ( .A(n8773), .ZN(n8782) );
  OAI211_X1 U10238 ( .C1(n8776), .C2(n8775), .A(n9379), .B(n8774), .ZN(n8781)
         );
  OAI211_X1 U10239 ( .C1(n8779), .C2(n8778), .A(n9383), .B(n8777), .ZN(n8780)
         );
  NAND3_X1 U10240 ( .A1(n8782), .A2(n8781), .A3(n8780), .ZN(P1_U3246) );
  AND2_X1 U10241 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8785) );
  NOR2_X1 U10242 ( .A1(n9389), .A2(n8783), .ZN(n8784) );
  AOI211_X1 U10243 ( .C1(n9305), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n8785), .B(
        n8784), .ZN(n8794) );
  OAI211_X1 U10244 ( .C1(n8788), .C2(n8787), .A(n9383), .B(n8786), .ZN(n8793)
         );
  OAI211_X1 U10245 ( .C1(n8791), .C2(n8790), .A(n9379), .B(n8789), .ZN(n8792)
         );
  NAND4_X1 U10246 ( .A1(n8795), .A2(n8794), .A3(n8793), .A4(n8792), .ZN(
        P1_U3247) );
  INV_X1 U10247 ( .A(n8813), .ZN(n8835) );
  OR2_X1 U10248 ( .A1(n8813), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U10249 ( .A1(n8813), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8796) );
  AND2_X1 U10250 ( .A1(n8841), .A2(n8796), .ZN(n8812) );
  XNOR2_X1 U10251 ( .A(n9367), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9365) );
  INV_X1 U10252 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U10253 ( .A1(n9346), .A2(n8798), .ZN(n8797) );
  OAI21_X1 U10254 ( .B1(n9346), .B2(n8798), .A(n8797), .ZN(n9339) );
  NAND2_X1 U10255 ( .A1(n8822), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8807) );
  INV_X1 U10256 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8799) );
  MUX2_X1 U10257 ( .A(n8799), .B(P1_REG1_REG_13__SCAN_IN), .S(n8822), .Z(n9324) );
  OR2_X1 U10258 ( .A1(n8821), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8805) );
  INV_X1 U10259 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8800) );
  MUX2_X1 U10260 ( .A(n8800), .B(P1_REG1_REG_10__SCAN_IN), .S(n8819), .Z(n9238) );
  OR2_X1 U10261 ( .A1(n8818), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U10262 ( .A1(n8802), .A2(n8801), .ZN(n9239) );
  NOR2_X1 U10263 ( .A1(n9238), .A2(n9239), .ZN(n9240) );
  AOI21_X1 U10264 ( .B1(n8819), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9240), .ZN(
        n9298) );
  INV_X1 U10265 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9570) );
  NOR2_X1 U10266 ( .A1(n9301), .A2(n9570), .ZN(n8803) );
  AOI21_X1 U10267 ( .B1(n9301), .B2(n9570), .A(n8803), .ZN(n9297) );
  NOR2_X1 U10268 ( .A1(n9298), .A2(n9297), .ZN(n9296) );
  AOI21_X1 U10269 ( .B1(n9301), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9296), .ZN(
        n9308) );
  INV_X1 U10270 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8804) );
  MUX2_X1 U10271 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n8804), .S(n8821), .Z(n9309) );
  NAND2_X1 U10272 ( .A1(n9308), .A2(n9309), .ZN(n9307) );
  NAND2_X1 U10273 ( .A1(n8805), .A2(n9307), .ZN(n9323) );
  NOR2_X1 U10274 ( .A1(n9324), .A2(n9323), .ZN(n9322) );
  INV_X1 U10275 ( .A(n9322), .ZN(n8806) );
  NAND2_X1 U10276 ( .A1(n8807), .A2(n8806), .ZN(n9338) );
  NAND2_X1 U10277 ( .A1(n9339), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U10278 ( .A1(n9346), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8808) );
  AND2_X1 U10279 ( .A1(n9337), .A2(n8808), .ZN(n8809) );
  NOR2_X1 U10280 ( .A1(n8809), .A2(n9359), .ZN(n8810) );
  INV_X1 U10281 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10101) );
  XNOR2_X1 U10282 ( .A(n8809), .B(n9359), .ZN(n9352) );
  NOR2_X1 U10283 ( .A1(n10101), .A2(n9352), .ZN(n9351) );
  NOR2_X1 U10284 ( .A1(n8810), .A2(n9351), .ZN(n9366) );
  NAND2_X1 U10285 ( .A1(n9365), .A2(n9366), .ZN(n9364) );
  OAI21_X1 U10286 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n8826), .A(n9364), .ZN(
        n8811) );
  NAND2_X1 U10287 ( .A1(n8812), .A2(n8811), .ZN(n8842) );
  OAI21_X1 U10288 ( .B1(n8812), .B2(n8811), .A(n8842), .ZN(n8830) );
  OR2_X1 U10289 ( .A1(n8813), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U10290 ( .A1(n8813), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8814) );
  AND2_X1 U10291 ( .A1(n8836), .A2(n8814), .ZN(n8828) );
  XNOR2_X1 U10292 ( .A(n9346), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9342) );
  INV_X1 U10293 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U10294 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9332), .B1(n8822), .B2(
        n10053), .ZN(n9328) );
  NOR2_X1 U10295 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n8821), .ZN(n8815) );
  AOI21_X1 U10296 ( .B1(n8821), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8815), .ZN(
        n9313) );
  NAND2_X1 U10297 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n8819), .ZN(n8816) );
  OAI21_X1 U10298 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n8819), .A(n8816), .ZN(
        n9245) );
  OAI21_X1 U10299 ( .B1(n8818), .B2(P1_REG2_REG_9__SCAN_IN), .A(n8817), .ZN(
        n9244) );
  NOR2_X1 U10300 ( .A1(n9245), .A2(n9244), .ZN(n9243) );
  NAND2_X1 U10301 ( .A1(n9301), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8820) );
  OAI21_X1 U10302 ( .B1(n9301), .B2(P1_REG2_REG_11__SCAN_IN), .A(n8820), .ZN(
        n9293) );
  OAI21_X1 U10303 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n8821), .A(n9311), .ZN(
        n9327) );
  NOR2_X1 U10304 ( .A1(n9328), .A2(n9327), .ZN(n9326) );
  NOR2_X1 U10305 ( .A1(n8823), .A2(n9359), .ZN(n8825) );
  INV_X1 U10306 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U10307 ( .A1(n10022), .A2(n9355), .ZN(n9354) );
  NOR2_X1 U10308 ( .A1(n8825), .A2(n9354), .ZN(n9371) );
  INV_X1 U10309 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U10310 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9367), .B1(n8826), .B2(
        n10008), .ZN(n9370) );
  NOR2_X1 U10311 ( .A1(n9371), .A2(n9370), .ZN(n9369) );
  OAI21_X1 U10312 ( .B1(n8828), .B2(n8827), .A(n8837), .ZN(n8829) );
  AOI22_X1 U10313 ( .A1(n9379), .A2(n8830), .B1(n9383), .B2(n8829), .ZN(n8834)
         );
  INV_X1 U10314 ( .A(n8831), .ZN(n8832) );
  AOI21_X1 U10315 ( .B1(n9305), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n8832), .ZN(
        n8833) );
  OAI211_X1 U10316 ( .C1(n8835), .C2(n9389), .A(n8834), .B(n8833), .ZN(
        P1_U3260) );
  NAND2_X1 U10317 ( .A1(n8843), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8839) );
  OR2_X1 U10318 ( .A1(n8843), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8838) );
  AND2_X1 U10319 ( .A1(n8839), .A2(n8838), .ZN(n9385) );
  NAND2_X1 U10320 ( .A1(n9382), .A2(n8839), .ZN(n8840) );
  XNOR2_X1 U10321 ( .A(n8840), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n8849) );
  INV_X1 U10322 ( .A(n8849), .ZN(n8848) );
  AND2_X1 U10323 ( .A1(n8842), .A2(n8841), .ZN(n9380) );
  NAND2_X1 U10324 ( .A1(n8843), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8845) );
  OR2_X1 U10325 ( .A1(n8843), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8844) );
  AND2_X1 U10326 ( .A1(n8845), .A2(n8844), .ZN(n9381) );
  NAND2_X1 U10327 ( .A1(n9380), .A2(n9381), .ZN(n9378) );
  NAND2_X1 U10328 ( .A1(n9378), .A2(n8845), .ZN(n8846) );
  XNOR2_X1 U10329 ( .A(n8846), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U10330 ( .A1(n9379), .A2(n8850), .ZN(n8847) );
  OAI211_X1 U10331 ( .C1(n9368), .C2(n8848), .A(n8847), .B(n9389), .ZN(n8852)
         );
  OAI22_X1 U10332 ( .A1(n9295), .A2(n8850), .B1(n8849), .B2(n9368), .ZN(n8851)
         );
  MUX2_X1 U10333 ( .A(n8852), .B(n8851), .S(n5549), .Z(n8853) );
  INV_X1 U10334 ( .A(n8853), .ZN(n8855) );
  NAND2_X1 U10335 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8854) );
  OAI211_X1 U10336 ( .C1(n10033), .C2(n9393), .A(n8855), .B(n8854), .ZN(
        P1_U3262) );
  INV_X1 U10337 ( .A(n9134), .ZN(n8911) );
  NAND2_X1 U10338 ( .A1(n9077), .A2(n9083), .ZN(n9078) );
  OR2_X2 U10339 ( .A1(n9078), .A2(n9182), .ZN(n9065) );
  OR2_X2 U10340 ( .A1(n9065), .A2(n9177), .ZN(n9051) );
  NAND2_X1 U10341 ( .A1(n9000), .A2(n9004), .ZN(n8994) );
  OR2_X2 U10342 ( .A1(n8994), .A2(n9152), .ZN(n8981) );
  NAND2_X1 U10343 ( .A1(n9128), .A2(n8907), .ZN(n8864) );
  INV_X1 U10344 ( .A(P1_B_REG_SCAN_IN), .ZN(n10050) );
  OR2_X1 U10345 ( .A1(n4421), .A2(n10050), .ZN(n8858) );
  NAND2_X1 U10346 ( .A1(n8859), .A2(n8858), .ZN(n8929) );
  OR2_X1 U10347 ( .A1(n8860), .A2(n8929), .ZN(n9126) );
  NOR2_X1 U10348 ( .A1(n9126), .A2(n9455), .ZN(n8867) );
  NOR2_X1 U10349 ( .A1(n8856), .A2(n9104), .ZN(n8862) );
  AOI211_X1 U10350 ( .C1(n9455), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8867), .B(
        n8862), .ZN(n8863) );
  OAI21_X1 U10351 ( .B1(n9119), .B2(n8871), .A(n8863), .ZN(P1_U3263) );
  OAI211_X1 U10352 ( .C1(n9128), .C2(n8907), .A(n9436), .B(n8864), .ZN(n9127)
         );
  INV_X1 U10353 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8865) );
  NOR2_X1 U10354 ( .A1(n9452), .A2(n8865), .ZN(n8866) );
  NOR2_X1 U10355 ( .A1(n8867), .A2(n8866), .ZN(n8870) );
  NAND2_X1 U10356 ( .A1(n8868), .A2(n9431), .ZN(n8869) );
  OAI211_X1 U10357 ( .C1(n9127), .C2(n8871), .A(n8870), .B(n8869), .ZN(
        P1_U3264) );
  NAND2_X1 U10358 ( .A1(n9192), .A2(n8875), .ZN(n8876) );
  INV_X1 U10359 ( .A(n9092), .ZN(n8879) );
  AOI21_X1 U10360 ( .B1(n9092), .B2(n9270), .A(n8877), .ZN(n8878) );
  NOR2_X1 U10361 ( .A1(n9182), .A2(n8885), .ZN(n8887) );
  INV_X1 U10362 ( .A(n9182), .ZN(n9070) );
  INV_X1 U10363 ( .A(n9177), .ZN(n9057) );
  NAND2_X1 U10364 ( .A1(n9043), .A2(n8889), .ZN(n8890) );
  NAND2_X1 U10365 ( .A1(n8891), .A2(n8890), .ZN(n9017) );
  NAND2_X1 U10366 ( .A1(n9030), .A2(n8892), .ZN(n8893) );
  NOR2_X1 U10367 ( .A1(n9161), .A2(n8895), .ZN(n8894) );
  NOR2_X1 U10368 ( .A1(n9152), .A2(n8897), .ZN(n8899) );
  OAI22_X1 U10369 ( .A1(n8976), .A2(n8899), .B1(n8898), .B2(n8986), .ZN(n8962)
         );
  NOR2_X1 U10370 ( .A1(n8966), .A2(n8901), .ZN(n8900) );
  NAND2_X1 U10371 ( .A1(n8966), .A2(n8901), .ZN(n8902) );
  AOI22_X1 U10372 ( .A1(n8933), .A2(n8923), .B1(n4643), .B2(n8926), .ZN(n8906)
         );
  XNOR2_X1 U10373 ( .A(n8906), .B(n8905), .ZN(n9131) );
  INV_X1 U10374 ( .A(n9131), .ZN(n8932) );
  AOI211_X1 U10375 ( .C1(n9134), .C2(n8908), .A(n9101), .B(n8907), .ZN(n9133)
         );
  AOI22_X1 U10376 ( .A1(n9455), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8909), .B2(
        n9447), .ZN(n8910) );
  OAI21_X1 U10377 ( .B1(n8911), .B2(n9104), .A(n8910), .ZN(n8912) );
  AOI21_X1 U10378 ( .B1(n9133), .B2(n9440), .A(n8912), .ZN(n8931) );
  NAND2_X1 U10379 ( .A1(n8914), .A2(n8913), .ZN(n9018) );
  INV_X1 U10380 ( .A(n8916), .ZN(n8917) );
  AOI21_X1 U10381 ( .B1(n8978), .B2(n8977), .A(n8920), .ZN(n8968) );
  NAND2_X1 U10382 ( .A1(n8968), .A2(n8969), .ZN(n8967) );
  NAND2_X1 U10383 ( .A1(n8967), .A2(n8921), .ZN(n8954) );
  NAND2_X1 U10384 ( .A1(n8953), .A2(n8922), .ZN(n8938) );
  NAND2_X1 U10385 ( .A1(n8938), .A2(n8939), .ZN(n8937) );
  NAND2_X1 U10386 ( .A1(n8937), .A2(n7464), .ZN(n8925) );
  NAND2_X1 U10387 ( .A1(n9132), .A2(n9452), .ZN(n8930) );
  OAI211_X1 U10388 ( .C1(n8932), .C2(n9086), .A(n8931), .B(n8930), .ZN(
        P1_U3356) );
  XNOR2_X1 U10389 ( .A(n8933), .B(n8939), .ZN(n9139) );
  AOI211_X1 U10390 ( .C1(n9136), .C2(n8947), .A(n9101), .B(n8934), .ZN(n9135)
         );
  AOI22_X1 U10391 ( .A1(n9455), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8935), .B2(
        n9447), .ZN(n8936) );
  OAI21_X1 U10392 ( .B1(n4643), .B2(n9104), .A(n8936), .ZN(n8944) );
  OAI21_X1 U10393 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8942) );
  INV_X1 U10394 ( .A(n8940), .ZN(n8941) );
  AOI21_X1 U10395 ( .B1(n8942), .B2(n9459), .A(n8941), .ZN(n9138) );
  NOR2_X1 U10396 ( .A1(n9138), .A2(n9455), .ZN(n8943) );
  AOI211_X1 U10397 ( .C1(n9440), .C2(n9135), .A(n8944), .B(n8943), .ZN(n8945)
         );
  OAI21_X1 U10398 ( .B1(n9139), .B2(n9086), .A(n8945), .ZN(P1_U3265) );
  XNOR2_X1 U10399 ( .A(n8946), .B(n8955), .ZN(n9144) );
  INV_X1 U10400 ( .A(n8963), .ZN(n8949) );
  INV_X1 U10401 ( .A(n8947), .ZN(n8948) );
  AOI211_X1 U10402 ( .C1(n9141), .C2(n8949), .A(n9101), .B(n8948), .ZN(n9140)
         );
  AOI22_X1 U10403 ( .A1(n9455), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9447), .B2(
        n8950), .ZN(n8951) );
  OAI21_X1 U10404 ( .B1(n8952), .B2(n9104), .A(n8951), .ZN(n8960) );
  OAI21_X1 U10405 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8958) );
  INV_X1 U10406 ( .A(n8956), .ZN(n8957) );
  AOI21_X1 U10407 ( .B1(n8958), .B2(n9459), .A(n8957), .ZN(n9143) );
  NOR2_X1 U10408 ( .A1(n9143), .A2(n9455), .ZN(n8959) );
  AOI211_X1 U10409 ( .C1(n9140), .C2(n9440), .A(n8960), .B(n8959), .ZN(n8961)
         );
  OAI21_X1 U10410 ( .B1(n9144), .B2(n9086), .A(n8961), .ZN(P1_U3266) );
  XOR2_X1 U10411 ( .A(n8969), .B(n8962), .Z(n9149) );
  AOI211_X1 U10412 ( .C1(n9146), .C2(n8981), .A(n9101), .B(n8963), .ZN(n9145)
         );
  AOI22_X1 U10413 ( .A1(n9455), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n8964), .B2(
        n9447), .ZN(n8965) );
  OAI21_X1 U10414 ( .B1(n8966), .B2(n9104), .A(n8965), .ZN(n8974) );
  OAI21_X1 U10415 ( .B1(n8969), .B2(n8968), .A(n8967), .ZN(n8972) );
  INV_X1 U10416 ( .A(n8970), .ZN(n8971) );
  AOI21_X1 U10417 ( .B1(n8972), .B2(n9459), .A(n8971), .ZN(n9148) );
  NOR2_X1 U10418 ( .A1(n9148), .A2(n9455), .ZN(n8973) );
  AOI211_X1 U10419 ( .C1(n9145), .C2(n9440), .A(n8974), .B(n8973), .ZN(n8975)
         );
  OAI21_X1 U10420 ( .B1(n9149), .B2(n9086), .A(n8975), .ZN(P1_U3267) );
  XNOR2_X1 U10421 ( .A(n8976), .B(n8977), .ZN(n9154) );
  XNOR2_X1 U10422 ( .A(n8978), .B(n8977), .ZN(n8980) );
  OAI21_X1 U10423 ( .B1(n8980), .B2(n9399), .A(n8979), .ZN(n9150) );
  INV_X1 U10424 ( .A(n8981), .ZN(n8982) );
  AOI211_X1 U10425 ( .C1(n9152), .C2(n8994), .A(n9101), .B(n8982), .ZN(n9151)
         );
  NAND2_X1 U10426 ( .A1(n9151), .A2(n9440), .ZN(n8985) );
  AOI22_X1 U10427 ( .A1(n9455), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n8983), .B2(
        n9447), .ZN(n8984) );
  OAI211_X1 U10428 ( .C1(n8986), .C2(n9104), .A(n8985), .B(n8984), .ZN(n8987)
         );
  AOI21_X1 U10429 ( .B1(n9150), .B2(n9452), .A(n8987), .ZN(n8988) );
  OAI21_X1 U10430 ( .B1(n9154), .B2(n9086), .A(n8988), .ZN(P1_U3268) );
  XNOR2_X1 U10431 ( .A(n8989), .B(n8990), .ZN(n9159) );
  XNOR2_X1 U10432 ( .A(n8991), .B(n8990), .ZN(n8993) );
  OAI21_X1 U10433 ( .B1(n8993), .B2(n9399), .A(n8992), .ZN(n9155) );
  INV_X1 U10434 ( .A(n8994), .ZN(n8995) );
  AOI211_X1 U10435 ( .C1(n9157), .C2(n8996), .A(n9101), .B(n8995), .ZN(n9156)
         );
  NAND2_X1 U10436 ( .A1(n9156), .A2(n9440), .ZN(n8999) );
  AOI22_X1 U10437 ( .A1(n9455), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n8997), .B2(
        n9447), .ZN(n8998) );
  OAI211_X1 U10438 ( .C1(n9000), .C2(n9104), .A(n8999), .B(n8998), .ZN(n9001)
         );
  AOI21_X1 U10439 ( .B1(n9155), .B2(n9452), .A(n9001), .ZN(n9002) );
  OAI21_X1 U10440 ( .B1(n9159), .B2(n9086), .A(n9002), .ZN(P1_U3269) );
  XNOR2_X1 U10441 ( .A(n9003), .B(n9010), .ZN(n9164) );
  AOI211_X1 U10442 ( .C1(n9161), .C2(n9024), .A(n9101), .B(n9004), .ZN(n9160)
         );
  AOI22_X1 U10443 ( .A1(n9455), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9005), .B2(
        n9447), .ZN(n9006) );
  OAI21_X1 U10444 ( .B1(n9007), .B2(n9104), .A(n9006), .ZN(n9015) );
  OAI21_X1 U10445 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(n9013) );
  INV_X1 U10446 ( .A(n9011), .ZN(n9012) );
  AOI21_X1 U10447 ( .B1(n9013), .B2(n9459), .A(n9012), .ZN(n9163) );
  NOR2_X1 U10448 ( .A1(n9163), .A2(n9455), .ZN(n9014) );
  AOI211_X1 U10449 ( .C1(n9160), .C2(n9440), .A(n9015), .B(n9014), .ZN(n9016)
         );
  OAI21_X1 U10450 ( .B1(n9164), .B2(n9086), .A(n9016), .ZN(P1_U3270) );
  XNOR2_X1 U10451 ( .A(n9017), .B(n9019), .ZN(n9169) );
  INV_X1 U10452 ( .A(n9018), .ZN(n9020) );
  OAI21_X1 U10453 ( .B1(n9020), .B2(n9019), .A(n9459), .ZN(n9023) );
  OAI21_X1 U10454 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9165) );
  INV_X1 U10455 ( .A(n9030), .ZN(n9167) );
  INV_X1 U10456 ( .A(n9039), .ZN(n9026) );
  INV_X1 U10457 ( .A(n9024), .ZN(n9025) );
  AOI211_X1 U10458 ( .C1(n9167), .C2(n9026), .A(n9101), .B(n9025), .ZN(n9166)
         );
  NAND2_X1 U10459 ( .A1(n9166), .A2(n9440), .ZN(n9029) );
  AOI22_X1 U10460 ( .A1(n9455), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9027), .B2(
        n9447), .ZN(n9028) );
  OAI211_X1 U10461 ( .C1(n9030), .C2(n9104), .A(n9029), .B(n9028), .ZN(n9031)
         );
  AOI21_X1 U10462 ( .B1(n9165), .B2(n9452), .A(n9031), .ZN(n9032) );
  OAI21_X1 U10463 ( .B1(n9169), .B2(n9086), .A(n9032), .ZN(P1_U3271) );
  XNOR2_X1 U10464 ( .A(n9033), .B(n9035), .ZN(n9174) );
  OAI21_X1 U10465 ( .B1(n9048), .B2(n9047), .A(n9034), .ZN(n9036) );
  XNOR2_X1 U10466 ( .A(n9036), .B(n9035), .ZN(n9038) );
  OAI21_X1 U10467 ( .B1(n9038), .B2(n9399), .A(n9037), .ZN(n9170) );
  AOI211_X1 U10468 ( .C1(n9172), .C2(n9051), .A(n9101), .B(n9039), .ZN(n9171)
         );
  NAND2_X1 U10469 ( .A1(n9171), .A2(n9440), .ZN(n9042) );
  AOI22_X1 U10470 ( .A1(n9455), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9040), .B2(
        n9447), .ZN(n9041) );
  OAI211_X1 U10471 ( .C1(n9043), .C2(n9104), .A(n9042), .B(n9041), .ZN(n9044)
         );
  AOI21_X1 U10472 ( .B1(n9170), .B2(n9452), .A(n9044), .ZN(n9045) );
  OAI21_X1 U10473 ( .B1(n9174), .B2(n9086), .A(n9045), .ZN(P1_U3272) );
  XNOR2_X1 U10474 ( .A(n9046), .B(n9047), .ZN(n9179) );
  XNOR2_X1 U10475 ( .A(n9048), .B(n9047), .ZN(n9050) );
  OAI21_X1 U10476 ( .B1(n9050), .B2(n9399), .A(n9049), .ZN(n9175) );
  INV_X1 U10477 ( .A(n9051), .ZN(n9052) );
  AOI211_X1 U10478 ( .C1(n9177), .C2(n9065), .A(n9101), .B(n9052), .ZN(n9176)
         );
  NAND2_X1 U10479 ( .A1(n9176), .A2(n9440), .ZN(n9056) );
  INV_X1 U10480 ( .A(n9053), .ZN(n9054) );
  AOI22_X1 U10481 ( .A1(n9455), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9054), .B2(
        n9447), .ZN(n9055) );
  OAI211_X1 U10482 ( .C1(n9057), .C2(n9104), .A(n9056), .B(n9055), .ZN(n9058)
         );
  AOI21_X1 U10483 ( .B1(n9175), .B2(n9452), .A(n9058), .ZN(n9059) );
  OAI21_X1 U10484 ( .B1(n9179), .B2(n9086), .A(n9059), .ZN(P1_U3273) );
  XOR2_X1 U10485 ( .A(n9062), .B(n9060), .Z(n9184) );
  XOR2_X1 U10486 ( .A(n9062), .B(n9061), .Z(n9064) );
  OAI21_X1 U10487 ( .B1(n9064), .B2(n9399), .A(n9063), .ZN(n9180) );
  INV_X1 U10488 ( .A(n9065), .ZN(n9066) );
  AOI211_X1 U10489 ( .C1(n9182), .C2(n9078), .A(n9101), .B(n9066), .ZN(n9181)
         );
  NAND2_X1 U10490 ( .A1(n9181), .A2(n9440), .ZN(n9069) );
  AOI22_X1 U10491 ( .A1(n9455), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9067), .B2(
        n9447), .ZN(n9068) );
  OAI211_X1 U10492 ( .C1(n9070), .C2(n9104), .A(n9069), .B(n9068), .ZN(n9071)
         );
  AOI21_X1 U10493 ( .B1(n9180), .B2(n9452), .A(n9071), .ZN(n9072) );
  OAI21_X1 U10494 ( .B1(n9184), .B2(n9086), .A(n9072), .ZN(P1_U3274) );
  XNOR2_X1 U10495 ( .A(n4499), .B(n9074), .ZN(n9189) );
  XOR2_X1 U10496 ( .A(n9074), .B(n9073), .Z(n9076) );
  OAI21_X1 U10497 ( .B1(n9076), .B2(n9399), .A(n9075), .ZN(n9185) );
  INV_X1 U10498 ( .A(n9077), .ZN(n9094) );
  INV_X1 U10499 ( .A(n9078), .ZN(n9079) );
  AOI211_X1 U10500 ( .C1(n9187), .C2(n9094), .A(n9101), .B(n9079), .ZN(n9186)
         );
  NAND2_X1 U10501 ( .A1(n9186), .A2(n9440), .ZN(n9082) );
  AOI22_X1 U10502 ( .A1(n9455), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9080), .B2(
        n9447), .ZN(n9081) );
  OAI211_X1 U10503 ( .C1(n9083), .C2(n9104), .A(n9082), .B(n9081), .ZN(n9084)
         );
  AOI21_X1 U10504 ( .B1(n9185), .B2(n9452), .A(n9084), .ZN(n9085) );
  OAI21_X1 U10505 ( .B1(n9189), .B2(n9086), .A(n9085), .ZN(P1_U3275) );
  AOI211_X1 U10506 ( .C1(n9093), .C2(n9088), .A(n9399), .B(n9087), .ZN(n9091)
         );
  INV_X1 U10507 ( .A(n9089), .ZN(n9090) );
  NOR2_X1 U10508 ( .A1(n9091), .A2(n9090), .ZN(n9269) );
  XNOR2_X1 U10509 ( .A(n9092), .B(n9093), .ZN(n9272) );
  NAND2_X1 U10510 ( .A1(n9272), .A2(n9441), .ZN(n9100) );
  OAI211_X1 U10511 ( .C1(n9270), .C2(n4492), .A(n9094), .B(n9436), .ZN(n9268)
         );
  INV_X1 U10512 ( .A(n9268), .ZN(n9098) );
  AOI22_X1 U10513 ( .A1(n9455), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9095), .B2(
        n9447), .ZN(n9096) );
  OAI21_X1 U10514 ( .B1(n9270), .B2(n9104), .A(n9096), .ZN(n9097) );
  AOI21_X1 U10515 ( .B1(n9098), .B2(n9440), .A(n9097), .ZN(n9099) );
  OAI211_X1 U10516 ( .C1(n9455), .C2(n9269), .A(n9100), .B(n9099), .ZN(
        P1_U3276) );
  AOI211_X1 U10517 ( .C1(n9192), .C2(n9102), .A(n9101), .B(n4492), .ZN(n9191)
         );
  AOI22_X1 U10518 ( .A1(n9455), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5023), .B2(
        n9447), .ZN(n9103) );
  OAI21_X1 U10519 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9117) );
  NAND2_X1 U10520 ( .A1(n9108), .A2(n9107), .ZN(n9190) );
  NAND3_X1 U10521 ( .A1(n9106), .A2(n9109), .A3(n9190), .ZN(n9115) );
  XNOR2_X1 U10522 ( .A(n9111), .B(n9110), .ZN(n9114) );
  INV_X1 U10523 ( .A(n9112), .ZN(n9113) );
  AOI21_X1 U10524 ( .B1(n9114), .B2(n9459), .A(n9113), .ZN(n9194) );
  AOI21_X1 U10525 ( .B1(n9115), .B2(n9194), .A(n9455), .ZN(n9116) );
  AOI211_X1 U10526 ( .C1(n9191), .C2(n9440), .A(n9117), .B(n9116), .ZN(n9118)
         );
  INV_X1 U10527 ( .A(n9118), .ZN(P1_U3277) );
  OAI211_X1 U10528 ( .C1(n8856), .C2(n9544), .A(n9119), .B(n9126), .ZN(n9204)
         );
  INV_X1 U10529 ( .A(n9120), .ZN(n9122) );
  NAND2_X1 U10530 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  MUX2_X1 U10531 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9204), .S(n9575), .Z(
        P1_U3553) );
  OAI211_X1 U10532 ( .C1(n9128), .C2(n9544), .A(n9127), .B(n9126), .ZN(n9205)
         );
  MUX2_X1 U10533 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9205), .S(n9575), .Z(
        P1_U3552) );
  OR2_X1 U10534 ( .A1(n9130), .A2(n9129), .ZN(n9509) );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9206), .S(n9575), .Z(
        P1_U3551) );
  AOI21_X1 U10536 ( .B1(n9507), .B2(n9136), .A(n9135), .ZN(n9137) );
  OAI211_X1 U10537 ( .C1(n9139), .C2(n9501), .A(n9138), .B(n9137), .ZN(n9207)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9207), .S(n9575), .Z(
        P1_U3550) );
  OAI211_X1 U10539 ( .C1(n9144), .C2(n9501), .A(n9143), .B(n9142), .ZN(n9208)
         );
  MUX2_X1 U10540 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9208), .S(n9575), .Z(
        P1_U3549) );
  AOI21_X1 U10541 ( .B1(n9507), .B2(n9146), .A(n9145), .ZN(n9147) );
  OAI211_X1 U10542 ( .C1(n9149), .C2(n9501), .A(n9148), .B(n9147), .ZN(n9209)
         );
  MUX2_X1 U10543 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9209), .S(n9575), .Z(
        P1_U3548) );
  AOI211_X1 U10544 ( .C1(n9507), .C2(n9152), .A(n9151), .B(n9150), .ZN(n9153)
         );
  OAI21_X1 U10545 ( .B1(n9154), .B2(n9501), .A(n9153), .ZN(n9210) );
  MUX2_X1 U10546 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9210), .S(n9575), .Z(
        P1_U3547) );
  AOI211_X1 U10547 ( .C1(n9507), .C2(n9157), .A(n9156), .B(n9155), .ZN(n9158)
         );
  OAI21_X1 U10548 ( .B1(n9159), .B2(n9501), .A(n9158), .ZN(n9211) );
  MUX2_X1 U10549 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9211), .S(n9575), .Z(
        P1_U3546) );
  AOI21_X1 U10550 ( .B1(n9507), .B2(n9161), .A(n9160), .ZN(n9162) );
  OAI211_X1 U10551 ( .C1(n9164), .C2(n9501), .A(n9163), .B(n9162), .ZN(n9212)
         );
  MUX2_X1 U10552 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9212), .S(n9575), .Z(
        P1_U3545) );
  AOI211_X1 U10553 ( .C1(n9507), .C2(n9167), .A(n9166), .B(n9165), .ZN(n9168)
         );
  OAI21_X1 U10554 ( .B1(n9169), .B2(n9501), .A(n9168), .ZN(n9213) );
  MUX2_X1 U10555 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9213), .S(n9575), .Z(
        P1_U3544) );
  AOI211_X1 U10556 ( .C1(n9507), .C2(n9172), .A(n9171), .B(n9170), .ZN(n9173)
         );
  OAI21_X1 U10557 ( .B1(n9174), .B2(n9501), .A(n9173), .ZN(n9214) );
  MUX2_X1 U10558 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9214), .S(n9575), .Z(
        P1_U3543) );
  AOI211_X1 U10559 ( .C1(n9507), .C2(n9177), .A(n9176), .B(n9175), .ZN(n9178)
         );
  OAI21_X1 U10560 ( .B1(n9179), .B2(n9501), .A(n9178), .ZN(n9215) );
  MUX2_X1 U10561 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9215), .S(n9575), .Z(
        P1_U3542) );
  AOI211_X1 U10562 ( .C1(n9507), .C2(n9182), .A(n9181), .B(n9180), .ZN(n9183)
         );
  OAI21_X1 U10563 ( .B1(n9184), .B2(n9501), .A(n9183), .ZN(n9216) );
  MUX2_X1 U10564 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9216), .S(n9575), .Z(
        P1_U3541) );
  AOI211_X1 U10565 ( .C1(n9507), .C2(n9187), .A(n9186), .B(n9185), .ZN(n9188)
         );
  OAI21_X1 U10566 ( .B1(n9189), .B2(n9501), .A(n9188), .ZN(n9217) );
  MUX2_X1 U10567 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9217), .S(n9575), .Z(
        P1_U3540) );
  NAND2_X1 U10568 ( .A1(n9190), .A2(n9541), .ZN(n9195) );
  AOI21_X1 U10569 ( .B1(n9507), .B2(n9192), .A(n9191), .ZN(n9193) );
  OAI211_X1 U10570 ( .C1(n9196), .C2(n9195), .A(n9194), .B(n9193), .ZN(n9218)
         );
  MUX2_X1 U10571 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9218), .S(n9575), .Z(
        P1_U3538) );
  AOI211_X1 U10572 ( .C1(n9507), .C2(n9199), .A(n9198), .B(n9197), .ZN(n9200)
         );
  OAI21_X1 U10573 ( .B1(n9201), .B2(n9501), .A(n9200), .ZN(n9219) );
  MUX2_X1 U10574 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9219), .S(n9575), .Z(
        P1_U3535) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9204), .S(n9553), .Z(
        P1_U3521) );
  MUX2_X1 U10576 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9205), .S(n9553), .Z(
        P1_U3520) );
  MUX2_X1 U10577 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9206), .S(n9553), .Z(
        P1_U3519) );
  MUX2_X1 U10578 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9207), .S(n9553), .Z(
        P1_U3518) );
  MUX2_X1 U10579 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9208), .S(n9553), .Z(
        P1_U3517) );
  MUX2_X1 U10580 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9209), .S(n9553), .Z(
        P1_U3516) );
  MUX2_X1 U10581 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9210), .S(n9553), .Z(
        P1_U3515) );
  MUX2_X1 U10582 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9211), .S(n9553), .Z(
        P1_U3514) );
  MUX2_X1 U10583 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9212), .S(n9553), .Z(
        P1_U3513) );
  MUX2_X1 U10584 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9213), .S(n9553), .Z(
        P1_U3512) );
  MUX2_X1 U10585 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9214), .S(n9553), .Z(
        P1_U3511) );
  MUX2_X1 U10586 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9215), .S(n9553), .Z(
        P1_U3510) );
  MUX2_X1 U10587 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9216), .S(n9553), .Z(
        P1_U3509) );
  MUX2_X1 U10588 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9217), .S(n9553), .Z(
        P1_U3507) );
  MUX2_X1 U10589 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9218), .S(n9553), .Z(
        P1_U3501) );
  MUX2_X1 U10590 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9219), .S(n9553), .Z(
        P1_U3492) );
  NOR2_X1 U10591 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n9222) );
  NAND4_X1 U10592 ( .A1(n9222), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .A4(n9221), .ZN(n9224) );
  OAI22_X1 U10593 ( .A1(n9220), .A2(n9224), .B1(n9223), .B2(n7620), .ZN(n9225)
         );
  AOI21_X1 U10594 ( .B1(n9227), .B2(n9226), .A(n9225), .ZN(n9228) );
  INV_X1 U10595 ( .A(n9228), .ZN(P1_U3324) );
  OAI222_X1 U10596 ( .A1(n7569), .A2(n9230), .B1(n4421), .B2(P1_U3086), .C1(
        n9229), .C2(n7620), .ZN(P1_U3328) );
  OAI222_X1 U10597 ( .A1(n7569), .A2(n9233), .B1(n9232), .B2(P1_U3086), .C1(
        n9231), .C2(n7620), .ZN(P1_U3329) );
  OAI222_X1 U10598 ( .A1(n7569), .A2(n9236), .B1(n9235), .B2(P1_U3086), .C1(
        n9234), .C2(n7620), .ZN(P1_U3330) );
  MUX2_X1 U10599 ( .A(n9237), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10600 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U10601 ( .A1(n9239), .A2(n9238), .ZN(n9242) );
  INV_X1 U10602 ( .A(n9240), .ZN(n9241) );
  NAND3_X1 U10603 ( .A1(n9379), .A2(n9242), .A3(n9241), .ZN(n9248) );
  AOI21_X1 U10604 ( .B1(n9245), .B2(n9244), .A(n9243), .ZN(n9246) );
  NAND2_X1 U10605 ( .A1(n9383), .A2(n9246), .ZN(n9247) );
  OAI211_X1 U10606 ( .C1(n9389), .C2(n9249), .A(n9248), .B(n9247), .ZN(n9250)
         );
  INV_X1 U10607 ( .A(n9250), .ZN(n9252) );
  OAI211_X1 U10608 ( .C1(n9393), .C2(n9253), .A(n9252), .B(n9251), .ZN(
        P1_U3253) );
  NOR2_X1 U10609 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10006), .ZN(n9303) );
  INV_X1 U10610 ( .A(n9303), .ZN(n9254) );
  OAI21_X1 U10611 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9263) );
  AOI21_X1 U10612 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(n9261) );
  NOR2_X1 U10613 ( .A1(n9261), .A2(n9260), .ZN(n9262) );
  AOI211_X1 U10614 ( .C1(n9264), .C2(n5768), .A(n9263), .B(n9262), .ZN(n9265)
         );
  OAI21_X1 U10615 ( .B1(n9267), .B2(n9266), .A(n9265), .ZN(P1_U3236) );
  OAI211_X1 U10616 ( .C1(n9270), .C2(n9544), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U10617 ( .B1(n9272), .B2(n9541), .A(n9271), .ZN(n9280) );
  INV_X1 U10618 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9273) );
  AOI22_X1 U10619 ( .A1(n9575), .A2(n9280), .B1(n9273), .B2(n9573), .ZN(
        P1_U3539) );
  OAI211_X1 U10620 ( .C1(n9276), .C2(n9544), .A(n9275), .B(n9274), .ZN(n9277)
         );
  AOI21_X1 U10621 ( .B1(n9278), .B2(n9541), .A(n9277), .ZN(n9282) );
  AOI22_X1 U10622 ( .A1(n9575), .A2(n9282), .B1(n10101), .B2(n9573), .ZN(
        P1_U3537) );
  INV_X1 U10623 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9279) );
  AOI22_X1 U10624 ( .A1(n9553), .A2(n9280), .B1(n9279), .B2(n9551), .ZN(
        P1_U3504) );
  INV_X1 U10625 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9281) );
  AOI22_X1 U10626 ( .A1(n9553), .A2(n9282), .B1(n9281), .B2(n9551), .ZN(
        P1_U3498) );
  XNOR2_X1 U10627 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10628 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10629 ( .A(n9283), .ZN(n9288) );
  INV_X1 U10630 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U10631 ( .A1(n4421), .A2(n9554), .ZN(n9286) );
  NAND2_X1 U10632 ( .A1(n9284), .A2(n9286), .ZN(n9285) );
  MUX2_X1 U10633 ( .A(n9286), .B(n9285), .S(P1_IR_REG_0__SCAN_IN), .Z(n9287)
         );
  NAND2_X1 U10634 ( .A1(n9288), .A2(n9287), .ZN(n9290) );
  AOI22_X1 U10635 ( .A1(n9305), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9289) );
  OAI21_X1 U10636 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(P1_U3243) );
  AOI211_X1 U10637 ( .C1(n9294), .C2(n9293), .A(n9292), .B(n9368), .ZN(n9300)
         );
  AOI211_X1 U10638 ( .C1(n9298), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9299)
         );
  AOI211_X1 U10639 ( .C1(n9347), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9302)
         );
  INV_X1 U10640 ( .A(n9302), .ZN(n9304) );
  AOI211_X1 U10641 ( .C1(n9305), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9304), .B(
        n9303), .ZN(n9306) );
  INV_X1 U10642 ( .A(n9306), .ZN(P1_U3254) );
  INV_X1 U10643 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9321) );
  OAI21_X1 U10644 ( .B1(n9309), .B2(n9308), .A(n9307), .ZN(n9310) );
  NAND2_X1 U10645 ( .A1(n9379), .A2(n9310), .ZN(n9316) );
  OAI21_X1 U10646 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9314) );
  NAND2_X1 U10647 ( .A1(n9383), .A2(n9314), .ZN(n9315) );
  OAI211_X1 U10648 ( .C1(n9389), .C2(n9317), .A(n9316), .B(n9315), .ZN(n9318)
         );
  INV_X1 U10649 ( .A(n9318), .ZN(n9320) );
  OAI211_X1 U10650 ( .C1(n9321), .C2(n9393), .A(n9320), .B(n9319), .ZN(
        P1_U3255) );
  INV_X1 U10651 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9336) );
  AOI21_X1 U10652 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9325) );
  NAND2_X1 U10653 ( .A1(n9379), .A2(n9325), .ZN(n9331) );
  AOI21_X1 U10654 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9329) );
  NAND2_X1 U10655 ( .A1(n9383), .A2(n9329), .ZN(n9330) );
  OAI211_X1 U10656 ( .C1(n9389), .C2(n9332), .A(n9331), .B(n9330), .ZN(n9333)
         );
  INV_X1 U10657 ( .A(n9333), .ZN(n9335) );
  OAI211_X1 U10658 ( .C1(n9393), .C2(n9336), .A(n9335), .B(n9334), .ZN(
        P1_U3256) );
  INV_X1 U10659 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9350) );
  OAI211_X1 U10660 ( .C1(n9339), .C2(n9338), .A(n9379), .B(n9337), .ZN(n9340)
         );
  INV_X1 U10661 ( .A(n9340), .ZN(n9345) );
  AOI211_X1 U10662 ( .C1(n9343), .C2(n9342), .A(n9341), .B(n9368), .ZN(n9344)
         );
  AOI211_X1 U10663 ( .C1(n9347), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9349)
         );
  NAND2_X1 U10664 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9348) );
  OAI211_X1 U10665 ( .C1(n9393), .C2(n9350), .A(n9349), .B(n9348), .ZN(
        P1_U3257) );
  INV_X1 U10666 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9363) );
  AOI21_X1 U10667 ( .B1(n9352), .B2(n10101), .A(n9351), .ZN(n9353) );
  NAND2_X1 U10668 ( .A1(n9379), .A2(n9353), .ZN(n9358) );
  AOI21_X1 U10669 ( .B1(n9355), .B2(n10022), .A(n9354), .ZN(n9356) );
  NAND2_X1 U10670 ( .A1(n9383), .A2(n9356), .ZN(n9357) );
  OAI211_X1 U10671 ( .C1(n9389), .C2(n9359), .A(n9358), .B(n9357), .ZN(n9360)
         );
  INV_X1 U10672 ( .A(n9360), .ZN(n9362) );
  OAI211_X1 U10673 ( .C1(n9363), .C2(n9393), .A(n9362), .B(n9361), .ZN(
        P1_U3258) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9377) );
  OAI21_X1 U10675 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9374) );
  NOR2_X1 U10676 ( .A1(n9389), .A2(n9367), .ZN(n9373) );
  AOI211_X1 U10677 ( .C1(n9371), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9372)
         );
  AOI211_X1 U10678 ( .C1(n9379), .C2(n9374), .A(n9373), .B(n9372), .ZN(n9376)
         );
  OAI211_X1 U10679 ( .C1(n9393), .C2(n9377), .A(n9376), .B(n9375), .ZN(
        P1_U3259) );
  OAI211_X1 U10680 ( .C1(n9381), .C2(n9380), .A(n9379), .B(n9378), .ZN(n9387)
         );
  OAI211_X1 U10681 ( .C1(n9385), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9386)
         );
  OAI211_X1 U10682 ( .C1(n9389), .C2(n9388), .A(n9387), .B(n9386), .ZN(n9390)
         );
  INV_X1 U10683 ( .A(n9390), .ZN(n9392) );
  NAND2_X1 U10684 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9391) );
  OAI211_X1 U10685 ( .C1(n9393), .C2(n9861), .A(n9392), .B(n9391), .ZN(
        P1_U3261) );
  XNOR2_X1 U10686 ( .A(n9394), .B(n9401), .ZN(n9549) );
  NAND2_X1 U10687 ( .A1(n9396), .A2(n9395), .ZN(n9400) );
  INV_X1 U10688 ( .A(n9397), .ZN(n9398) );
  AOI211_X1 U10689 ( .C1(n9401), .C2(n9400), .A(n9399), .B(n9398), .ZN(n9404)
         );
  INV_X1 U10690 ( .A(n9402), .ZN(n9403) );
  AOI211_X1 U10691 ( .C1(n9549), .C2(n9513), .A(n9404), .B(n9403), .ZN(n9546)
         );
  AOI222_X1 U10692 ( .A1(n9406), .A2(n9431), .B1(n9405), .B2(n9447), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(n9455), .ZN(n9411) );
  OAI211_X1 U10693 ( .C1(n9408), .C2(n9545), .A(n9436), .B(n9407), .ZN(n9543)
         );
  INV_X1 U10694 ( .A(n9543), .ZN(n9409) );
  AOI22_X1 U10695 ( .A1(n9549), .A2(n9424), .B1(n9440), .B2(n9409), .ZN(n9410)
         );
  OAI211_X1 U10696 ( .C1(n9455), .C2(n9546), .A(n9411), .B(n9410), .ZN(
        P1_U3279) );
  OAI21_X1 U10697 ( .B1(n4941), .B2(n9413), .A(n9412), .ZN(n9418) );
  XNOR2_X1 U10698 ( .A(n9414), .B(n4941), .ZN(n9421) );
  NOR2_X1 U10699 ( .A1(n9421), .A2(n9415), .ZN(n9416) );
  AOI211_X1 U10700 ( .C1(n9418), .C2(n9459), .A(n9417), .B(n9416), .ZN(n9516)
         );
  AOI222_X1 U10701 ( .A1(n9420), .A2(n9431), .B1(n9419), .B2(n9447), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n9455), .ZN(n9426) );
  INV_X1 U10702 ( .A(n9421), .ZN(n9519) );
  OAI211_X1 U10703 ( .C1(n4639), .C2(n9515), .A(n9436), .B(n9422), .ZN(n9514)
         );
  INV_X1 U10704 ( .A(n9514), .ZN(n9423) );
  AOI22_X1 U10705 ( .A1(n9519), .A2(n9424), .B1(n9440), .B2(n9423), .ZN(n9425)
         );
  OAI211_X1 U10706 ( .C1(n9455), .C2(n9516), .A(n9426), .B(n9425), .ZN(
        P1_U3285) );
  XNOR2_X1 U10707 ( .A(n9427), .B(n9434), .ZN(n9429) );
  AOI21_X1 U10708 ( .B1(n9429), .B2(n9459), .A(n9428), .ZN(n9485) );
  AOI222_X1 U10709 ( .A1(n9432), .A2(n9431), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9455), .C1(n9447), .C2(n9430), .ZN(n9443) );
  XNOR2_X1 U10710 ( .A(n9433), .B(n9434), .ZN(n9488) );
  INV_X1 U10711 ( .A(n9435), .ZN(n9437) );
  OAI211_X1 U10712 ( .C1(n9484), .C2(n9438), .A(n9437), .B(n9436), .ZN(n9483)
         );
  INV_X1 U10713 ( .A(n9483), .ZN(n9439) );
  AOI22_X1 U10714 ( .A1(n9488), .A2(n9441), .B1(n9440), .B2(n9439), .ZN(n9442)
         );
  OAI211_X1 U10715 ( .C1(n9455), .C2(n9485), .A(n9443), .B(n9442), .ZN(
        P1_U3289) );
  INV_X1 U10716 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9454) );
  INV_X1 U10717 ( .A(n9444), .ZN(n9451) );
  NAND2_X1 U10718 ( .A1(n9446), .A2(n9445), .ZN(n9460) );
  NAND2_X1 U10719 ( .A1(n9447), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9448) );
  OAI211_X1 U10720 ( .C1(n9449), .C2(n9460), .A(n9461), .B(n9448), .ZN(n9450)
         );
  AOI21_X1 U10721 ( .B1(n9458), .B2(n9451), .A(n9450), .ZN(n9453) );
  AOI22_X1 U10722 ( .A1(n9455), .A2(n9454), .B1(n9453), .B2(n9452), .ZN(
        P1_U3293) );
  AND2_X1 U10723 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9457), .ZN(P1_U3294) );
  AND2_X1 U10724 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9457), .ZN(P1_U3295) );
  AND2_X1 U10725 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9457), .ZN(P1_U3296) );
  AND2_X1 U10726 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9457), .ZN(P1_U3297) );
  AND2_X1 U10727 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9457), .ZN(P1_U3298) );
  INV_X1 U10728 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U10729 ( .A1(n9456), .A2(n9942), .ZN(P1_U3299) );
  INV_X1 U10730 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U10731 ( .A1(n9456), .A2(n10067), .ZN(P1_U3300) );
  AND2_X1 U10732 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9457), .ZN(P1_U3301) );
  AND2_X1 U10733 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9457), .ZN(P1_U3302) );
  INV_X1 U10734 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10124) );
  NOR2_X1 U10735 ( .A1(n9456), .A2(n10124), .ZN(P1_U3303) );
  INV_X1 U10736 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U10737 ( .A1(n9456), .A2(n10116), .ZN(P1_U3304) );
  AND2_X1 U10738 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9457), .ZN(P1_U3305) );
  AND2_X1 U10739 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9457), .ZN(P1_U3306) );
  AND2_X1 U10740 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9457), .ZN(P1_U3307) );
  AND2_X1 U10741 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9457), .ZN(P1_U3308) );
  AND2_X1 U10742 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9457), .ZN(P1_U3309) );
  AND2_X1 U10743 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9457), .ZN(P1_U3310) );
  AND2_X1 U10744 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9457), .ZN(P1_U3311) );
  AND2_X1 U10745 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9457), .ZN(P1_U3312) );
  INV_X1 U10746 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U10747 ( .A1(n9456), .A2(n9984), .ZN(P1_U3313) );
  AND2_X1 U10748 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9457), .ZN(P1_U3314) );
  AND2_X1 U10749 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9457), .ZN(P1_U3315) );
  AND2_X1 U10750 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9457), .ZN(P1_U3316) );
  AND2_X1 U10751 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9457), .ZN(P1_U3317) );
  AND2_X1 U10752 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9457), .ZN(P1_U3318) );
  AND2_X1 U10753 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9457), .ZN(P1_U3319) );
  AND2_X1 U10754 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9457), .ZN(P1_U3320) );
  INV_X1 U10755 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U10756 ( .A1(n9456), .A2(n10009), .ZN(P1_U3321) );
  AND2_X1 U10757 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9457), .ZN(P1_U3322) );
  AND2_X1 U10758 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9457), .ZN(P1_U3323) );
  OAI21_X1 U10759 ( .B1(n9541), .B2(n9459), .A(n9458), .ZN(n9462) );
  AND3_X1 U10760 ( .A1(n9462), .A2(n9461), .A3(n9460), .ZN(n9555) );
  INV_X1 U10761 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U10762 ( .A1(n9553), .A2(n9555), .B1(n10005), .B2(n9551), .ZN(
        P1_U3453) );
  INV_X1 U10763 ( .A(n9509), .ZN(n9550) );
  OAI21_X1 U10764 ( .B1(n9464), .B2(n9544), .A(n9463), .ZN(n9465) );
  AOI21_X1 U10765 ( .B1(n9466), .B2(n9550), .A(n9465), .ZN(n9467) );
  AND2_X1 U10766 ( .A1(n9468), .A2(n9467), .ZN(n9556) );
  INV_X1 U10767 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U10768 ( .A1(n9553), .A2(n9556), .B1(n9469), .B2(n9551), .ZN(
        P1_U3456) );
  INV_X1 U10769 ( .A(n9470), .ZN(n9475) );
  OAI21_X1 U10770 ( .B1(n9472), .B2(n9544), .A(n9471), .ZN(n9474) );
  AOI211_X1 U10771 ( .C1(n9475), .C2(n9541), .A(n9474), .B(n9473), .ZN(n9558)
         );
  INV_X1 U10772 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U10773 ( .A1(n9553), .A2(n9558), .B1(n9476), .B2(n9551), .ZN(
        P1_U3459) );
  AOI21_X1 U10774 ( .B1(n9507), .B2(n9478), .A(n9477), .ZN(n9479) );
  OAI211_X1 U10775 ( .C1(n9481), .C2(n9501), .A(n9480), .B(n9479), .ZN(n9482)
         );
  INV_X1 U10776 ( .A(n9482), .ZN(n9559) );
  INV_X1 U10777 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U10778 ( .A1(n9553), .A2(n9559), .B1(n10068), .B2(n9551), .ZN(
        P1_U3462) );
  OAI21_X1 U10779 ( .B1(n9484), .B2(n9544), .A(n9483), .ZN(n9487) );
  INV_X1 U10780 ( .A(n9485), .ZN(n9486) );
  AOI211_X1 U10781 ( .C1(n9541), .C2(n9488), .A(n9487), .B(n9486), .ZN(n9561)
         );
  INV_X1 U10782 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9489) );
  AOI22_X1 U10783 ( .A1(n9553), .A2(n9561), .B1(n9489), .B2(n9551), .ZN(
        P1_U3465) );
  AND2_X1 U10784 ( .A1(n9490), .A2(n9541), .ZN(n9494) );
  OAI21_X1 U10785 ( .B1(n9492), .B2(n9544), .A(n9491), .ZN(n9493) );
  NOR3_X1 U10786 ( .A1(n9495), .A2(n9494), .A3(n9493), .ZN(n9562) );
  INV_X1 U10787 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U10788 ( .A1(n9553), .A2(n9562), .B1(n10047), .B2(n9551), .ZN(
        P1_U3468) );
  AOI21_X1 U10789 ( .B1(n9507), .B2(n9497), .A(n9496), .ZN(n9498) );
  OAI211_X1 U10790 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9502)
         );
  INV_X1 U10791 ( .A(n9502), .ZN(n9564) );
  INV_X1 U10792 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9503) );
  AOI22_X1 U10793 ( .A1(n9553), .A2(n9564), .B1(n9503), .B2(n9551), .ZN(
        P1_U3471) );
  INV_X1 U10794 ( .A(n9510), .ZN(n9512) );
  AOI211_X1 U10795 ( .C1(n9507), .C2(n9506), .A(n9505), .B(n9504), .ZN(n9508)
         );
  OAI21_X1 U10796 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9511) );
  AOI21_X1 U10797 ( .B1(n9513), .B2(n9512), .A(n9511), .ZN(n9565) );
  INV_X1 U10798 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U10799 ( .A1(n9553), .A2(n9565), .B1(n9988), .B2(n9551), .ZN(
        P1_U3474) );
  OAI21_X1 U10800 ( .B1(n9515), .B2(n9544), .A(n9514), .ZN(n9518) );
  INV_X1 U10801 ( .A(n9516), .ZN(n9517) );
  AOI211_X1 U10802 ( .C1(n9550), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9567)
         );
  INV_X1 U10803 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U10804 ( .A1(n9553), .A2(n9567), .B1(n10153), .B2(n9551), .ZN(
        P1_U3477) );
  OAI21_X1 U10805 ( .B1(n9521), .B2(n9544), .A(n9520), .ZN(n9523) );
  AOI211_X1 U10806 ( .C1(n9541), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9568)
         );
  INV_X1 U10807 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U10808 ( .A1(n9553), .A2(n9568), .B1(n9944), .B2(n9551), .ZN(
        P1_U3480) );
  OAI211_X1 U10809 ( .C1(n9527), .C2(n9544), .A(n9526), .B(n9525), .ZN(n9528)
         );
  AOI21_X1 U10810 ( .B1(n9541), .B2(n9529), .A(n9528), .ZN(n9569) );
  INV_X1 U10811 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9530) );
  AOI22_X1 U10812 ( .A1(n9553), .A2(n9569), .B1(n9530), .B2(n9551), .ZN(
        P1_U3483) );
  OAI21_X1 U10813 ( .B1(n9532), .B2(n9544), .A(n9531), .ZN(n9533) );
  AOI21_X1 U10814 ( .B1(n9534), .B2(n9550), .A(n9533), .ZN(n9535) );
  AND2_X1 U10815 ( .A1(n9536), .A2(n9535), .ZN(n9571) );
  INV_X1 U10816 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10023) );
  AOI22_X1 U10817 ( .A1(n9553), .A2(n9571), .B1(n10023), .B2(n9551), .ZN(
        P1_U3486) );
  OAI21_X1 U10818 ( .B1(n9538), .B2(n9544), .A(n9537), .ZN(n9539) );
  AOI211_X1 U10819 ( .C1(n9542), .C2(n9541), .A(n9540), .B(n9539), .ZN(n9572)
         );
  INV_X1 U10820 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U10821 ( .A1(n9553), .A2(n9572), .B1(n10119), .B2(n9551), .ZN(
        P1_U3489) );
  OAI21_X1 U10822 ( .B1(n9545), .B2(n9544), .A(n9543), .ZN(n9548) );
  INV_X1 U10823 ( .A(n9546), .ZN(n9547) );
  AOI211_X1 U10824 ( .C1(n9550), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9574)
         );
  INV_X1 U10825 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10826 ( .A1(n9553), .A2(n9574), .B1(n9552), .B2(n9551), .ZN(
        P1_U3495) );
  AOI22_X1 U10827 ( .A1(n9575), .A2(n9555), .B1(n9554), .B2(n9573), .ZN(
        P1_U3522) );
  AOI22_X1 U10828 ( .A1(n9575), .A2(n9556), .B1(n10181), .B2(n9573), .ZN(
        P1_U3523) );
  INV_X1 U10829 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10830 ( .A1(n9575), .A2(n9558), .B1(n9557), .B2(n9573), .ZN(
        P1_U3524) );
  AOI22_X1 U10831 ( .A1(n9575), .A2(n9559), .B1(n6448), .B2(n9573), .ZN(
        P1_U3525) );
  AOI22_X1 U10832 ( .A1(n9575), .A2(n9561), .B1(n9560), .B2(n9573), .ZN(
        P1_U3526) );
  AOI22_X1 U10833 ( .A1(n9575), .A2(n9562), .B1(n6452), .B2(n9573), .ZN(
        P1_U3527) );
  AOI22_X1 U10834 ( .A1(n9575), .A2(n9564), .B1(n9563), .B2(n9573), .ZN(
        P1_U3528) );
  AOI22_X1 U10835 ( .A1(n9575), .A2(n9565), .B1(n6455), .B2(n9573), .ZN(
        P1_U3529) );
  AOI22_X1 U10836 ( .A1(n9575), .A2(n9567), .B1(n9566), .B2(n9573), .ZN(
        P1_U3530) );
  AOI22_X1 U10837 ( .A1(n9575), .A2(n9568), .B1(n10031), .B2(n9573), .ZN(
        P1_U3531) );
  AOI22_X1 U10838 ( .A1(n9575), .A2(n9569), .B1(n8800), .B2(n9573), .ZN(
        P1_U3532) );
  AOI22_X1 U10839 ( .A1(n9575), .A2(n9571), .B1(n9570), .B2(n9573), .ZN(
        P1_U3533) );
  AOI22_X1 U10840 ( .A1(n9575), .A2(n9572), .B1(n8804), .B2(n9573), .ZN(
        P1_U3534) );
  AOI22_X1 U10841 ( .A1(n9575), .A2(n9574), .B1(n8798), .B2(n9573), .ZN(
        P1_U3536) );
  INV_X1 U10842 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9595) );
  XOR2_X1 U10843 ( .A(n9577), .B(n9576), .Z(n9593) );
  OAI21_X1 U10844 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(n9588) );
  INV_X1 U10845 ( .A(n9581), .ZN(n9583) );
  NAND3_X1 U10846 ( .A1(n9584), .A2(n9583), .A3(n9582), .ZN(n9585) );
  AOI21_X1 U10847 ( .B1(n9586), .B2(n9585), .A(n10220), .ZN(n9587) );
  AOI21_X1 U10848 ( .B1(n10223), .B2(n9588), .A(n9587), .ZN(n9590) );
  OAI211_X1 U10849 ( .C1(n9754), .C2(n9591), .A(n9590), .B(n9589), .ZN(n9592)
         );
  AOI21_X1 U10850 ( .B1(n9593), .B2(n10207), .A(n9592), .ZN(n9594) );
  OAI21_X1 U10851 ( .B1(n10217), .B2(n9595), .A(n9594), .ZN(P2_U3186) );
  INV_X1 U10852 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9613) );
  AOI211_X1 U10853 ( .C1(n9599), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9611)
         );
  NOR2_X1 U10854 ( .A1(n9754), .A2(n9600), .ZN(n9609) );
  XOR2_X1 U10855 ( .A(n9601), .B(P2_REG1_REG_5__SCAN_IN), .Z(n9606) );
  INV_X1 U10856 ( .A(n9602), .ZN(n9603) );
  AOI21_X1 U10857 ( .B1(n5880), .B2(n9604), .A(n9603), .ZN(n9605) );
  OAI22_X1 U10858 ( .A1(n9607), .A2(n9606), .B1(n9605), .B2(n10220), .ZN(n9608) );
  NOR4_X1 U10859 ( .A1(n9611), .A2(n9610), .A3(n9609), .A4(n9608), .ZN(n9612)
         );
  OAI21_X1 U10860 ( .B1(n10217), .B2(n9613), .A(n9612), .ZN(P2_U3187) );
  AOI22_X1 U10861 ( .A1(n9614), .A2(n10209), .B1(P2_ADDR_REG_9__SCAN_IN), .B2(
        n9740), .ZN(n9628) );
  OAI21_X1 U10862 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9621) );
  OAI21_X1 U10863 ( .B1(n9619), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9618), .ZN(
        n9620) );
  AOI22_X1 U10864 ( .A1(n9621), .A2(n10207), .B1(n10223), .B2(n9620), .ZN(
        n9627) );
  AOI21_X1 U10865 ( .B1(n5946), .B2(n9623), .A(n9622), .ZN(n9624) );
  OR2_X1 U10866 ( .A1(n9624), .A2(n10220), .ZN(n9625) );
  NAND4_X1 U10867 ( .A1(n9628), .A2(n9627), .A3(n9626), .A4(n9625), .ZN(
        P2_U3191) );
  AOI22_X1 U10868 ( .A1(n9629), .A2(n10209), .B1(n9740), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n9645) );
  OAI21_X1 U10869 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9637) );
  OAI21_X1 U10870 ( .B1(n9635), .B2(n9634), .A(n9633), .ZN(n9636) );
  AOI22_X1 U10871 ( .A1(n9637), .A2(n10223), .B1(n10207), .B2(n9636), .ZN(
        n9644) );
  AOI21_X1 U10872 ( .B1(n9640), .B2(n9639), .A(n9638), .ZN(n9641) );
  OR2_X1 U10873 ( .A1(n9641), .A2(n10220), .ZN(n9642) );
  NAND4_X1 U10874 ( .A1(n9645), .A2(n9644), .A3(n9643), .A4(n9642), .ZN(
        P2_U3192) );
  AOI22_X1 U10875 ( .A1(n9646), .A2(n10209), .B1(n9740), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n9660) );
  OAI21_X1 U10876 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9648), .A(n9647), .ZN(
        n9653) );
  OAI21_X1 U10877 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9652) );
  AOI22_X1 U10878 ( .A1(n9653), .A2(n10223), .B1(n10207), .B2(n9652), .ZN(
        n9659) );
  AOI21_X1 U10879 ( .B1(n9655), .B2(n5978), .A(n9654), .ZN(n9656) );
  OR2_X1 U10880 ( .A1(n10220), .A2(n9656), .ZN(n9657) );
  NAND4_X1 U10881 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(
        P2_U3193) );
  AOI22_X1 U10882 ( .A1(n9661), .A2(n10209), .B1(n9740), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9678) );
  OAI21_X1 U10883 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9669) );
  OAI21_X1 U10884 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9668) );
  AOI22_X1 U10885 ( .A1(n9669), .A2(n10223), .B1(n10207), .B2(n9668), .ZN(
        n9677) );
  INV_X1 U10886 ( .A(n9670), .ZN(n9676) );
  AOI21_X1 U10887 ( .B1(n9673), .B2(n9672), .A(n9671), .ZN(n9674) );
  OR2_X1 U10888 ( .A1(n9674), .A2(n10220), .ZN(n9675) );
  NAND4_X1 U10889 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(
        P2_U3194) );
  AOI22_X1 U10890 ( .A1(n9679), .A2(n10209), .B1(n9740), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9693) );
  OAI21_X1 U10891 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9681), .A(n9680), .ZN(
        n9686) );
  OAI21_X1 U10892 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9685) );
  AOI22_X1 U10893 ( .A1(n9686), .A2(n10223), .B1(n10207), .B2(n9685), .ZN(
        n9692) );
  NAND2_X1 U10894 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n9691) );
  AOI21_X1 U10895 ( .B1(n9688), .B2(n6010), .A(n9687), .ZN(n9689) );
  OR2_X1 U10896 ( .A1(n10220), .A2(n9689), .ZN(n9690) );
  NAND4_X1 U10897 ( .A1(n9693), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(
        P2_U3195) );
  AOI22_X1 U10898 ( .A1(n9740), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n9694), .B2(
        n10209), .ZN(n9710) );
  XNOR2_X1 U10899 ( .A(n9696), .B(n9695), .ZN(n9701) );
  OAI21_X1 U10900 ( .B1(n9699), .B2(n9698), .A(n9697), .ZN(n9700) );
  AOI22_X1 U10901 ( .A1(n9701), .A2(n10223), .B1(n10207), .B2(n9700), .ZN(
        n9709) );
  NAND2_X1 U10902 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9708) );
  AOI21_X1 U10903 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9703), .A(n9702), .ZN(
        n9705) );
  XOR2_X1 U10904 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND2_X1 U10905 ( .A1(n9706), .A2(n9749), .ZN(n9707) );
  NAND4_X1 U10906 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(
        P2_U3196) );
  AOI21_X1 U10907 ( .B1(n9740), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n9711), .ZN(
        n9722) );
  OAI21_X1 U10908 ( .B1(n9713), .B2(P2_REG1_REG_15__SCAN_IN), .A(n9712), .ZN(
        n9720) );
  OAI21_X1 U10909 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n9715), .A(n9714), .ZN(
        n9719) );
  XNOR2_X1 U10910 ( .A(n9717), .B(n9716), .ZN(n9718) );
  AOI222_X1 U10911 ( .A1(n9720), .A2(n10223), .B1(n9749), .B2(n9719), .C1(
        n9718), .C2(n10207), .ZN(n9721) );
  OAI211_X1 U10912 ( .C1(n9754), .C2(n9723), .A(n9722), .B(n9721), .ZN(
        P2_U3197) );
  AOI21_X1 U10913 ( .B1(n9740), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9724), .ZN(
        n9737) );
  OAI21_X1 U10914 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9735) );
  XNOR2_X1 U10915 ( .A(n9729), .B(n9728), .ZN(n9734) );
  OAI21_X1 U10916 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  AOI222_X1 U10917 ( .A1(n9735), .A2(n10223), .B1(n10207), .B2(n9734), .C1(
        n9749), .C2(n9733), .ZN(n9736) );
  OAI211_X1 U10918 ( .C1(n9754), .C2(n9738), .A(n9737), .B(n9736), .ZN(
        P2_U3198) );
  AOI21_X1 U10919 ( .B1(n9740), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9739), .ZN(
        n9752) );
  OAI21_X1 U10920 ( .B1(n9742), .B2(P2_REG1_REG_17__SCAN_IN), .A(n9741), .ZN(
        n9750) );
  OAI21_X1 U10921 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9744), .A(n9743), .ZN(
        n9748) );
  XNOR2_X1 U10922 ( .A(n9746), .B(n9745), .ZN(n9747) );
  AOI222_X1 U10923 ( .A1(n9750), .A2(n10223), .B1(n9749), .B2(n9748), .C1(
        n9747), .C2(n10207), .ZN(n9751) );
  OAI211_X1 U10924 ( .C1(n9754), .C2(n9753), .A(n9752), .B(n9751), .ZN(
        P2_U3199) );
  XNOR2_X1 U10925 ( .A(n9755), .B(n9757), .ZN(n9781) );
  XNOR2_X1 U10926 ( .A(n9756), .B(n9757), .ZN(n9763) );
  AOI22_X1 U10927 ( .A1(n8352), .A2(n9760), .B1(n9759), .B2(n9758), .ZN(n9761)
         );
  OAI21_X1 U10928 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  AOI21_X1 U10929 ( .B1(n9765), .B2(n9781), .A(n9764), .ZN(n9778) );
  NOR2_X1 U10930 ( .A1(n9766), .A2(n9821), .ZN(n9780) );
  INV_X1 U10931 ( .A(n9767), .ZN(n9769) );
  AOI22_X1 U10932 ( .A1(n9780), .A2(n9769), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9768), .ZN(n9772) );
  AOI22_X1 U10933 ( .A1(n9781), .A2(n9770), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n9773), .ZN(n9771) );
  OAI221_X1 U10934 ( .B1(n9773), .B2(n9778), .C1(n9773), .C2(n9772), .A(n9771), 
        .ZN(P2_U3231) );
  NOR2_X1 U10935 ( .A1(n9774), .A2(n9821), .ZN(n9776) );
  AOI211_X1 U10936 ( .C1(n9794), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9836)
         );
  AOI22_X1 U10937 ( .A1(n9835), .A2(n5807), .B1(n9836), .B2(n9833), .ZN(
        P2_U3393) );
  INV_X1 U10938 ( .A(n9778), .ZN(n9779) );
  AOI211_X1 U10939 ( .C1(n9781), .C2(n9794), .A(n9780), .B(n9779), .ZN(n9837)
         );
  AOI22_X1 U10940 ( .A1(n9835), .A2(n5839), .B1(n9837), .B2(n9833), .ZN(
        P2_U3396) );
  OAI21_X1 U10941 ( .B1(n9783), .B2(n9821), .A(n9782), .ZN(n9784) );
  AOI21_X1 U10942 ( .B1(n9819), .B2(n9785), .A(n9784), .ZN(n9839) );
  AOI22_X1 U10943 ( .A1(n9835), .A2(n5855), .B1(n9839), .B2(n9833), .ZN(
        P2_U3399) );
  OAI21_X1 U10944 ( .B1(n9787), .B2(n9821), .A(n9786), .ZN(n9788) );
  AOI21_X1 U10945 ( .B1(n9789), .B2(n9819), .A(n9788), .ZN(n9840) );
  AOI22_X1 U10946 ( .A1(n9835), .A2(n5872), .B1(n9840), .B2(n9833), .ZN(
        P2_U3402) );
  NOR2_X1 U10947 ( .A1(n9790), .A2(n9821), .ZN(n9792) );
  AOI211_X1 U10948 ( .C1(n9794), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9841)
         );
  AOI22_X1 U10949 ( .A1(n9835), .A2(n5885), .B1(n9841), .B2(n9833), .ZN(
        P2_U3405) );
  NOR2_X1 U10950 ( .A1(n9795), .A2(n9821), .ZN(n9797) );
  AOI211_X1 U10951 ( .C1(n9798), .C2(n9819), .A(n9797), .B(n9796), .ZN(n9843)
         );
  AOI22_X1 U10952 ( .A1(n9835), .A2(n5899), .B1(n9843), .B2(n9833), .ZN(
        P2_U3408) );
  OAI22_X1 U10953 ( .A1(n9800), .A2(n9808), .B1(n9799), .B2(n9821), .ZN(n9801)
         );
  NOR2_X1 U10954 ( .A1(n9802), .A2(n9801), .ZN(n9844) );
  AOI22_X1 U10955 ( .A1(n9835), .A2(n5919), .B1(n9844), .B2(n9833), .ZN(
        P2_U3411) );
  OAI21_X1 U10956 ( .B1(n9804), .B2(n9821), .A(n9803), .ZN(n9805) );
  AOI21_X1 U10957 ( .B1(n9819), .B2(n9806), .A(n9805), .ZN(n9845) );
  AOI22_X1 U10958 ( .A1(n9835), .A2(n5934), .B1(n9845), .B2(n9833), .ZN(
        P2_U3414) );
  INV_X1 U10959 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9812) );
  OAI22_X1 U10960 ( .A1(n9809), .A2(n9808), .B1(n9807), .B2(n9821), .ZN(n9810)
         );
  NOR2_X1 U10961 ( .A1(n9811), .A2(n9810), .ZN(n9846) );
  AOI22_X1 U10962 ( .A1(n9835), .A2(n9812), .B1(n9846), .B2(n9833), .ZN(
        P2_U3417) );
  INV_X1 U10963 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U10964 ( .A1(n9813), .A2(n9819), .ZN(n9816) );
  NAND2_X1 U10965 ( .A1(n9814), .A2(n9832), .ZN(n9815) );
  AND3_X1 U10966 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9847) );
  AOI22_X1 U10967 ( .A1(n9835), .A2(n9818), .B1(n9847), .B2(n9833), .ZN(
        P2_U3420) );
  INV_X1 U10968 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9826) );
  NAND2_X1 U10969 ( .A1(n9820), .A2(n9819), .ZN(n9824) );
  OR2_X1 U10970 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  AOI22_X1 U10971 ( .A1(n9835), .A2(n9826), .B1(n9848), .B2(n9833), .ZN(
        P2_U3423) );
  INV_X1 U10972 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9834) );
  NOR2_X1 U10973 ( .A1(n9828), .A2(n9827), .ZN(n9830) );
  AOI211_X1 U10974 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9850)
         );
  AOI22_X1 U10975 ( .A1(n9835), .A2(n9834), .B1(n9850), .B2(n9833), .ZN(
        P2_U3426) );
  AOI22_X1 U10976 ( .A1(n9851), .A2(n9836), .B1(n5808), .B2(n9849), .ZN(
        P2_U3460) );
  AOI22_X1 U10977 ( .A1(n9851), .A2(n9837), .B1(n6653), .B2(n9849), .ZN(
        P2_U3461) );
  INV_X1 U10978 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U10979 ( .A1(n9851), .A2(n9839), .B1(n9838), .B2(n9849), .ZN(
        P2_U3462) );
  AOI22_X1 U10980 ( .A1(n9851), .A2(n9840), .B1(n6751), .B2(n9849), .ZN(
        P2_U3463) );
  INV_X1 U10981 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U10982 ( .A1(n9851), .A2(n9841), .B1(n9959), .B2(n9849), .ZN(
        P2_U3464) );
  AOI22_X1 U10983 ( .A1(n9851), .A2(n9843), .B1(n9842), .B2(n9849), .ZN(
        P2_U3465) );
  AOI22_X1 U10984 ( .A1(n9851), .A2(n9844), .B1(n6976), .B2(n9849), .ZN(
        P2_U3466) );
  AOI22_X1 U10985 ( .A1(n9851), .A2(n9845), .B1(n6973), .B2(n9849), .ZN(
        P2_U3467) );
  AOI22_X1 U10986 ( .A1(n9851), .A2(n9846), .B1(n5947), .B2(n9849), .ZN(
        P2_U3468) );
  AOI22_X1 U10987 ( .A1(n9851), .A2(n9847), .B1(n5963), .B2(n9849), .ZN(
        P2_U3469) );
  AOI22_X1 U10988 ( .A1(n9851), .A2(n9848), .B1(n5979), .B2(n9849), .ZN(
        P2_U3470) );
  AOI22_X1 U10989 ( .A1(n9851), .A2(n9850), .B1(n5993), .B2(n9849), .ZN(
        P2_U3471) );
  OAI222_X1 U10990 ( .A1(n9856), .A2(n9855), .B1(n9856), .B2(n9854), .C1(n9853), .C2(n9852), .ZN(ADD_1068_U5) );
  AOI21_X1 U10991 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(ADD_1068_U46) );
  OAI21_X1 U10992 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9863) );
  XNOR2_X1 U10993 ( .A(n9863), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U10994 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(ADD_1068_U56) );
  OAI21_X1 U10995 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(ADD_1068_U57) );
  OAI21_X1 U10996 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(ADD_1068_U58) );
  OAI21_X1 U10997 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(ADD_1068_U59) );
  OAI21_X1 U10998 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(ADD_1068_U60) );
  OAI21_X1 U10999 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(ADD_1068_U61) );
  OAI21_X1 U11000 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(ADD_1068_U62) );
  OAI21_X1 U11001 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(ADD_1068_U63) );
  NAND4_X1 U11002 ( .A1(keyinput44), .A2(keyinput40), .A3(keyinput59), .A4(
        keyinput68), .ZN(n9888) );
  NOR3_X1 U11003 ( .A1(keyinput66), .A2(keyinput113), .A3(n9888), .ZN(n9903)
         );
  NAND2_X1 U11004 ( .A1(keyinput114), .A2(keyinput73), .ZN(n9889) );
  NOR3_X1 U11005 ( .A1(keyinput78), .A2(keyinput115), .A3(n9889), .ZN(n9890)
         );
  NAND3_X1 U11006 ( .A1(keyinput5), .A2(keyinput77), .A3(n9890), .ZN(n9900) );
  INV_X1 U11007 ( .A(keyinput48), .ZN(n9891) );
  NOR4_X1 U11008 ( .A1(keyinput87), .A2(keyinput112), .A3(keyinput123), .A4(
        n9891), .ZN(n9898) );
  NAND2_X1 U11009 ( .A1(keyinput95), .A2(keyinput80), .ZN(n9892) );
  NOR3_X1 U11010 ( .A1(keyinput16), .A2(keyinput83), .A3(n9892), .ZN(n9897) );
  NAND2_X1 U11011 ( .A1(keyinput13), .A2(keyinput124), .ZN(n9893) );
  NOR3_X1 U11012 ( .A1(keyinput121), .A2(keyinput4), .A3(n9893), .ZN(n9896) );
  NAND2_X1 U11013 ( .A1(keyinput14), .A2(keyinput107), .ZN(n9894) );
  NOR3_X1 U11014 ( .A1(keyinput47), .A2(keyinput45), .A3(n9894), .ZN(n9895) );
  NAND4_X1 U11015 ( .A1(n9898), .A2(n9897), .A3(n9896), .A4(n9895), .ZN(n9899)
         );
  NOR4_X1 U11016 ( .A1(keyinput104), .A2(keyinput9), .A3(n9900), .A4(n9899), 
        .ZN(n9902) );
  INV_X1 U11017 ( .A(keyinput99), .ZN(n9901) );
  NAND4_X1 U11018 ( .A1(keyinput90), .A2(n9903), .A3(n9902), .A4(n9901), .ZN(
        n9914) );
  NAND4_X1 U11019 ( .A1(keyinput2), .A2(keyinput55), .A3(keyinput54), .A4(
        keyinput111), .ZN(n9913) );
  NAND4_X1 U11020 ( .A1(keyinput50), .A2(keyinput71), .A3(keyinput42), .A4(
        keyinput67), .ZN(n9912) );
  NAND4_X1 U11021 ( .A1(keyinput28), .A2(keyinput12), .A3(keyinput116), .A4(
        keyinput64), .ZN(n9904) );
  NOR3_X1 U11022 ( .A1(keyinput110), .A2(keyinput63), .A3(n9904), .ZN(n9910)
         );
  NAND4_X1 U11023 ( .A1(keyinput70), .A2(keyinput74), .A3(keyinput86), .A4(
        keyinput91), .ZN(n9908) );
  NAND4_X1 U11024 ( .A1(keyinput94), .A2(keyinput127), .A3(keyinput75), .A4(
        keyinput119), .ZN(n9907) );
  NAND4_X1 U11025 ( .A1(keyinput81), .A2(keyinput65), .A3(keyinput89), .A4(
        keyinput118), .ZN(n9906) );
  NAND4_X1 U11026 ( .A1(keyinput41), .A2(keyinput105), .A3(keyinput21), .A4(
        keyinput17), .ZN(n9905) );
  NOR4_X1 U11027 ( .A1(n9908), .A2(n9907), .A3(n9906), .A4(n9905), .ZN(n9909)
         );
  NAND4_X1 U11028 ( .A1(keyinput32), .A2(keyinput84), .A3(n9910), .A4(n9909), 
        .ZN(n9911) );
  NOR4_X1 U11029 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n10201)
         );
  INV_X1 U11030 ( .A(keyinput61), .ZN(n9915) );
  NAND4_X1 U11031 ( .A1(keyinput46), .A2(keyinput3), .A3(keyinput56), .A4(
        n9915), .ZN(n9921) );
  NAND4_X1 U11032 ( .A1(keyinput85), .A2(keyinput125), .A3(keyinput60), .A4(
        keyinput88), .ZN(n9920) );
  NOR3_X1 U11033 ( .A1(keyinput24), .A2(keyinput79), .A3(keyinput7), .ZN(n9916) );
  NAND2_X1 U11034 ( .A1(keyinput126), .A2(n9916), .ZN(n9919) );
  INV_X1 U11035 ( .A(keyinput69), .ZN(n9917) );
  NAND4_X1 U11036 ( .A1(keyinput122), .A2(keyinput23), .A3(keyinput25), .A4(
        n9917), .ZN(n9918) );
  OR4_X1 U11037 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(n9940)
         );
  NAND2_X1 U11038 ( .A1(keyinput11), .A2(keyinput30), .ZN(n9922) );
  NOR3_X1 U11039 ( .A1(keyinput109), .A2(keyinput100), .A3(n9922), .ZN(n9928)
         );
  NAND2_X1 U11040 ( .A1(keyinput82), .A2(keyinput102), .ZN(n9923) );
  NOR3_X1 U11041 ( .A1(keyinput6), .A2(keyinput15), .A3(n9923), .ZN(n9927) );
  NOR4_X1 U11042 ( .A1(keyinput10), .A2(keyinput62), .A3(keyinput108), .A4(
        keyinput49), .ZN(n9926) );
  NAND2_X1 U11043 ( .A1(keyinput101), .A2(keyinput51), .ZN(n9924) );
  NOR3_X1 U11044 ( .A1(keyinput43), .A2(keyinput58), .A3(n9924), .ZN(n9925) );
  NAND4_X1 U11045 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n9939)
         );
  NOR4_X1 U11046 ( .A1(keyinput27), .A2(keyinput31), .A3(keyinput34), .A4(
        keyinput35), .ZN(n9932) );
  NOR4_X1 U11047 ( .A1(keyinput29), .A2(keyinput1), .A3(keyinput93), .A4(
        keyinput26), .ZN(n9931) );
  NOR4_X1 U11048 ( .A1(keyinput22), .A2(keyinput98), .A3(keyinput103), .A4(
        keyinput106), .ZN(n9930) );
  NOR4_X1 U11049 ( .A1(keyinput38), .A2(keyinput39), .A3(keyinput18), .A4(
        keyinput19), .ZN(n9929) );
  NAND4_X1 U11050 ( .A1(n9932), .A2(n9931), .A3(n9930), .A4(n9929), .ZN(n9938)
         );
  NOR4_X1 U11051 ( .A1(keyinput36), .A2(keyinput20), .A3(keyinput8), .A4(
        keyinput0), .ZN(n9936) );
  NOR4_X1 U11052 ( .A1(keyinput52), .A2(keyinput72), .A3(keyinput76), .A4(
        keyinput92), .ZN(n9935) );
  NOR4_X1 U11053 ( .A1(keyinput37), .A2(keyinput33), .A3(keyinput117), .A4(
        keyinput97), .ZN(n9934) );
  NOR4_X1 U11054 ( .A1(keyinput96), .A2(keyinput120), .A3(keyinput57), .A4(
        keyinput53), .ZN(n9933) );
  NAND4_X1 U11055 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(n9937)
         );
  NOR4_X1 U11056 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), .ZN(n10200)
         );
  AOI22_X1 U11057 ( .A1(n9942), .A2(keyinput76), .B1(keyinput117), .B2(n5919), 
        .ZN(n9941) );
  OAI221_X1 U11058 ( .B1(n9942), .B2(keyinput76), .C1(n5919), .C2(keyinput117), 
        .A(n9941), .ZN(n9953) );
  AOI22_X1 U11059 ( .A1(n9945), .A2(keyinput52), .B1(keyinput119), .B2(n9944), 
        .ZN(n9943) );
  OAI221_X1 U11060 ( .B1(n9945), .B2(keyinput52), .C1(n9944), .C2(keyinput119), 
        .A(n9943), .ZN(n9952) );
  INV_X1 U11061 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9946) );
  XOR2_X1 U11062 ( .A(n9946), .B(keyinput32), .Z(n9950) );
  XNOR2_X1 U11063 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput116), .ZN(n9949) );
  XNOR2_X1 U11064 ( .A(P2_REG1_REG_25__SCAN_IN), .B(keyinput91), .ZN(n9948) );
  XNOR2_X1 U11065 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput110), .ZN(n9947)
         );
  NAND4_X1 U11066 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n9951)
         );
  NOR3_X1 U11067 ( .A1(n9953), .A2(n9952), .A3(n9951), .ZN(n9998) );
  INV_X1 U11068 ( .A(SI_10_), .ZN(n9956) );
  AOI22_X1 U11069 ( .A1(n9956), .A2(keyinput72), .B1(keyinput17), .B2(n9955), 
        .ZN(n9954) );
  OAI221_X1 U11070 ( .B1(n9956), .B2(keyinput72), .C1(n9955), .C2(keyinput17), 
        .A(n9954), .ZN(n9969) );
  INV_X1 U11071 ( .A(keyinput120), .ZN(n9958) );
  AOI22_X1 U11072 ( .A1(n9959), .A2(keyinput19), .B1(P1_ADDR_REG_9__SCAN_IN), 
        .B2(n9958), .ZN(n9957) );
  OAI221_X1 U11073 ( .B1(n9959), .B2(keyinput19), .C1(n9958), .C2(
        P1_ADDR_REG_9__SCAN_IN), .A(n9957), .ZN(n9968) );
  INV_X1 U11074 ( .A(keyinput127), .ZN(n9961) );
  AOI22_X1 U11075 ( .A1(n9962), .A2(keyinput63), .B1(P2_ADDR_REG_6__SCAN_IN), 
        .B2(n9961), .ZN(n9960) );
  OAI221_X1 U11076 ( .B1(n9962), .B2(keyinput63), .C1(n9961), .C2(
        P2_ADDR_REG_6__SCAN_IN), .A(n9960), .ZN(n9967) );
  AOI22_X1 U11077 ( .A1(n9965), .A2(keyinput39), .B1(keyinput118), .B2(n9964), 
        .ZN(n9963) );
  OAI221_X1 U11078 ( .B1(n9965), .B2(keyinput39), .C1(n9964), .C2(keyinput118), 
        .A(n9963), .ZN(n9966) );
  NOR4_X1 U11079 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9997)
         );
  INV_X1 U11080 ( .A(keyinput0), .ZN(n9971) );
  AOI22_X1 U11081 ( .A1(n8096), .A2(keyinput106), .B1(P1_ADDR_REG_1__SCAN_IN), 
        .B2(n9971), .ZN(n9970) );
  OAI221_X1 U11082 ( .B1(n8096), .B2(keyinput106), .C1(n9971), .C2(
        P1_ADDR_REG_1__SCAN_IN), .A(n9970), .ZN(n9982) );
  INV_X1 U11083 ( .A(keyinput57), .ZN(n9973) );
  AOI22_X1 U11084 ( .A1(n5375), .A2(keyinput64), .B1(P2_ADDR_REG_9__SCAN_IN), 
        .B2(n9973), .ZN(n9972) );
  OAI221_X1 U11085 ( .B1(n5375), .B2(keyinput64), .C1(n9973), .C2(
        P2_ADDR_REG_9__SCAN_IN), .A(n9972), .ZN(n9981) );
  AOI22_X1 U11086 ( .A1(n9976), .A2(keyinput27), .B1(n9975), .B2(keyinput34), 
        .ZN(n9974) );
  OAI221_X1 U11087 ( .B1(n9976), .B2(keyinput27), .C1(n9975), .C2(keyinput34), 
        .A(n9974), .ZN(n9980) );
  XNOR2_X1 U11088 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput71), .ZN(n9978) );
  XNOR2_X1 U11089 ( .A(keyinput20), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U11090 ( .A1(n9978), .A2(n9977), .ZN(n9979) );
  NOR4_X1 U11091 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n9996)
         );
  AOI22_X1 U11092 ( .A1(n9984), .A2(keyinput37), .B1(n5756), .B2(keyinput111), 
        .ZN(n9983) );
  OAI221_X1 U11093 ( .B1(n9984), .B2(keyinput37), .C1(n5756), .C2(keyinput111), 
        .A(n9983), .ZN(n9994) );
  AOI22_X1 U11094 ( .A1(P2_U3151), .A2(keyinput42), .B1(keyinput75), .B2(n9986), .ZN(n9985) );
  OAI221_X1 U11095 ( .B1(P2_U3151), .B2(keyinput42), .C1(n9986), .C2(
        keyinput75), .A(n9985), .ZN(n9993) );
  AOI22_X1 U11096 ( .A1(n9988), .A2(keyinput1), .B1(n5153), .B2(keyinput12), 
        .ZN(n9987) );
  OAI221_X1 U11097 ( .B1(n9988), .B2(keyinput1), .C1(n5153), .C2(keyinput12), 
        .A(n9987), .ZN(n9992) );
  AOI22_X1 U11098 ( .A1(n5934), .A2(keyinput41), .B1(n9990), .B2(keyinput89), 
        .ZN(n9989) );
  OAI221_X1 U11099 ( .B1(n5934), .B2(keyinput41), .C1(n9990), .C2(keyinput89), 
        .A(n9989), .ZN(n9991) );
  NOR4_X1 U11100 ( .A1(n9994), .A2(n9993), .A3(n9992), .A4(n9991), .ZN(n9995)
         );
  NAND4_X1 U11101 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n10199) );
  INV_X1 U11102 ( .A(keyinput97), .ZN(n10000) );
  OAI22_X1 U11103 ( .A1(n7118), .A2(keyinput8), .B1(n10000), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n9999) );
  AOI221_X1 U11104 ( .B1(n7118), .B2(keyinput8), .C1(P1_ADDR_REG_0__SCAN_IN), 
        .C2(n10000), .A(n9999), .ZN(n10013) );
  INV_X1 U11105 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10002) );
  OAI22_X1 U11106 ( .A1(n10003), .A2(keyinput2), .B1(n10002), .B2(keyinput65), 
        .ZN(n10001) );
  AOI221_X1 U11107 ( .B1(n10003), .B2(keyinput2), .C1(keyinput65), .C2(n10002), 
        .A(n10001), .ZN(n10012) );
  OAI22_X1 U11108 ( .A1(n10006), .A2(keyinput92), .B1(n10005), .B2(keyinput33), 
        .ZN(n10004) );
  AOI221_X1 U11109 ( .B1(n10006), .B2(keyinput92), .C1(keyinput33), .C2(n10005), .A(n10004), .ZN(n10011) );
  OAI22_X1 U11110 ( .A1(n10009), .A2(keyinput67), .B1(n10008), .B2(keyinput105), .ZN(n10007) );
  AOI221_X1 U11111 ( .B1(n10009), .B2(keyinput67), .C1(keyinput105), .C2(
        n10008), .A(n10007), .ZN(n10010) );
  NAND4_X1 U11112 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n10065) );
  XOR2_X1 U11113 ( .A(P2_B_REG_SCAN_IN), .B(keyinput29), .Z(n10020) );
  XNOR2_X1 U11114 ( .A(n10014), .B(keyinput18), .ZN(n10019) );
  INV_X1 U11115 ( .A(keyinput96), .ZN(n10015) );
  XNOR2_X1 U11116 ( .A(n10015), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n10018) );
  XNOR2_X1 U11117 ( .A(n10016), .B(keyinput74), .ZN(n10017) );
  NOR4_X1 U11118 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10029) );
  OAI22_X1 U11119 ( .A1(n10023), .A2(keyinput36), .B1(n10022), .B2(keyinput55), 
        .ZN(n10021) );
  AOI221_X1 U11120 ( .B1(n10023), .B2(keyinput36), .C1(keyinput55), .C2(n10022), .A(n10021), .ZN(n10028) );
  INV_X1 U11121 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10026) );
  INV_X1 U11122 ( .A(keyinput54), .ZN(n10025) );
  OAI22_X1 U11123 ( .A1(n10026), .A2(keyinput98), .B1(n10025), .B2(
        P1_ADDR_REG_15__SCAN_IN), .ZN(n10024) );
  AOI221_X1 U11124 ( .B1(n10026), .B2(keyinput98), .C1(P1_ADDR_REG_15__SCAN_IN), .C2(n10025), .A(n10024), .ZN(n10027) );
  NAND3_X1 U11125 ( .A1(n10029), .A2(n10028), .A3(n10027), .ZN(n10064) );
  OAI22_X1 U11126 ( .A1(n10031), .A2(keyinput38), .B1(n5993), .B2(keyinput50), 
        .ZN(n10030) );
  AOI221_X1 U11127 ( .B1(n10031), .B2(keyinput38), .C1(keyinput50), .C2(n5993), 
        .A(n10030), .ZN(n10044) );
  XNOR2_X1 U11128 ( .A(n10032), .B(keyinput21), .ZN(n10038) );
  XOR2_X1 U11129 ( .A(P1_REG0_REG_22__SCAN_IN), .B(keyinput86), .Z(n10037) );
  XNOR2_X1 U11130 ( .A(n10033), .B(keyinput84), .ZN(n10036) );
  XNOR2_X1 U11131 ( .A(n10034), .B(keyinput35), .ZN(n10035) );
  NOR4_X1 U11132 ( .A1(n10038), .A2(n10037), .A3(n10036), .A4(n10035), .ZN(
        n10043) );
  INV_X1 U11133 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10041) );
  OAI22_X1 U11134 ( .A1(n10041), .A2(keyinput26), .B1(n10040), .B2(keyinput103), .ZN(n10039) );
  AOI221_X1 U11135 ( .B1(n10041), .B2(keyinput26), .C1(keyinput103), .C2(
        n10040), .A(n10039), .ZN(n10042) );
  NAND3_X1 U11136 ( .A1(n10044), .A2(n10043), .A3(n10042), .ZN(n10063) );
  INV_X1 U11137 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10046) );
  OAI22_X1 U11138 ( .A1(n10047), .A2(keyinput22), .B1(n10046), .B2(keyinput70), 
        .ZN(n10045) );
  AOI221_X1 U11139 ( .B1(n10047), .B2(keyinput22), .C1(keyinput70), .C2(n10046), .A(n10045), .ZN(n10061) );
  INV_X1 U11140 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10049) );
  OAI22_X1 U11141 ( .A1(n10050), .A2(keyinput94), .B1(n10049), .B2(keyinput81), 
        .ZN(n10048) );
  AOI221_X1 U11142 ( .B1(n10050), .B2(keyinput94), .C1(keyinput81), .C2(n10049), .A(n10048), .ZN(n10060) );
  INV_X1 U11143 ( .A(keyinput31), .ZN(n10052) );
  OAI22_X1 U11144 ( .A1(n10053), .A2(keyinput28), .B1(n10052), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n10051) );
  AOI221_X1 U11145 ( .B1(n10053), .B2(keyinput28), .C1(P2_REG2_REG_28__SCAN_IN), .C2(n10052), .A(n10051), .ZN(n10059) );
  XNOR2_X1 U11146 ( .A(n10054), .B(keyinput93), .ZN(n10057) );
  XNOR2_X1 U11147 ( .A(n10055), .B(keyinput53), .ZN(n10056) );
  NOR2_X1 U11148 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  NAND4_X1 U11149 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10062) );
  NOR4_X1 U11150 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10197) );
  AOI22_X1 U11151 ( .A1(n10068), .A2(keyinput10), .B1(n10067), .B2(keyinput62), 
        .ZN(n10066) );
  OAI221_X1 U11152 ( .B1(n10068), .B2(keyinput10), .C1(n10067), .C2(keyinput62), .A(n10066), .ZN(n10079) );
  AOI22_X1 U11153 ( .A1(n10071), .A2(keyinput43), .B1(n10070), .B2(keyinput51), 
        .ZN(n10069) );
  OAI221_X1 U11154 ( .B1(n10071), .B2(keyinput43), .C1(n10070), .C2(keyinput51), .A(n10069), .ZN(n10078) );
  INV_X1 U11155 ( .A(keyinput101), .ZN(n10072) );
  XNOR2_X1 U11156 ( .A(n10072), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n10077) );
  XNOR2_X1 U11157 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput58), .ZN(n10075) );
  XNOR2_X1 U11158 ( .A(P2_REG0_REG_30__SCAN_IN), .B(keyinput49), .ZN(n10074)
         );
  XNOR2_X1 U11159 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput108), .ZN(n10073)
         );
  NAND3_X1 U11160 ( .A1(n10075), .A2(n10074), .A3(n10073), .ZN(n10076) );
  NOR4_X1 U11161 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10196) );
  AOI22_X1 U11162 ( .A1(n10082), .A2(keyinput109), .B1(n10081), .B2(keyinput11), .ZN(n10080) );
  OAI221_X1 U11163 ( .B1(n10082), .B2(keyinput109), .C1(n10081), .C2(
        keyinput11), .A(n10080), .ZN(n10083) );
  INV_X1 U11164 ( .A(n10083), .ZN(n10096) );
  AOI22_X1 U11165 ( .A1(n10086), .A2(keyinput6), .B1(n10085), .B2(keyinput82), 
        .ZN(n10084) );
  OAI221_X1 U11166 ( .B1(n10086), .B2(keyinput6), .C1(n10085), .C2(keyinput82), 
        .A(n10084), .ZN(n10087) );
  INV_X1 U11167 ( .A(n10087), .ZN(n10095) );
  XNOR2_X1 U11168 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput102), .ZN(n10090)
         );
  XNOR2_X1 U11169 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput100), .ZN(n10089)
         );
  XNOR2_X1 U11170 ( .A(keyinput15), .B(P1_REG0_REG_17__SCAN_IN), .ZN(n10088)
         );
  AND3_X1 U11171 ( .A1(n10090), .A2(n10089), .A3(n10088), .ZN(n10094) );
  INV_X1 U11172 ( .A(keyinput30), .ZN(n10091) );
  XNOR2_X1 U11173 ( .A(n10092), .B(n10091), .ZN(n10093) );
  AND4_X1 U11174 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10195) );
  AOI22_X1 U11175 ( .A1(n10098), .A2(keyinput66), .B1(keyinput113), .B2(n5978), 
        .ZN(n10097) );
  OAI221_X1 U11176 ( .B1(n10098), .B2(keyinput66), .C1(n5978), .C2(keyinput113), .A(n10097), .ZN(n10111) );
  AOI22_X1 U11177 ( .A1(n10101), .A2(keyinput90), .B1(keyinput99), .B2(n10100), 
        .ZN(n10099) );
  OAI221_X1 U11178 ( .B1(n10101), .B2(keyinput90), .C1(n10100), .C2(keyinput99), .A(n10099), .ZN(n10110) );
  INV_X1 U11179 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10104) );
  INV_X1 U11180 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11181 ( .A1(n10104), .A2(keyinput59), .B1(keyinput68), .B2(n10103), 
        .ZN(n10102) );
  OAI221_X1 U11182 ( .B1(n10104), .B2(keyinput59), .C1(n10103), .C2(keyinput68), .A(n10102), .ZN(n10109) );
  AOI22_X1 U11183 ( .A1(n10107), .A2(keyinput44), .B1(n10106), .B2(keyinput40), 
        .ZN(n10105) );
  OAI221_X1 U11184 ( .B1(n10107), .B2(keyinput44), .C1(n10106), .C2(keyinput40), .A(n10105), .ZN(n10108) );
  NOR4_X1 U11185 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10193) );
  INV_X1 U11186 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10114) );
  OAI22_X1 U11187 ( .A1(n10114), .A2(keyinput122), .B1(n10113), .B2(keyinput69), .ZN(n10112) );
  AOI221_X1 U11188 ( .B1(n10114), .B2(keyinput122), .C1(keyinput69), .C2(
        n10113), .A(n10112), .ZN(n10147) );
  AOI22_X1 U11189 ( .A1(n10117), .A2(keyinput87), .B1(n10116), .B2(keyinput123), .ZN(n10115) );
  OAI221_X1 U11190 ( .B1(n10117), .B2(keyinput87), .C1(n10116), .C2(
        keyinput123), .A(n10115), .ZN(n10122) );
  AOI22_X1 U11191 ( .A1(n10120), .A2(keyinput3), .B1(n10119), .B2(keyinput56), 
        .ZN(n10118) );
  OAI221_X1 U11192 ( .B1(n10120), .B2(keyinput3), .C1(n10119), .C2(keyinput56), 
        .A(n10118), .ZN(n10121) );
  NOR2_X1 U11193 ( .A1(n10122), .A2(n10121), .ZN(n10146) );
  INV_X1 U11194 ( .A(keyinput77), .ZN(n10123) );
  XNOR2_X1 U11195 ( .A(n10124), .B(n10123), .ZN(n10135) );
  XNOR2_X1 U11196 ( .A(P1_REG3_REG_17__SCAN_IN), .B(keyinput88), .ZN(n10128)
         );
  XNOR2_X1 U11197 ( .A(P1_REG0_REG_16__SCAN_IN), .B(keyinput79), .ZN(n10127)
         );
  XNOR2_X1 U11198 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput16), .ZN(n10126) );
  XNOR2_X1 U11199 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput5), .ZN(n10125) );
  NAND4_X1 U11200 ( .A1(n10128), .A2(n10127), .A3(n10126), .A4(n10125), .ZN(
        n10133) );
  XNOR2_X1 U11201 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput124), .ZN(n10131) );
  XNOR2_X1 U11202 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput60), .ZN(n10130)
         );
  XNOR2_X1 U11203 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput126), .ZN(n10129) );
  NAND3_X1 U11204 ( .A1(n10131), .A2(n10130), .A3(n10129), .ZN(n10132) );
  NOR2_X1 U11205 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  AND2_X1 U11206 ( .A1(n10135), .A2(n10134), .ZN(n10145) );
  INV_X1 U11207 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U11208 ( .A1(n6180), .A2(keyinput24), .B1(n10137), .B2(keyinput7), 
        .ZN(n10136) );
  OAI221_X1 U11209 ( .B1(n6180), .B2(keyinput24), .C1(n10137), .C2(keyinput7), 
        .A(n10136), .ZN(n10143) );
  XNOR2_X1 U11210 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput107), .ZN(n10141) );
  XNOR2_X1 U11211 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput80), .ZN(n10140) );
  XNOR2_X1 U11212 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput13), .ZN(n10139) );
  XNOR2_X1 U11213 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput47), .ZN(n10138) );
  NAND4_X1 U11214 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10142) );
  NOR2_X1 U11215 ( .A1(n10143), .A2(n10142), .ZN(n10144) );
  AND4_X1 U11216 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10192) );
  INV_X1 U11217 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10150) );
  OAI22_X1 U11218 ( .A1(n10150), .A2(keyinput23), .B1(n10149), .B2(keyinput25), 
        .ZN(n10148) );
  AOI221_X1 U11219 ( .B1(n10150), .B2(keyinput23), .C1(keyinput25), .C2(n10149), .A(n10148), .ZN(n10191) );
  AOI22_X1 U11220 ( .A1(n10153), .A2(keyinput78), .B1(n10152), .B2(keyinput73), 
        .ZN(n10151) );
  OAI221_X1 U11221 ( .B1(n10153), .B2(keyinput78), .C1(n10152), .C2(keyinput73), .A(n10151), .ZN(n10158) );
  INV_X1 U11222 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10156) );
  INV_X1 U11223 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11224 ( .A1(n10156), .A2(keyinput48), .B1(keyinput112), .B2(n10155), .ZN(n10154) );
  OAI221_X1 U11225 ( .B1(n10156), .B2(keyinput48), .C1(n10155), .C2(
        keyinput112), .A(n10154), .ZN(n10157) );
  NOR2_X1 U11226 ( .A1(n10158), .A2(n10157), .ZN(n10166) );
  AOI22_X1 U11227 ( .A1(n10161), .A2(keyinput61), .B1(keyinput46), .B2(n10160), 
        .ZN(n10159) );
  OAI221_X1 U11228 ( .B1(n10161), .B2(keyinput61), .C1(n10160), .C2(keyinput46), .A(n10159), .ZN(n10164) );
  INV_X1 U11229 ( .A(keyinput4), .ZN(n10162) );
  XNOR2_X1 U11230 ( .A(n10162), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U11231 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  AND2_X1 U11232 ( .A1(n10166), .A2(n10165), .ZN(n10189) );
  AOI22_X1 U11233 ( .A1(n10168), .A2(keyinput85), .B1(keyinput125), .B2(n8331), 
        .ZN(n10167) );
  OAI221_X1 U11234 ( .B1(n10168), .B2(keyinput85), .C1(n8331), .C2(keyinput125), .A(n10167), .ZN(n10173) );
  INV_X1 U11235 ( .A(keyinput83), .ZN(n10170) );
  AOI22_X1 U11236 ( .A1(n10171), .A2(keyinput95), .B1(P1_ADDR_REG_6__SCAN_IN), 
        .B2(n10170), .ZN(n10169) );
  OAI221_X1 U11237 ( .B1(n10171), .B2(keyinput95), .C1(n10170), .C2(
        P1_ADDR_REG_6__SCAN_IN), .A(n10169), .ZN(n10172) );
  NOR2_X1 U11238 ( .A1(n10173), .A2(n10172), .ZN(n10188) );
  INV_X1 U11239 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U11240 ( .A1(n10175), .A2(keyinput114), .B1(keyinput115), .B2(n6733), .ZN(n10174) );
  OAI221_X1 U11241 ( .B1(n10175), .B2(keyinput114), .C1(n6733), .C2(
        keyinput115), .A(n10174), .ZN(n10179) );
  AOI22_X1 U11242 ( .A1(n10177), .A2(keyinput104), .B1(keyinput9), .B2(n6009), 
        .ZN(n10176) );
  OAI221_X1 U11243 ( .B1(n10177), .B2(keyinput104), .C1(n6009), .C2(keyinput9), 
        .A(n10176), .ZN(n10178) );
  NOR2_X1 U11244 ( .A1(n10179), .A2(n10178), .ZN(n10187) );
  XNOR2_X1 U11245 ( .A(n10183), .B(keyinput121), .ZN(n10184) );
  NOR2_X1 U11246 ( .A1(n10185), .A2(n10184), .ZN(n10186) );
  AND4_X1 U11247 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10190) );
  AND4_X1 U11248 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10194) );
  NAND4_X1 U11249 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  AOI211_X1 U11250 ( .C1(n10201), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10224) );
  OAI21_X1 U11251 ( .B1(n10204), .B2(n10203), .A(n10202), .ZN(n10222) );
  INV_X1 U11252 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10216) );
  XNOR2_X1 U11253 ( .A(n10206), .B(n10205), .ZN(n10210) );
  INV_X1 U11254 ( .A(n10210), .ZN(n10208) );
  NAND2_X1 U11255 ( .A1(n10208), .A2(n10207), .ZN(n10213) );
  AOI21_X1 U11256 ( .B1(n10210), .B2(P2_U3893), .A(n10209), .ZN(n10212) );
  MUX2_X1 U11257 ( .A(n10213), .B(n10212), .S(n10211), .Z(n10215) );
  NAND2_X1 U11258 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n10214)
         );
  OAI211_X1 U11259 ( .C1(n10217), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n10221) );
  OAI21_X1 U11260 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(ADD_1068_U50) );
  OAI21_X1 U11261 ( .B1(n10230), .B2(n10229), .A(n10228), .ZN(ADD_1068_U51) );
  OAI21_X1 U11262 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(ADD_1068_U47) );
  OAI21_X1 U11263 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(ADD_1068_U49) );
  OAI21_X1 U11264 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(ADD_1068_U48) );
  AOI21_X1 U11265 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(ADD_1068_U54) );
  AOI21_X1 U11266 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(ADD_1068_U53) );
  OAI21_X1 U11267 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(ADD_1068_U52) );
  NOR2_X2 U4923 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5208) );
  CLKBUF_X2 U4933 ( .A(n5850), .Z(n4415) );
  NAND2_X1 U4935 ( .A1(n6720), .A2(n7121), .ZN(n9452) );
  OR2_X1 U4974 ( .A1(n6647), .A2(P2_U3151), .ZN(n10253) );
endmodule

