

module b15_C_SARLock_k_128_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025;

  OR2_X1 U3568 ( .A1(n5366), .A2(n5590), .ZN(n3123) );
  NOR2_X1 U3569 ( .A1(n5336), .A2(n3776), .ZN(n3779) );
  NAND2_X1 U3571 ( .A1(n5062), .A2(n3727), .ZN(n5094) );
  OR2_X1 U3572 ( .A1(n4026), .A2(n5429), .ZN(n4027) );
  NAND2_X1 U3573 ( .A1(n3683), .A2(n3682), .ZN(n4507) );
  CLKBUF_X2 U3574 ( .A(n3331), .Z(n4317) );
  CLKBUF_X2 U3575 ( .A(n3247), .Z(n4307) );
  CLKBUF_X2 U3576 ( .A(n3234), .Z(n3120) );
  CLKBUF_X2 U3577 ( .A(n3213), .Z(n4316) );
  CLKBUF_X2 U3578 ( .A(n3364), .Z(n3121) );
  NAND2_X1 U3579 ( .A1(n3262), .A2(n3261), .ZN(n3635) );
  CLKBUF_X2 U3580 ( .A(n3350), .Z(n4178) );
  CLKBUF_X2 U3581 ( .A(n3348), .Z(n4284) );
  NAND4_X2 U3582 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3277)
         );
  AND2_X2 U3583 ( .A1(n4563), .A2(n4375), .ZN(n3213) );
  INV_X1 U3584 ( .A(n3597), .ZN(n3612) );
  INV_X1 U3585 ( .A(n5223), .ZN(n5164) );
  NAND2_X1 U3587 ( .A1(n5091), .A2(n5162), .ZN(n5161) );
  CLKBUF_X2 U3588 ( .A(n3316), .Z(n4559) );
  OR2_X1 U3589 ( .A1(n4210), .A2(n5306), .ZN(n4231) );
  NAND2_X1 U3590 ( .A1(n3932), .A2(n3931), .ZN(n4470) );
  AND2_X1 U3592 ( .A1(n3139), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4381)
         );
  INV_X1 U3593 ( .A(n5590), .ZN(n6105) );
  NAND2_X1 U3594 ( .A1(n5342), .A2(n5341), .ZN(n5471) );
  NAND2_X2 U3595 ( .A1(n3288), .A2(n3780), .ZN(n3293) );
  AND4_X2 U3596 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3253)
         );
  NOR2_X4 U3597 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4374) );
  AND2_X1 U3598 ( .A1(n4563), .A2(n4375), .ZN(n3119) );
  NAND2_X2 U3599 ( .A1(n3259), .A2(n3780), .ZN(n3232) );
  NAND2_X2 U3600 ( .A1(n3165), .A2(n3260), .ZN(n3259) );
  AND4_X2 U3601 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3163)
         );
  AND2_X2 U3602 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n3140), .ZN(n3148)
         );
  AND4_X2 U3603 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3164)
         );
  INV_X1 U3604 ( .A(n5802), .ZN(n6696) );
  NOR2_X2 U3605 ( .A1(n5276), .A2(n5389), .ZN(n5309) );
  NAND2_X2 U3606 ( .A1(n3164), .A2(n3163), .ZN(n3260) );
  XNOR2_X2 U3607 ( .A(n3456), .B(n6167), .ZN(n6091) );
  XNOR2_X2 U3608 ( .A(n3502), .B(n3480), .ZN(n3896) );
  NAND2_X2 U3609 ( .A1(n3455), .A2(n3454), .ZN(n3456) );
  NAND2_X2 U3610 ( .A1(n5294), .A2(n5293), .ZN(n5577) );
  XNOR2_X2 U3611 ( .A(n3428), .B(n3429), .ZN(n4398) );
  NAND2_X2 U3612 ( .A1(n3303), .A2(n3326), .ZN(n3428) );
  NAND2_X1 U3613 ( .A1(n5561), .A2(n3571), .ZN(n5593) );
  AND2_X1 U3614 ( .A1(n5309), .A2(n4195), .ZN(n5499) );
  NAND2_X1 U3615 ( .A1(n4785), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U3616 ( .A1(n3517), .A2(n3518), .ZN(n3536) );
  AND2_X1 U3617 ( .A1(n3403), .A2(n3419), .ZN(n4462) );
  CLKBUF_X1 U3618 ( .A(n4584), .Z(n6210) );
  NAND2_X1 U3619 ( .A1(n3427), .A2(n3426), .ZN(n3458) );
  XNOR2_X1 U3621 ( .A(n3411), .B(n3410), .ZN(n3907) );
  OR2_X1 U3622 ( .A1(n4857), .A2(n3602), .ZN(n3400) );
  XNOR2_X1 U3623 ( .A(n3408), .B(n3407), .ZN(n3411) );
  NAND2_X1 U3624 ( .A1(n3344), .A2(n3343), .ZN(n3409) );
  OR2_X1 U3625 ( .A1(n3405), .A2(n3404), .ZN(n3408) );
  CLKBUF_X1 U3626 ( .A(n4367), .Z(n6004) );
  INV_X1 U3627 ( .A(n4505), .ZN(n3683) );
  OAI211_X1 U3628 ( .C1(n3299), .C2(n3287), .A(n3300), .B(n3298), .ZN(n3327)
         );
  NAND2_X1 U3629 ( .A1(n3677), .A2(n3676), .ZN(n4505) );
  NOR2_X2 U3630 ( .A1(n6733), .A2(n4027), .ZN(n4073) );
  CLKBUF_X1 U3631 ( .A(n3654), .Z(n5910) );
  INV_X1 U3632 ( .A(n4504), .ZN(n3682) );
  NOR2_X1 U3633 ( .A1(n4368), .A2(n5097), .ZN(n3781) );
  INV_X1 U3634 ( .A(n3636), .ZN(n3414) );
  CLKBUF_X1 U3635 ( .A(n3277), .Z(n4605) );
  BUF_X2 U3636 ( .A(n3288), .Z(n4615) );
  OR2_X2 U3637 ( .A1(n3203), .A2(n3202), .ZN(n5098) );
  INV_X1 U3638 ( .A(n3788), .ZN(n4621) );
  AND4_X1 U3639 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3231)
         );
  AND4_X1 U3640 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n3228)
         );
  AND4_X1 U3641 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3230)
         );
  AND4_X1 U3642 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3229)
         );
  OR2_X2 U3643 ( .A1(n6574), .A2(n6401), .ZN(n5590) );
  BUF_X2 U3644 ( .A(n3309), .Z(n4305) );
  BUF_X2 U3645 ( .A(n3310), .Z(n4260) );
  AND2_X2 U3646 ( .A1(n6972), .A2(n4594), .ZN(n6677) );
  OR2_X2 U3647 ( .A1(n4792), .A2(n4793), .ZN(n4854) );
  XNOR2_X1 U3648 ( .A(n3330), .B(n3329), .ZN(n4367) );
  OAI22_X2 U3650 ( .A1(n5559), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5571), .B2(n5297), .ZN(n5298) );
  AND2_X4 U3651 ( .A1(n5482), .A2(n5476), .ZN(n5478) );
  NOR2_X4 U3652 ( .A1(n5494), .A2(n5481), .ZN(n5482) );
  OR2_X2 U3653 ( .A1(n5500), .A2(n5493), .ZN(n5494) );
  NOR2_X4 U3654 ( .A1(n4507), .A2(n4499), .ZN(n4652) );
  AND2_X2 U3655 ( .A1(n4855), .A2(n4809), .ZN(n5062) );
  NOR2_X2 U3656 ( .A1(n4854), .A2(n4853), .ZN(n4855) );
  OR2_X1 U3658 ( .A1(n3342), .A2(n3341), .ZN(n3412) );
  NAND2_X1 U3659 ( .A1(n3585), .A2(n4643), .ZN(n3597) );
  NAND2_X1 U3660 ( .A1(n3437), .A2(n3436), .ZN(n3620) );
  NOR2_X1 U3661 ( .A1(n6525), .A2(n6972), .ZN(n4296) );
  NAND2_X1 U3662 ( .A1(n3979), .A2(n3978), .ZN(n4783) );
  INV_X1 U3663 ( .A(n4790), .ZN(n3978) );
  INV_X1 U3664 ( .A(n4774), .ZN(n3979) );
  NAND2_X1 U3665 ( .A1(n5516), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4228) );
  OR2_X1 U3666 ( .A1(n4419), .A2(n5917), .ZN(n4439) );
  NAND2_X1 U3667 ( .A1(n3780), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3437) );
  CLKBUF_X1 U3668 ( .A(n3655), .Z(n3631) );
  NOR2_X2 U3669 ( .A1(n5490), .A2(n5484), .ZN(n5485) );
  NOR2_X1 U3670 ( .A1(n5117), .A2(n6557), .ZN(n5116) );
  NOR2_X1 U3671 ( .A1(n3290), .A2(n6972), .ZN(n3585) );
  AND2_X1 U3672 ( .A1(n3620), .A2(n3539), .ZN(n3518) );
  NOR2_X2 U3673 ( .A1(n3502), .A2(n3506), .ZN(n3517) );
  AND2_X1 U3674 ( .A1(n4420), .A2(n5098), .ZN(n3262) );
  NAND2_X1 U3675 ( .A1(n3302), .A2(n3124), .ZN(n3326) );
  INV_X1 U3676 ( .A(n3300), .ZN(n3302) );
  BUF_X1 U3677 ( .A(n3304), .Z(n3431) );
  AND2_X2 U3678 ( .A1(n4374), .A2(n4562), .ZN(n3219) );
  AOI22_X1 U3679 ( .A1(n3213), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U3680 ( .A1(n3309), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3161) );
  BUF_X1 U3681 ( .A(n3259), .Z(n4420) );
  NAND2_X1 U3682 ( .A1(n5274), .A2(n5277), .ZN(n5276) );
  AND2_X1 U3683 ( .A1(n4771), .A2(n3895), .ZN(n3961) );
  INV_X1 U3684 ( .A(n3766), .ZN(n3759) );
  OR2_X1 U3685 ( .A1(n3375), .A2(n3374), .ZN(n3413) );
  NAND2_X1 U3686 ( .A1(n4367), .A2(n6972), .ZN(n3344) );
  INV_X1 U3687 ( .A(n3260), .ZN(n3912) );
  AND2_X2 U3688 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4375) );
  OR2_X1 U3689 ( .A1(n6661), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4337) );
  INV_X1 U3690 ( .A(n3290), .ZN(n3256) );
  AND2_X1 U3691 ( .A1(n3290), .A2(n3655), .ZN(n5171) );
  NAND2_X1 U3692 ( .A1(n4300), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4342)
         );
  OR2_X1 U3693 ( .A1(n4237), .A2(n4236), .ZN(n5492) );
  INV_X1 U3694 ( .A(n4439), .ZN(n4491) );
  OR2_X1 U3695 ( .A1(n5617), .A2(n5703), .ZN(n5293) );
  OR2_X1 U3696 ( .A1(n5603), .A2(n7008), .ZN(n5265) );
  AND2_X1 U3697 ( .A1(n5603), .A2(n7008), .ZN(n5266) );
  AND2_X1 U3698 ( .A1(n5103), .A2(n3555), .ZN(n3556) );
  NOR2_X1 U3699 ( .A1(n3795), .A2(n3794), .ZN(n4417) );
  OAI21_X1 U3700 ( .B1(n4439), .B2(n3653), .A(n3652), .ZN(n3806) );
  NAND2_X1 U3701 ( .A1(n3382), .A2(n3381), .ZN(n3405) );
  AND2_X1 U3702 ( .A1(n3626), .A2(n3625), .ZN(n4419) );
  INV_X1 U3703 ( .A(n4857), .ZN(n6323) );
  AND2_X1 U3704 ( .A1(n6557), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6553) );
  INV_X1 U3705 ( .A(n5981), .ZN(n6002) );
  OR2_X1 U3706 ( .A1(n6675), .A2(n5115), .ZN(n6011) );
  INV_X1 U3707 ( .A(n5505), .ZN(n5511) );
  XNOR2_X1 U3708 ( .A(n3779), .B(n3778), .ZN(n5328) );
  INV_X1 U3709 ( .A(n3817), .ZN(n3819) );
  AND2_X1 U3710 ( .A1(n5657), .A2(n3803), .ZN(n5644) );
  NOR2_X1 U3711 ( .A1(n5682), .A2(n3813), .ZN(n5664) );
  CLKBUF_X1 U3712 ( .A(n4398), .Z(n5178) );
  NOR2_X1 U3713 ( .A1(n3355), .A2(n3354), .ZN(n3357) );
  INV_X1 U3714 ( .A(n3349), .ZN(n3355) );
  NAND2_X1 U3715 ( .A1(n4308), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3356)
         );
  NAND2_X1 U3716 ( .A1(n3267), .A2(n3663), .ZN(n3279) );
  CLKBUF_X1 U3717 ( .A(n3365), .Z(n4315) );
  OR2_X1 U3718 ( .A1(n3516), .A2(n3515), .ZN(n3539) );
  OR2_X1 U3719 ( .A1(n3491), .A2(n3490), .ZN(n3524) );
  NOR2_X1 U3720 ( .A1(n3665), .A2(n5223), .ZN(n3671) );
  OR2_X1 U3721 ( .A1(n6688), .A2(n4333), .ZN(n4191) );
  NOR2_X1 U3722 ( .A1(n5218), .A2(n5285), .ZN(n5274) );
  NAND2_X1 U3723 ( .A1(n5203), .A2(n4113), .ZN(n5218) );
  INV_X1 U3724 ( .A(n5219), .ZN(n4113) );
  NOR2_X2 U3725 ( .A1(n5161), .A2(n5205), .ZN(n5203) );
  NOR2_X2 U3726 ( .A1(n4783), .A2(n4784), .ZN(n4785) );
  XNOR2_X1 U3727 ( .A(n3536), .B(n3535), .ZN(n3826) );
  AND2_X1 U3728 ( .A1(n4657), .A2(n4656), .ZN(n3960) );
  AND2_X1 U3729 ( .A1(n5603), .A2(n6913), .ZN(n3576) );
  CLKBUF_X1 U3730 ( .A(n3671), .Z(n3755) );
  INV_X1 U3731 ( .A(n3635), .ZN(n3638) );
  INV_X1 U3732 ( .A(n3541), .ZN(n3548) );
  NAND2_X1 U3734 ( .A1(n3327), .A2(n3326), .ZN(n3330) );
  AND2_X1 U3735 ( .A1(n3619), .A2(n3618), .ZN(n3644) );
  OR2_X1 U3736 ( .A1(n3617), .A2(n3616), .ZN(n3619) );
  OR2_X1 U3737 ( .A1(n3597), .A2(n3602), .ZN(n3624) );
  AOI21_X1 U3738 ( .B1(n3431), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3308), 
        .ZN(n3429) );
  OR2_X1 U3739 ( .A1(n6400), .A2(n4585), .ZN(n6354) );
  AND4_X1 U3740 ( .A1(n3238), .A2(n3237), .A3(n3236), .A4(n3235), .ZN(n3255)
         );
  AND4_X1 U3741 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3254)
         );
  BUF_X2 U3742 ( .A(n3182), .Z(n3288) );
  AOI22_X1 U3743 ( .A1(n3365), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U3744 ( .A1(n3449), .A2(n3448), .ZN(n4663) );
  NAND2_X1 U3745 ( .A1(n4554), .A2(n6972), .ZN(n3449) );
  INV_X1 U3746 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6539) );
  CLKBUF_X1 U3747 ( .A(n4350), .Z(n4437) );
  NAND2_X1 U3748 ( .A1(n5320), .A2(n5124), .ZN(n5962) );
  AND2_X1 U3749 ( .A1(n4432), .A2(n5126), .ZN(n6023) );
  AND2_X1 U3750 ( .A1(n5799), .A2(n4299), .ZN(n4211) );
  CLKBUF_X1 U3751 ( .A(n5488), .Z(n5489) );
  OR2_X1 U3752 ( .A1(n4190), .A2(n5565), .ZN(n4210) );
  AND2_X1 U3753 ( .A1(n4148), .A2(n4147), .ZN(n5277) );
  BUF_X1 U3754 ( .A(n5276), .Z(n5388) );
  CLKBUF_X1 U3755 ( .A(n5274), .Z(n5275) );
  NAND2_X1 U3756 ( .A1(n4110), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4127)
         );
  CLKBUF_X1 U3757 ( .A(n5218), .Z(n5284) );
  AND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4092), .ZN(n4110)
         );
  CLKBUF_X1 U3759 ( .A(n5203), .Z(n5204) );
  NOR2_X1 U3760 ( .A1(n4074), .A2(n5609), .ZN(n4075) );
  INV_X1 U3761 ( .A(n4073), .ZN(n4074) );
  NAND2_X1 U3762 ( .A1(n4075), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4091)
         );
  AND2_X1 U3764 ( .A1(n4042), .A2(n4041), .ZN(n5066) );
  NAND2_X1 U3765 ( .A1(n4021), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4026)
         );
  AND3_X1 U3766 ( .A1(n4025), .A2(n4024), .A3(n4023), .ZN(n4993) );
  INV_X1 U3767 ( .A(n4994), .ZN(n5067) );
  CLKBUF_X1 U3768 ( .A(n4785), .Z(n4786) );
  NAND2_X1 U3769 ( .A1(n3980), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3981)
         );
  NOR2_X1 U3770 ( .A1(n6943), .A2(n3981), .ZN(n4021) );
  AND2_X1 U3771 ( .A1(n3877), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3847)
         );
  NOR2_X1 U3772 ( .A1(n6794), .A2(n3878), .ZN(n3877) );
  OR2_X1 U3773 ( .A1(n4798), .A2(n4799), .ZN(n4900) );
  NOR2_X1 U3774 ( .A1(n3955), .A2(n5154), .ZN(n3827) );
  CLKBUF_X1 U3775 ( .A(n4655), .Z(n4770) );
  NOR2_X1 U3776 ( .A1(n3936), .A2(n3900), .ZN(n3945) );
  INV_X1 U3777 ( .A(n3922), .ZN(n3937) );
  NAND2_X1 U3778 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3937), .ZN(n3936)
         );
  NAND2_X1 U3779 ( .A1(n3392), .A2(n3391), .ZN(n6104) );
  NAND2_X1 U3780 ( .A1(n3766), .A2(n5164), .ZN(n4478) );
  AND2_X1 U3781 ( .A1(n5339), .A2(n5164), .ZN(n5336) );
  NOR2_X1 U3782 ( .A1(n5356), .A2(n3801), .ZN(n5331) );
  AND2_X1 U3783 ( .A1(n5393), .A2(n5299), .ZN(n5502) );
  NAND2_X1 U3784 ( .A1(n5502), .A2(n5501), .ZN(n5500) );
  NOR2_X2 U3785 ( .A1(n5394), .A2(n5395), .ZN(n5393) );
  OR2_X1 U3786 ( .A1(n5617), .A2(n6702), .ZN(n5292) );
  NAND2_X1 U3787 ( .A1(n4778), .A2(n4779), .ZN(n4792) );
  OR2_X1 U3788 ( .A1(n5603), .A2(n3554), .ZN(n5103) );
  OR2_X1 U3789 ( .A1(n5603), .A2(n5079), .ZN(n5054) );
  AND2_X1 U3790 ( .A1(n3707), .A2(n3706), .ZN(n5042) );
  INV_X1 U3791 ( .A(n4474), .ZN(n3676) );
  INV_X1 U3792 ( .A(n4475), .ZN(n3677) );
  AND2_X1 U3793 ( .A1(n3681), .A2(n3680), .ZN(n4504) );
  AND2_X1 U3794 ( .A1(n5253), .A2(n3805), .ZN(n5693) );
  XNOR2_X1 U3795 ( .A(n4575), .B(n5725), .ZN(n4554) );
  NAND2_X1 U3796 ( .A1(n3632), .A2(n3631), .ZN(n3654) );
  INV_X1 U3797 ( .A(n5989), .ZN(n6325) );
  OR2_X1 U3798 ( .A1(n6354), .A2(n6323), .ZN(n6332) );
  OR2_X1 U3799 ( .A1(n4747), .A2(n6353), .ZN(n4744) );
  OR2_X1 U3800 ( .A1(n4662), .A2(n4585), .ZN(n4747) );
  BUF_X1 U3801 ( .A(n3260), .Z(n4626) );
  INV_X1 U3802 ( .A(n6685), .ZN(n5977) );
  INV_X1 U3803 ( .A(n6000), .ZN(n6692) );
  AND2_X1 U3805 ( .A1(n5172), .A2(n5802), .ZN(n5981) );
  INV_X1 U3806 ( .A(n5507), .ZN(n5512) );
  NAND2_X1 U3807 ( .A1(n4426), .A2(n4425), .ZN(n5505) );
  OR2_X1 U3808 ( .A1(n5475), .A2(n5360), .ZN(n5361) );
  NOR2_X1 U3809 ( .A1(n6023), .A2(n6677), .ZN(n6039) );
  INV_X1 U3810 ( .A(n6071), .ZN(n4551) );
  XNOR2_X1 U3811 ( .A(n4344), .B(n4343), .ZN(n5117) );
  OR2_X1 U3812 ( .A1(n4342), .A2(n4341), .ZN(n4344) );
  INV_X1 U3813 ( .A(n5535), .ZN(n5832) );
  OR2_X1 U3814 ( .A1(n5486), .A2(n5485), .ZN(n5783) );
  INV_X1 U3815 ( .A(n6110), .ZN(n5622) );
  AND2_X1 U3816 ( .A1(n5924), .A2(n4338), .ZN(n6099) );
  AND2_X1 U3817 ( .A1(n5664), .A2(n3815), .ZN(n5657) );
  OR2_X1 U3818 ( .A1(n5670), .A2(n3816), .ZN(n5661) );
  OR2_X1 U3819 ( .A1(n3800), .A2(n5863), .ZN(n5682) );
  CLKBUF_X1 U3820 ( .A(n5286), .Z(n5288) );
  CLKBUF_X1 U3821 ( .A(n5263), .Z(n5264) );
  CLKBUF_X1 U3822 ( .A(n5245), .Z(n5247) );
  INV_X1 U3823 ( .A(n5881), .ZN(n6190) );
  NAND2_X2 U3824 ( .A1(n3394), .A2(n3130), .ZN(n4857) );
  INV_X1 U3825 ( .A(n3405), .ZN(n3394) );
  CLKBUF_X1 U3826 ( .A(n6324), .Z(n6447) );
  CLKBUF_X1 U3827 ( .A(n4554), .Z(n5989) );
  INV_X1 U3828 ( .A(n6352), .ZN(n6311) );
  AND2_X1 U3829 ( .A1(n6451), .A2(n6450), .ZN(n6519) );
  INV_X2 U3830 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6972) );
  INV_X1 U3831 ( .A(n4397), .ZN(n6558) );
  INV_X1 U3832 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U3833 ( .A1(n3821), .A2(n3820), .ZN(n3822) );
  NOR2_X1 U3834 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  NAND2_X1 U3835 ( .A1(n5362), .A2(n5361), .ZN(n5366) );
  XOR2_X1 U3836 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5332), .Z(n3122) );
  OR2_X1 U3837 ( .A1(n3301), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3124)
         );
  NAND2_X1 U3838 ( .A1(n3536), .A2(n3547), .ZN(n3558) );
  INV_X1 U3839 ( .A(n3558), .ZN(n5296) );
  BUF_X2 U3840 ( .A(n3460), .Z(n4177) );
  INV_X1 U3841 ( .A(n5580), .ZN(n6193) );
  NOR2_X2 U3842 ( .A1(n6595), .A2(n6684), .ZN(n6638) );
  NOR3_X4 U3843 ( .A1(n6289), .A2(n6323), .A3(n4585), .ZN(n6267) );
  AND2_X1 U3844 ( .A1(n5046), .A2(n3709), .ZN(n4778) );
  OR2_X2 U3845 ( .A1(n3192), .A2(n3191), .ZN(n3663) );
  AND2_X2 U3846 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4562) );
  OR2_X1 U3847 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3125)
         );
  AND4_X1 U3848 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3126)
         );
  OR2_X1 U3849 ( .A1(n3293), .A2(n5122), .ZN(n3127) );
  AND4_X1 U3850 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3128)
         );
  AND4_X1 U3851 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3129)
         );
  OR2_X1 U3852 ( .A1(n3393), .A2(n3133), .ZN(n3130) );
  OR2_X1 U3853 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3131)
         );
  AND4_X1 U3854 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3132)
         );
  AND2_X1 U3855 ( .A1(n3377), .A2(n3376), .ZN(n3133) );
  INV_X1 U3856 ( .A(n5319), .ZN(n3395) );
  OR2_X1 U3857 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3134)
         );
  OR2_X1 U3858 ( .A1(n5617), .A2(n6760), .ZN(n3135) );
  OR2_X1 U3859 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3136)
         );
  AND2_X1 U3860 ( .A1(n5359), .A2(n5630), .ZN(n3137) );
  INV_X1 U3861 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3900) );
  OR2_X1 U3862 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3138)
         );
  INV_X1 U3863 ( .A(n5204), .ZN(n5220) );
  CLKBUF_X1 U3864 ( .A(n4375), .Z(n4376) );
  AND2_X1 U3865 ( .A1(n3258), .A2(n3257), .ZN(n3283) );
  NAND2_X1 U3866 ( .A1(n3633), .A2(n5319), .ZN(n3258) );
  NOR2_X1 U3867 ( .A1(n3635), .A2(n3263), .ZN(n3264) );
  AND2_X1 U3868 ( .A1(n6355), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3594)
         );
  OR2_X1 U3869 ( .A1(n3470), .A2(n3469), .ZN(n3525) );
  OR2_X1 U3870 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  AOI22_X1 U3871 ( .A1(n3331), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3119), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U3872 ( .A1(n3612), .A2(n4493), .ZN(n3268) );
  INV_X1 U3873 ( .A(n3182), .ZN(n3165) );
  NAND2_X1 U3874 ( .A1(n3357), .A2(n3356), .ZN(n3363) );
  OR2_X1 U3875 ( .A1(n3293), .A2(n4626), .ZN(n3261) );
  AOI22_X1 U3876 ( .A1(n3348), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U3877 ( .A1(n3297), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3300) );
  OR2_X1 U3878 ( .A1(n3405), .A2(n3387), .ZN(n3388) );
  AOI22_X1 U3879 ( .A1(n3331), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3156) );
  OR2_X1 U3880 ( .A1(n3363), .A2(n3362), .ZN(n3541) );
  NOR2_X1 U3881 ( .A1(n3322), .A2(n3321), .ZN(n3450) );
  OR2_X1 U3882 ( .A1(n5603), .A2(n6117), .ZN(n3555) );
  NAND2_X1 U3883 ( .A1(n3663), .A2(n3788), .ZN(n3636) );
  XNOR2_X1 U3884 ( .A(n3494), .B(n3503), .ZN(n3944) );
  INV_X1 U3885 ( .A(n4301), .ZN(n4300) );
  INV_X1 U3886 ( .A(n4277), .ZN(n4275) );
  INV_X1 U3887 ( .A(n4091), .ZN(n4092) );
  INV_X1 U3888 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6794) );
  AND2_X1 U3889 ( .A1(n5603), .A2(n6117), .ZN(n3557) );
  BUF_X1 U3890 ( .A(n3328), .Z(n3329) );
  INV_X1 U3891 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3287) );
  NAND2_X1 U3892 ( .A1(n3133), .A2(n3393), .ZN(n3381) );
  OR2_X1 U3893 ( .A1(n3447), .A2(n3446), .ZN(n3473) );
  AND2_X1 U3894 ( .A1(n4370), .A2(n5122), .ZN(n4350) );
  INV_X1 U3895 ( .A(n3277), .ZN(n3655) );
  INV_X1 U3896 ( .A(n4296), .ZN(n4330) );
  INV_X1 U3897 ( .A(n5066), .ZN(n4043) );
  NAND2_X1 U3898 ( .A1(n3670), .A2(n3669), .ZN(n4475) );
  NOR2_X1 U3899 ( .A1(n4621), .A2(n3663), .ZN(n4422) );
  NAND2_X1 U3900 ( .A1(n3288), .A2(n3912), .ZN(n3267) );
  NAND2_X1 U3901 ( .A1(n4275), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4301)
         );
  NOR2_X1 U3902 ( .A1(n4127), .A2(n6790), .ZN(n4145) );
  AND2_X1 U3903 ( .A1(n4077), .A2(n4076), .ZN(n5162) );
  AND2_X1 U3904 ( .A1(n3847), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3962)
         );
  NAND2_X1 U3905 ( .A1(n3832), .A2(n3831), .ZN(n4771) );
  NAND2_X1 U3906 ( .A1(n5329), .A2(n5546), .ZN(n5356) );
  OAI21_X1 U3907 ( .B1(n5104), .B2(n3557), .A(n3556), .ZN(n5184) );
  OR2_X1 U3908 ( .A1(n3655), .A2(n3290), .ZN(n3665) );
  OR2_X1 U3909 ( .A1(n3624), .A2(n3623), .ZN(n3625) );
  AND2_X1 U3910 ( .A1(n4665), .A2(n6447), .ZN(n6206) );
  XNOR2_X1 U3911 ( .A(n3458), .B(n4663), .ZN(n3933) );
  NAND2_X1 U3912 ( .A1(n3435), .A2(n3434), .ZN(n5725) );
  NOR2_X1 U3913 ( .A1(n4231), .A2(n5796), .ZN(n4232) );
  AND2_X1 U3914 ( .A1(n5117), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5118) );
  AND2_X1 U3915 ( .A1(n6011), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5320) );
  INV_X1 U3916 ( .A(n4428), .ZN(n4424) );
  INV_X1 U3917 ( .A(n5311), .ZN(n4195) );
  AND2_X1 U3918 ( .A1(n4658), .A2(n3960), .ZN(n4655) );
  OR2_X1 U3919 ( .A1(n4254), .A2(n6762), .ZN(n4277) );
  NAND2_X1 U3920 ( .A1(n4145), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4190)
         );
  OR2_X1 U3921 ( .A1(n5603), .A2(n3570), .ZN(n3571) );
  INV_X1 U3922 ( .A(n5296), .ZN(n5603) );
  AND2_X1 U3923 ( .A1(n3962), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3980)
         );
  INV_X1 U3924 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5154) );
  INV_X1 U3925 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3818) );
  AOI21_X1 U3927 ( .B1(n5593), .B2(n3575), .A(n3574), .ZN(n5553) );
  INV_X1 U3928 ( .A(n5296), .ZN(n5617) );
  NOR2_X1 U3929 ( .A1(n5617), .A2(n5197), .ZN(n5188) );
  INV_X1 U3930 ( .A(n3665), .ZN(n4428) );
  NAND2_X1 U3931 ( .A1(n3400), .A2(n3399), .ZN(n4509) );
  INV_X1 U3932 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3139) );
  OR3_X1 U3933 ( .A1(n6289), .A2(n4857), .A3(n4585), .ZN(n6275) );
  INV_X1 U3934 ( .A(n4663), .ZN(n4664) );
  INV_X1 U3935 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6534) );
  OR2_X1 U3936 ( .A1(n4747), .A2(n6323), .ZN(n6516) );
  NAND2_X1 U3937 ( .A1(n4232), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4254)
         );
  NOR2_X1 U3938 ( .A1(n5962), .A2(n5315), .ZN(n5942) );
  AND2_X1 U3939 ( .A1(n5320), .A2(n5131), .ZN(n6686) );
  AND2_X1 U3940 ( .A1(n5320), .A2(n5121), .ZN(n6000) );
  AND2_X1 U3941 ( .A1(n6011), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6685) );
  OR2_X1 U3942 ( .A1(n5336), .A2(n5335), .ZN(n5342) );
  INV_X1 U3943 ( .A(n5098), .ZN(n5516) );
  AND2_X1 U3944 ( .A1(n5515), .A2(n5100), .ZN(n6020) );
  INV_X1 U3945 ( .A(n5515), .ZN(n6019) );
  INV_X1 U3946 ( .A(n3290), .ZN(n5122) );
  INV_X1 U3947 ( .A(n6060), .ZN(n6072) );
  OR2_X1 U3948 ( .A1(n5616), .A2(n5602), .ZN(n5851) );
  OR2_X1 U3949 ( .A1(n4900), .A2(n4899), .ZN(n5040) );
  NAND2_X1 U3950 ( .A1(n3827), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3878)
         );
  NAND2_X1 U3951 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3945), .ZN(n3955)
         );
  NAND2_X1 U3952 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3922) );
  BUF_X1 U3953 ( .A(n5329), .Z(n5547) );
  NOR2_X1 U3954 ( .A1(n7008), .A2(n5908), .ZN(n5892) );
  INV_X1 U3955 ( .A(n6193), .ZN(n6178) );
  INV_X1 U3956 ( .A(n6195), .ZN(n6180) );
  NOR2_X1 U3957 ( .A1(n6942), .A2(n4419), .ZN(n4397) );
  INV_X1 U3958 ( .A(n5004), .ZN(n5036) );
  INV_X1 U3959 ( .A(n4907), .ZN(n6233) );
  INV_X1 U3960 ( .A(n6280), .ZN(n6313) );
  INV_X1 U3961 ( .A(n6332), .ZN(n6389) );
  INV_X1 U3962 ( .A(n4863), .ZN(n6390) );
  INV_X1 U3963 ( .A(n6326), .ZN(n4820) );
  INV_X1 U3964 ( .A(n6516), .ZN(n4764) );
  INV_X1 U3965 ( .A(n4944), .ZN(n4988) );
  INV_X1 U3966 ( .A(n4705), .ZN(n4735) );
  INV_X1 U3967 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6557) );
  INV_X1 U3968 ( .A(n6686), .ZN(n5811) );
  NAND2_X1 U3969 ( .A1(n6011), .A2(n5116), .ZN(n5802) );
  INV_X1 U3970 ( .A(n5509), .ZN(n5514) );
  NAND2_X1 U3971 ( .A1(n6052), .A2(n4492), .ZN(n5515) );
  INV_X1 U3972 ( .A(n6023), .ZN(n6051) );
  NAND2_X1 U3973 ( .A1(n4491), .A2(n4430), .ZN(n6060) );
  OR2_X1 U3974 ( .A1(n6099), .A2(n4511), .ZN(n6110) );
  NAND2_X1 U3975 ( .A1(n4491), .A2(n4351), .ZN(n5924) );
  INV_X1 U3976 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6355) );
  INV_X1 U3977 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6397) );
  OR2_X1 U3978 ( .A1(n6289), .A2(n6396), .ZN(n6352) );
  OR2_X1 U3979 ( .A1(n6400), .A2(n4906), .ZN(n6440) );
  OR2_X1 U3980 ( .A1(n6400), .A2(n6396), .ZN(n6523) );
  OR2_X1 U3981 ( .A1(n4747), .A2(n4857), .ZN(n4992) );
  OAI21_X1 U3982 ( .B1(n3823), .B2(n5881), .A(n3822), .ZN(U2987) );
  AND2_X2 U3983 ( .A1(n4381), .A2(n4562), .ZN(n3336) );
  INV_X1 U3984 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3935) );
  AND2_X2 U3985 ( .A1(n3935), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3146)
         );
  AND2_X2 U3986 ( .A1(n3146), .A2(n4374), .ZN(n3309) );
  AOI22_X1 U3987 ( .A1(n3336), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3145) );
  INV_X1 U3988 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3140) );
  AND2_X2 U3989 ( .A1(n3148), .A2(n4381), .ZN(n3348) );
  INV_X1 U3990 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3141) );
  AND2_X2 U3991 ( .A1(n3141), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3147)
         );
  AND2_X2 U3992 ( .A1(n3146), .A2(n3147), .ZN(n3247) );
  AOI22_X1 U3993 ( .A1(n3348), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3144) );
  NOR2_X4 U3994 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4563) );
  AND2_X2 U3995 ( .A1(n4381), .A2(n4563), .ZN(n3460) );
  AND2_X2 U3996 ( .A1(n4374), .A2(n4563), .ZN(n3310) );
  AOI22_X1 U3997 ( .A1(n3460), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3143) );
  AND2_X2 U3998 ( .A1(n3148), .A2(n4375), .ZN(n3365) );
  AND2_X2 U3999 ( .A1(n4562), .A2(n4375), .ZN(n3316) );
  AOI22_X1 U4000 ( .A1(n3365), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3142) );
  NAND4_X1 U4001 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3154)
         );
  AND2_X2 U4002 ( .A1(n3148), .A2(n4374), .ZN(n3350) );
  AND2_X2 U4003 ( .A1(n3147), .A2(n4563), .ZN(n3234) );
  AOI22_X1 U4004 ( .A1(n3350), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3152) );
  AND2_X2 U4005 ( .A1(n4381), .A2(n3146), .ZN(n3364) );
  AND2_X2 U4006 ( .A1(n3147), .A2(n4562), .ZN(n3193) );
  AOI22_X1 U4007 ( .A1(n3364), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3151) );
  AND2_X2 U4008 ( .A1(n3146), .A2(n4375), .ZN(n3218) );
  AOI22_X1 U4009 ( .A1(n3218), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3150) );
  AND2_X2 U4010 ( .A1(n3148), .A2(n3147), .ZN(n3331) );
  NAND4_X1 U4011 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3153)
         );
  OR2_X2 U4012 ( .A1(n3154), .A2(n3153), .ZN(n3182) );
  AOI22_X1 U4013 ( .A1(n3364), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4014 ( .A1(n3350), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4015 ( .A1(n3460), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4016 ( .A1(n3348), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4017 ( .A1(n3364), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4018 ( .A1(n3309), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4019 ( .A1(n3350), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4020 ( .A1(n3460), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4021 ( .A1(n3348), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4022 ( .A1(n3331), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4023 ( .A1(n3213), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4024 ( .A1(n3218), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3170) );
  AND2_X2 U4025 ( .A1(n3129), .A2(n3132), .ZN(n3780) );
  AOI22_X1 U4026 ( .A1(n3364), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3193), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4027 ( .A1(n3460), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4028 ( .A1(n3213), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4029 ( .A1(n3350), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4030 ( .A1(n3247), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4031 ( .A1(n3309), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4032 ( .A1(n3331), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3178) );
  AND2_X2 U4033 ( .A1(n3128), .A2(n3126), .ZN(n3788) );
  NAND2_X1 U4034 ( .A1(n3232), .A2(n4621), .ZN(n3204) );
  AOI22_X1 U4035 ( .A1(n3331), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4036 ( .A1(n3348), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3185) );
  BUF_X2 U4037 ( .A(n3219), .Z(n3315) );
  AOI22_X1 U4038 ( .A1(n3218), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4039 ( .A1(n3213), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4040 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3192)
         );
  BUF_X2 U4041 ( .A(n3193), .Z(n3208) );
  AOI22_X1 U4042 ( .A1(n3350), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4043 ( .A1(n3309), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4044 ( .A1(n3364), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4045 ( .A1(n3460), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3187) );
  NAND4_X1 U4046 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3191)
         );
  AOI22_X1 U4047 ( .A1(n3309), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4048 ( .A1(n3364), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4049 ( .A1(n3350), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4050 ( .A1(n3460), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3194) );
  NAND4_X1 U4051 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3203)
         );
  AOI22_X1 U4052 ( .A1(n3331), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4053 ( .A1(n3348), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4054 ( .A1(n3218), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3315), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4055 ( .A1(n3213), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3198) );
  NAND4_X1 U4056 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3202)
         );
  AND3_X2 U4057 ( .A1(n3204), .A2(n3279), .A3(n5098), .ZN(n3207) );
  NAND2_X1 U4058 ( .A1(n3259), .A2(n3788), .ZN(n3205) );
  MUX2_X2 U4059 ( .A(n3232), .B(n3205), .S(n3260), .Z(n3206) );
  NAND2_X2 U4060 ( .A1(n3207), .A2(n3206), .ZN(n3294) );
  NAND2_X1 U4061 ( .A1(n3309), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4062 ( .A1(n3350), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4063 ( .A1(n3234), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4064 ( .A1(n3208), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3209)
         );
  NAND2_X1 U4065 ( .A1(n3331), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3217)
         );
  NAND2_X1 U4066 ( .A1(n3365), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4067 ( .A1(n3316), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4068 ( .A1(n3213), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4069 ( .A1(n3247), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4070 ( .A1(n3348), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4071 ( .A1(n3218), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4072 ( .A1(n3219), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4073 ( .A1(n3364), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4074 ( .A1(n3336), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4075 ( .A1(n3460), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4076 ( .A1(n3310), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3224) );
  AND4_X4 U4077 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3290)
         );
  NAND2_X1 U4078 ( .A1(n3294), .A2(n3290), .ZN(n3265) );
  INV_X1 U4079 ( .A(n3232), .ZN(n3233) );
  NAND2_X2 U4080 ( .A1(n3233), .A2(n5098), .ZN(n3633) );
  NAND2_X1 U4081 ( .A1(n3336), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3238)
         );
  NAND2_X1 U4082 ( .A1(n3350), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U4083 ( .A1(n3309), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3236) );
  NAND2_X1 U4084 ( .A1(n3234), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4085 ( .A1(n3365), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3242)
         );
  NAND2_X1 U4086 ( .A1(n3348), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4087 ( .A1(n3218), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4088 ( .A1(n3316), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3239)
         );
  NAND2_X1 U4089 ( .A1(n3364), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4090 ( .A1(n3460), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U4091 ( .A1(n3208), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3244)
         );
  NAND2_X1 U4092 ( .A1(n3310), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4093 ( .A1(n3331), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3251)
         );
  NAND2_X1 U4094 ( .A1(n3247), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4095 ( .A1(n3315), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3249)
         );
  NAND2_X1 U4096 ( .A1(n3213), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3248) );
  AND4_X2 U4097 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3252)
         );
  AND2_X2 U4098 ( .A1(n3256), .A2(n3655), .ZN(n5319) );
  NAND2_X2 U4099 ( .A1(n3277), .A2(n3663), .ZN(n3661) );
  OR2_X1 U4100 ( .A1(n3293), .A2(n3661), .ZN(n3257) );
  INV_X1 U4101 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6595) );
  INV_X1 U4102 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U4103 ( .A1(n6584), .A2(n6595), .ZN(n6585) );
  AOI21_X1 U4104 ( .B1(n6595), .B2(n6584), .A(n6585), .ZN(n3627) );
  NOR2_X1 U4105 ( .A1(n3277), .A2(n3627), .ZN(n3291) );
  NAND2_X1 U4106 ( .A1(n3290), .A2(n3277), .ZN(n5176) );
  OAI211_X1 U4107 ( .C1(n3291), .C2(n4615), .A(n3414), .B(n5176), .ZN(n3263)
         );
  NAND3_X1 U4108 ( .A1(n3265), .A2(n3283), .A3(n3264), .ZN(n3266) );
  NAND2_X1 U4109 ( .A1(n3266), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3269) );
  INV_X2 U4110 ( .A(n3780), .ZN(n4643) );
  NAND2_X2 U4111 ( .A1(n3269), .A2(n3268), .ZN(n3304) );
  NAND2_X1 U4112 ( .A1(n3304), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3274) );
  INV_X1 U4113 ( .A(n6553), .ZN(n3271) );
  NAND2_X1 U4114 ( .A1(n6942), .A2(n6557), .ZN(n6661) );
  INV_X1 U4115 ( .A(n4337), .ZN(n3270) );
  MUX2_X1 U4116 ( .A(n3271), .B(n3270), .S(n6355), .Z(n3272) );
  INV_X1 U4117 ( .A(n3272), .ZN(n3273) );
  NAND2_X1 U4118 ( .A1(n3274), .A2(n3273), .ZN(n3347) );
  INV_X1 U4119 ( .A(n3293), .ZN(n3656) );
  OAI22_X1 U4120 ( .A1(n3656), .A2(n5176), .B1(n3290), .B2(n3788), .ZN(n3275)
         );
  AOI21_X1 U4121 ( .B1(n3294), .B2(n5171), .A(n3275), .ZN(n3792) );
  NAND2_X1 U4122 ( .A1(n4493), .A2(n4643), .ZN(n3276) );
  NAND2_X1 U4123 ( .A1(n3276), .A2(n3663), .ZN(n3278) );
  OAI21_X1 U4124 ( .B1(n3635), .B2(n3278), .A(n4605), .ZN(n3282) );
  NOR2_X1 U4125 ( .A1(n6661), .A2(n6972), .ZN(n6567) );
  NAND2_X1 U4126 ( .A1(n5319), .A2(n3279), .ZN(n3281) );
  AND4_X1 U4127 ( .A1(n3912), .A2(n3290), .A3(n4643), .A4(n5098), .ZN(n3280)
         );
  NAND2_X1 U4128 ( .A1(n3280), .A2(n4422), .ZN(n4557) );
  NAND4_X1 U4129 ( .A1(n3282), .A2(n6567), .A3(n3281), .A4(n4557), .ZN(n3285)
         );
  INV_X1 U4130 ( .A(n3283), .ZN(n3284) );
  NOR2_X1 U4131 ( .A1(n3285), .A2(n3284), .ZN(n3286) );
  NAND2_X1 U4132 ( .A1(n3792), .A2(n3286), .ZN(n3345) );
  AND2_X2 U4133 ( .A1(n3347), .A2(n3345), .ZN(n3328) );
  INV_X1 U4134 ( .A(n3304), .ZN(n3299) );
  INV_X1 U4135 ( .A(n3288), .ZN(n5099) );
  NAND3_X1 U4136 ( .A1(n5171), .A2(n4422), .A3(n5099), .ZN(n4368) );
  NAND2_X1 U4137 ( .A1(n4626), .A2(n5098), .ZN(n5097) );
  INV_X1 U4138 ( .A(n3781), .ZN(n3296) );
  NAND2_X1 U4139 ( .A1(n3414), .A2(n5099), .ZN(n3289) );
  NOR2_X2 U4140 ( .A1(n3633), .A2(n3289), .ZN(n4370) );
  INV_X1 U4141 ( .A(n3291), .ZN(n3292) );
  NAND2_X1 U4142 ( .A1(n4350), .A2(n3292), .ZN(n3295) );
  NOR2_X2 U4143 ( .A1(n3294), .A2(n3127), .ZN(n3632) );
  NAND3_X1 U4144 ( .A1(n3296), .A2(n3295), .A3(n3654), .ZN(n3297) );
  XNOR2_X1 U4145 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6320) );
  OAI22_X1 U4146 ( .A1(n4337), .A2(n6320), .B1(n6553), .B2(n6534), .ZN(n3301)
         );
  INV_X1 U4147 ( .A(n3301), .ZN(n3298) );
  NAND2_X1 U4148 ( .A1(n3328), .A2(n3327), .ZN(n3303) );
  AND2_X1 U4149 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4150 ( .A1(n3305), .A2(n6539), .ZN(n6398) );
  INV_X1 U4151 ( .A(n3305), .ZN(n3306) );
  NAND2_X1 U4152 ( .A1(n3306), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3307) );
  AND2_X1 U4153 ( .A1(n6398), .A2(n3307), .ZN(n4708) );
  OAI22_X1 U4154 ( .A1(n4708), .A2(n4337), .B1(n6553), .B2(n6539), .ZN(n3308)
         );
  AOI22_X1 U4155 ( .A1(n4305), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3314) );
  BUF_X2 U4156 ( .A(n3336), .Z(n4313) );
  AOI22_X1 U4157 ( .A1(n3121), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3313) );
  BUF_X2 U4158 ( .A(n3208), .Z(n4306) );
  AOI22_X1 U4159 ( .A1(n4178), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4160 ( .A1(n4177), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4161 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3322)
         );
  AOI22_X1 U4163 ( .A1(n4317), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4164 ( .A1(n4284), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3319) );
  BUF_X2 U4165 ( .A(n3218), .Z(n4314) );
  BUF_X2 U4166 ( .A(n3315), .Z(n4308) );
  AOI22_X1 U4167 ( .A1(n4314), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3318) );
  INV_X1 U4168 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U4169 ( .A1(n4316), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4170 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3321)
         );
  NOR2_X1 U4171 ( .A1(n3437), .A2(n3450), .ZN(n3323) );
  AOI21_X2 U4172 ( .B1(n4398), .B2(n6972), .A(n3323), .ZN(n3325) );
  INV_X1 U4173 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6937) );
  NAND2_X1 U4174 ( .A1(n3290), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3436) );
  OAI22_X1 U4175 ( .A1(n3597), .A2(n6937), .B1(n3450), .B2(n3436), .ZN(n3324)
         );
  XNOR2_X2 U4176 ( .A(n3325), .B(n3324), .ZN(n3427) );
  AOI22_X1 U4177 ( .A1(n4305), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4178 ( .A1(n4317), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4179 ( .A1(n4284), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4180 ( .A1(n3121), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3332) );
  NAND4_X1 U4181 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3342)
         );
  AOI22_X1 U4182 ( .A1(n4178), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4183 ( .A1(n4177), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4184 ( .A1(n4314), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4185 ( .A1(n4316), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4186 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3341)
         );
  INV_X1 U4187 ( .A(n3412), .ZN(n3383) );
  OR2_X1 U4188 ( .A1(n3437), .A2(n3383), .ZN(n3343) );
  INV_X1 U4189 ( .A(n3345), .ZN(n3346) );
  XNOR2_X1 U4190 ( .A(n3347), .B(n3346), .ZN(n3914) );
  NAND2_X1 U4191 ( .A1(n3914), .A2(n6972), .ZN(n3382) );
  INV_X1 U4192 ( .A(n3437), .ZN(n3377) );
  AOI22_X1 U4193 ( .A1(n4284), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4194 ( .A1(n4178), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4195 ( .A1(n4313), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4196 ( .A1(n4315), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3351)
         );
  NAND3_X1 U4197 ( .A1(n3353), .A2(n3352), .A3(n3351), .ZN(n3354) );
  AOI22_X1 U4198 ( .A1(n4317), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4199 ( .A1(n3120), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4200 ( .A1(n3121), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4201 ( .A1(n4316), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3358) );
  NAND4_X1 U4202 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3362)
         );
  AOI22_X1 U4203 ( .A1(n3121), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4204 ( .A1(n4284), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4205 ( .A1(n4285), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4206 ( .A1(n3120), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4207 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3375)
         );
  AOI22_X1 U4208 ( .A1(n4178), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4209 ( .A1(n4313), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4210 ( .A1(n4317), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4211 ( .A1(n4316), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3370) );
  NAND4_X1 U4212 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3374)
         );
  XNOR2_X1 U4213 ( .A(n3548), .B(n3413), .ZN(n3376) );
  NAND2_X1 U4214 ( .A1(n3290), .A2(n3413), .ZN(n3378) );
  OAI211_X1 U4215 ( .C1(n3548), .C2(n4643), .A(STATE2_REG_0__SCAN_IN), .B(
        n3378), .ZN(n3379) );
  AOI21_X1 U4216 ( .B1(n3612), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n3379), 
        .ZN(n3380) );
  INV_X1 U4217 ( .A(n3380), .ZN(n3393) );
  NOR2_X1 U4218 ( .A1(n3437), .A2(n3548), .ZN(n3404) );
  NAND2_X1 U4219 ( .A1(n3612), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3386) );
  OAI22_X1 U4220 ( .A1(n3437), .A2(n3541), .B1(n3436), .B2(n3383), .ZN(n3384)
         );
  INV_X1 U4221 ( .A(n3384), .ZN(n3385) );
  NAND2_X1 U4222 ( .A1(n3386), .A2(n3385), .ZN(n3406) );
  OR2_X1 U4223 ( .A1(n3404), .A2(n3406), .ZN(n3387) );
  AND2_X2 U4224 ( .A1(n3409), .A2(n3388), .ZN(n3426) );
  INV_X1 U4225 ( .A(n3426), .ZN(n3389) );
  XNOR2_X1 U4226 ( .A(n3427), .B(n3389), .ZN(n3905) );
  NAND2_X1 U4227 ( .A1(n4615), .A2(n4605), .ZN(n3602) );
  INV_X1 U4228 ( .A(n3602), .ZN(n3537) );
  NAND2_X1 U4229 ( .A1(n3905), .A2(n3537), .ZN(n3392) );
  NAND2_X1 U4230 ( .A1(n3412), .A2(n3413), .ZN(n3451) );
  XNOR2_X1 U4231 ( .A(n3451), .B(n3450), .ZN(n3390) );
  AND2_X1 U4232 ( .A1(n3290), .A2(n3663), .ZN(n3396) );
  AOI21_X1 U4233 ( .B1(n3390), .B2(n5319), .A(n3396), .ZN(n3391) );
  NAND2_X1 U4234 ( .A1(n6104), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3421)
         );
  INV_X1 U4235 ( .A(n3396), .ZN(n3397) );
  OAI21_X1 U4236 ( .B1(n3395), .B2(n3413), .A(n3397), .ZN(n3398) );
  INV_X1 U4237 ( .A(n3398), .ZN(n3399) );
  NAND2_X1 U4238 ( .A1(n4509), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3401)
         );
  INV_X1 U4239 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U4240 ( .A1(n3401), .A2(n4464), .ZN(n3403) );
  AND2_X1 U4241 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4242 ( .A1(n4509), .A2(n3402), .ZN(n3419) );
  INV_X1 U4243 ( .A(n3406), .ZN(n3407) );
  INV_X1 U4244 ( .A(n3409), .ZN(n3410) );
  NAND2_X1 U4245 ( .A1(n3907), .A2(n3537), .ZN(n3418) );
  OAI21_X1 U4246 ( .B1(n3413), .B2(n3412), .A(n3451), .ZN(n3415) );
  OAI211_X1 U4247 ( .C1(n3415), .C2(n3395), .A(n3414), .B(n4615), .ZN(n3416)
         );
  INV_X1 U4248 ( .A(n3416), .ZN(n3417) );
  NAND2_X1 U4249 ( .A1(n3418), .A2(n3417), .ZN(n4463) );
  INV_X1 U4250 ( .A(n3419), .ZN(n3420) );
  AOI21_X2 U4251 ( .B1(n4462), .B2(n4463), .A(n3420), .ZN(n6101) );
  NAND2_X1 U4252 ( .A1(n3421), .A2(n6101), .ZN(n3425) );
  INV_X1 U4253 ( .A(n6104), .ZN(n3423) );
  INV_X1 U4254 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4255 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  AND2_X1 U4256 ( .A1(n3425), .A2(n3424), .ZN(n6093) );
  INV_X1 U4257 ( .A(n3429), .ZN(n3430) );
  NAND2_X1 U4258 ( .A1(n3428), .A2(n3430), .ZN(n4575) );
  NAND2_X1 U4259 ( .A1(n3431), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3435) );
  NOR3_X1 U4260 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6539), .A3(n6534), 
        .ZN(n6288) );
  NAND2_X1 U4261 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6288), .ZN(n6282) );
  NAND2_X1 U4262 ( .A1(n6397), .A2(n6282), .ZN(n3432) );
  NOR3_X1 U4263 ( .A1(n6397), .A2(n6539), .A3(n6534), .ZN(n4947) );
  NAND2_X1 U4264 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4947), .ZN(n4645) );
  NAND2_X1 U4265 ( .A1(n3432), .A2(n4645), .ZN(n4703) );
  OAI22_X1 U4266 ( .A1(n4337), .A2(n4703), .B1(n6553), .B2(n6397), .ZN(n3433)
         );
  INV_X1 U4267 ( .A(n3433), .ZN(n3434) );
  AOI22_X1 U4268 ( .A1(n4305), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4269 ( .A1(n3121), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4270 ( .A1(n4178), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4271 ( .A1(n4177), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3438) );
  NAND4_X1 U4272 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n3447)
         );
  AOI22_X1 U4273 ( .A1(n4317), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4274 ( .A1(n4284), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4275 ( .A1(n4314), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4276 ( .A1(n4316), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4277 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3446)
         );
  AOI22_X1 U4278 ( .A1(n3612), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3620), 
        .B2(n3473), .ZN(n3448) );
  NAND2_X1 U4279 ( .A1(n3933), .A2(n3537), .ZN(n3455) );
  NAND2_X1 U4280 ( .A1(n3451), .A2(n3450), .ZN(n3474) );
  INV_X1 U4281 ( .A(n3473), .ZN(n3452) );
  XNOR2_X1 U4282 ( .A(n3474), .B(n3452), .ZN(n3453) );
  NAND2_X1 U4283 ( .A1(n3453), .A2(n5319), .ZN(n3454) );
  INV_X1 U4284 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U4285 ( .A1(n6093), .A2(n6091), .ZN(n6092) );
  NAND2_X1 U4286 ( .A1(n3456), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3457)
         );
  NAND2_X1 U4287 ( .A1(n6092), .A2(n3457), .ZN(n4694) );
  INV_X1 U4288 ( .A(n3458), .ZN(n3459) );
  NAND2_X2 U4289 ( .A1(n3459), .A2(n4663), .ZN(n3502) );
  NAND2_X1 U4290 ( .A1(n3612), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4291 ( .A1(n4305), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4292 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4313), .B1(n3121), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4293 ( .A1(n4178), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4294 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4177), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3461) );
  NAND4_X1 U4295 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3470)
         );
  AOI22_X1 U4296 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4285), .B1(n4317), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4297 ( .A1(n4284), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4298 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4314), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4299 ( .A1(n4316), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4300 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3469)
         );
  NAND2_X1 U4301 ( .A1(n3620), .A2(n3525), .ZN(n3471) );
  NAND2_X1 U4302 ( .A1(n3472), .A2(n3471), .ZN(n3480) );
  NAND2_X1 U4303 ( .A1(n3896), .A2(n3537), .ZN(n3477) );
  NAND2_X1 U4304 ( .A1(n3474), .A2(n3473), .ZN(n3527) );
  XNOR2_X1 U4305 ( .A(n3527), .B(n3525), .ZN(n3475) );
  NAND2_X1 U4306 ( .A1(n3475), .A2(n5319), .ZN(n3476) );
  NAND2_X1 U4307 ( .A1(n3477), .A2(n3476), .ZN(n3478) );
  INV_X1 U4308 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6757) );
  XNOR2_X1 U4309 ( .A(n3478), .B(n6757), .ZN(n4691) );
  NAND2_X1 U4310 ( .A1(n4694), .A2(n4691), .ZN(n4692) );
  NAND2_X1 U4311 ( .A1(n3478), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3479)
         );
  NAND2_X1 U4312 ( .A1(n4692), .A2(n3479), .ZN(n6083) );
  INV_X1 U4313 ( .A(n3502), .ZN(n3481) );
  INV_X1 U4314 ( .A(n3480), .ZN(n3504) );
  NAND2_X1 U4315 ( .A1(n3481), .A2(n3480), .ZN(n3494) );
  NAND2_X1 U4316 ( .A1(n3612), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4317 ( .A1(n4305), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4318 ( .A1(n3121), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4319 ( .A1(n4178), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3483) );
  INV_X1 U4320 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U4321 ( .A1(n4177), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3482) );
  NAND4_X1 U4322 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(n3491)
         );
  AOI22_X1 U4323 ( .A1(n4317), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4324 ( .A1(n4284), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4325 ( .A1(n4314), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4326 ( .A1(n4316), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3486) );
  NAND4_X1 U4327 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3490)
         );
  NAND2_X1 U4328 ( .A1(n3620), .A2(n3524), .ZN(n3492) );
  NAND2_X1 U4329 ( .A1(n3493), .A2(n3492), .ZN(n3503) );
  NAND2_X1 U4330 ( .A1(n3944), .A2(n3537), .ZN(n3499) );
  INV_X1 U4331 ( .A(n3525), .ZN(n3495) );
  OR2_X1 U4332 ( .A1(n3527), .A2(n3495), .ZN(n3496) );
  XNOR2_X1 U4333 ( .A(n3496), .B(n3524), .ZN(n3497) );
  NAND2_X1 U4334 ( .A1(n3497), .A2(n5319), .ZN(n3498) );
  NAND2_X1 U4335 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  INV_X1 U4336 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U4337 ( .A(n3500), .B(n5077), .ZN(n6085) );
  NAND2_X1 U4338 ( .A1(n6083), .A2(n6085), .ZN(n6084) );
  NAND2_X1 U4339 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3501)
         );
  NAND2_X1 U4340 ( .A1(n6084), .A2(n3501), .ZN(n4815) );
  INV_X1 U4341 ( .A(n3503), .ZN(n3505) );
  AOI22_X1 U4342 ( .A1(n4305), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4343 ( .A1(n3121), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4344 ( .A1(n4178), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4345 ( .A1(n4177), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4346 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3516)
         );
  AOI22_X1 U4347 ( .A1(n4317), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4348 ( .A1(n4284), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4349 ( .A1(n4314), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4350 ( .A1(n4316), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4351 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3515)
         );
  INV_X1 U4352 ( .A(n3517), .ZN(n3523) );
  INV_X1 U4353 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3520) );
  INV_X1 U4354 ( .A(n3518), .ZN(n3519) );
  OAI21_X1 U4355 ( .B1(n3597), .B2(n3520), .A(n3519), .ZN(n3521) );
  INV_X1 U4356 ( .A(n3521), .ZN(n3522) );
  NAND2_X1 U4357 ( .A1(n3523), .A2(n3522), .ZN(n3952) );
  NAND3_X1 U4358 ( .A1(n3536), .A2(n3537), .A3(n3952), .ZN(n3530) );
  NAND2_X1 U4359 ( .A1(n3525), .A2(n3524), .ZN(n3526) );
  OR2_X1 U4360 ( .A1(n3527), .A2(n3526), .ZN(n3538) );
  XNOR2_X1 U4361 ( .A(n3538), .B(n3539), .ZN(n3528) );
  NAND2_X1 U4362 ( .A1(n3528), .A2(n5319), .ZN(n3529) );
  NAND2_X1 U4363 ( .A1(n3530), .A2(n3529), .ZN(n3531) );
  INV_X1 U4364 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U4365 ( .A(n3531), .B(n5078), .ZN(n4813) );
  NAND2_X1 U4366 ( .A1(n4815), .A2(n4813), .ZN(n4814) );
  NAND2_X1 U4367 ( .A1(n3531), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3532)
         );
  NAND2_X1 U4368 ( .A1(n4814), .A2(n3532), .ZN(n6075) );
  INV_X1 U4369 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4370 ( .A1(n3620), .A2(n3541), .ZN(n3533) );
  OAI21_X1 U4371 ( .B1(n3597), .B2(n3534), .A(n3533), .ZN(n3535) );
  NAND2_X1 U4372 ( .A1(n3826), .A2(n3537), .ZN(n3544) );
  INV_X1 U4373 ( .A(n3538), .ZN(n3540) );
  NAND2_X1 U4374 ( .A1(n3540), .A2(n3539), .ZN(n3549) );
  XNOR2_X1 U4375 ( .A(n3549), .B(n3541), .ZN(n3542) );
  NAND2_X1 U4376 ( .A1(n3542), .A2(n5319), .ZN(n3543) );
  NAND2_X1 U4377 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  INV_X1 U4378 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U4379 ( .A(n3545), .B(n6723), .ZN(n6077) );
  NAND2_X1 U4380 ( .A1(n6075), .A2(n6077), .ZN(n6076) );
  NAND2_X1 U4381 ( .A1(n3545), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3546)
         );
  NAND2_X1 U4382 ( .A1(n6076), .A2(n3546), .ZN(n4893) );
  NOR2_X1 U4383 ( .A1(n3602), .A2(n3548), .ZN(n3547) );
  OR3_X1 U4384 ( .A1(n3549), .A2(n3548), .A3(n3395), .ZN(n3550) );
  NAND2_X1 U4385 ( .A1(n3558), .A2(n3550), .ZN(n3551) );
  INV_X1 U4386 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U4387 ( .A(n3551), .B(n6135), .ZN(n4892) );
  NAND2_X1 U4388 ( .A1(n4893), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U4389 ( .A1(n3551), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3552)
         );
  NAND2_X1 U4390 ( .A1(n4891), .A2(n3552), .ZN(n5052) );
  INV_X1 U4391 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U4392 ( .A1(n5617), .A2(n5079), .ZN(n5053) );
  NAND2_X1 U4393 ( .A1(n5052), .A2(n5053), .ZN(n3553) );
  NAND2_X1 U4394 ( .A1(n3553), .A2(n5054), .ZN(n5071) );
  INV_X1 U4395 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3554) );
  NAND2_X1 U4396 ( .A1(n5603), .A2(n3554), .ZN(n5070) );
  NAND2_X1 U4397 ( .A1(n5071), .A2(n5070), .ZN(n5104) );
  INV_X1 U4398 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6117) );
  INV_X1 U4399 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U4400 ( .A1(n5617), .A2(n5197), .ZN(n5186) );
  OAI21_X1 U4401 ( .B1(n5184), .B2(n5188), .A(n5186), .ZN(n5245) );
  XNOR2_X1 U4402 ( .A(n5617), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5246)
         );
  NAND2_X1 U4403 ( .A1(n5245), .A2(n5246), .ZN(n3561) );
  INV_X1 U4404 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4405 ( .A1(n5603), .A2(n3559), .ZN(n3560) );
  NAND2_X1 U4406 ( .A1(n3561), .A2(n3560), .ZN(n5263) );
  INV_X1 U4407 ( .A(n5263), .ZN(n3563) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n7008) );
  INV_X1 U4409 ( .A(n5266), .ZN(n3562) );
  NAND2_X1 U4410 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  NAND2_X1 U4411 ( .A1(n3564), .A2(n5265), .ZN(n5286) );
  INV_X1 U4412 ( .A(n5286), .ZN(n3565) );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6760) );
  NAND2_X1 U4414 ( .A1(n3565), .A2(n3135), .ZN(n5599) );
  NAND2_X1 U4415 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3784) );
  AND2_X1 U4416 ( .A1(n5603), .A2(n3784), .ZN(n3566) );
  INV_X1 U4417 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3569) );
  AND2_X1 U4418 ( .A1(n5603), .A2(n3569), .ZN(n5602) );
  NOR2_X1 U4419 ( .A1(n3566), .A2(n5602), .ZN(n3567) );
  NAND2_X1 U4420 ( .A1(n5603), .A2(n6760), .ZN(n5600) );
  AND2_X1 U4421 ( .A1(n3567), .A2(n5600), .ZN(n3568) );
  NAND2_X1 U4422 ( .A1(n5599), .A2(n3568), .ZN(n5561) );
  INV_X1 U4423 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5690) );
  INV_X1 U4424 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5865) );
  AND3_X1 U4425 ( .A1(n5690), .A2(n3569), .A3(n5865), .ZN(n3570) );
  AND2_X1 U4426 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5697) );
  AND2_X1 U4427 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5674) );
  AND2_X1 U4428 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3815) );
  NAND3_X1 U4429 ( .A1(n5697), .A2(n5674), .A3(n3815), .ZN(n3572) );
  NAND2_X1 U4430 ( .A1(n5617), .A2(n3572), .ZN(n3575) );
  NOR2_X1 U4431 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5302) );
  NOR2_X1 U4432 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5698) );
  NOR2_X1 U4433 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5673) );
  AND3_X1 U4434 ( .A1(n5302), .A2(n5698), .A3(n5673), .ZN(n3573) );
  NOR2_X1 U4435 ( .A1(n5617), .A2(n3573), .ZN(n3574) );
  XNOR2_X1 U4436 ( .A(n3558), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5554)
         );
  AND2_X2 U4437 ( .A1(n5553), .A2(n5554), .ZN(n3577) );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6913) );
  NOR2_X2 U4439 ( .A1(n3577), .A2(n3576), .ZN(n5329) );
  INV_X1 U4440 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5530) );
  NOR2_X1 U4441 ( .A1(n5296), .A2(n5530), .ZN(n5546) );
  AND2_X1 U4442 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U4443 ( .A1(n5628), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3801) );
  NOR2_X1 U4444 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3578)
         );
  AND2_X1 U4445 ( .A1(n3577), .A2(n3578), .ZN(n5531) );
  NOR4_X1 U4446 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4447 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n5531), .B2(n3579), .ZN(n3580) );
  XNOR2_X1 U4448 ( .A(n3580), .B(n3818), .ZN(n3823) );
  XNOR2_X1 U4449 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3593) );
  XOR2_X1 U4450 ( .A(n3593), .B(n3594), .Z(n3641) );
  INV_X1 U4451 ( .A(n3620), .ZN(n3581) );
  OAI21_X1 U4452 ( .B1(n3581), .B2(n3631), .A(n4615), .ZN(n3590) );
  INV_X1 U4453 ( .A(n3594), .ZN(n3583) );
  INV_X1 U4454 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3917) );
  NAND2_X1 U4455 ( .A1(n3917), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4456 ( .A1(n3583), .A2(n3582), .ZN(n3586) );
  INV_X1 U4457 ( .A(n3586), .ZN(n3584) );
  NAND2_X1 U4458 ( .A1(n3620), .A2(n3584), .ZN(n3588) );
  OAI21_X1 U4459 ( .B1(n3656), .B2(n3586), .A(n3585), .ZN(n3587) );
  OAI21_X1 U4460 ( .B1(n3290), .B2(n4615), .A(n3631), .ZN(n3603) );
  AOI22_X1 U4461 ( .A1(n3624), .A2(n3588), .B1(n3587), .B2(n3603), .ZN(n3589)
         );
  OAI21_X1 U4462 ( .B1(n3590), .B2(n3641), .A(n3589), .ZN(n3592) );
  NAND3_X1 U4463 ( .A1(n3590), .A2(STATE2_REG_0__SCAN_IN), .A3(n3641), .ZN(
        n3591) );
  OAI211_X1 U4464 ( .C1(n3641), .C2(n3624), .A(n3592), .B(n3591), .ZN(n3607)
         );
  XNOR2_X1 U4465 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4466 ( .A1(n3594), .A2(n3593), .ZN(n3596) );
  NAND2_X1 U4467 ( .A1(n6534), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3595) );
  NAND2_X1 U4468 ( .A1(n3596), .A2(n3595), .ZN(n3599) );
  XOR2_X1 U4469 ( .A(n3598), .B(n3599), .Z(n3642) );
  NAND2_X1 U4470 ( .A1(n3620), .A2(n3642), .ZN(n3604) );
  OAI211_X1 U4471 ( .C1(n3597), .C2(n3642), .A(n3604), .B(n3603), .ZN(n3606)
         );
  XNOR2_X1 U4472 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3608) );
  NAND2_X1 U4473 ( .A1(n3599), .A2(n3598), .ZN(n3601) );
  NAND2_X1 U4474 ( .A1(n6539), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4475 ( .A1(n3601), .A2(n3600), .ZN(n3609) );
  XOR2_X1 U4476 ( .A(n3608), .B(n3609), .Z(n3640) );
  OAI22_X1 U4477 ( .A1(n3604), .A2(n3603), .B1(n3640), .B2(n3602), .ZN(n3605)
         );
  AOI21_X1 U4478 ( .B1(n3607), .B2(n3606), .A(n3605), .ZN(n3614) );
  NAND2_X1 U4479 ( .A1(n3609), .A2(n3608), .ZN(n3611) );
  NAND2_X1 U4480 ( .A1(n6397), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4481 ( .A1(n3611), .A2(n3610), .ZN(n3617) );
  INV_X1 U4482 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U4483 ( .A1(n4577), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3618) );
  OR2_X1 U4484 ( .A1(n3617), .A2(n3618), .ZN(n3645) );
  AOI21_X1 U4485 ( .B1(n3640), .B2(n3645), .A(n3612), .ZN(n3613) );
  OAI22_X1 U4486 ( .A1(n3614), .A2(n3613), .B1(n3624), .B2(n3645), .ZN(n3615)
         );
  AOI21_X1 U4487 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6972), .A(n3615), 
        .ZN(n3622) );
  INV_X1 U4488 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6983) );
  AND2_X1 U4489 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6983), .ZN(n3616)
         );
  NAND2_X1 U4490 ( .A1(n3620), .A2(n3644), .ZN(n3621) );
  NAND2_X1 U4491 ( .A1(n3622), .A2(n3621), .ZN(n3626) );
  INV_X1 U4492 ( .A(n3644), .ZN(n3623) );
  AND2_X1 U4493 ( .A1(n6553), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6566) );
  INV_X1 U4494 ( .A(n6566), .ZN(n5917) );
  INV_X1 U4495 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U4496 ( .A1(n3627), .A2(n6588), .ZN(n6583) );
  NAND2_X1 U4497 ( .A1(n3631), .A2(n6583), .ZN(n5123) );
  INV_X1 U4498 ( .A(READY_N), .ZN(n6892) );
  NAND3_X1 U4499 ( .A1(n4370), .A2(n5123), .A3(n6892), .ZN(n3628) );
  NAND3_X1 U4500 ( .A1(n3628), .A2(n5122), .A3(n5097), .ZN(n3629) );
  NAND2_X1 U4501 ( .A1(n3629), .A2(n3788), .ZN(n3653) );
  NAND2_X1 U4502 ( .A1(n4643), .A2(n5098), .ZN(n3630) );
  OR2_X1 U4503 ( .A1(n4493), .A2(n3630), .ZN(n6525) );
  NOR2_X1 U4504 ( .A1(n6525), .A2(n3631), .ZN(n3793) );
  NAND2_X1 U4505 ( .A1(n4419), .A2(n3793), .ZN(n3650) );
  INV_X1 U4506 ( .A(n3632), .ZN(n4353) );
  NAND2_X1 U4507 ( .A1(n3633), .A2(n5122), .ZN(n3634) );
  MUX2_X1 U4508 ( .A(n3395), .B(n3634), .S(n4493), .Z(n3791) );
  AOI21_X1 U4509 ( .B1(n6525), .B2(n3290), .A(n3636), .ZN(n3637) );
  AND2_X1 U4510 ( .A1(n3638), .A2(n3637), .ZN(n3657) );
  NAND2_X1 U4511 ( .A1(n3791), .A2(n3657), .ZN(n3639) );
  NAND2_X1 U4512 ( .A1(n4353), .A2(n3639), .ZN(n4388) );
  NAND2_X1 U4513 ( .A1(n4605), .A2(n6583), .ZN(n3648) );
  AND3_X1 U4514 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(n3643) );
  OR2_X1 U4515 ( .A1(n3644), .A2(n3643), .ZN(n3646) );
  NAND2_X1 U4516 ( .A1(n3646), .A2(n3645), .ZN(n4352) );
  INV_X1 U4517 ( .A(n4352), .ZN(n3647) );
  NOR2_X1 U4518 ( .A1(READY_N), .A2(n3647), .ZN(n4485) );
  NAND3_X1 U4519 ( .A1(n3648), .A2(n4485), .A3(n4621), .ZN(n3649) );
  NAND3_X1 U4520 ( .A1(n3650), .A2(n4388), .A3(n3649), .ZN(n3651) );
  NAND2_X1 U4521 ( .A1(n3651), .A2(n6566), .ZN(n3652) );
  AOI22_X1 U4522 ( .A1(n4370), .A2(n4428), .B1(n3781), .B2(n4643), .ZN(n3659)
         );
  AND2_X1 U4523 ( .A1(n3657), .A2(n5171), .ZN(n4490) );
  INV_X1 U4524 ( .A(n4490), .ZN(n3658) );
  AND2_X1 U4525 ( .A1(n3657), .A2(n3656), .ZN(n4351) );
  INV_X1 U4526 ( .A(n4351), .ZN(n6545) );
  NAND4_X1 U4527 ( .A1(n5910), .A2(n3659), .A3(n3658), .A4(n6545), .ZN(n3660)
         );
  NAND2_X1 U4528 ( .A1(n3806), .A2(n3660), .ZN(n5881) );
  INV_X2 U4529 ( .A(n3661), .ZN(n5223) );
  INV_X1 U4530 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3662) );
  NAND2_X1 U4531 ( .A1(n3671), .A2(n3662), .ZN(n3667) );
  OR2_X2 U4532 ( .A1(n3663), .A2(n3290), .ZN(n3766) );
  NAND2_X1 U4533 ( .A1(n3661), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3664)
         );
  OAI211_X1 U4534 ( .C1(n3665), .C2(EBX_REG_1__SCAN_IN), .A(n3766), .B(n3664), 
        .ZN(n3666) );
  NAND2_X1 U4535 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  INV_X1 U4536 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5212) );
  OAI22_X1 U4537 ( .A1(n3766), .A2(n5212), .B1(n3661), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4479) );
  XNOR2_X1 U4538 ( .A(n3668), .B(n4479), .ZN(n4427) );
  NAND2_X1 U4539 ( .A1(n4427), .A2(n4428), .ZN(n3670) );
  INV_X1 U4540 ( .A(n3668), .ZN(n3669) );
  INV_X1 U4541 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6986) );
  NAND2_X1 U4542 ( .A1(n3755), .A2(n6986), .ZN(n3675) );
  INV_X1 U4543 ( .A(n4428), .ZN(n3673) );
  INV_X2 U4544 ( .A(n5223), .ZN(n5340) );
  NAND2_X1 U4545 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3672)
         );
  OAI211_X1 U4546 ( .C1(n3673), .C2(EBX_REG_2__SCAN_IN), .A(n3766), .B(n3672), 
        .ZN(n3674) );
  NAND2_X1 U4547 ( .A1(n3675), .A2(n3674), .ZN(n4474) );
  INV_X1 U4548 ( .A(EBX_REG_3__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4549 ( .A1(n5223), .A2(n3678), .ZN(n3681) );
  NAND2_X1 U4550 ( .A1(n3766), .A2(n6167), .ZN(n3679) );
  OAI211_X1 U4551 ( .C1(n3673), .C2(EBX_REG_3__SCAN_IN), .A(n3679), .B(n5340), 
        .ZN(n3680) );
  INV_X1 U4552 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U4553 ( .A1(n3755), .A2(n3684), .ZN(n3687) );
  NAND2_X1 U4554 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3685)
         );
  OAI211_X1 U4555 ( .C1(n4424), .C2(EBX_REG_4__SCAN_IN), .A(n3766), .B(n3685), 
        .ZN(n3686) );
  NAND2_X1 U4556 ( .A1(n3687), .A2(n3686), .ZN(n4499) );
  NAND2_X1 U4557 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3689)
         );
  NOR2_X1 U4558 ( .A1(n4424), .A2(EBX_REG_5__SCAN_IN), .ZN(n3688) );
  MUX2_X1 U4559 ( .A(n3689), .B(n5164), .S(n3688), .Z(n3692) );
  NAND2_X1 U4560 ( .A1(n3759), .A2(n4424), .ZN(n3731) );
  NAND2_X1 U4561 ( .A1(n3759), .A2(EBX_REG_5__SCAN_IN), .ZN(n3690) );
  AND2_X1 U4562 ( .A1(n3731), .A2(n3690), .ZN(n3691) );
  NAND2_X1 U4563 ( .A1(n3692), .A2(n3691), .ZN(n4651) );
  NAND2_X1 U4564 ( .A1(n4652), .A2(n4651), .ZN(n4671) );
  INV_X1 U4565 ( .A(n3755), .ZN(n3764) );
  MUX2_X1 U4566 ( .A(n3764), .B(n5340), .S(EBX_REG_6__SCAN_IN), .Z(n3693) );
  NAND2_X1 U4567 ( .A1(n3693), .A2(n3131), .ZN(n4670) );
  OR2_X2 U4568 ( .A1(n4671), .A2(n4670), .ZN(n4801) );
  NAND2_X1 U4569 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3695)
         );
  NOR2_X1 U4570 ( .A1(n4424), .A2(EBX_REG_7__SCAN_IN), .ZN(n3694) );
  MUX2_X1 U4571 ( .A(n3695), .B(n5340), .S(n3694), .Z(n3698) );
  NAND2_X1 U4572 ( .A1(n3759), .A2(EBX_REG_7__SCAN_IN), .ZN(n3696) );
  AND2_X1 U4573 ( .A1(n3731), .A2(n3696), .ZN(n3697) );
  NAND2_X1 U4574 ( .A1(n3698), .A2(n3697), .ZN(n4803) );
  INV_X1 U4575 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U4576 ( .A1(n3755), .A2(n5450), .ZN(n3701) );
  NAND2_X1 U4577 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3699)
         );
  OAI211_X1 U4578 ( .C1(n4424), .C2(EBX_REG_8__SCAN_IN), .A(n3766), .B(n3699), 
        .ZN(n3700) );
  AND2_X1 U4579 ( .A1(n3701), .A2(n3700), .ZN(n4802) );
  NAND2_X1 U4580 ( .A1(n4803), .A2(n4802), .ZN(n3702) );
  NOR2_X4 U4581 ( .A1(n4801), .A2(n3702), .ZN(n5046) );
  NAND2_X1 U4582 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3704)
         );
  NOR2_X1 U4583 ( .A1(n4424), .A2(EBX_REG_9__SCAN_IN), .ZN(n3703) );
  MUX2_X1 U4584 ( .A(n3704), .B(n5164), .S(n3703), .Z(n3707) );
  NAND2_X1 U4585 ( .A1(n3759), .A2(EBX_REG_9__SCAN_IN), .ZN(n3705) );
  AND2_X1 U4586 ( .A1(n3731), .A2(n3705), .ZN(n3706) );
  MUX2_X1 U4587 ( .A(n3764), .B(n5164), .S(EBX_REG_10__SCAN_IN), .Z(n3708) );
  NAND2_X1 U4588 ( .A1(n3708), .A2(n3134), .ZN(n5043) );
  NOR2_X1 U4589 ( .A1(n5042), .A2(n5043), .ZN(n3709) );
  INV_X1 U4590 ( .A(EBX_REG_11__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4591 ( .A1(n5223), .A2(n3710), .ZN(n3713) );
  NAND2_X1 U4592 ( .A1(n3766), .A2(n6117), .ZN(n3711) );
  OAI211_X1 U4593 ( .C1(n4424), .C2(EBX_REG_11__SCAN_IN), .A(n3711), .B(n5164), 
        .ZN(n3712) );
  NAND2_X1 U4594 ( .A1(n3713), .A2(n3712), .ZN(n4779) );
  MUX2_X1 U4595 ( .A(n3764), .B(n5340), .S(EBX_REG_12__SCAN_IN), .Z(n3714) );
  NAND2_X1 U4596 ( .A1(n3714), .A2(n3138), .ZN(n4793) );
  NAND2_X1 U4597 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3716) );
  NOR2_X1 U4598 ( .A1(n4424), .A2(EBX_REG_13__SCAN_IN), .ZN(n3715) );
  MUX2_X1 U4599 ( .A(n3716), .B(n5164), .S(n3715), .Z(n3718) );
  NAND2_X1 U4600 ( .A1(n3759), .A2(EBX_REG_13__SCAN_IN), .ZN(n3717) );
  AND3_X1 U4601 ( .A1(n3718), .A2(n3731), .A3(n3717), .ZN(n4853) );
  INV_X1 U4602 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U4603 ( .A1(n3755), .A2(n6803), .ZN(n3721) );
  NAND2_X1 U4604 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3719) );
  OAI211_X1 U4605 ( .C1(n4424), .C2(EBX_REG_14__SCAN_IN), .A(n3766), .B(n3719), 
        .ZN(n3720) );
  AND2_X1 U4606 ( .A1(n3721), .A2(n3720), .ZN(n4809) );
  NAND2_X1 U4607 ( .A1(n4478), .A2(EBX_REG_15__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4608 ( .A1(n4424), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4609 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  XNOR2_X1 U4610 ( .A(n3724), .B(n5223), .ZN(n4998) );
  MUX2_X1 U4611 ( .A(n3764), .B(n5164), .S(EBX_REG_16__SCAN_IN), .Z(n3726) );
  INV_X1 U4612 ( .A(n4478), .ZN(n3770) );
  NAND2_X1 U4613 ( .A1(n3770), .A2(n3569), .ZN(n3725) );
  NAND2_X1 U4614 ( .A1(n3726), .A2(n3725), .ZN(n5063) );
  NOR2_X1 U4615 ( .A1(n4998), .A2(n5063), .ZN(n3727) );
  NAND2_X1 U4616 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3729) );
  NOR2_X1 U4617 ( .A1(n4424), .A2(EBX_REG_17__SCAN_IN), .ZN(n3728) );
  MUX2_X1 U4618 ( .A(n3729), .B(n5164), .S(n3728), .Z(n3732) );
  NAND2_X1 U4619 ( .A1(n3759), .A2(EBX_REG_17__SCAN_IN), .ZN(n3730) );
  AND3_X1 U4620 ( .A1(n3732), .A2(n3731), .A3(n3730), .ZN(n5095) );
  OR2_X2 U4621 ( .A1(n5094), .A2(n5095), .ZN(n5167) );
  INV_X1 U4622 ( .A(EBX_REG_19__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4623 ( .A1(n3755), .A2(n3733), .ZN(n3736) );
  NAND2_X1 U4624 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3734) );
  OAI211_X1 U4625 ( .C1(n4424), .C2(EBX_REG_19__SCAN_IN), .A(n3766), .B(n3734), 
        .ZN(n3735) );
  NAND2_X1 U4626 ( .A1(n3736), .A2(n3735), .ZN(n5208) );
  OR2_X2 U4627 ( .A1(n5167), .A2(n5208), .ZN(n5222) );
  NAND2_X1 U4628 ( .A1(n4478), .A2(EBX_REG_18__SCAN_IN), .ZN(n3738) );
  NAND2_X1 U4629 ( .A1(n4424), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3737) );
  AND2_X1 U4630 ( .A1(n3738), .A2(n3737), .ZN(n5165) );
  INV_X1 U4631 ( .A(n5165), .ZN(n5224) );
  OAI22_X1 U4632 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4424), .ZN(n5225) );
  MUX2_X1 U4633 ( .A(n5340), .B(n5165), .S(n5225), .Z(n3739) );
  OAI21_X1 U4634 ( .B1(n5223), .B2(n5224), .A(n3739), .ZN(n3740) );
  NOR2_X2 U4635 ( .A1(n5222), .A2(n3740), .ZN(n5282) );
  INV_X1 U4636 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U4637 ( .A1(n3755), .A2(n5402), .ZN(n3743) );
  NAND2_X1 U4638 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3741) );
  OAI211_X1 U4639 ( .C1(n4424), .C2(EBX_REG_21__SCAN_IN), .A(n3766), .B(n3741), 
        .ZN(n3742) );
  AND2_X1 U4640 ( .A1(n3743), .A2(n3742), .ZN(n5281) );
  NAND2_X1 U4641 ( .A1(n5282), .A2(n5281), .ZN(n5278) );
  NAND2_X1 U4642 ( .A1(n3759), .A2(EBX_REG_22__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4643 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3745) );
  NOR2_X1 U4644 ( .A1(n4424), .A2(EBX_REG_22__SCAN_IN), .ZN(n3744) );
  MUX2_X1 U4645 ( .A(n3745), .B(n5164), .S(n3744), .Z(n3746) );
  AND2_X1 U4646 ( .A1(n3747), .A2(n3746), .ZN(n5279) );
  OR2_X2 U4647 ( .A1(n5278), .A2(n5279), .ZN(n5394) );
  INV_X1 U4648 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U4649 ( .A1(n3755), .A2(n6956), .ZN(n3750) );
  NAND2_X1 U4650 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3748) );
  OAI211_X1 U4651 ( .C1(n4424), .C2(EBX_REG_23__SCAN_IN), .A(n3766), .B(n3748), 
        .ZN(n3749) );
  NAND2_X1 U4652 ( .A1(n3750), .A2(n3749), .ZN(n5395) );
  INV_X1 U4653 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U4654 ( .A1(n5223), .A2(n5506), .ZN(n3754) );
  INV_X1 U4655 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3751) );
  NAND2_X1 U4656 ( .A1(n3766), .A2(n3751), .ZN(n3752) );
  OAI211_X1 U4657 ( .C1(n4424), .C2(EBX_REG_24__SCAN_IN), .A(n3752), .B(n5164), 
        .ZN(n3753) );
  NAND2_X1 U4658 ( .A1(n3754), .A2(n3753), .ZN(n5299) );
  INV_X1 U4659 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U4660 ( .A1(n3755), .A2(n5807), .ZN(n3758) );
  NAND2_X1 U4661 ( .A1(n5164), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3756) );
  OAI211_X1 U4662 ( .C1(n4424), .C2(EBX_REG_25__SCAN_IN), .A(n3766), .B(n3756), 
        .ZN(n3757) );
  AND2_X1 U4663 ( .A1(n3758), .A2(n3757), .ZN(n5501) );
  NAND2_X1 U4664 ( .A1(n3759), .A2(EBX_REG_26__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4665 ( .A1(n5340), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3761) );
  NOR2_X1 U4666 ( .A1(n3673), .A2(EBX_REG_26__SCAN_IN), .ZN(n3760) );
  MUX2_X1 U4667 ( .A(n3761), .B(n5340), .S(n3760), .Z(n3762) );
  AND2_X1 U4668 ( .A1(n3763), .A2(n3762), .ZN(n5493) );
  MUX2_X1 U4669 ( .A(n3764), .B(n5164), .S(EBX_REG_27__SCAN_IN), .Z(n3765) );
  NAND2_X1 U4670 ( .A1(n3765), .A2(n3125), .ZN(n5481) );
  INV_X1 U4671 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6748) );
  NAND2_X1 U4672 ( .A1(n5223), .A2(n6748), .ZN(n3769) );
  INV_X1 U4673 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U4674 ( .A1(n3766), .A2(n5533), .ZN(n3767) );
  OAI211_X1 U4675 ( .C1(n4424), .C2(EBX_REG_28__SCAN_IN), .A(n3767), .B(n5164), 
        .ZN(n3768) );
  NAND2_X1 U4676 ( .A1(n3769), .A2(n3768), .ZN(n5476) );
  INV_X1 U4677 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5627) );
  INV_X1 U4678 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U4679 ( .A1(n3770), .A2(n5627), .B1(n4428), .B2(n6895), .ZN(n3771)
         );
  NAND2_X1 U4680 ( .A1(n5478), .A2(n3771), .ZN(n5339) );
  INV_X1 U4681 ( .A(n3771), .ZN(n3772) );
  MUX2_X1 U4682 ( .A(EBX_REG_29__SCAN_IN), .B(n3772), .S(n5340), .Z(n5369) );
  NAND2_X1 U4683 ( .A1(n4478), .A2(EBX_REG_30__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U4684 ( .A1(n3673), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4685 ( .A1(n3774), .A2(n3773), .ZN(n5337) );
  NOR2_X1 U4686 ( .A1(n5369), .A2(n5337), .ZN(n3775) );
  AND2_X1 U4687 ( .A1(n5478), .A2(n3775), .ZN(n3776) );
  OAI22_X1 U4688 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4424), .ZN(n3777) );
  INV_X1 U4689 ( .A(n3777), .ZN(n3778) );
  NAND2_X1 U4690 ( .A1(n4370), .A2(n5319), .ZN(n6555) );
  NAND2_X1 U4691 ( .A1(n3781), .A2(n3780), .ZN(n3782) );
  NAND2_X1 U4692 ( .A1(n6555), .A2(n3782), .ZN(n3783) );
  NAND2_X1 U4693 ( .A1(n3806), .A2(n3783), .ZN(n6195) );
  NOR2_X1 U4694 ( .A1(n4337), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U4695 ( .A1(n6178), .A2(REIP_REG_31__SCAN_IN), .ZN(n4346) );
  INV_X1 U4696 ( .A(n5697), .ZN(n3800) );
  INV_X1 U4697 ( .A(n3784), .ZN(n3804) );
  NOR2_X1 U4698 ( .A1(n5197), .A2(n6117), .ZN(n5252) );
  INV_X1 U4699 ( .A(n5252), .ZN(n5257) );
  NOR2_X1 U4700 ( .A1(n3559), .A2(n5257), .ZN(n5254) );
  AND2_X1 U4701 ( .A1(n3632), .A2(n4605), .ZN(n6529) );
  NAND2_X1 U4702 ( .A1(n3806), .A2(n6529), .ZN(n5253) );
  NAND4_X1 U4703 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U4704 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3785) );
  OR2_X1 U4705 ( .A1(n6161), .A2(n3785), .ZN(n5075) );
  NOR2_X1 U4706 ( .A1(n6135), .A2(n6723), .ZN(n6130) );
  NAND2_X1 U4707 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5080) );
  INV_X1 U4708 ( .A(n5080), .ZN(n3786) );
  NAND2_X1 U4709 ( .A1(n6130), .A2(n3786), .ZN(n3796) );
  NOR2_X1 U4710 ( .A1(n5075), .A2(n3796), .ZN(n5195) );
  INV_X1 U4711 ( .A(n5195), .ZN(n3798) );
  INV_X1 U4712 ( .A(n5097), .ZN(n3897) );
  NAND2_X1 U4713 ( .A1(n4478), .A2(n3636), .ZN(n3787) );
  OR2_X1 U4714 ( .A1(n5176), .A2(n4621), .ZN(n4387) );
  OAI211_X1 U4715 ( .C1(n3788), .C2(n3897), .A(n3787), .B(n4387), .ZN(n3789)
         );
  AOI21_X1 U4716 ( .B1(n3635), .B2(n5223), .A(n3789), .ZN(n3790) );
  AND3_X1 U4717 ( .A1(n3792), .A2(n3791), .A3(n3790), .ZN(n4372) );
  NAND2_X1 U4718 ( .A1(n4372), .A2(n4557), .ZN(n3795) );
  NAND2_X1 U4719 ( .A1(n3806), .A2(n3795), .ZN(n3805) );
  NOR2_X1 U4720 ( .A1(n3798), .A2(n3805), .ZN(n3797) );
  INV_X1 U4721 ( .A(n3793), .ZN(n3794) );
  NAND2_X1 U4722 ( .A1(n3806), .A2(n4417), .ZN(n6187) );
  NAND2_X1 U4723 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U4724 ( .A1(n3422), .A2(n6188), .ZN(n6189) );
  NAND3_X1 U4725 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6189), .ZN(n5076) );
  NOR2_X1 U4726 ( .A1(n6187), .A2(n5076), .ZN(n6158) );
  NAND3_X1 U4727 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6158), .ZN(n5074) );
  NOR2_X1 U4728 ( .A1(n3796), .A2(n5074), .ZN(n5194) );
  AOI21_X1 U4729 ( .B1(n3797), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5194), 
        .ZN(n5903) );
  OAI21_X1 U4730 ( .B1(n5253), .B2(n3798), .A(n5903), .ZN(n5196) );
  NAND2_X1 U4731 ( .A1(n5254), .A2(n5196), .ZN(n5908) );
  NAND3_X1 U4732 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5892), .ZN(n5876) );
  INV_X1 U4733 ( .A(n5876), .ZN(n3799) );
  NAND2_X1 U4734 ( .A1(n3804), .A2(n3799), .ZN(n5863) );
  INV_X1 U4735 ( .A(n5674), .ZN(n3813) );
  AND2_X1 U4736 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3803) );
  INV_X1 U4737 ( .A(n3801), .ZN(n5344) );
  NAND4_X1 U4738 ( .A1(n5644), .A2(n5344), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n3818), .ZN(n3802) );
  OAI211_X1 U4739 ( .C1(n5328), .C2(n6195), .A(n4346), .B(n3802), .ZN(n3821)
         );
  NAND2_X1 U4740 ( .A1(n5693), .A2(n6187), .ZN(n5878) );
  INV_X1 U4741 ( .A(n5878), .ZN(n6151) );
  INV_X1 U4742 ( .A(n3803), .ZN(n5651) );
  NAND2_X1 U4743 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U4744 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5254), .ZN(n5877) );
  NOR2_X1 U4745 ( .A1(n5885), .A2(n5877), .ZN(n3807) );
  NAND2_X1 U4746 ( .A1(n5194), .A2(n3807), .ZN(n5689) );
  NAND2_X1 U4747 ( .A1(n3804), .A2(n5697), .ZN(n3808) );
  INV_X1 U4748 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U4749 ( .A1(n6187), .A2(n3805), .ZN(n5256) );
  AND2_X1 U4750 ( .A1(n4406), .A2(n5256), .ZN(n5704) );
  NOR2_X1 U4751 ( .A1(n3806), .A2(n6178), .ZN(n5709) );
  NOR2_X1 U4752 ( .A1(n5704), .A2(n5709), .ZN(n6146) );
  NAND2_X1 U4753 ( .A1(n6187), .A2(n6146), .ZN(n5688) );
  OAI21_X1 U4754 ( .B1(n5689), .B2(n3808), .A(n5688), .ZN(n3812) );
  AND2_X1 U4755 ( .A1(n5195), .A2(n3807), .ZN(n5692) );
  INV_X1 U4756 ( .A(n3808), .ZN(n3809) );
  AND2_X1 U4757 ( .A1(n5692), .A2(n3809), .ZN(n3810) );
  OR2_X1 U4758 ( .A1(n5693), .A2(n3810), .ZN(n3811) );
  NAND2_X1 U4759 ( .A1(n3812), .A2(n3811), .ZN(n5685) );
  AND2_X1 U4760 ( .A1(n5878), .A2(n3813), .ZN(n3814) );
  OR2_X1 U4761 ( .A1(n5685), .A2(n3814), .ZN(n5670) );
  INV_X1 U4762 ( .A(n5253), .ZN(n5710) );
  NOR2_X1 U4763 ( .A1(n5710), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4465)
         );
  NOR2_X1 U4764 ( .A1(n5693), .A2(n4465), .ZN(n6186) );
  INV_X1 U4765 ( .A(n6186), .ZN(n6160) );
  AOI21_X1 U4766 ( .B1(n6187), .B2(n6160), .A(n3815), .ZN(n3816) );
  AOI21_X1 U4767 ( .B1(n5878), .B2(n5651), .A(n5661), .ZN(n5636) );
  OAI21_X1 U4768 ( .B1(n5628), .B2(n6151), .A(n5636), .ZN(n5633) );
  AOI21_X1 U4769 ( .B1(n5627), .B2(n5878), .A(n5633), .ZN(n5333) );
  OAI21_X1 U4770 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6151), .A(n5333), 
        .ZN(n3817) );
  INV_X1 U4771 ( .A(n3823), .ZN(n3825) );
  INV_X1 U4772 ( .A(n5924), .ZN(n3824) );
  NAND2_X1 U4773 ( .A1(n3825), .A2(n3824), .ZN(n4349) );
  INV_X2 U4774 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6568) );
  NOR2_X2 U4775 ( .A1(n4626), .A2(n6568), .ZN(n4018) );
  NAND2_X1 U4776 ( .A1(n3826), .A2(n4018), .ZN(n3832) );
  OR2_X1 U4777 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4333) );
  OAI21_X1 U4778 ( .B1(n3827), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3878), 
        .ZN(n6082) );
  INV_X1 U4779 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4780 ( .A1(n6568), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4038) );
  INV_X1 U4781 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3828) );
  OAI22_X1 U4782 ( .A1(n4228), .A2(n3829), .B1(n4038), .B2(n3828), .ZN(n3830)
         );
  AOI21_X1 U4783 ( .B1(n4299), .B2(n6082), .A(n3830), .ZN(n3831) );
  AOI22_X1 U4784 ( .A1(n4305), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4785 ( .A1(n4284), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4786 ( .A1(n4307), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4787 ( .A1(n4178), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4788 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AOI22_X1 U4789 ( .A1(n3121), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4790 ( .A1(n4317), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4315), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4791 ( .A1(n4260), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4792 ( .A1(n4316), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4793 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4794 ( .A1(n3842), .A2(n3841), .ZN(n3846) );
  INV_X1 U4795 ( .A(n4018), .ZN(n3845) );
  XNOR2_X1 U4796 ( .A(n3962), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5140)
         );
  NAND2_X1 U4797 ( .A1(n5140), .A2(n4299), .ZN(n3844) );
  INV_X2 U4798 ( .A(n4228), .ZN(n4335) );
  INV_X1 U4799 ( .A(n4038), .ZN(n4334) );
  AOI22_X1 U4800 ( .A1(n4335), .A2(EAX_REG_11__SCAN_IN), .B1(n4334), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3843) );
  OAI211_X1 U4801 ( .C1(n3846), .C2(n3845), .A(n3844), .B(n3843), .ZN(n4776)
         );
  XOR2_X1 U4802 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3847), .Z(n5965) );
  INV_X1 U4803 ( .A(n5965), .ZN(n3862) );
  INV_X1 U4804 ( .A(n4333), .ZN(n4299) );
  AOI22_X1 U4805 ( .A1(n4178), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4806 ( .A1(n4177), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4807 ( .A1(n4305), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4808 ( .A1(n4316), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4809 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AOI22_X1 U4810 ( .A1(n4317), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4811 ( .A1(n4313), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4812 ( .A1(n4284), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4813 ( .A1(n4307), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4814 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  OAI21_X1 U4815 ( .B1(n3857), .B2(n3856), .A(n4018), .ZN(n3860) );
  NAND2_X1 U4816 ( .A1(n4335), .A2(EAX_REG_10__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4817 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3858)
         );
  NAND3_X1 U4818 ( .A1(n3860), .A2(n3859), .A3(n3858), .ZN(n3861) );
  AOI21_X1 U4819 ( .B1(n3862), .B2(n4299), .A(n3861), .ZN(n5041) );
  XNOR2_X1 U4820 ( .A(n3877), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5119) );
  AOI22_X1 U4821 ( .A1(n3121), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4822 ( .A1(n4305), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4823 ( .A1(n4314), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4824 ( .A1(n4285), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4825 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3872)
         );
  AOI22_X1 U4826 ( .A1(n4313), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4827 ( .A1(n4178), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4828 ( .A1(n4284), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4829 ( .A1(n4317), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4830 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  OAI21_X1 U4831 ( .B1(n3872), .B2(n3871), .A(n4018), .ZN(n3875) );
  NAND2_X1 U4832 ( .A1(n4335), .A2(EAX_REG_9__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4833 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3873)
         );
  NAND3_X1 U4834 ( .A1(n3875), .A2(n3874), .A3(n3873), .ZN(n3876) );
  AOI21_X1 U4835 ( .B1(n5119), .B2(n4299), .A(n3876), .ZN(n4899) );
  OR2_X1 U4836 ( .A1(n5041), .A2(n4899), .ZN(n3894) );
  AOI21_X1 U4837 ( .B1(n6794), .B2(n3878), .A(n3877), .ZN(n4894) );
  OR2_X1 U4838 ( .A1(n4894), .A2(n4333), .ZN(n3893) );
  AOI22_X1 U4839 ( .A1(n4178), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4840 ( .A1(n3121), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4841 ( .A1(n4284), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4842 ( .A1(n4317), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4843 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3888)
         );
  AOI22_X1 U4844 ( .A1(n3120), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4845 ( .A1(n4313), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4846 ( .A1(n4314), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4847 ( .A1(n4285), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4848 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3887)
         );
  OAI21_X1 U4849 ( .B1(n3888), .B2(n3887), .A(n4018), .ZN(n3891) );
  NAND2_X1 U4850 ( .A1(n4335), .A2(EAX_REG_8__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4851 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3889)
         );
  AND3_X1 U4852 ( .A1(n3891), .A2(n3890), .A3(n3889), .ZN(n3892) );
  AND2_X1 U4853 ( .A1(n3893), .A2(n3892), .ZN(n4799) );
  NOR2_X1 U4854 ( .A1(n3894), .A2(n4799), .ZN(n4772) );
  AND2_X1 U4855 ( .A1(n4776), .A2(n4772), .ZN(n3895) );
  NAND2_X1 U4856 ( .A1(n3896), .A2(n4018), .ZN(n3904) );
  NAND2_X1 U4857 ( .A1(n3897), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3940) );
  INV_X1 U4858 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6353) );
  OAI21_X1 U4859 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6353), .A(n6568), 
        .ZN(n3899) );
  NAND2_X1 U4860 ( .A1(n4335), .A2(EAX_REG_4__SCAN_IN), .ZN(n3898) );
  OAI211_X1 U4861 ( .C1(n3940), .C2(n4577), .A(n3899), .B(n3898), .ZN(n3902)
         );
  AOI21_X1 U4862 ( .B1(n3936), .B2(n3900), .A(n3945), .ZN(n5458) );
  NAND2_X1 U4863 ( .A1(n5458), .A2(n4299), .ZN(n3901) );
  NAND2_X1 U4864 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  NAND2_X1 U4865 ( .A1(n3904), .A2(n3903), .ZN(n4497) );
  BUF_X1 U4866 ( .A(n3905), .Z(n4584) );
  NAND2_X1 U4867 ( .A1(n4584), .A2(n4018), .ZN(n3906) );
  NAND2_X1 U4868 ( .A1(n3906), .A2(n4038), .ZN(n4473) );
  NAND2_X1 U4869 ( .A1(n3907), .A2(n4018), .ZN(n3911) );
  AOI22_X1 U4870 ( .A1(n4335), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6568), .ZN(n3909) );
  INV_X1 U4871 ( .A(n3940), .ZN(n3921) );
  NAND2_X1 U4872 ( .A1(n3921), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3908) );
  AND2_X1 U4873 ( .A1(n3909), .A2(n3908), .ZN(n3910) );
  NAND2_X1 U4874 ( .A1(n3911), .A2(n3910), .ZN(n4414) );
  NAND2_X1 U4875 ( .A1(n4857), .A2(n3912), .ZN(n3913) );
  NAND2_X1 U4876 ( .A1(n3913), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U4877 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6568), .ZN(n3916)
         );
  NAND2_X1 U4878 ( .A1(n4335), .A2(EAX_REG_0__SCAN_IN), .ZN(n3915) );
  OAI211_X1 U4879 ( .C1(n3940), .C2(n3917), .A(n3916), .B(n3915), .ZN(n3918)
         );
  AOI21_X1 U4880 ( .B1(n6528), .B2(n4018), .A(n3918), .ZN(n4481) );
  OR2_X1 U4881 ( .A1(n4482), .A2(n4481), .ZN(n4484) );
  INV_X1 U4882 ( .A(n4481), .ZN(n3919) );
  OR2_X1 U4883 ( .A1(n3919), .A2(n4333), .ZN(n3920) );
  NAND2_X1 U4884 ( .A1(n4484), .A2(n3920), .ZN(n4413) );
  NAND2_X1 U4885 ( .A1(n4414), .A2(n4413), .ZN(n4416) );
  NAND2_X1 U4886 ( .A1(n3921), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3927) );
  OAI21_X1 U4887 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3922), .ZN(n6109) );
  NAND2_X1 U4888 ( .A1(n6109), .A2(n4299), .ZN(n3924) );
  NAND2_X1 U4889 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3923)
         );
  NAND2_X1 U4890 ( .A1(n3924), .A2(n3923), .ZN(n3925) );
  AOI21_X1 U4891 ( .B1(n4335), .B2(EAX_REG_2__SCAN_IN), .A(n3925), .ZN(n3926)
         );
  AND2_X1 U4892 ( .A1(n3927), .A2(n3926), .ZN(n3928) );
  NAND2_X1 U4893 ( .A1(n4416), .A2(n3928), .ZN(n4472) );
  NAND2_X1 U4894 ( .A1(n4473), .A2(n4472), .ZN(n3932) );
  INV_X1 U4895 ( .A(n4416), .ZN(n3930) );
  INV_X1 U4896 ( .A(n3928), .ZN(n3929) );
  NAND2_X1 U4897 ( .A1(n3930), .A2(n3929), .ZN(n3931) );
  BUF_X1 U4898 ( .A(n3933), .Z(n3934) );
  NAND2_X1 U4899 ( .A1(n3934), .A2(n4018), .ZN(n3943) );
  OAI21_X1 U4900 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3937), .A(n3936), 
        .ZN(n6098) );
  AOI22_X1 U4901 ( .A1(n6098), .A2(n4299), .B1(n4334), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3939) );
  NAND2_X1 U4902 ( .A1(n4335), .A2(EAX_REG_3__SCAN_IN), .ZN(n3938) );
  OAI211_X1 U4903 ( .C1(n3940), .C2(n3935), .A(n3939), .B(n3938), .ZN(n3941)
         );
  INV_X1 U4904 ( .A(n3941), .ZN(n3942) );
  NAND2_X1 U4905 ( .A1(n3943), .A2(n3942), .ZN(n4502) );
  AND3_X2 U4906 ( .A1(n4497), .A2(n4470), .A3(n4502), .ZN(n4658) );
  NAND2_X1 U4907 ( .A1(n3944), .A2(n4018), .ZN(n3951) );
  INV_X1 U4908 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3948) );
  NAND2_X1 U4909 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3947)
         );
  OAI21_X1 U4910 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3945), .A(n3955), 
        .ZN(n6090) );
  NAND2_X1 U4911 ( .A1(n6090), .A2(n4299), .ZN(n3946) );
  OAI211_X1 U4912 ( .C1(n4228), .C2(n3948), .A(n3947), .B(n3946), .ZN(n3949)
         );
  INV_X1 U4913 ( .A(n3949), .ZN(n3950) );
  NAND2_X1 U4914 ( .A1(n3951), .A2(n3950), .ZN(n4657) );
  NAND2_X1 U4915 ( .A1(n3952), .A2(n4018), .ZN(n3959) );
  INV_X1 U4916 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3954) );
  OAI21_X1 U4917 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6353), .A(n6568), 
        .ZN(n3953) );
  OAI21_X1 U4918 ( .B1(n4228), .B2(n3954), .A(n3953), .ZN(n3957) );
  XOR2_X1 U4919 ( .A(n5154), .B(n3955), .Z(n5158) );
  NAND2_X1 U4920 ( .A1(n5158), .A2(n4299), .ZN(n3956) );
  NAND2_X1 U4921 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  NAND2_X1 U4922 ( .A1(n3959), .A2(n3958), .ZN(n4656) );
  NAND2_X1 U4923 ( .A1(n3961), .A2(n4655), .ZN(n4774) );
  XOR2_X1 U4924 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3980), .Z(n5954) );
  INV_X1 U4925 ( .A(n5954), .ZN(n3977) );
  AOI22_X1 U4926 ( .A1(n4178), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4927 ( .A1(n3121), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4928 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4285), .B1(n4307), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4929 ( .A1(n4313), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U4930 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3972)
         );
  AOI22_X1 U4931 ( .A1(n4284), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4932 ( .A1(n4305), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4933 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4317), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4934 ( .A1(n4316), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3967) );
  NAND4_X1 U4935 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3971)
         );
  OAI21_X1 U4936 ( .B1(n3972), .B2(n3971), .A(n4018), .ZN(n3975) );
  NAND2_X1 U4937 ( .A1(n4335), .A2(EAX_REG_12__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4938 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3973)
         );
  NAND3_X1 U4939 ( .A1(n3975), .A2(n3974), .A3(n3973), .ZN(n3976) );
  AOI21_X1 U4940 ( .B1(n3977), .B2(n4299), .A(n3976), .ZN(n4790) );
  INV_X1 U4941 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U4942 ( .A1(n3981), .A2(n6943), .ZN(n3983) );
  INV_X1 U4943 ( .A(n4021), .ZN(n3982) );
  NAND2_X1 U4944 ( .A1(n3983), .A2(n3982), .ZN(n5441) );
  AOI22_X1 U4945 ( .A1(n4178), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4946 ( .A1(n3121), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4947 ( .A1(n4305), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4948 ( .A1(n4315), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U4949 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3993)
         );
  AOI22_X1 U4950 ( .A1(n4317), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4951 ( .A1(n4177), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4952 ( .A1(n4284), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4953 ( .A1(n4316), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4954 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3992)
         );
  OAI21_X1 U4955 ( .B1(n3993), .B2(n3992), .A(n4018), .ZN(n3995) );
  NAND2_X1 U4956 ( .A1(n4335), .A2(EAX_REG_13__SCAN_IN), .ZN(n3994) );
  AOI21_X1 U4957 ( .B1(n5441), .B2(n4299), .A(n3996), .ZN(n4784) );
  INV_X1 U4958 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U4959 ( .A(n5232), .B(n4021), .ZN(n5270) );
  AOI22_X1 U4960 ( .A1(n4305), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4961 ( .A1(n4284), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4962 ( .A1(n4178), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4963 ( .A1(n4316), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4964 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4006)
         );
  AOI22_X1 U4965 ( .A1(n3121), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4966 ( .A1(n4307), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4967 ( .A1(n4177), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4968 ( .A1(n4317), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4969 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  OR2_X1 U4970 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  AOI22_X1 U4971 ( .A1(n4018), .A2(n4007), .B1(n4334), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U4972 ( .A1(n4335), .A2(EAX_REG_14__SCAN_IN), .ZN(n4008) );
  OAI211_X1 U4973 ( .C1(n5270), .C2(n4333), .A(n4009), .B(n4008), .ZN(n4808)
         );
  AOI22_X1 U4974 ( .A1(n4178), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4975 ( .A1(n4305), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4976 ( .A1(n4285), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4977 ( .A1(n4317), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4978 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4020)
         );
  AOI22_X1 U4979 ( .A1(n3121), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4980 ( .A1(n4313), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4981 ( .A1(n4284), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4982 ( .A1(n4307), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4983 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4019)
         );
  OAI21_X1 U4984 ( .B1(n4020), .B2(n4019), .A(n4018), .ZN(n4025) );
  INV_X1 U4985 ( .A(n4026), .ZN(n4022) );
  XNOR2_X1 U4986 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4022), .ZN(n5430)
         );
  AOI22_X1 U4987 ( .A1(n4299), .A2(n5430), .B1(n4334), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U4988 ( .A1(n4335), .A2(EAX_REG_15__SCAN_IN), .ZN(n4023) );
  NOR2_X2 U4989 ( .A1(n4807), .A2(n4993), .ZN(n4994) );
  INV_X1 U4990 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6733) );
  INV_X1 U4991 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5429) );
  AOI21_X1 U4992 ( .B1(n6733), .B2(n4027), .A(n4073), .ZN(n5621) );
  OR2_X1 U4993 ( .A1(n5621), .A2(n4333), .ZN(n4042) );
  AOI22_X1 U4994 ( .A1(n4284), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4995 ( .A1(n4307), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4996 ( .A1(n4313), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4997 ( .A1(n4317), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U4998 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4037)
         );
  AOI22_X1 U4999 ( .A1(n4178), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5000 ( .A1(n4177), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5001 ( .A1(n4260), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5002 ( .A1(n4285), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U5003 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4036)
         );
  OR2_X1 U5004 ( .A1(n4037), .A2(n4036), .ZN(n4040) );
  INV_X1 U5005 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4451) );
  OAI22_X1 U5006 ( .A1(n4228), .A2(n4451), .B1(n4038), .B2(n6733), .ZN(n4039)
         );
  AOI21_X1 U5007 ( .B1(n4296), .B2(n4040), .A(n4039), .ZN(n4041) );
  AND2_X2 U5008 ( .A1(n4994), .A2(n4043), .ZN(n5068) );
  XNOR2_X1 U5009 ( .A(n4073), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5607)
         );
  NAND2_X1 U5010 ( .A1(n5607), .A2(n4299), .ZN(n4058) );
  AOI22_X1 U5011 ( .A1(n4313), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5012 ( .A1(n4177), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5013 ( .A1(n4285), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5014 ( .A1(n4317), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U5015 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4053)
         );
  AOI22_X1 U5016 ( .A1(n4178), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U5017 ( .A1(n3121), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U5018 ( .A1(n4284), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5019 ( .A1(n4314), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U5020 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4052)
         );
  NOR2_X1 U5021 ( .A1(n4053), .A2(n4052), .ZN(n4055) );
  AOI22_X1 U5022 ( .A1(n4335), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6568), .ZN(n4054) );
  OAI21_X1 U5023 ( .B1(n4330), .B2(n4055), .A(n4054), .ZN(n4056) );
  NAND2_X1 U5024 ( .A1(n4056), .A2(n4333), .ZN(n4057) );
  NAND2_X1 U5025 ( .A1(n4058), .A2(n4057), .ZN(n5092) );
  AND2_X2 U5026 ( .A1(n5068), .A2(n5092), .ZN(n5091) );
  AOI22_X1 U5027 ( .A1(n4305), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5028 ( .A1(n4315), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5029 ( .A1(n4307), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5030 ( .A1(n4317), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5031 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4068)
         );
  AOI22_X1 U5032 ( .A1(n4178), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5033 ( .A1(n3121), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5034 ( .A1(n4284), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5035 ( .A1(n4308), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5036 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR2_X1 U5037 ( .A1(n4068), .A2(n4067), .ZN(n4072) );
  OAI21_X1 U5038 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6353), .A(n6568), 
        .ZN(n4069) );
  INV_X1 U5039 ( .A(n4069), .ZN(n4070) );
  AOI21_X1 U5040 ( .B1(n4335), .B2(EAX_REG_18__SCAN_IN), .A(n4070), .ZN(n4071)
         );
  OAI21_X1 U5041 ( .B1(n4330), .B2(n4072), .A(n4071), .ZN(n4077) );
  INV_X1 U5042 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5609) );
  OAI21_X1 U5043 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4075), .A(n4091), 
        .ZN(n5949) );
  OR2_X1 U5044 ( .A1(n4333), .A2(n5949), .ZN(n4076) );
  AOI22_X1 U5045 ( .A1(n4305), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5046 ( .A1(n3121), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5047 ( .A1(n4178), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5048 ( .A1(n4177), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4078) );
  NAND4_X1 U5049 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .ZN(n4087)
         );
  AOI22_X1 U5050 ( .A1(n4317), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5051 ( .A1(n4284), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5052 ( .A1(n4314), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5053 ( .A1(n4316), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5054 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4086)
         );
  NOR2_X1 U5055 ( .A1(n4087), .A2(n4086), .ZN(n4090) );
  INV_X1 U5056 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6804) );
  AOI21_X1 U5057 ( .B1(n6804), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4088) );
  AOI21_X1 U5058 ( .B1(n4335), .B2(EAX_REG_19__SCAN_IN), .A(n4088), .ZN(n4089)
         );
  OAI21_X1 U5059 ( .B1(n4330), .B2(n4090), .A(n4089), .ZN(n4095) );
  NOR2_X1 U5060 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4092), .ZN(n4093)
         );
  NOR2_X1 U5061 ( .A1(n4110), .A2(n4093), .ZN(n5594) );
  NAND2_X1 U5062 ( .A1(n5594), .A2(n4299), .ZN(n4094) );
  NAND2_X1 U5063 ( .A1(n4095), .A2(n4094), .ZN(n5205) );
  AOI22_X1 U5064 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3121), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5065 ( .A1(n4178), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5066 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n4177), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5067 ( .A1(n4317), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4096) );
  NAND4_X1 U5068 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4105)
         );
  AOI22_X1 U5069 ( .A1(n4284), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5070 ( .A1(n4305), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5071 ( .A1(n4314), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5072 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4315), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4100) );
  NAND4_X1 U5073 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104)
         );
  NOR2_X1 U5074 ( .A1(n4105), .A2(n4104), .ZN(n4109) );
  NAND2_X1 U5075 ( .A1(n6568), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4106)
         );
  NAND2_X1 U5076 ( .A1(n4333), .A2(n4106), .ZN(n4107) );
  AOI21_X1 U5077 ( .B1(n4335), .B2(EAX_REG_20__SCAN_IN), .A(n4107), .ZN(n4108)
         );
  OAI21_X1 U5078 ( .B1(n4330), .B2(n4109), .A(n4108), .ZN(n4112) );
  OAI21_X1 U5079 ( .B1(n4110), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4127), 
        .ZN(n5824) );
  OR2_X1 U5080 ( .A1(n5824), .A2(n4333), .ZN(n4111) );
  NAND2_X1 U5081 ( .A1(n4112), .A2(n4111), .ZN(n5219) );
  AOI22_X1 U5082 ( .A1(n4178), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5083 ( .A1(n4284), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5084 ( .A1(n4307), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5085 ( .A1(n4308), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4114) );
  NAND4_X1 U5086 ( .A1(n4117), .A2(n4116), .A3(n4115), .A4(n4114), .ZN(n4123)
         );
  AOI22_X1 U5087 ( .A1(n3121), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5088 ( .A1(n3120), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5089 ( .A1(n4285), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5090 ( .A1(n4317), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4118) );
  NAND4_X1 U5091 ( .A1(n4121), .A2(n4120), .A3(n4119), .A4(n4118), .ZN(n4122)
         );
  NOR2_X1 U5092 ( .A1(n4123), .A2(n4122), .ZN(n4126) );
  INV_X1 U5093 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6790) );
  OAI21_X1 U5094 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6790), .A(n4333), .ZN(
        n4124) );
  AOI21_X1 U5095 ( .B1(n4335), .B2(EAX_REG_21__SCAN_IN), .A(n4124), .ZN(n4125)
         );
  OAI21_X1 U5096 ( .B1(n4330), .B2(n4126), .A(n4125), .ZN(n4130) );
  AND2_X1 U5097 ( .A1(n4127), .A2(n6790), .ZN(n4128) );
  NOR2_X1 U5098 ( .A1(n4145), .A2(n4128), .ZN(n5579) );
  NAND2_X1 U5099 ( .A1(n5579), .A2(n4299), .ZN(n4129) );
  NAND2_X1 U5100 ( .A1(n4130), .A2(n4129), .ZN(n5285) );
  AOI22_X1 U5101 ( .A1(n3121), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5102 ( .A1(n4178), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5103 ( .A1(n4307), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5104 ( .A1(n4285), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4131) );
  NAND4_X1 U5105 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4140)
         );
  AOI22_X1 U5106 ( .A1(n4284), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5107 ( .A1(n4305), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5108 ( .A1(n4177), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5109 ( .A1(n4317), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5110 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4139)
         );
  NOR2_X1 U5111 ( .A1(n4140), .A2(n4139), .ZN(n4144) );
  NAND2_X1 U5112 ( .A1(n6568), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4141)
         );
  NAND2_X1 U5113 ( .A1(n4333), .A2(n4141), .ZN(n4142) );
  AOI21_X1 U5114 ( .B1(n4335), .B2(EAX_REG_22__SCAN_IN), .A(n4142), .ZN(n4143)
         );
  OAI21_X1 U5115 ( .B1(n4330), .B2(n4144), .A(n4143), .ZN(n4148) );
  OR2_X1 U5116 ( .A1(n4145), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4146)
         );
  AND2_X1 U5117 ( .A1(n4190), .A2(n4146), .ZN(n5817) );
  NAND2_X1 U5118 ( .A1(n5817), .A2(n4299), .ZN(n4147) );
  AOI22_X1 U5119 ( .A1(n4305), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5120 ( .A1(n3121), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5121 ( .A1(n4178), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5122 ( .A1(n4177), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U5123 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4158)
         );
  AOI22_X1 U5124 ( .A1(n4317), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5125 ( .A1(n4284), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5126 ( .A1(n4314), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5127 ( .A1(n4316), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4153) );
  NAND4_X1 U5128 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157)
         );
  NOR2_X1 U5129 ( .A1(n4158), .A2(n4157), .ZN(n4176) );
  AOI22_X1 U5130 ( .A1(n4178), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5131 ( .A1(n4177), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4315), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5132 ( .A1(n4313), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5133 ( .A1(n4317), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4159) );
  NAND4_X1 U5134 ( .A1(n4162), .A2(n4161), .A3(n4160), .A4(n4159), .ZN(n4168)
         );
  AOI22_X1 U5135 ( .A1(n3121), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5136 ( .A1(n4307), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5137 ( .A1(n4284), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5138 ( .A1(n4308), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U5139 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4167)
         );
  NOR2_X1 U5140 ( .A1(n4168), .A2(n4167), .ZN(n4175) );
  XOR2_X1 U5141 ( .A(n4176), .B(n4175), .Z(n4169) );
  NAND2_X1 U5142 ( .A1(n4169), .A2(n4296), .ZN(n4172) );
  INV_X1 U5143 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5565) );
  OAI21_X1 U5144 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5565), .A(n4333), .ZN(
        n4170) );
  AOI21_X1 U5145 ( .B1(n4335), .B2(EAX_REG_23__SCAN_IN), .A(n4170), .ZN(n4171)
         );
  NAND2_X1 U5146 ( .A1(n4172), .A2(n4171), .ZN(n4174) );
  XNOR2_X1 U5147 ( .A(n4190), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5563)
         );
  NAND2_X1 U5148 ( .A1(n5563), .A2(n4299), .ZN(n4173) );
  NAND2_X1 U5149 ( .A1(n4174), .A2(n4173), .ZN(n5389) );
  OR2_X1 U5150 ( .A1(n4176), .A2(n4175), .ZN(n4197) );
  AOI22_X1 U5151 ( .A1(n4178), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5152 ( .A1(n4284), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5153 ( .A1(n4307), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5154 ( .A1(n4313), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4179) );
  NAND4_X1 U5155 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4188)
         );
  INV_X1 U5156 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6957) );
  AOI22_X1 U5157 ( .A1(n4317), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4285), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U5158 ( .A1(n4308), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4316), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5159 ( .A1(n3120), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U5160 ( .A1(n3121), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4183) );
  NAND4_X1 U5161 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4187)
         );
  NOR2_X1 U5162 ( .A1(n4188), .A2(n4187), .ZN(n4196) );
  INV_X1 U5163 ( .A(n4196), .ZN(n4189) );
  XNOR2_X1 U5164 ( .A(n4197), .B(n4189), .ZN(n4194) );
  INV_X1 U5165 ( .A(EAX_REG_24__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U5166 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4192)
         );
  XNOR2_X1 U5167 ( .A(n4210), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6688)
         );
  OAI211_X1 U5168 ( .C1(n4228), .C2(n7002), .A(n4192), .B(n4191), .ZN(n4193)
         );
  AOI21_X1 U5169 ( .B1(n4194), .B2(n4296), .A(n4193), .ZN(n5311) );
  OR2_X1 U5170 ( .A1(n4197), .A2(n4196), .ZN(n4214) );
  AOI22_X1 U5171 ( .A1(n4284), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5172 ( .A1(n4305), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5173 ( .A1(n4314), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5174 ( .A1(n4316), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4198) );
  NAND4_X1 U5175 ( .A1(n4201), .A2(n4200), .A3(n4199), .A4(n4198), .ZN(n4207)
         );
  AOI22_X1 U5176 ( .A1(n3121), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5177 ( .A1(n4317), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4315), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5178 ( .A1(n4178), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5179 ( .A1(n4307), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U5180 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4206)
         );
  NOR2_X1 U5181 ( .A1(n4207), .A2(n4206), .ZN(n4215) );
  XOR2_X1 U5182 ( .A(n4214), .B(n4215), .Z(n4208) );
  NAND2_X1 U5183 ( .A1(n4208), .A2(n4296), .ZN(n4213) );
  INV_X1 U5184 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5796) );
  OAI21_X1 U5185 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5796), .A(n4333), .ZN(
        n4209) );
  AOI21_X1 U5186 ( .B1(n4335), .B2(EAX_REG_25__SCAN_IN), .A(n4209), .ZN(n4212)
         );
  INV_X1 U5187 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5306) );
  XNOR2_X1 U5188 ( .A(n4231), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5799)
         );
  AOI21_X1 U5189 ( .B1(n4213), .B2(n4212), .A(n4211), .ZN(n5498) );
  NAND2_X1 U5190 ( .A1(n5499), .A2(n5498), .ZN(n5488) );
  NOR2_X1 U5191 ( .A1(n4215), .A2(n4214), .ZN(n4239) );
  AOI22_X1 U5192 ( .A1(n4305), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5193 ( .A1(n3121), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5194 ( .A1(n4178), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5195 ( .A1(n4177), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4216) );
  NAND4_X1 U5196 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4225)
         );
  AOI22_X1 U5197 ( .A1(n4317), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4315), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U5198 ( .A1(n4284), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5199 ( .A1(n4314), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5200 ( .A1(n4316), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4220) );
  NAND4_X1 U5201 ( .A1(n4223), .A2(n4222), .A3(n4221), .A4(n4220), .ZN(n4224)
         );
  OR2_X1 U5202 ( .A1(n4225), .A2(n4224), .ZN(n4238) );
  INV_X1 U5203 ( .A(n4238), .ZN(n4226) );
  XNOR2_X1 U5204 ( .A(n4239), .B(n4226), .ZN(n4230) );
  INV_X1 U5205 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U5206 ( .A1(n6568), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4227)
         );
  OAI211_X1 U5207 ( .C1(n4228), .C2(n4447), .A(n4333), .B(n4227), .ZN(n4229)
         );
  AOI21_X1 U5208 ( .B1(n4230), .B2(n4296), .A(n4229), .ZN(n4237) );
  INV_X1 U5209 ( .A(n4232), .ZN(n4234) );
  INV_X1 U5210 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U5211 ( .A1(n4234), .A2(n4233), .ZN(n4235) );
  NAND2_X1 U5212 ( .A1(n4254), .A2(n4235), .ZN(n5795) );
  NOR2_X1 U5213 ( .A1(n5795), .A2(n4333), .ZN(n4236) );
  OR2_X2 U5214 ( .A1(n5488), .A2(n5492), .ZN(n5490) );
  NAND2_X1 U5215 ( .A1(n4239), .A2(n4238), .ZN(n4258) );
  AOI22_X1 U5216 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4284), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5217 ( .A1(n4178), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5218 ( .A1(n4317), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5219 ( .A1(n3213), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4240) );
  NAND4_X1 U5220 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4249)
         );
  AOI22_X1 U5221 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4177), .B1(n4313), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U5222 ( .A1(n4285), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U5223 ( .A1(n4305), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U5224 ( .A1(n4307), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4244) );
  NAND4_X1 U5225 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4248)
         );
  NOR2_X1 U5226 ( .A1(n4249), .A2(n4248), .ZN(n4259) );
  XOR2_X1 U5227 ( .A(n4258), .B(n4259), .Z(n4250) );
  NAND2_X1 U5228 ( .A1(n4250), .A2(n4296), .ZN(n4253) );
  INV_X1 U5229 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6762) );
  OAI21_X1 U5230 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6762), .A(n4333), .ZN(
        n4251) );
  AOI21_X1 U5231 ( .B1(n4335), .B2(EAX_REG_27__SCAN_IN), .A(n4251), .ZN(n4252)
         );
  NAND2_X1 U5232 ( .A1(n4253), .A2(n4252), .ZN(n4257) );
  NAND2_X1 U5233 ( .A1(n4254), .A2(n6762), .ZN(n4255) );
  AND2_X1 U5234 ( .A1(n4277), .A2(n4255), .ZN(n5778) );
  NAND2_X1 U5235 ( .A1(n5778), .A2(n4299), .ZN(n4256) );
  NAND2_X1 U5236 ( .A1(n4257), .A2(n4256), .ZN(n5484) );
  NOR2_X1 U5237 ( .A1(n4259), .A2(n4258), .ZN(n4283) );
  AOI22_X1 U5238 ( .A1(n4305), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U5239 ( .A1(n3121), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U5240 ( .A1(n4178), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U5241 ( .A1(n4177), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4261) );
  NAND4_X1 U5242 ( .A1(n4264), .A2(n4263), .A3(n4262), .A4(n4261), .ZN(n4270)
         );
  AOI22_X1 U5243 ( .A1(n4317), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4315), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5244 ( .A1(n4284), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5245 ( .A1(n4314), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U5246 ( .A1(n3213), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4265) );
  NAND4_X1 U5247 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4269)
         );
  OR2_X1 U5248 ( .A1(n4270), .A2(n4269), .ZN(n4282) );
  INV_X1 U5249 ( .A(n4282), .ZN(n4271) );
  XNOR2_X1 U5250 ( .A(n4283), .B(n4271), .ZN(n4272) );
  NAND2_X1 U5251 ( .A1(n4272), .A2(n4296), .ZN(n4281) );
  NAND2_X1 U5252 ( .A1(n6568), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4273)
         );
  NAND2_X1 U5253 ( .A1(n4333), .A2(n4273), .ZN(n4274) );
  AOI21_X1 U5254 ( .B1(n4335), .B2(EAX_REG_28__SCAN_IN), .A(n4274), .ZN(n4280)
         );
  INV_X1 U5255 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U5256 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  NAND2_X1 U5257 ( .A1(n4301), .A2(n4278), .ZN(n5769) );
  NOR2_X1 U5258 ( .A1(n5769), .A2(n4333), .ZN(n4279) );
  AOI21_X1 U5259 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(n5473) );
  AND2_X2 U5260 ( .A1(n5485), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U5261 ( .A1(n4283), .A2(n4282), .ZN(n4324) );
  AOI22_X1 U5262 ( .A1(n4178), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4289) );
  AOI22_X1 U5263 ( .A1(n4284), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4307), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4288) );
  AOI22_X1 U5264 ( .A1(n4177), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4287) );
  AOI22_X1 U5265 ( .A1(n4285), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4286) );
  NAND4_X1 U5266 ( .A1(n4289), .A2(n4288), .A3(n4287), .A4(n4286), .ZN(n4295)
         );
  AOI22_X1 U5267 ( .A1(n4313), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4305), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U5268 ( .A1(n3121), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U5269 ( .A1(n4314), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4308), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U5270 ( .A1(n4317), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4290) );
  NAND4_X1 U5271 ( .A1(n4293), .A2(n4292), .A3(n4291), .A4(n4290), .ZN(n4294)
         );
  NOR2_X1 U5272 ( .A1(n4295), .A2(n4294), .ZN(n4325) );
  XOR2_X1 U5273 ( .A(n4324), .B(n4325), .Z(n4297) );
  NAND2_X1 U5274 ( .A1(n4297), .A2(n4296), .ZN(n4304) );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U5276 ( .A1(n6706), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4298) );
  AOI211_X1 U5277 ( .C1(n4335), .C2(EAX_REG_29__SCAN_IN), .A(n4299), .B(n4298), 
        .ZN(n4303) );
  NAND2_X1 U5278 ( .A1(n4301), .A2(n6706), .ZN(n4302) );
  AND2_X1 U5279 ( .A1(n4342), .A2(n4302), .ZN(n5370) );
  AOI22_X1 U5280 ( .A1(n4304), .A2(n4303), .B1(n4299), .B2(n5370), .ZN(n5360)
         );
  INV_X1 U5282 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4341) );
  XNOR2_X1 U5283 ( .A(n4342), .B(n4341), .ZN(n5379) );
  AOI22_X1 U5284 ( .A1(n4305), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U5285 ( .A1(n3460), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4306), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U5286 ( .A1(n4307), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4260), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4310) );
  AOI22_X1 U5287 ( .A1(n4308), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4309) );
  NAND4_X1 U5288 ( .A1(n4312), .A2(n4311), .A3(n4310), .A4(n4309), .ZN(n4323)
         );
  AOI22_X1 U5289 ( .A1(n4178), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4313), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U5290 ( .A1(n4284), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U5291 ( .A1(n4315), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4314), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U5292 ( .A1(n4317), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4318) );
  NAND4_X1 U5293 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4322)
         );
  NOR2_X1 U5294 ( .A1(n4323), .A2(n4322), .ZN(n4327) );
  NOR2_X1 U5295 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  XOR2_X1 U5296 ( .A(n4327), .B(n4326), .Z(n4331) );
  AOI21_X1 U5297 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6568), .A(n4299), 
        .ZN(n4329) );
  NAND2_X1 U5298 ( .A1(n4335), .A2(EAX_REG_30__SCAN_IN), .ZN(n4328) );
  OAI211_X1 U5299 ( .C1(n4331), .C2(n4330), .A(n4329), .B(n4328), .ZN(n4332)
         );
  OAI21_X1 U5300 ( .B1(n4333), .B2(n5379), .A(n4332), .ZN(n5350) );
  AOI22_X1 U5301 ( .A1(n4335), .A2(EAX_REG_31__SCAN_IN), .B1(n4334), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4336) );
  XNOR2_X2 U5302 ( .A(n5349), .B(n4336), .ZN(n5517) );
  AND2_X1 U5303 ( .A1(n6972), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5304 ( .A1(n5112), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6574) );
  NOR2_X1 U5305 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6324) );
  INV_X1 U5306 ( .A(n6324), .ZN(n6401) );
  NAND2_X1 U5307 ( .A1(n6401), .A2(n4337), .ZN(n6676) );
  NAND2_X1 U5308 ( .A1(n6676), .A2(n6972), .ZN(n4338) );
  NAND2_X1 U5309 ( .A1(n6972), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U5310 ( .A1(n6353), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4339) );
  AND2_X1 U5311 ( .A1(n4340), .A2(n4339), .ZN(n4511) );
  INV_X1 U5312 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5313 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4345)
         );
  OAI211_X1 U5314 ( .C1(n6110), .C2(n5117), .A(n4346), .B(n4345), .ZN(n4347)
         );
  AOI21_X1 U5315 ( .B1(n5517), .B2(n6105), .A(n4347), .ZN(n4348) );
  NAND2_X1 U5316 ( .A1(n4349), .A2(n4348), .ZN(U2955) );
  INV_X1 U5317 ( .A(n4419), .ZN(n4356) );
  AND2_X1 U5318 ( .A1(n3632), .A2(n4352), .ZN(n4360) );
  OAI22_X1 U5319 ( .A1(n4356), .A2(n5171), .B1(n4437), .B2(n4360), .ZN(n5918)
         );
  NAND2_X1 U5320 ( .A1(n3395), .A2(n5176), .ZN(n4363) );
  AOI21_X1 U5321 ( .B1(n4363), .B2(n6583), .A(READY_N), .ZN(n6678) );
  NOR2_X1 U5322 ( .A1(n5918), .A2(n6678), .ZN(n6543) );
  NOR2_X1 U5323 ( .A1(n6543), .A2(n5917), .ZN(n5926) );
  INV_X1 U5324 ( .A(MORE_REG_SCAN_IN), .ZN(n6736) );
  NOR3_X1 U5325 ( .A1(n4490), .A2(n4351), .A3(n4437), .ZN(n4354) );
  OAI22_X1 U5326 ( .A1(n4356), .A2(n4354), .B1(n4353), .B2(n4352), .ZN(n4355)
         );
  AOI21_X1 U5327 ( .B1(n4417), .B2(n4356), .A(n4355), .ZN(n6546) );
  INV_X1 U5328 ( .A(n6546), .ZN(n4357) );
  NAND2_X1 U5329 ( .A1(n5926), .A2(n4357), .ZN(n4358) );
  OAI21_X1 U5330 ( .B1(n5926), .B2(n6736), .A(n4358), .ZN(U3471) );
  NAND2_X1 U5331 ( .A1(n4491), .A2(n4437), .ZN(n4362) );
  NAND2_X1 U5332 ( .A1(n6447), .A2(n6557), .ZN(n4359) );
  NAND2_X1 U5333 ( .A1(n4362), .A2(n4359), .ZN(n5766) );
  NAND2_X1 U5334 ( .A1(n4360), .A2(n6566), .ZN(n5767) );
  INV_X1 U5335 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n4361) );
  NAND2_X1 U5336 ( .A1(n5767), .A2(n4361), .ZN(n4365) );
  NAND2_X1 U5337 ( .A1(n4362), .A2(n5767), .ZN(n6675) );
  NAND2_X1 U5338 ( .A1(n6675), .A2(n4363), .ZN(n4364) );
  OAI21_X1 U5339 ( .B1(n5766), .B2(n4365), .A(n4364), .ZN(n4366) );
  INV_X1 U5340 ( .A(n4366), .ZN(U3474) );
  INV_X1 U5341 ( .A(n4368), .ZN(n4369) );
  NOR2_X1 U5342 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  AND2_X1 U5343 ( .A1(n5910), .A2(n4371), .ZN(n4373) );
  NAND2_X1 U5344 ( .A1(n4373), .A2(n4372), .ZN(n6527) );
  NAND2_X1 U5345 ( .A1(n6004), .A2(n6527), .ZN(n4380) );
  INV_X1 U5346 ( .A(n4374), .ZN(n4574) );
  INV_X1 U5347 ( .A(n4376), .ZN(n4407) );
  NAND2_X1 U5348 ( .A1(n4574), .A2(n4407), .ZN(n4377) );
  NOR2_X1 U5349 ( .A1(n6525), .A2(n4377), .ZN(n4378) );
  AOI21_X1 U5350 ( .B1(n6529), .B2(n3287), .A(n4378), .ZN(n4379) );
  NAND2_X1 U5351 ( .A1(n4380), .A2(n4379), .ZN(n6531) );
  INV_X1 U5352 ( .A(n6661), .ZN(n5912) );
  AOI22_X1 U5353 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3818), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4464), .ZN(n4405) );
  NOR2_X1 U5354 ( .A1(n6557), .A2(n4406), .ZN(n4382) );
  AOI222_X1 U5355 ( .A1(n6531), .A2(n5912), .B1(n4405), .B2(n4382), .C1(n4381), 
        .C2(n4397), .ZN(n4396) );
  INV_X1 U5356 ( .A(n6583), .ZN(n5126) );
  NAND2_X1 U5357 ( .A1(n6529), .A2(n5126), .ZN(n4384) );
  NAND2_X1 U5358 ( .A1(n4437), .A2(n5123), .ZN(n4383) );
  NAND2_X1 U5359 ( .A1(n4384), .A2(n4383), .ZN(n4385) );
  AOI21_X1 U5360 ( .B1(n4385), .B2(n6892), .A(n4490), .ZN(n4386) );
  OR2_X1 U5361 ( .A1(n4419), .A2(n4386), .ZN(n4393) );
  NAND2_X1 U5362 ( .A1(n4419), .A2(n4417), .ZN(n4392) );
  INV_X1 U5363 ( .A(n4485), .ZN(n4389) );
  OAI211_X1 U5364 ( .C1(n5910), .C2(n4389), .A(n4388), .B(n4387), .ZN(n4390)
         );
  INV_X1 U5365 ( .A(n4390), .ZN(n4391) );
  NAND3_X1 U5366 ( .A1(n4393), .A2(n4392), .A3(n4391), .ZN(n6532) );
  INV_X1 U5367 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5925) );
  NOR2_X1 U5368 ( .A1(n6568), .A2(n6557), .ZN(n4594) );
  NAND2_X1 U5369 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4594), .ZN(n6652) );
  NOR2_X1 U5370 ( .A1(n5925), .A2(n6652), .ZN(n4394) );
  AOI21_X1 U5371 ( .B1(n6566), .B2(n6532), .A(n4394), .ZN(n5915) );
  NAND2_X1 U5372 ( .A1(n6972), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U5373 ( .A1(n5915), .A2(n6653), .ZN(n6659) );
  INV_X1 U5374 ( .A(n6659), .ZN(n4410) );
  NOR2_X1 U5375 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6558), .ZN(n6655)
         );
  OAI21_X1 U5376 ( .B1(n4410), .B2(n6655), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4395) );
  OAI21_X1 U5377 ( .B1(n4396), .B2(n4410), .A(n4395), .ZN(U3460) );
  AOI21_X1 U5378 ( .B1(n4397), .B2(n4407), .A(n4410), .ZN(n4412) );
  NAND2_X1 U5379 ( .A1(n5178), .A2(n6527), .ZN(n4404) );
  OR2_X1 U5380 ( .A1(n4417), .A2(n4490), .ZN(n4567) );
  XNOR2_X1 U5381 ( .A(n4376), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4402)
         );
  XNOR2_X1 U5382 ( .A(n3287), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4399)
         );
  NAND2_X1 U5383 ( .A1(n6529), .A2(n4399), .ZN(n4400) );
  OAI21_X1 U5384 ( .B1(n4402), .B2(n4557), .A(n4400), .ZN(n4401) );
  AOI21_X1 U5385 ( .B1(n4567), .B2(n4402), .A(n4401), .ZN(n4403) );
  NAND2_X1 U5386 ( .A1(n4404), .A2(n4403), .ZN(n4553) );
  NOR3_X1 U5387 ( .A1(n6557), .A2(n4406), .A3(n4405), .ZN(n4409) );
  NOR3_X1 U5388 ( .A1(n4407), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6558), 
        .ZN(n4408) );
  AOI211_X1 U5389 ( .C1(n4553), .C2(n5912), .A(n4409), .B(n4408), .ZN(n4411)
         );
  OAI22_X1 U5390 ( .A1(n4412), .A2(n3140), .B1(n4411), .B2(n4410), .ZN(U3459)
         );
  OR2_X1 U5391 ( .A1(n4414), .A2(n4413), .ZN(n4415) );
  AND2_X1 U5392 ( .A1(n4416), .A2(n4415), .ZN(n6001) );
  INV_X1 U5393 ( .A(n6001), .ZN(n4699) );
  AND2_X1 U5394 ( .A1(n4417), .A2(n6566), .ZN(n4418) );
  NAND2_X1 U5395 ( .A1(n4419), .A2(n4418), .ZN(n4426) );
  INV_X1 U5396 ( .A(n4420), .ZN(n4423) );
  NOR2_X1 U5397 ( .A1(n4643), .A2(n5917), .ZN(n4421) );
  NAND4_X1 U5398 ( .A1(n4423), .A2(n5516), .A3(n4422), .A4(n4421), .ZN(n4486)
         );
  OR2_X1 U5399 ( .A1(n4486), .A2(n4424), .ZN(n4425) );
  NAND2_X1 U5400 ( .A1(n5505), .A2(n5098), .ZN(n5228) );
  NAND2_X1 U5401 ( .A1(n5505), .A2(n5516), .ZN(n5507) );
  XNOR2_X1 U5402 ( .A(n4427), .B(n4428), .ZN(n4468) );
  AOI22_X1 U5403 ( .A1(n5512), .A2(n4468), .B1(n5511), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4429) );
  OAI21_X1 U5404 ( .B1(n4699), .B2(n5228), .A(n4429), .ZN(U2858) );
  INV_X1 U5405 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4434) );
  INV_X1 U5406 ( .A(n6555), .ZN(n4430) );
  NAND2_X1 U5407 ( .A1(n4491), .A2(n6529), .ZN(n4431) );
  NAND2_X1 U5408 ( .A1(n6060), .A2(n4431), .ZN(n4432) );
  NAND2_X1 U5409 ( .A1(n6023), .A2(n5122), .ZN(n4686) );
  AOI22_X1 U5410 ( .A1(DATAO_REG_23__SCAN_IN), .A2(n6039), .B1(
        UWORD_REG_7__SCAN_IN), .B2(n6677), .ZN(n4433) );
  OAI21_X1 U5411 ( .B1(n4434), .B2(n4686), .A(n4433), .ZN(U2900) );
  AOI22_X1 U5412 ( .A1(DATAO_REG_16__SCAN_IN), .A2(n6039), .B1(
        UWORD_REG_0__SCAN_IN), .B2(n6677), .ZN(n4435) );
  OAI21_X1 U5413 ( .B1(n4451), .B2(n4686), .A(n4435), .ZN(U2907) );
  INV_X1 U5414 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U5415 ( .A1(DATAO_REG_25__SCAN_IN), .A2(n6039), .B1(
        UWORD_REG_9__SCAN_IN), .B2(n6677), .ZN(n4436) );
  OAI21_X1 U5416 ( .B1(n6707), .B2(n4686), .A(n4436), .ZN(U2898) );
  INV_X1 U5417 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4442) );
  NAND2_X1 U5418 ( .A1(n4437), .A2(n6892), .ZN(n4438) );
  NOR2_X1 U5419 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  NOR2_X2 U5420 ( .A1(n6072), .A2(n4440), .ZN(n6071) );
  NAND2_X1 U5421 ( .A1(n6071), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4441) );
  NAND2_X1 U5422 ( .A1(n4440), .A2(n4605), .ZN(n6052) );
  INV_X1 U5423 ( .A(DATAI_10_), .ZN(n5049) );
  OR2_X1 U5424 ( .A1(n6052), .A2(n5049), .ZN(n4445) );
  OAI211_X1 U5425 ( .C1(n6060), .C2(n4442), .A(n4441), .B(n4445), .ZN(U2949)
         );
  INV_X1 U5426 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U5427 ( .A1(n6071), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4443) );
  INV_X1 U5428 ( .A(DATAI_0_), .ZN(n4702) );
  OR2_X1 U5429 ( .A1(n6052), .A2(n4702), .ZN(n4449) );
  OAI211_X1 U5430 ( .C1(n6060), .C2(n4444), .A(n4443), .B(n4449), .ZN(U2939)
         );
  NAND2_X1 U5431 ( .A1(n6071), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4446) );
  OAI211_X1 U5432 ( .C1(n6060), .C2(n4447), .A(n4446), .B(n4445), .ZN(U2934)
         );
  INV_X1 U5433 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5434 ( .A1(n6071), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4448) );
  INV_X1 U5435 ( .A(DATAI_2_), .ZN(n4496) );
  OR2_X1 U5436 ( .A1(n6052), .A2(n4496), .ZN(n4452) );
  OAI211_X1 U5437 ( .C1(n6060), .C2(n4678), .A(n4448), .B(n4452), .ZN(U2926)
         );
  NAND2_X1 U5438 ( .A1(n6071), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4450) );
  OAI211_X1 U5439 ( .C1(n6060), .C2(n4451), .A(n4450), .B(n4449), .ZN(U2924)
         );
  INV_X1 U5440 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U5441 ( .A1(n6071), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4453) );
  OAI211_X1 U5442 ( .C1(n6060), .C2(n4454), .A(n4453), .B(n4452), .ZN(U2941)
         );
  AOI22_X1 U5443 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4455) );
  OAI21_X1 U5444 ( .B1(n4447), .B2(n4686), .A(n4455), .ZN(U2897) );
  INV_X1 U5445 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U5446 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4456) );
  OAI21_X1 U5447 ( .B1(n4457), .B2(n4686), .A(n4456), .ZN(U2901) );
  AOI22_X1 U5448 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5449 ( .B1(n7002), .B2(n4686), .A(n4458), .ZN(U2899) );
  INV_X1 U5450 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6780) );
  AOI22_X1 U5451 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4459) );
  OAI21_X1 U5452 ( .B1(n6780), .B2(n4686), .A(n4459), .ZN(U2895) );
  INV_X1 U5453 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U5454 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4460) );
  OAI21_X1 U5455 ( .B1(n4461), .B2(n4686), .A(n4460), .ZN(U2894) );
  XNOR2_X1 U5456 ( .A(n4462), .B(n4463), .ZN(n4593) );
  NAND2_X1 U5457 ( .A1(n5580), .A2(REIP_REG_1__SCAN_IN), .ZN(n4589) );
  OAI21_X1 U5458 ( .B1(n6146), .B2(n4464), .A(n4589), .ZN(n4467) );
  NOR3_X1 U5459 ( .A1(n6151), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4465), 
        .ZN(n4466) );
  AOI211_X1 U5460 ( .C1(n6180), .C2(n4468), .A(n4467), .B(n4466), .ZN(n4469)
         );
  OAI21_X1 U5461 ( .B1(n4593), .B2(n5881), .A(n4469), .ZN(U3017) );
  INV_X1 U5462 ( .A(n4470), .ZN(n4471) );
  OAI21_X1 U5463 ( .B1(n4473), .B2(n4472), .A(n4471), .ZN(n6100) );
  INV_X1 U5464 ( .A(n5228), .ZN(n5509) );
  NAND2_X1 U5465 ( .A1(n4475), .A2(n4474), .ZN(n4476) );
  AND2_X1 U5466 ( .A1(n4505), .A2(n4476), .ZN(n6192) );
  AOI22_X1 U5467 ( .A1(n5512), .A2(n6192), .B1(n5511), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4477) );
  OAI21_X1 U5468 ( .B1(n6100), .B2(n5514), .A(n4477), .ZN(U2857) );
  NOR2_X1 U5469 ( .A1(n4478), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4480)
         );
  OR2_X1 U5470 ( .A1(n4480), .A2(n4479), .ZN(n5706) );
  NAND2_X1 U5471 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  NAND2_X1 U5472 ( .A1(n4484), .A2(n4483), .ZN(n5217) );
  OAI222_X1 U5473 ( .A1(n5706), .A2(n5507), .B1(n5505), .B2(n5212), .C1(n5217), 
        .C2(n5514), .ZN(U2859) );
  NAND2_X1 U5474 ( .A1(n6566), .A2(n4485), .ZN(n4488) );
  INV_X1 U5475 ( .A(n5171), .ZN(n4487) );
  OAI22_X1 U5476 ( .A1(n5910), .A2(n4488), .B1(n4487), .B2(n4486), .ZN(n4489)
         );
  AOI21_X1 U5477 ( .B1(n4491), .B2(n4490), .A(n4489), .ZN(n4492) );
  NAND2_X1 U5478 ( .A1(n4493), .A2(n5098), .ZN(n4494) );
  NAND2_X1 U5479 ( .A1(n5515), .A2(n4494), .ZN(n5831) );
  INV_X1 U5480 ( .A(n4494), .ZN(n4495) );
  NAND2_X1 U5481 ( .A1(n5515), .A2(n4495), .ZN(n5050) );
  OAI222_X1 U5482 ( .A1(n6100), .A2(n5831), .B1(n5050), .B2(n4496), .C1(n5515), 
        .C2(n4454), .ZN(U2889) );
  AOI21_X1 U5483 ( .B1(n4470), .B2(n4502), .A(n4497), .ZN(n4498) );
  OR2_X1 U5484 ( .A1(n4498), .A2(n4658), .ZN(n5470) );
  AND2_X1 U5485 ( .A1(n4507), .A2(n4499), .ZN(n4500) );
  NOR2_X1 U5486 ( .A1(n4652), .A2(n4500), .ZN(n6170) );
  AOI22_X1 U5487 ( .A1(n5512), .A2(n6170), .B1(n5511), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4501) );
  OAI21_X1 U5488 ( .B1(n5470), .B2(n5514), .A(n4501), .ZN(U2855) );
  INV_X1 U5489 ( .A(n4502), .ZN(n4503) );
  XNOR2_X1 U5490 ( .A(n4503), .B(n4470), .ZN(n6095) );
  INV_X1 U5491 ( .A(n6095), .ZN(n4701) );
  NAND2_X1 U5492 ( .A1(n4505), .A2(n4504), .ZN(n4506) );
  AND2_X1 U5493 ( .A1(n4507), .A2(n4506), .ZN(n6179) );
  AOI22_X1 U5494 ( .A1(n5512), .A2(n6179), .B1(n5511), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4508) );
  OAI21_X1 U5495 ( .B1(n4701), .B2(n5228), .A(n4508), .ZN(U2856) );
  XOR2_X1 U5496 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n4509), .Z(n5708) );
  NAND2_X1 U5497 ( .A1(n6178), .A2(REIP_REG_0__SCAN_IN), .ZN(n5705) );
  OAI21_X1 U5498 ( .B1(n5217), .B2(n5590), .A(n5705), .ZN(n4513) );
  INV_X1 U5499 ( .A(n6099), .ZN(n5610) );
  INV_X1 U5500 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4510) );
  AOI21_X1 U5501 ( .B1(n5610), .B2(n4511), .A(n4510), .ZN(n4512) );
  AOI211_X1 U5502 ( .C1(n3824), .C2(n5708), .A(n4513), .B(n4512), .ZN(n4514)
         );
  INV_X1 U5503 ( .A(n4514), .ZN(U2986) );
  INV_X1 U5504 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4516) );
  INV_X1 U5505 ( .A(DATAI_6_), .ZN(n4660) );
  NOR2_X1 U5506 ( .A1(n6052), .A2(n4660), .ZN(n4530) );
  AOI21_X1 U5507 ( .B1(n6072), .B2(EAX_REG_6__SCAN_IN), .A(n4530), .ZN(n4515)
         );
  OAI21_X1 U5508 ( .B1(n4551), .B2(n4516), .A(n4515), .ZN(U2945) );
  INV_X1 U5509 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n4518) );
  INV_X1 U5510 ( .A(DATAI_14_), .ZN(n6973) );
  NOR2_X1 U5511 ( .A1(n6052), .A2(n6973), .ZN(n4525) );
  AOI21_X1 U5512 ( .B1(n6072), .B2(EAX_REG_30__SCAN_IN), .A(n4525), .ZN(n4517)
         );
  OAI21_X1 U5513 ( .B1(n4551), .B2(n4518), .A(n4517), .ZN(U2938) );
  INV_X1 U5514 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4520) );
  INV_X1 U5515 ( .A(DATAI_7_), .ZN(n4768) );
  NOR2_X1 U5516 ( .A1(n6052), .A2(n4768), .ZN(n4538) );
  AOI21_X1 U5517 ( .B1(n6072), .B2(EAX_REG_7__SCAN_IN), .A(n4538), .ZN(n4519)
         );
  OAI21_X1 U5518 ( .B1(n4551), .B2(n4520), .A(n4519), .ZN(U2946) );
  INV_X1 U5519 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4522) );
  INV_X1 U5520 ( .A(DATAI_1_), .ZN(n4698) );
  NOR2_X1 U5521 ( .A1(n6052), .A2(n4698), .ZN(n4547) );
  AOI21_X1 U5522 ( .B1(n6072), .B2(EAX_REG_1__SCAN_IN), .A(n4547), .ZN(n4521)
         );
  OAI21_X1 U5523 ( .B1(n4551), .B2(n4522), .A(n4521), .ZN(U2940) );
  INV_X1 U5524 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4524) );
  INV_X1 U5525 ( .A(DATAI_4_), .ZN(n4690) );
  NOR2_X1 U5526 ( .A1(n6052), .A2(n4690), .ZN(n4541) );
  AOI21_X1 U5527 ( .B1(n6072), .B2(EAX_REG_4__SCAN_IN), .A(n4541), .ZN(n4523)
         );
  OAI21_X1 U5528 ( .B1(n4551), .B2(n4524), .A(n4523), .ZN(U2943) );
  INV_X1 U5529 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n4527) );
  AOI21_X1 U5530 ( .B1(n6072), .B2(EAX_REG_14__SCAN_IN), .A(n4525), .ZN(n4526)
         );
  OAI21_X1 U5531 ( .B1(n4551), .B2(n4527), .A(n4526), .ZN(U2953) );
  INV_X1 U5532 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4529) );
  INV_X1 U5533 ( .A(DATAI_5_), .ZN(n4688) );
  NOR2_X1 U5534 ( .A1(n6052), .A2(n4688), .ZN(n4544) );
  AOI21_X1 U5535 ( .B1(n6072), .B2(EAX_REG_21__SCAN_IN), .A(n4544), .ZN(n4528)
         );
  OAI21_X1 U5536 ( .B1(n4551), .B2(n4529), .A(n4528), .ZN(U2929) );
  INV_X1 U5537 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4532) );
  AOI21_X1 U5538 ( .B1(n6072), .B2(EAX_REG_22__SCAN_IN), .A(n4530), .ZN(n4531)
         );
  OAI21_X1 U5539 ( .B1(n4551), .B2(n4532), .A(n4531), .ZN(U2930) );
  INV_X1 U5540 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4534) );
  INV_X1 U5541 ( .A(DATAI_3_), .ZN(n4700) );
  NOR2_X1 U5542 ( .A1(n6052), .A2(n4700), .ZN(n4535) );
  AOI21_X1 U5543 ( .B1(n6072), .B2(EAX_REG_3__SCAN_IN), .A(n4535), .ZN(n4533)
         );
  OAI21_X1 U5544 ( .B1(n4551), .B2(n4534), .A(n4533), .ZN(U2942) );
  INV_X1 U5545 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4537) );
  AOI21_X1 U5546 ( .B1(n6072), .B2(EAX_REG_19__SCAN_IN), .A(n4535), .ZN(n4536)
         );
  OAI21_X1 U5547 ( .B1(n4551), .B2(n4537), .A(n4536), .ZN(U2927) );
  INV_X1 U5548 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4540) );
  AOI21_X1 U5549 ( .B1(n6072), .B2(EAX_REG_23__SCAN_IN), .A(n4538), .ZN(n4539)
         );
  OAI21_X1 U5550 ( .B1(n4551), .B2(n4540), .A(n4539), .ZN(U2931) );
  INV_X1 U5551 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4543) );
  AOI21_X1 U5552 ( .B1(n6072), .B2(EAX_REG_20__SCAN_IN), .A(n4541), .ZN(n4542)
         );
  OAI21_X1 U5553 ( .B1(n4551), .B2(n4543), .A(n4542), .ZN(U2928) );
  INV_X1 U5554 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4546) );
  AOI21_X1 U5555 ( .B1(n6072), .B2(EAX_REG_5__SCAN_IN), .A(n4544), .ZN(n4545)
         );
  OAI21_X1 U5556 ( .B1(n4551), .B2(n4546), .A(n4545), .ZN(U2944) );
  INV_X1 U5557 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4549) );
  AOI21_X1 U5558 ( .B1(n6072), .B2(EAX_REG_17__SCAN_IN), .A(n4547), .ZN(n4548)
         );
  OAI21_X1 U5559 ( .B1(n4551), .B2(n4549), .A(n4548), .ZN(U2925) );
  INV_X1 U5560 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4552) );
  INV_X1 U5561 ( .A(DATAI_15_), .ZN(n4997) );
  INV_X1 U5562 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4550) );
  OAI222_X1 U5563 ( .A1(n4552), .A2(n4551), .B1(n6052), .B2(n4997), .C1(n4550), 
        .C2(n6060), .ZN(U2954) );
  MUX2_X1 U5564 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4553), .S(n6532), 
        .Z(n6538) );
  INV_X1 U5565 ( .A(n6527), .ZN(n4570) );
  NAND2_X1 U5566 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4555) );
  INV_X1 U5567 ( .A(n4555), .ZN(n4556) );
  MUX2_X1 U5568 ( .A(n4556), .B(n4555), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4561) );
  INV_X1 U5569 ( .A(n4557), .ZN(n4560) );
  AOI21_X1 U5570 ( .B1(n4376), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4558) );
  NOR2_X1 U5571 ( .A1(n4559), .A2(n4558), .ZN(n5720) );
  AOI22_X1 U5572 ( .A1(n6529), .A2(n4561), .B1(n4560), .B2(n5720), .ZN(n4569)
         );
  INV_X1 U5573 ( .A(n4562), .ZN(n4566) );
  INV_X1 U5574 ( .A(n4563), .ZN(n4564) );
  MUX2_X1 U5575 ( .A(n4564), .B(n3935), .S(n4376), .Z(n4565) );
  NAND3_X1 U5576 ( .A1(n4567), .A2(n4566), .A3(n4565), .ZN(n4568) );
  OAI211_X1 U5577 ( .C1(n6325), .C2(n4570), .A(n4569), .B(n4568), .ZN(n5719)
         );
  MUX2_X1 U5578 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5719), .S(n6532), 
        .Z(n6540) );
  NAND3_X1 U5579 ( .A1(n6538), .A2(n6540), .A3(n6557), .ZN(n4573) );
  NAND2_X1 U5580 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5925), .ZN(n4578) );
  INV_X1 U5581 ( .A(n4578), .ZN(n4571) );
  NAND2_X1 U5582 ( .A1(n4562), .A2(n4571), .ZN(n4572) );
  NAND2_X1 U5583 ( .A1(n4573), .A2(n4572), .ZN(n6549) );
  NAND2_X1 U5584 ( .A1(n6549), .A2(n4574), .ZN(n4596) );
  INV_X1 U5585 ( .A(n5725), .ZN(n6449) );
  OR2_X1 U5586 ( .A1(n4575), .A2(n6449), .ZN(n4576) );
  XNOR2_X1 U5587 ( .A(n4576), .B(n4577), .ZN(n5909) );
  OAI22_X1 U5588 ( .A1(n6532), .A2(n4577), .B1(n5910), .B2(n5909), .ZN(n4580)
         );
  NOR2_X1 U5589 ( .A1(n4577), .A2(n4578), .ZN(n4579) );
  AOI21_X1 U5590 ( .B1(n4580), .B2(n6557), .A(n4579), .ZN(n6547) );
  AND2_X1 U5591 ( .A1(n6547), .A2(n5925), .ZN(n4581) );
  NAND2_X1 U5592 ( .A1(n4596), .A2(n4581), .ZN(n4583) );
  INV_X1 U5593 ( .A(n6652), .ZN(n4582) );
  NOR2_X1 U5594 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6679) );
  OAI21_X1 U5595 ( .B1(n6679), .B2(n4594), .A(n6558), .ZN(n4603) );
  NAND2_X1 U5596 ( .A1(n6972), .A2(n4603), .ZN(n6326) );
  AOI21_X1 U5597 ( .B1(n4583), .B2(n4582), .A(n4820), .ZN(n5717) );
  NAND2_X1 U5598 ( .A1(n4585), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U5599 ( .A(n6210), .B(n6203), .ZN(n4586) );
  NAND2_X1 U5600 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6942), .ZN(n4661) );
  AOI22_X1 U5601 ( .A1(n4586), .A2(n6447), .B1(n5178), .B2(n4661), .ZN(n4588)
         );
  NAND2_X1 U5602 ( .A1(n5717), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4587) );
  OAI21_X1 U5603 ( .B1(n5717), .B2(n4588), .A(n4587), .ZN(U3463) );
  NAND2_X1 U5604 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4590)
         );
  OAI211_X1 U5605 ( .C1(n6110), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4590), 
        .B(n4589), .ZN(n4591) );
  AOI21_X1 U5606 ( .B1(n6105), .B2(n6001), .A(n4591), .ZN(n4592) );
  OAI21_X1 U5607 ( .B1(n4593), .B2(n5924), .A(n4592), .ZN(U2985) );
  INV_X1 U5608 ( .A(n5717), .ZN(n6202) );
  AND2_X1 U5609 ( .A1(n6547), .A2(n4594), .ZN(n4595) );
  NAND2_X1 U5610 ( .A1(n4596), .A2(n4595), .ZN(n6565) );
  INV_X1 U5611 ( .A(n6565), .ZN(n4598) );
  INV_X1 U5612 ( .A(n6528), .ZN(n5001) );
  INV_X1 U5613 ( .A(n4661), .ZN(n5716) );
  OAI22_X1 U5614 ( .A1(n4857), .A2(n6401), .B1(n5001), .B2(n5716), .ZN(n4597)
         );
  OAI21_X1 U5615 ( .B1(n4598), .B2(n4597), .A(n6202), .ZN(n4599) );
  OAI21_X1 U5616 ( .B1(n6202), .B2(n6355), .A(n4599), .ZN(U3465) );
  NAND2_X1 U5617 ( .A1(n6210), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5618 ( .A1(n4585), .A2(n4857), .ZN(n4906) );
  OR2_X1 U5619 ( .A1(n4662), .A2(n4906), .ZN(n4944) );
  INV_X1 U5620 ( .A(DATAI_25_), .ZN(n4600) );
  NOR2_X1 U5621 ( .A1(n5590), .A2(n4600), .ZN(n6367) );
  INV_X1 U5622 ( .A(n6367), .ZN(n6466) );
  INV_X1 U5623 ( .A(DATAI_17_), .ZN(n4601) );
  NOR2_X1 U5624 ( .A1(n5590), .A2(n4601), .ZN(n6414) );
  NAND2_X1 U5625 ( .A1(n4585), .A2(n6323), .ZN(n6396) );
  OR2_X1 U5626 ( .A1(n4662), .A2(n6396), .ZN(n4705) );
  NAND2_X1 U5627 ( .A1(DATAI_1_), .A2(n4820), .ZN(n6295) );
  NAND2_X1 U5628 ( .A1(n5989), .A2(n6528), .ZN(n6358) );
  NAND2_X1 U5629 ( .A1(n5178), .A2(n6004), .ZN(n4953) );
  OR2_X1 U5630 ( .A1(n6358), .A2(n4953), .ZN(n4602) );
  NAND2_X1 U5631 ( .A1(n4602), .A2(n4645), .ZN(n4608) );
  AOI22_X1 U5632 ( .A1(n4608), .A2(n6324), .B1(n4947), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4646) );
  INV_X1 U5633 ( .A(n6653), .ZN(n4604) );
  AND2_X1 U5634 ( .A1(n4604), .A2(n4603), .ZN(n4644) );
  NAND2_X1 U5635 ( .A1(n4644), .A2(n4605), .ZN(n4968) );
  OAI22_X1 U5636 ( .A1(n6295), .A2(n4646), .B1(n4645), .B2(n4968), .ZN(n4606)
         );
  AOI21_X1 U5637 ( .B1(n6414), .B2(n4735), .A(n4606), .ZN(n4613) );
  AOI21_X1 U5638 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6355), .A(n6326), .ZN(
        n6406) );
  INV_X1 U5639 ( .A(n4662), .ZN(n4607) );
  AOI21_X1 U5640 ( .B1(n4607), .B2(n4585), .A(n5590), .ZN(n4610) );
  AND2_X1 U5641 ( .A1(n6447), .A2(n6353), .ZN(n6248) );
  INV_X1 U5642 ( .A(n4608), .ZN(n4609) );
  OAI21_X1 U5643 ( .B1(n4610), .B2(n6248), .A(n4609), .ZN(n4611) );
  OAI211_X1 U5644 ( .C1(n4947), .C2(n6447), .A(n6406), .B(n4611), .ZN(n4648)
         );
  NAND2_X1 U5645 ( .A1(n4648), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4612)
         );
  OAI211_X1 U5646 ( .C1(n4944), .C2(n6466), .A(n4613), .B(n4612), .ZN(U3141)
         );
  NAND2_X1 U5647 ( .A1(n6105), .A2(DATAI_29_), .ZN(n6503) );
  INV_X1 U5648 ( .A(DATAI_21_), .ZN(n4614) );
  NOR2_X1 U5649 ( .A1(n5590), .A2(n4614), .ZN(n6427) );
  NAND2_X1 U5650 ( .A1(DATAI_5_), .A2(n4820), .ZN(n6307) );
  NAND2_X1 U5651 ( .A1(n4644), .A2(n4615), .ZN(n4949) );
  OAI22_X1 U5652 ( .A1(n6307), .A2(n4646), .B1(n4645), .B2(n4949), .ZN(n4616)
         );
  AOI21_X1 U5653 ( .B1(n6427), .B2(n4735), .A(n4616), .ZN(n4618) );
  NAND2_X1 U5654 ( .A1(n4648), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4617)
         );
  OAI211_X1 U5655 ( .C1(n4944), .C2(n6503), .A(n4618), .B(n4617), .ZN(U3145)
         );
  INV_X1 U5656 ( .A(DATAI_26_), .ZN(n4619) );
  NOR2_X1 U5657 ( .A1(n5590), .A2(n4619), .ZN(n6370) );
  INV_X1 U5658 ( .A(n6370), .ZN(n6479) );
  INV_X1 U5659 ( .A(DATAI_18_), .ZN(n4620) );
  NOR2_X1 U5660 ( .A1(n5590), .A2(n4620), .ZN(n6417) );
  NAND2_X1 U5661 ( .A1(DATAI_2_), .A2(n4820), .ZN(n6298) );
  NAND2_X1 U5662 ( .A1(n4644), .A2(n4621), .ZN(n4972) );
  OAI22_X1 U5663 ( .A1(n6298), .A2(n4646), .B1(n4645), .B2(n4972), .ZN(n4622)
         );
  AOI21_X1 U5664 ( .B1(n6417), .B2(n4735), .A(n4622), .ZN(n4624) );
  NAND2_X1 U5665 ( .A1(n4648), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4623)
         );
  OAI211_X1 U5666 ( .C1(n4944), .C2(n6479), .A(n4624), .B(n4623), .ZN(U3142)
         );
  INV_X1 U5667 ( .A(DATAI_30_), .ZN(n6781) );
  NOR2_X1 U5668 ( .A1(n5590), .A2(n6781), .ZN(n6383) );
  INV_X1 U5669 ( .A(n6383), .ZN(n6511) );
  INV_X1 U5670 ( .A(DATAI_22_), .ZN(n4625) );
  NOR2_X1 U5671 ( .A1(n5590), .A2(n4625), .ZN(n6430) );
  NAND2_X1 U5672 ( .A1(DATAI_6_), .A2(n4820), .ZN(n6310) );
  NAND2_X1 U5673 ( .A1(n4644), .A2(n4626), .ZN(n4960) );
  OAI22_X1 U5674 ( .A1(n6310), .A2(n4646), .B1(n4645), .B2(n4960), .ZN(n4627)
         );
  AOI21_X1 U5675 ( .B1(n6430), .B2(n4735), .A(n4627), .ZN(n4629) );
  NAND2_X1 U5676 ( .A1(n4648), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4628)
         );
  OAI211_X1 U5677 ( .C1(n4944), .C2(n6511), .A(n4629), .B(n4628), .ZN(U3146)
         );
  NAND2_X1 U5678 ( .A1(n6105), .A2(DATAI_24_), .ZN(n6458) );
  INV_X1 U5679 ( .A(DATAI_16_), .ZN(n4630) );
  NOR2_X1 U5680 ( .A1(n5590), .A2(n4630), .ZN(n6364) );
  NAND2_X1 U5681 ( .A1(DATAI_0_), .A2(n4820), .ZN(n6292) );
  NAND2_X1 U5682 ( .A1(n4644), .A2(n5122), .ZN(n4964) );
  OAI22_X1 U5683 ( .A1(n6292), .A2(n4646), .B1(n4645), .B2(n4964), .ZN(n4631)
         );
  AOI21_X1 U5684 ( .B1(n6364), .B2(n4735), .A(n4631), .ZN(n4633) );
  NAND2_X1 U5685 ( .A1(n4648), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4632)
         );
  OAI211_X1 U5686 ( .C1(n4944), .C2(n6458), .A(n4633), .B(n4632), .ZN(U3140)
         );
  NAND2_X1 U5687 ( .A1(n6105), .A2(DATAI_27_), .ZN(n6487) );
  INV_X1 U5688 ( .A(DATAI_19_), .ZN(n4634) );
  NOR2_X1 U5689 ( .A1(n5590), .A2(n4634), .ZN(n6373) );
  NAND2_X1 U5690 ( .A1(DATAI_3_), .A2(n4820), .ZN(n6301) );
  NAND2_X1 U5691 ( .A1(n4644), .A2(n3663), .ZN(n4980) );
  OAI22_X1 U5692 ( .A1(n6301), .A2(n4646), .B1(n4645), .B2(n4980), .ZN(n4635)
         );
  AOI21_X1 U5693 ( .B1(n6373), .B2(n4735), .A(n4635), .ZN(n4637) );
  NAND2_X1 U5694 ( .A1(n4648), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4636)
         );
  OAI211_X1 U5695 ( .C1(n4944), .C2(n6487), .A(n4637), .B(n4636), .ZN(U3143)
         );
  INV_X1 U5696 ( .A(DATAI_31_), .ZN(n6775) );
  NOR2_X1 U5697 ( .A1(n5590), .A2(n6775), .ZN(n6388) );
  INV_X1 U5698 ( .A(n6388), .ZN(n6524) );
  INV_X1 U5699 ( .A(DATAI_23_), .ZN(n4638) );
  NOR2_X1 U5700 ( .A1(n5590), .A2(n4638), .ZN(n6433) );
  NAND2_X1 U5701 ( .A1(DATAI_7_), .A2(n4820), .ZN(n6317) );
  NAND2_X1 U5702 ( .A1(n4644), .A2(n5098), .ZN(n4985) );
  OAI22_X1 U5703 ( .A1(n6317), .A2(n4646), .B1(n4645), .B2(n4985), .ZN(n4639)
         );
  AOI21_X1 U5704 ( .B1(n6433), .B2(n4735), .A(n4639), .ZN(n4641) );
  NAND2_X1 U5705 ( .A1(n4648), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4640)
         );
  OAI211_X1 U5706 ( .C1(n4944), .C2(n6524), .A(n4641), .B(n4640), .ZN(U3147)
         );
  NAND2_X1 U5707 ( .A1(n6105), .A2(DATAI_28_), .ZN(n6495) );
  INV_X1 U5708 ( .A(DATAI_20_), .ZN(n4642) );
  NOR2_X1 U5709 ( .A1(n5590), .A2(n4642), .ZN(n6424) );
  NAND2_X1 U5710 ( .A1(DATAI_4_), .A2(n4820), .ZN(n6304) );
  NAND2_X1 U5711 ( .A1(n4644), .A2(n4643), .ZN(n4976) );
  OAI22_X1 U5712 ( .A1(n6304), .A2(n4646), .B1(n4645), .B2(n4976), .ZN(n4647)
         );
  AOI21_X1 U5713 ( .B1(n6424), .B2(n4735), .A(n4647), .ZN(n4650) );
  NAND2_X1 U5714 ( .A1(n4648), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4649)
         );
  OAI211_X1 U5715 ( .C1(n4944), .C2(n6495), .A(n4650), .B(n4649), .ZN(U3144)
         );
  OAI21_X1 U5716 ( .B1(n4652), .B2(n4651), .A(n4671), .ZN(n6159) );
  INV_X1 U5717 ( .A(n4657), .ZN(n4653) );
  XNOR2_X1 U5718 ( .A(n4653), .B(n4658), .ZN(n6087) );
  INV_X1 U5719 ( .A(n6087), .ZN(n4689) );
  INV_X1 U5720 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4654) );
  OAI222_X1 U5721 ( .A1(n6159), .A2(n5507), .B1(n5228), .B2(n4689), .C1(n4654), 
        .C2(n5505), .ZN(U2854) );
  AOI21_X1 U5722 ( .B1(n4658), .B2(n4657), .A(n4656), .ZN(n4659) );
  OR2_X1 U5723 ( .A1(n4770), .A2(n4659), .ZN(n5160) );
  OAI222_X1 U5724 ( .A1(n5160), .A2(n5831), .B1(n5050), .B2(n4660), .C1(n5515), 
        .C2(n3954), .ZN(U2885) );
  NAND2_X1 U5725 ( .A1(n5989), .A2(n4661), .ZN(n4667) );
  INV_X1 U5726 ( .A(n6210), .ZN(n6204) );
  NAND2_X1 U5727 ( .A1(n6204), .A2(n3934), .ZN(n6400) );
  NAND2_X1 U5728 ( .A1(n6210), .A2(n4664), .ZN(n6289) );
  OR2_X1 U5729 ( .A1(n6289), .A2(n6203), .ZN(n6281) );
  NAND3_X1 U5730 ( .A1(n4744), .A2(n6400), .A3(n6281), .ZN(n4665) );
  NOR2_X1 U5731 ( .A1(n5717), .A2(n6206), .ZN(n4666) );
  NAND2_X1 U5732 ( .A1(n4667), .A2(n4666), .ZN(n4668) );
  AOI21_X1 U5733 ( .B1(n3934), .B2(n6248), .A(n4668), .ZN(n4669) );
  AOI21_X1 U5734 ( .B1(n5717), .B2(n6397), .A(n4669), .ZN(U3462) );
  NAND2_X1 U5735 ( .A1(n4671), .A2(n4670), .ZN(n4672) );
  NAND2_X1 U5736 ( .A1(n4801), .A2(n4672), .ZN(n6142) );
  INV_X1 U5737 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4673) );
  OAI222_X1 U5738 ( .A1(n6142), .A2(n5507), .B1(n5505), .B2(n4673), .C1(n5514), 
        .C2(n5160), .ZN(U2853) );
  INV_X1 U5739 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U5740 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4674) );
  OAI21_X1 U5741 ( .B1(n6743), .B2(n4686), .A(n4674), .ZN(U2893) );
  INV_X1 U5742 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5743 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4675) );
  OAI21_X1 U5744 ( .B1(n4676), .B2(n4686), .A(n4675), .ZN(U2904) );
  AOI22_X1 U5745 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4677) );
  OAI21_X1 U5746 ( .B1(n4678), .B2(n4686), .A(n4677), .ZN(U2905) );
  INV_X1 U5747 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5748 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4679) );
  OAI21_X1 U5749 ( .B1(n4680), .B2(n4686), .A(n4679), .ZN(U2906) );
  INV_X1 U5750 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5751 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4681) );
  OAI21_X1 U5752 ( .B1(n4682), .B2(n4686), .A(n4681), .ZN(U2903) );
  INV_X1 U5753 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5754 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4683) );
  OAI21_X1 U5755 ( .B1(n4684), .B2(n4686), .A(n4683), .ZN(U2896) );
  INV_X1 U5756 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5757 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4685) );
  OAI21_X1 U5758 ( .B1(n4687), .B2(n4686), .A(n4685), .ZN(U2902) );
  OAI222_X1 U5759 ( .A1(n5831), .A2(n4689), .B1(n5050), .B2(n4688), .C1(n5515), 
        .C2(n3948), .ZN(U2886) );
  INV_X1 U5760 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6043) );
  OAI222_X1 U5761 ( .A1(n5831), .A2(n5470), .B1(n5515), .B2(n6043), .C1(n5050), 
        .C2(n4690), .ZN(U2887) );
  CLKBUF_X1 U5762 ( .A(n4692), .Z(n4693) );
  OAI21_X1 U5763 ( .B1(n4694), .B2(n4691), .A(n4693), .ZN(n6171) );
  NAND2_X1 U5764 ( .A1(n5580), .A2(REIP_REG_4__SCAN_IN), .ZN(n6168) );
  OAI21_X1 U5765 ( .B1(n5610), .B2(n3900), .A(n6168), .ZN(n4696) );
  NOR2_X1 U5766 ( .A1(n5470), .A2(n5590), .ZN(n4695) );
  AOI211_X1 U5767 ( .C1(n5622), .C2(n5458), .A(n4696), .B(n4695), .ZN(n4697)
         );
  OAI21_X1 U5768 ( .B1(n5924), .B2(n6171), .A(n4697), .ZN(U2982) );
  INV_X1 U5769 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6048) );
  OAI222_X1 U5770 ( .A1(n4699), .A2(n5831), .B1(n5050), .B2(n4698), .C1(n5515), 
        .C2(n6048), .ZN(U2890) );
  INV_X1 U5771 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6045) );
  OAI222_X1 U5772 ( .A1(n4701), .A2(n5831), .B1(n5050), .B2(n4700), .C1(n5515), 
        .C2(n6045), .ZN(U2888) );
  OAI222_X1 U5773 ( .A1(n5217), .A2(n5831), .B1(n5050), .B2(n4702), .C1(n5515), 
        .C2(n4444), .ZN(U2891) );
  NOR3_X1 U5774 ( .A1(n3934), .A2(n6210), .A3(n4585), .ZN(n4905) );
  NAND2_X1 U5775 ( .A1(n4905), .A2(n4857), .ZN(n5004) );
  INV_X1 U5776 ( .A(n6414), .ZN(n6468) );
  NAND3_X1 U5777 ( .A1(n6397), .A2(n6539), .A3(n6534), .ZN(n5006) );
  OR2_X1 U5778 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5006), .ZN(n4732)
         );
  NOR2_X1 U5779 ( .A1(n4708), .A2(n6568), .ZN(n6327) );
  INV_X1 U5780 ( .A(n4703), .ZN(n6321) );
  INV_X1 U5781 ( .A(n6320), .ZN(n4823) );
  NOR2_X1 U5782 ( .A1(n6321), .A2(n4823), .ZN(n6240) );
  OAI21_X1 U5783 ( .B1(n6240), .B2(n6568), .A(n4820), .ZN(n6244) );
  AOI211_X1 U5784 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4732), .A(n6327), .B(
        n6244), .ZN(n4707) );
  INV_X1 U5785 ( .A(n6248), .ZN(n4908) );
  OAI21_X1 U5786 ( .B1(n4905), .B2(n6401), .A(n4908), .ZN(n5007) );
  OR2_X1 U5787 ( .A1(n5178), .A2(n6004), .ZN(n6357) );
  INV_X1 U5788 ( .A(n6357), .ZN(n4704) );
  NAND2_X1 U5789 ( .A1(n4704), .A2(n6325), .ZN(n5002) );
  OAI211_X1 U5790 ( .C1(n6248), .C2(n4705), .A(n5007), .B(n5002), .ZN(n4706)
         );
  NAND2_X1 U5791 ( .A1(n4707), .A2(n4706), .ZN(n4731) );
  NAND2_X1 U5792 ( .A1(n4731), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4712) );
  INV_X1 U5793 ( .A(n5002), .ZN(n4709) );
  AND2_X1 U5794 ( .A1(n4708), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6442) );
  AOI22_X1 U5795 ( .A1(n4709), .A2(n6324), .B1(n6442), .B2(n6240), .ZN(n4733)
         );
  OAI22_X1 U5796 ( .A1(n6295), .A2(n4733), .B1(n4968), .B2(n4732), .ZN(n4710)
         );
  AOI21_X1 U5797 ( .B1(n6367), .B2(n4735), .A(n4710), .ZN(n4711) );
  OAI211_X1 U5798 ( .C1(n5004), .C2(n6468), .A(n4712), .B(n4711), .ZN(U3021)
         );
  INV_X1 U5799 ( .A(n6373), .ZN(n6482) );
  NAND2_X1 U5800 ( .A1(n4731), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4715) );
  INV_X1 U5801 ( .A(n6487), .ZN(n6420) );
  OAI22_X1 U5802 ( .A1(n6301), .A2(n4733), .B1(n4980), .B2(n4732), .ZN(n4713)
         );
  AOI21_X1 U5803 ( .B1(n6420), .B2(n4735), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5804 ( .C1(n5004), .C2(n6482), .A(n4715), .B(n4714), .ZN(U3023)
         );
  INV_X1 U5805 ( .A(n6433), .ZN(n6517) );
  NAND2_X1 U5806 ( .A1(n4731), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4718) );
  OAI22_X1 U5807 ( .A1(n6317), .A2(n4733), .B1(n4985), .B2(n4732), .ZN(n4716)
         );
  AOI21_X1 U5808 ( .B1(n6388), .B2(n4735), .A(n4716), .ZN(n4717) );
  OAI211_X1 U5809 ( .C1(n5004), .C2(n6517), .A(n4718), .B(n4717), .ZN(U3027)
         );
  INV_X1 U5810 ( .A(n6417), .ZN(n6474) );
  NAND2_X1 U5811 ( .A1(n4731), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4721) );
  OAI22_X1 U5812 ( .A1(n6298), .A2(n4733), .B1(n4972), .B2(n4732), .ZN(n4719)
         );
  AOI21_X1 U5813 ( .B1(n6370), .B2(n4735), .A(n4719), .ZN(n4720) );
  OAI211_X1 U5814 ( .C1(n5004), .C2(n6474), .A(n4721), .B(n4720), .ZN(U3022)
         );
  INV_X1 U5815 ( .A(n6364), .ZN(n6460) );
  NAND2_X1 U5816 ( .A1(n4731), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4724) );
  INV_X1 U5817 ( .A(n6458), .ZN(n6399) );
  OAI22_X1 U5818 ( .A1(n6292), .A2(n4733), .B1(n4964), .B2(n4732), .ZN(n4722)
         );
  AOI21_X1 U5819 ( .B1(n6399), .B2(n4735), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5820 ( .C1(n5004), .C2(n6460), .A(n4724), .B(n4723), .ZN(U3020)
         );
  INV_X1 U5821 ( .A(n6430), .ZN(n6506) );
  NAND2_X1 U5822 ( .A1(n4731), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4727) );
  OAI22_X1 U5823 ( .A1(n6310), .A2(n4733), .B1(n4960), .B2(n4732), .ZN(n4725)
         );
  AOI21_X1 U5824 ( .B1(n6383), .B2(n4735), .A(n4725), .ZN(n4726) );
  OAI211_X1 U5825 ( .C1(n5004), .C2(n6506), .A(n4727), .B(n4726), .ZN(U3026)
         );
  INV_X1 U5826 ( .A(n6424), .ZN(n6490) );
  NAND2_X1 U5827 ( .A1(n4731), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4730) );
  INV_X1 U5828 ( .A(n6495), .ZN(n6377) );
  OAI22_X1 U5829 ( .A1(n6304), .A2(n4733), .B1(n4976), .B2(n4732), .ZN(n4728)
         );
  AOI21_X1 U5830 ( .B1(n6377), .B2(n4735), .A(n4728), .ZN(n4729) );
  OAI211_X1 U5831 ( .C1(n5004), .C2(n6490), .A(n4730), .B(n4729), .ZN(U3024)
         );
  INV_X1 U5832 ( .A(n6427), .ZN(n6498) );
  NAND2_X1 U5833 ( .A1(n4731), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4737) );
  INV_X1 U5834 ( .A(n6503), .ZN(n6380) );
  OAI22_X1 U5835 ( .A1(n6307), .A2(n4733), .B1(n4949), .B2(n4732), .ZN(n4734)
         );
  AOI21_X1 U5836 ( .B1(n6380), .B2(n4735), .A(n4734), .ZN(n4736) );
  OAI211_X1 U5837 ( .C1(n5004), .C2(n6498), .A(n4737), .B(n4736), .ZN(U3025)
         );
  NAND2_X1 U5838 ( .A1(n4771), .A2(n4770), .ZN(n4798) );
  OR2_X1 U5839 ( .A1(n4771), .A2(n4770), .ZN(n4738) );
  AND2_X1 U5840 ( .A1(n4798), .A2(n4738), .ZN(n6079) );
  INV_X1 U5841 ( .A(n6079), .ZN(n4769) );
  XNOR2_X1 U5842 ( .A(n4801), .B(n4803), .ZN(n6136) );
  AOI22_X1 U5843 ( .A1(n5512), .A2(n6136), .B1(EBX_REG_7__SCAN_IN), .B2(n5511), 
        .ZN(n4739) );
  OAI21_X1 U5844 ( .B1(n4769), .B2(n5228), .A(n4739), .ZN(U2852) );
  NAND3_X1 U5845 ( .A1(n6534), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6441) );
  INV_X1 U5846 ( .A(n6441), .ZN(n4743) );
  INV_X1 U5847 ( .A(n6358), .ZN(n4741) );
  INV_X1 U5848 ( .A(n6004), .ZN(n5715) );
  NAND2_X1 U5849 ( .A1(n5178), .A2(n5715), .ZN(n6454) );
  INV_X1 U5850 ( .A(n6454), .ZN(n4740) );
  NOR2_X1 U5851 ( .A1(n6355), .A2(n6441), .ZN(n4765) );
  AOI21_X1 U5852 ( .B1(n4741), .B2(n4740), .A(n4765), .ZN(n4746) );
  NAND3_X1 U5853 ( .A1(n6324), .A2(n4746), .A3(n4744), .ZN(n4742) );
  OAI211_X1 U5854 ( .C1(n6447), .C2(n4743), .A(n6406), .B(n4742), .ZN(n4763)
         );
  INV_X1 U5855 ( .A(n6298), .ZN(n6473) );
  NAND2_X1 U5856 ( .A1(n6447), .A2(n4744), .ZN(n4745) );
  OAI22_X1 U5857 ( .A1(n4746), .A2(n4745), .B1(n6568), .B2(n6441), .ZN(n4762)
         );
  AOI22_X1 U5858 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4763), .B1(n6473), 
        .B2(n4762), .ZN(n4749) );
  INV_X1 U5859 ( .A(n4972), .ZN(n6472) );
  AOI22_X1 U5860 ( .A1(n6472), .A2(n4765), .B1(n4764), .B2(n6370), .ZN(n4748)
         );
  OAI211_X1 U5861 ( .C1(n6474), .C2(n4992), .A(n4749), .B(n4748), .ZN(U3126)
         );
  INV_X1 U5862 ( .A(n6304), .ZN(n6489) );
  AOI22_X1 U5863 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4763), .B1(n6489), 
        .B2(n4762), .ZN(n4751) );
  INV_X1 U5864 ( .A(n4976), .ZN(n6488) );
  AOI22_X1 U5865 ( .A1(n6488), .A2(n4765), .B1(n4764), .B2(n6377), .ZN(n4750)
         );
  OAI211_X1 U5866 ( .C1(n6490), .C2(n4992), .A(n4751), .B(n4750), .ZN(U3128)
         );
  INV_X1 U5867 ( .A(n6292), .ZN(n6457) );
  AOI22_X1 U5868 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4763), .B1(n6457), 
        .B2(n4762), .ZN(n4753) );
  INV_X1 U5869 ( .A(n4964), .ZN(n6456) );
  AOI22_X1 U5870 ( .A1(n6456), .A2(n4765), .B1(n4764), .B2(n6399), .ZN(n4752)
         );
  OAI211_X1 U5871 ( .C1(n6460), .C2(n4992), .A(n4753), .B(n4752), .ZN(U3124)
         );
  INV_X1 U5872 ( .A(n6295), .ZN(n6465) );
  AOI22_X1 U5873 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4763), .B1(n6465), 
        .B2(n4762), .ZN(n4755) );
  INV_X1 U5874 ( .A(n4968), .ZN(n6464) );
  AOI22_X1 U5875 ( .A1(n6464), .A2(n4765), .B1(n4764), .B2(n6367), .ZN(n4754)
         );
  OAI211_X1 U5876 ( .C1(n6468), .C2(n4992), .A(n4755), .B(n4754), .ZN(U3125)
         );
  INV_X1 U5877 ( .A(n6307), .ZN(n6497) );
  AOI22_X1 U5878 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4763), .B1(n6497), 
        .B2(n4762), .ZN(n4757) );
  INV_X1 U5879 ( .A(n4949), .ZN(n6496) );
  AOI22_X1 U5880 ( .A1(n6496), .A2(n4765), .B1(n4764), .B2(n6380), .ZN(n4756)
         );
  OAI211_X1 U5881 ( .C1(n6498), .C2(n4992), .A(n4757), .B(n4756), .ZN(U3129)
         );
  INV_X1 U5882 ( .A(n6317), .ZN(n6515) );
  AOI22_X1 U5883 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4763), .B1(n6515), 
        .B2(n4762), .ZN(n4759) );
  INV_X1 U5884 ( .A(n4985), .ZN(n6513) );
  AOI22_X1 U5885 ( .A1(n6513), .A2(n4765), .B1(n4764), .B2(n6388), .ZN(n4758)
         );
  OAI211_X1 U5886 ( .C1(n6517), .C2(n4992), .A(n4759), .B(n4758), .ZN(U3131)
         );
  INV_X1 U5887 ( .A(n6310), .ZN(n6505) );
  AOI22_X1 U5888 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4763), .B1(n6505), 
        .B2(n4762), .ZN(n4761) );
  INV_X1 U5889 ( .A(n4960), .ZN(n6504) );
  AOI22_X1 U5890 ( .A1(n6504), .A2(n4765), .B1(n4764), .B2(n6383), .ZN(n4760)
         );
  OAI211_X1 U5891 ( .C1(n6506), .C2(n4992), .A(n4761), .B(n4760), .ZN(U3130)
         );
  INV_X1 U5892 ( .A(n6301), .ZN(n6481) );
  AOI22_X1 U5893 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4763), .B1(n6481), 
        .B2(n4762), .ZN(n4767) );
  INV_X1 U5894 ( .A(n4980), .ZN(n6480) );
  AOI22_X1 U5895 ( .A1(n6480), .A2(n4765), .B1(n4764), .B2(n6420), .ZN(n4766)
         );
  OAI211_X1 U5896 ( .C1(n6482), .C2(n4992), .A(n4767), .B(n4766), .ZN(U3127)
         );
  OAI222_X1 U5897 ( .A1(n4769), .A2(n5831), .B1(n5050), .B2(n4768), .C1(n5515), 
        .C2(n3829), .ZN(U2884) );
  AND2_X1 U5898 ( .A1(n4771), .A2(n4770), .ZN(n4773) );
  AND2_X1 U5899 ( .A1(n4773), .A2(n4772), .ZN(n5039) );
  CLKBUF_X1 U5900 ( .A(n4774), .Z(n4775) );
  OAI21_X1 U5901 ( .B1(n5039), .B2(n4776), .A(n4775), .ZN(n5151) );
  INV_X1 U5902 ( .A(n5050), .ZN(n4902) );
  AOI22_X1 U5903 ( .A1(n4902), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6019), .ZN(n4777) );
  OAI21_X1 U5904 ( .B1(n5151), .B2(n5831), .A(n4777), .ZN(U2880) );
  OR2_X1 U5905 ( .A1(n4778), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5906 ( .A1(n4792), .A2(n4780), .ZN(n6112) );
  INV_X1 U5907 ( .A(n6112), .ZN(n4781) );
  AOI22_X1 U5908 ( .A1(n5512), .A2(n4781), .B1(n5511), .B2(EBX_REG_11__SCAN_IN), .ZN(n4782) );
  OAI21_X1 U5909 ( .B1(n5151), .B2(n5228), .A(n4782), .ZN(U2848) );
  AND2_X1 U5910 ( .A1(n4783), .A2(n4784), .ZN(n4787) );
  OR2_X1 U5911 ( .A1(n4787), .A2(n4786), .ZN(n5248) );
  AOI22_X1 U5912 ( .A1(n4902), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6019), .ZN(n4788) );
  OAI21_X1 U5913 ( .B1(n5248), .B2(n5831), .A(n4788), .ZN(U2878) );
  INV_X1 U5914 ( .A(n4783), .ZN(n4789) );
  AOI21_X1 U5915 ( .B1(n4790), .B2(n4775), .A(n4789), .ZN(n5955) );
  INV_X1 U5916 ( .A(n5955), .ZN(n4796) );
  INV_X1 U5917 ( .A(n4854), .ZN(n4791) );
  AOI21_X1 U5918 ( .B1(n4793), .B2(n4792), .A(n4791), .ZN(n5952) );
  AOI22_X1 U5919 ( .A1(n5952), .A2(n5512), .B1(EBX_REG_12__SCAN_IN), .B2(n5511), .ZN(n4794) );
  OAI21_X1 U5920 ( .B1(n4796), .B2(n5228), .A(n4794), .ZN(U2847) );
  AOI22_X1 U5921 ( .A1(n4902), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6019), .ZN(n4795) );
  OAI21_X1 U5922 ( .B1(n4796), .B2(n5831), .A(n4795), .ZN(U2879) );
  INV_X1 U5923 ( .A(n4900), .ZN(n4797) );
  AOI21_X1 U5924 ( .B1(n4799), .B2(n4798), .A(n4797), .ZN(n4897) );
  INV_X1 U5925 ( .A(n4897), .ZN(n5457) );
  AOI22_X1 U5926 ( .A1(n4902), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6019), .ZN(n4800) );
  OAI21_X1 U5927 ( .B1(n5457), .B2(n5831), .A(n4800), .ZN(U2883) );
  INV_X1 U5928 ( .A(n4801), .ZN(n4804) );
  AOI21_X1 U5929 ( .B1(n4804), .B2(n4803), .A(n4802), .ZN(n4805) );
  OR2_X1 U5930 ( .A1(n4805), .A2(n5046), .ZN(n5452) );
  INV_X1 U5931 ( .A(n5452), .ZN(n6128) );
  AOI22_X1 U5932 ( .A1(n5512), .A2(n6128), .B1(n5511), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4806) );
  OAI21_X1 U5933 ( .B1(n5457), .B2(n5228), .A(n4806), .ZN(U2851) );
  OAI21_X1 U5934 ( .B1(n4786), .B2(n4808), .A(n4807), .ZN(n5273) );
  NOR2_X1 U5935 ( .A1(n4855), .A2(n4809), .ZN(n4810) );
  OR2_X1 U5936 ( .A1(n5062), .A2(n4810), .ZN(n5897) );
  OAI22_X1 U5937 ( .A1(n5897), .A2(n5507), .B1(n6803), .B2(n5505), .ZN(n4811)
         );
  INV_X1 U5938 ( .A(n4811), .ZN(n4812) );
  OAI21_X1 U5939 ( .B1(n5273), .B2(n5228), .A(n4812), .ZN(U2845) );
  OAI21_X1 U5940 ( .B1(n4815), .B2(n4813), .A(n4814), .ZN(n6152) );
  NAND2_X1 U5941 ( .A1(n5580), .A2(REIP_REG_6__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U5942 ( .B1(n5610), .B2(n5154), .A(n6143), .ZN(n4817) );
  NOR2_X1 U5943 ( .A1(n5160), .A2(n5590), .ZN(n4816) );
  AOI211_X1 U5944 ( .C1(n5622), .C2(n5158), .A(n4817), .B(n4816), .ZN(n4818)
         );
  OAI21_X1 U5945 ( .B1(n5924), .B2(n6152), .A(n4818), .ZN(U2980) );
  OR2_X1 U5946 ( .A1(n6289), .A2(n4906), .ZN(n6280) );
  NAND3_X1 U5947 ( .A1(n6280), .A2(n6447), .A3(n6275), .ZN(n4819) );
  NOR2_X1 U5948 ( .A1(n4953), .A2(n5725), .ZN(n6283) );
  AOI21_X1 U5949 ( .B1(n4819), .B2(n4908), .A(n6283), .ZN(n4822) );
  OAI21_X1 U5950 ( .B1(n4823), .B2(n6568), .A(n4820), .ZN(n4954) );
  AND2_X1 U5951 ( .A1(n6355), .A2(n6288), .ZN(n6272) );
  INV_X1 U5952 ( .A(n6442), .ZN(n6322) );
  OAI211_X1 U5953 ( .C1(n6272), .C2(n6942), .A(n6322), .B(n6397), .ZN(n4821)
         );
  NOR3_X2 U5954 ( .A1(n4822), .A2(n4954), .A3(n4821), .ZN(n6274) );
  INV_X1 U5955 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4828) );
  OR2_X1 U5956 ( .A1(n5989), .A2(n6401), .ZN(n6242) );
  NAND3_X1 U5957 ( .A1(n6327), .A2(n4823), .A3(n6397), .ZN(n4824) );
  OAI21_X1 U5958 ( .B1(n6242), .B2(n4953), .A(n4824), .ZN(n6273) );
  AOI22_X1 U5959 ( .A1(n6505), .A2(n6273), .B1(n6504), .B2(n6272), .ZN(n4825)
         );
  OAI21_X1 U5960 ( .B1(n6511), .B2(n6275), .A(n4825), .ZN(n4826) );
  AOI21_X1 U5961 ( .B1(n6430), .B2(n6313), .A(n4826), .ZN(n4827) );
  OAI21_X1 U5962 ( .B1(n6274), .B2(n4828), .A(n4827), .ZN(U3074) );
  INV_X1 U5963 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4832) );
  AOI22_X1 U5964 ( .A1(n6489), .A2(n6273), .B1(n6488), .B2(n6272), .ZN(n4829)
         );
  OAI21_X1 U5965 ( .B1(n6495), .B2(n6275), .A(n4829), .ZN(n4830) );
  AOI21_X1 U5966 ( .B1(n6424), .B2(n6313), .A(n4830), .ZN(n4831) );
  OAI21_X1 U5967 ( .B1(n6274), .B2(n4832), .A(n4831), .ZN(U3072) );
  INV_X1 U5968 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5969 ( .A1(n6515), .A2(n6273), .B1(n6513), .B2(n6272), .ZN(n4833)
         );
  OAI21_X1 U5970 ( .B1(n6524), .B2(n6275), .A(n4833), .ZN(n4834) );
  AOI21_X1 U5971 ( .B1(n6433), .B2(n6313), .A(n4834), .ZN(n4835) );
  OAI21_X1 U5972 ( .B1(n6274), .B2(n4836), .A(n4835), .ZN(U3075) );
  INV_X1 U5973 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U5974 ( .A1(n6497), .A2(n6273), .B1(n6496), .B2(n6272), .ZN(n4837)
         );
  OAI21_X1 U5975 ( .B1(n6503), .B2(n6275), .A(n4837), .ZN(n4838) );
  AOI21_X1 U5976 ( .B1(n6427), .B2(n6313), .A(n4838), .ZN(n4839) );
  OAI21_X1 U5977 ( .B1(n6274), .B2(n4840), .A(n4839), .ZN(U3073) );
  INV_X1 U5978 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U5979 ( .A1(n6473), .A2(n6273), .B1(n6472), .B2(n6272), .ZN(n4841)
         );
  OAI21_X1 U5980 ( .B1(n6479), .B2(n6275), .A(n4841), .ZN(n4842) );
  AOI21_X1 U5981 ( .B1(n6417), .B2(n6313), .A(n4842), .ZN(n4843) );
  OAI21_X1 U5982 ( .B1(n6274), .B2(n4844), .A(n4843), .ZN(U3070) );
  INV_X1 U5983 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U5984 ( .A1(n6481), .A2(n6273), .B1(n6480), .B2(n6272), .ZN(n4845)
         );
  OAI21_X1 U5985 ( .B1(n6487), .B2(n6275), .A(n4845), .ZN(n4846) );
  AOI21_X1 U5986 ( .B1(n6373), .B2(n6313), .A(n4846), .ZN(n4847) );
  OAI21_X1 U5987 ( .B1(n6274), .B2(n4848), .A(n4847), .ZN(U3071) );
  INV_X1 U5988 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U5989 ( .A1(n6465), .A2(n6273), .B1(n6464), .B2(n6272), .ZN(n4849)
         );
  OAI21_X1 U5990 ( .B1(n6466), .B2(n6275), .A(n4849), .ZN(n4850) );
  AOI21_X1 U5991 ( .B1(n6414), .B2(n6313), .A(n4850), .ZN(n4851) );
  OAI21_X1 U5992 ( .B1(n6274), .B2(n4852), .A(n4851), .ZN(U3069) );
  AND2_X1 U5993 ( .A1(n4854), .A2(n4853), .ZN(n4856) );
  OR2_X1 U5994 ( .A1(n4856), .A2(n4855), .ZN(n5437) );
  INV_X1 U5995 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5438) );
  OAI222_X1 U5996 ( .A1(n5437), .A2(n5507), .B1(n5505), .B2(n5438), .C1(n5514), 
        .C2(n5248), .ZN(U2846) );
  OR2_X1 U5997 ( .A1(n6354), .A2(n4857), .ZN(n4863) );
  AOI21_X1 U5998 ( .B1(n4863), .B2(n6440), .A(n6353), .ZN(n4858) );
  NOR2_X1 U5999 ( .A1(n4858), .A2(n6401), .ZN(n4861) );
  NOR2_X1 U6000 ( .A1(n5178), .A2(n5715), .ZN(n4910) );
  AND2_X1 U6001 ( .A1(n4910), .A2(n5989), .ZN(n6404) );
  NOR3_X1 U6002 ( .A1(n6322), .A2(n6397), .A3(n6320), .ZN(n4859) );
  AOI21_X1 U6003 ( .B1(n4861), .B2(n6404), .A(n4859), .ZN(n4890) );
  NOR2_X1 U6004 ( .A1(n6327), .A2(n4954), .ZN(n4913) );
  INV_X1 U6005 ( .A(n6404), .ZN(n4860) );
  NAND3_X1 U6006 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6539), .ZN(n6409) );
  OR2_X1 U6007 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6409), .ZN(n4886)
         );
  AOI22_X1 U6008 ( .A1(n4861), .A2(n4860), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4886), .ZN(n4862) );
  OAI211_X1 U6009 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6568), .A(n4913), .B(n4862), .ZN(n4885) );
  NAND2_X1 U6010 ( .A1(n4885), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4866)
         );
  OAI22_X1 U6011 ( .A1(n4972), .A2(n4886), .B1(n6440), .B2(n6474), .ZN(n4864)
         );
  AOI21_X1 U6012 ( .B1(n6390), .B2(n6370), .A(n4864), .ZN(n4865) );
  OAI211_X1 U6013 ( .C1(n4890), .C2(n6298), .A(n4866), .B(n4865), .ZN(U3102)
         );
  NAND2_X1 U6014 ( .A1(n4885), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4869)
         );
  OAI22_X1 U6015 ( .A1(n4968), .A2(n4886), .B1(n6440), .B2(n6468), .ZN(n4867)
         );
  AOI21_X1 U6016 ( .B1(n6390), .B2(n6367), .A(n4867), .ZN(n4868) );
  OAI211_X1 U6017 ( .C1(n4890), .C2(n6295), .A(n4869), .B(n4868), .ZN(U3101)
         );
  NAND2_X1 U6018 ( .A1(n4885), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4872)
         );
  OAI22_X1 U6019 ( .A1(n4985), .A2(n4886), .B1(n6440), .B2(n6517), .ZN(n4870)
         );
  AOI21_X1 U6020 ( .B1(n6390), .B2(n6388), .A(n4870), .ZN(n4871) );
  OAI211_X1 U6021 ( .C1(n4890), .C2(n6317), .A(n4872), .B(n4871), .ZN(U3107)
         );
  NAND2_X1 U6022 ( .A1(n4885), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4875)
         );
  OAI22_X1 U6023 ( .A1(n4960), .A2(n4886), .B1(n6440), .B2(n6506), .ZN(n4873)
         );
  AOI21_X1 U6024 ( .B1(n6390), .B2(n6383), .A(n4873), .ZN(n4874) );
  OAI211_X1 U6025 ( .C1(n4890), .C2(n6310), .A(n4875), .B(n4874), .ZN(U3106)
         );
  NAND2_X1 U6026 ( .A1(n4885), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4878)
         );
  OAI22_X1 U6027 ( .A1(n4949), .A2(n4886), .B1(n6440), .B2(n6498), .ZN(n4876)
         );
  AOI21_X1 U6028 ( .B1(n6390), .B2(n6380), .A(n4876), .ZN(n4877) );
  OAI211_X1 U6029 ( .C1(n4890), .C2(n6307), .A(n4878), .B(n4877), .ZN(U3105)
         );
  NAND2_X1 U6030 ( .A1(n4885), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4881)
         );
  OAI22_X1 U6031 ( .A1(n4976), .A2(n4886), .B1(n6440), .B2(n6490), .ZN(n4879)
         );
  AOI21_X1 U6032 ( .B1(n6390), .B2(n6377), .A(n4879), .ZN(n4880) );
  OAI211_X1 U6033 ( .C1(n4890), .C2(n6304), .A(n4881), .B(n4880), .ZN(U3104)
         );
  NAND2_X1 U6034 ( .A1(n4885), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4884)
         );
  OAI22_X1 U6035 ( .A1(n4980), .A2(n4886), .B1(n6440), .B2(n6482), .ZN(n4882)
         );
  AOI21_X1 U6036 ( .B1(n6390), .B2(n6420), .A(n4882), .ZN(n4883) );
  OAI211_X1 U6037 ( .C1(n4890), .C2(n6301), .A(n4884), .B(n4883), .ZN(U3103)
         );
  NAND2_X1 U6038 ( .A1(n4885), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4889)
         );
  OAI22_X1 U6039 ( .A1(n4964), .A2(n4886), .B1(n6440), .B2(n6460), .ZN(n4887)
         );
  AOI21_X1 U6040 ( .B1(n6390), .B2(n6399), .A(n4887), .ZN(n4888) );
  OAI211_X1 U6041 ( .C1(n4890), .C2(n6292), .A(n4889), .B(n4888), .ZN(U3100)
         );
  OAI21_X1 U6042 ( .B1(n4893), .B2(n4892), .A(n4891), .ZN(n6129) );
  INV_X1 U6043 ( .A(n4894), .ZN(n5451) );
  NAND2_X1 U6044 ( .A1(n6178), .A2(REIP_REG_8__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U6045 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4895)
         );
  OAI211_X1 U6046 ( .C1(n6110), .C2(n5451), .A(n6126), .B(n4895), .ZN(n4896)
         );
  AOI21_X1 U6047 ( .B1(n4897), .B2(n6105), .A(n4896), .ZN(n4898) );
  OAI21_X1 U6048 ( .B1(n6129), .B2(n5924), .A(n4898), .ZN(U2978) );
  INV_X1 U6049 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6026) );
  OAI222_X1 U6050 ( .A1(n5273), .A2(n5831), .B1(n5050), .B2(n6973), .C1(n5515), 
        .C2(n6026), .ZN(U2877) );
  NAND2_X1 U6051 ( .A1(n4900), .A2(n4899), .ZN(n4901) );
  NAND2_X1 U6052 ( .A1(n5040), .A2(n4901), .ZN(n5139) );
  AOI22_X1 U6053 ( .A1(n4902), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6019), .ZN(n4903) );
  OAI21_X1 U6054 ( .B1(n5139), .B2(n5831), .A(n4903), .ZN(U2882) );
  XNOR2_X1 U6055 ( .A(n5046), .B(n5042), .ZN(n6120) );
  AOI22_X1 U6056 ( .A1(n5512), .A2(n6120), .B1(EBX_REG_9__SCAN_IN), .B2(n5511), 
        .ZN(n4904) );
  OAI21_X1 U6057 ( .B1(n5139), .B2(n5228), .A(n4904), .ZN(U2850) );
  NAND2_X1 U6058 ( .A1(n4905), .A2(n6323), .ZN(n5034) );
  NAND3_X1 U6059 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6397), .A3(n6539), .ZN(n6211) );
  NOR2_X1 U6060 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6211), .ZN(n4916)
         );
  INV_X1 U6061 ( .A(n5034), .ZN(n4909) );
  OR3_X1 U6062 ( .A1(n3934), .A2(n6210), .A3(n4906), .ZN(n4907) );
  OAI21_X1 U6063 ( .B1(n4909), .B2(n6233), .A(n4908), .ZN(n4912) );
  AND2_X1 U6064 ( .A1(n4910), .A2(n6325), .ZN(n6207) );
  INV_X1 U6065 ( .A(n6207), .ZN(n4911) );
  NAND2_X1 U6066 ( .A1(n4912), .A2(n4911), .ZN(n4914) );
  OAI221_X1 U6067 ( .B1(n4916), .B2(n6942), .C1(n4916), .C2(n4914), .A(n4913), 
        .ZN(n4938) );
  NAND2_X1 U6068 ( .A1(n4938), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4919) );
  NOR3_X1 U6069 ( .A1(n6322), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6320), 
        .ZN(n4915) );
  AOI21_X1 U6070 ( .B1(n6207), .B2(n6324), .A(n4915), .ZN(n4940) );
  INV_X1 U6071 ( .A(n4916), .ZN(n4939) );
  OAI22_X1 U6072 ( .A1(n6295), .A2(n4940), .B1(n4968), .B2(n4939), .ZN(n4917)
         );
  AOI21_X1 U6073 ( .B1(n6414), .B2(n6233), .A(n4917), .ZN(n4918) );
  OAI211_X1 U6074 ( .C1(n5034), .C2(n6466), .A(n4919), .B(n4918), .ZN(U3037)
         );
  NAND2_X1 U6075 ( .A1(n4938), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4922) );
  OAI22_X1 U6076 ( .A1(n6317), .A2(n4940), .B1(n4985), .B2(n4939), .ZN(n4920)
         );
  AOI21_X1 U6077 ( .B1(n6433), .B2(n6233), .A(n4920), .ZN(n4921) );
  OAI211_X1 U6078 ( .C1(n5034), .C2(n6524), .A(n4922), .B(n4921), .ZN(U3043)
         );
  NAND2_X1 U6079 ( .A1(n4938), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4925) );
  OAI22_X1 U6080 ( .A1(n6298), .A2(n4940), .B1(n4972), .B2(n4939), .ZN(n4923)
         );
  AOI21_X1 U6081 ( .B1(n6417), .B2(n6233), .A(n4923), .ZN(n4924) );
  OAI211_X1 U6082 ( .C1(n5034), .C2(n6479), .A(n4925), .B(n4924), .ZN(U3038)
         );
  NAND2_X1 U6083 ( .A1(n4938), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4928) );
  OAI22_X1 U6084 ( .A1(n6292), .A2(n4940), .B1(n4964), .B2(n4939), .ZN(n4926)
         );
  AOI21_X1 U6085 ( .B1(n6364), .B2(n6233), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6086 ( .C1(n6458), .C2(n5034), .A(n4928), .B(n4927), .ZN(U3036)
         );
  NAND2_X1 U6087 ( .A1(n4938), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6088 ( .A1(n6301), .A2(n4940), .B1(n4980), .B2(n4939), .ZN(n4929)
         );
  AOI21_X1 U6089 ( .B1(n6373), .B2(n6233), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6090 ( .C1(n5034), .C2(n6487), .A(n4931), .B(n4930), .ZN(U3039)
         );
  NAND2_X1 U6091 ( .A1(n4938), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6092 ( .A1(n6304), .A2(n4940), .B1(n4976), .B2(n4939), .ZN(n4932)
         );
  AOI21_X1 U6093 ( .B1(n6424), .B2(n6233), .A(n4932), .ZN(n4933) );
  OAI211_X1 U6094 ( .C1(n5034), .C2(n6495), .A(n4934), .B(n4933), .ZN(U3040)
         );
  NAND2_X1 U6095 ( .A1(n4938), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4937) );
  OAI22_X1 U6096 ( .A1(n6307), .A2(n4940), .B1(n4949), .B2(n4939), .ZN(n4935)
         );
  AOI21_X1 U6097 ( .B1(n6427), .B2(n6233), .A(n4935), .ZN(n4936) );
  OAI211_X1 U6098 ( .C1(n5034), .C2(n6503), .A(n4937), .B(n4936), .ZN(U3041)
         );
  NAND2_X1 U6099 ( .A1(n4938), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4943) );
  OAI22_X1 U6100 ( .A1(n6310), .A2(n4940), .B1(n4960), .B2(n4939), .ZN(n4941)
         );
  AOI21_X1 U6101 ( .B1(n6430), .B2(n6233), .A(n4941), .ZN(n4942) );
  OAI211_X1 U6102 ( .C1(n5034), .C2(n6511), .A(n4943), .B(n4942), .ZN(U3042)
         );
  NOR2_X1 U6103 ( .A1(n6325), .A2(n6401), .ZN(n6319) );
  INV_X1 U6104 ( .A(n4953), .ZN(n4946) );
  INV_X1 U6105 ( .A(n6327), .ZN(n6453) );
  NOR3_X1 U6106 ( .A1(n6453), .A2(n6397), .A3(n6320), .ZN(n4945) );
  AOI21_X1 U6107 ( .B1(n6319), .B2(n4946), .A(n4945), .ZN(n4986) );
  INV_X1 U6108 ( .A(n4947), .ZN(n4948) );
  NOR2_X1 U6109 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4948), .ZN(n4957)
         );
  INV_X1 U6110 ( .A(n4957), .ZN(n4984) );
  OAI22_X1 U6111 ( .A1(n6307), .A2(n4986), .B1(n4949), .B2(n4984), .ZN(n4950)
         );
  AOI21_X1 U6112 ( .B1(n6427), .B2(n4988), .A(n4950), .ZN(n4959) );
  INV_X1 U6113 ( .A(n4992), .ZN(n4951) );
  OAI21_X1 U6114 ( .B1(n4951), .B2(n4988), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4952) );
  NAND3_X1 U6115 ( .A1(n4953), .A2(n6447), .A3(n4952), .ZN(n4956) );
  NOR3_X1 U6116 ( .A1(n4954), .A2(n6397), .A3(n6442), .ZN(n4955) );
  OAI211_X1 U6117 ( .C1(n4957), .C2(n6942), .A(n4956), .B(n4955), .ZN(n4989)
         );
  NAND2_X1 U6118 ( .A1(n4989), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4958)
         );
  OAI211_X1 U6119 ( .C1(n4992), .C2(n6503), .A(n4959), .B(n4958), .ZN(U3137)
         );
  OAI22_X1 U6120 ( .A1(n6310), .A2(n4986), .B1(n4960), .B2(n4984), .ZN(n4961)
         );
  AOI21_X1 U6121 ( .B1(n6430), .B2(n4988), .A(n4961), .ZN(n4963) );
  NAND2_X1 U6122 ( .A1(n4989), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4962)
         );
  OAI211_X1 U6123 ( .C1(n4992), .C2(n6511), .A(n4963), .B(n4962), .ZN(U3138)
         );
  OAI22_X1 U6124 ( .A1(n6292), .A2(n4986), .B1(n4964), .B2(n4984), .ZN(n4965)
         );
  AOI21_X1 U6125 ( .B1(n6364), .B2(n4988), .A(n4965), .ZN(n4967) );
  NAND2_X1 U6126 ( .A1(n4989), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4966)
         );
  OAI211_X1 U6127 ( .C1(n4992), .C2(n6458), .A(n4967), .B(n4966), .ZN(U3132)
         );
  OAI22_X1 U6128 ( .A1(n6295), .A2(n4986), .B1(n4968), .B2(n4984), .ZN(n4969)
         );
  AOI21_X1 U6129 ( .B1(n6414), .B2(n4988), .A(n4969), .ZN(n4971) );
  NAND2_X1 U6130 ( .A1(n4989), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4970)
         );
  OAI211_X1 U6131 ( .C1(n4992), .C2(n6466), .A(n4971), .B(n4970), .ZN(U3133)
         );
  OAI22_X1 U6132 ( .A1(n6298), .A2(n4986), .B1(n4972), .B2(n4984), .ZN(n4973)
         );
  AOI21_X1 U6133 ( .B1(n6417), .B2(n4988), .A(n4973), .ZN(n4975) );
  NAND2_X1 U6134 ( .A1(n4989), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4974)
         );
  OAI211_X1 U6135 ( .C1(n4992), .C2(n6479), .A(n4975), .B(n4974), .ZN(U3134)
         );
  OAI22_X1 U6136 ( .A1(n6304), .A2(n4986), .B1(n4976), .B2(n4984), .ZN(n4977)
         );
  AOI21_X1 U6137 ( .B1(n6424), .B2(n4988), .A(n4977), .ZN(n4979) );
  NAND2_X1 U6138 ( .A1(n4989), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4978)
         );
  OAI211_X1 U6139 ( .C1(n4992), .C2(n6495), .A(n4979), .B(n4978), .ZN(U3136)
         );
  OAI22_X1 U6140 ( .A1(n6301), .A2(n4986), .B1(n4980), .B2(n4984), .ZN(n4981)
         );
  AOI21_X1 U6141 ( .B1(n6373), .B2(n4988), .A(n4981), .ZN(n4983) );
  NAND2_X1 U6142 ( .A1(n4989), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4982)
         );
  OAI211_X1 U6143 ( .C1(n4992), .C2(n6487), .A(n4983), .B(n4982), .ZN(U3135)
         );
  OAI22_X1 U6144 ( .A1(n6317), .A2(n4986), .B1(n4985), .B2(n4984), .ZN(n4987)
         );
  AOI21_X1 U6145 ( .B1(n6433), .B2(n4988), .A(n4987), .ZN(n4991) );
  NAND2_X1 U6146 ( .A1(n4989), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4990)
         );
  OAI211_X1 U6147 ( .C1(n4992), .C2(n6524), .A(n4991), .B(n4990), .ZN(U3139)
         );
  INV_X1 U6148 ( .A(n4807), .ZN(n4996) );
  INV_X1 U6149 ( .A(n4993), .ZN(n4995) );
  OAI21_X1 U6150 ( .B1(n4996), .B2(n4995), .A(n5067), .ZN(n5435) );
  OAI222_X1 U6151 ( .A1(n5831), .A2(n5435), .B1(n5050), .B2(n4997), .C1(n5515), 
        .C2(n4550), .ZN(U2876) );
  INV_X1 U6152 ( .A(n4998), .ZN(n5061) );
  XNOR2_X1 U6153 ( .A(n5062), .B(n5061), .ZN(n5889) );
  INV_X1 U6154 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4999) );
  OAI222_X1 U6155 ( .A1(n5514), .A2(n5435), .B1(n5507), .B2(n5889), .C1(n4999), 
        .C2(n5505), .ZN(U2844) );
  NOR2_X1 U6156 ( .A1(n6355), .A2(n5006), .ZN(n5032) );
  INV_X1 U6157 ( .A(n5032), .ZN(n5000) );
  OAI21_X1 U6158 ( .B1(n5002), .B2(n5001), .A(n5000), .ZN(n5005) );
  INV_X1 U6159 ( .A(n5006), .ZN(n5003) );
  AOI22_X1 U6160 ( .A1(n5007), .A2(n5005), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5003), .ZN(n5038) );
  INV_X1 U6161 ( .A(n5005), .ZN(n5008) );
  AOI22_X1 U6162 ( .A1(n5008), .A2(n5007), .B1(n5006), .B2(n6401), .ZN(n5009)
         );
  NAND2_X1 U6163 ( .A1(n6406), .A2(n5009), .ZN(n5031) );
  AOI22_X1 U6164 ( .A1(n6464), .A2(n5032), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5031), .ZN(n5010) );
  OAI21_X1 U6165 ( .B1(n6468), .B2(n5034), .A(n5010), .ZN(n5011) );
  AOI21_X1 U6166 ( .B1(n6367), .B2(n5036), .A(n5011), .ZN(n5012) );
  OAI21_X1 U6167 ( .B1(n5038), .B2(n6295), .A(n5012), .ZN(U3029) );
  AOI22_X1 U6168 ( .A1(n6496), .A2(n5032), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5031), .ZN(n5013) );
  OAI21_X1 U6169 ( .B1(n6498), .B2(n5034), .A(n5013), .ZN(n5014) );
  AOI21_X1 U6170 ( .B1(n6380), .B2(n5036), .A(n5014), .ZN(n5015) );
  OAI21_X1 U6171 ( .B1(n5038), .B2(n6307), .A(n5015), .ZN(U3033) );
  AOI22_X1 U6172 ( .A1(n6472), .A2(n5032), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5031), .ZN(n5016) );
  OAI21_X1 U6173 ( .B1(n6474), .B2(n5034), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6174 ( .B1(n6370), .B2(n5036), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6175 ( .B1(n5038), .B2(n6298), .A(n5018), .ZN(U3030) );
  AOI22_X1 U6176 ( .A1(n6488), .A2(n5032), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5031), .ZN(n5019) );
  OAI21_X1 U6177 ( .B1(n6490), .B2(n5034), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6178 ( .B1(n6377), .B2(n5036), .A(n5020), .ZN(n5021) );
  OAI21_X1 U6179 ( .B1(n5038), .B2(n6304), .A(n5021), .ZN(U3032) );
  AOI22_X1 U6180 ( .A1(n6513), .A2(n5032), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5031), .ZN(n5022) );
  OAI21_X1 U6181 ( .B1(n6517), .B2(n5034), .A(n5022), .ZN(n5023) );
  AOI21_X1 U6182 ( .B1(n6388), .B2(n5036), .A(n5023), .ZN(n5024) );
  OAI21_X1 U6183 ( .B1(n5038), .B2(n6317), .A(n5024), .ZN(U3035) );
  AOI22_X1 U6184 ( .A1(n6504), .A2(n5032), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5031), .ZN(n5025) );
  OAI21_X1 U6185 ( .B1(n6506), .B2(n5034), .A(n5025), .ZN(n5026) );
  AOI21_X1 U6186 ( .B1(n6383), .B2(n5036), .A(n5026), .ZN(n5027) );
  OAI21_X1 U6187 ( .B1(n5038), .B2(n6310), .A(n5027), .ZN(U3034) );
  AOI22_X1 U6188 ( .A1(n6480), .A2(n5032), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5031), .ZN(n5028) );
  OAI21_X1 U6189 ( .B1(n6482), .B2(n5034), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6190 ( .B1(n6420), .B2(n5036), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6191 ( .B1(n5038), .B2(n6301), .A(n5030), .ZN(U3031) );
  AOI22_X1 U6192 ( .A1(n6456), .A2(n5032), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5031), .ZN(n5033) );
  OAI21_X1 U6193 ( .B1(n6460), .B2(n5034), .A(n5033), .ZN(n5035) );
  AOI21_X1 U6194 ( .B1(n6399), .B2(n5036), .A(n5035), .ZN(n5037) );
  OAI21_X1 U6195 ( .B1(n5038), .B2(n6292), .A(n5037), .ZN(U3028) );
  AOI21_X1 U6196 ( .B1(n5041), .B2(n5040), .A(n5039), .ZN(n5966) );
  INV_X1 U6197 ( .A(n5966), .ZN(n5051) );
  INV_X1 U6198 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5048) );
  INV_X1 U6199 ( .A(n5042), .ZN(n5045) );
  INV_X1 U6200 ( .A(n5043), .ZN(n5044) );
  AOI21_X1 U6201 ( .B1(n5046), .B2(n5045), .A(n5044), .ZN(n5047) );
  OR2_X1 U6202 ( .A1(n4778), .A2(n5047), .ZN(n5082) );
  OAI222_X1 U6203 ( .A1(n5051), .A2(n5514), .B1(n5505), .B2(n5048), .C1(n5082), 
        .C2(n5507), .ZN(U2849) );
  OAI222_X1 U6204 ( .A1(n5051), .A2(n5831), .B1(n5050), .B2(n5049), .C1(n5515), 
        .C2(n4442), .ZN(U2881) );
  CLKBUF_X1 U6205 ( .A(n5052), .Z(n5056) );
  NAND2_X1 U6206 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  XNOR2_X1 U6207 ( .A(n5056), .B(n5055), .ZN(n6122) );
  NAND2_X1 U6208 ( .A1(n6122), .A2(n3824), .ZN(n5060) );
  INV_X1 U6209 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U6210 ( .A1(n6193), .A2(n5057), .ZN(n6119) );
  NOR2_X1 U6211 ( .A1(n6110), .A2(n5119), .ZN(n5058) );
  AOI211_X1 U6212 ( .C1(n6099), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6119), 
        .B(n5058), .ZN(n5059) );
  OAI211_X1 U6213 ( .C1(n5590), .C2(n5139), .A(n5060), .B(n5059), .ZN(U2977)
         );
  INV_X1 U6214 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6215 ( .A1(n5062), .A2(n5061), .ZN(n5064) );
  NAND2_X1 U6216 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NAND2_X1 U6217 ( .A1(n5065), .A2(n5094), .ZN(n5880) );
  AND2_X1 U6218 ( .A1(n5067), .A2(n5066), .ZN(n5069) );
  OR2_X1 U6219 ( .A1(n5069), .A2(n5068), .ZN(n6015) );
  OAI222_X1 U6220 ( .A1(n5417), .A2(n5505), .B1(n5507), .B2(n5880), .C1(n6015), 
        .C2(n5514), .ZN(U2843) );
  NAND2_X1 U6221 ( .A1(n5103), .A2(n5070), .ZN(n5073) );
  CLKBUF_X1 U6222 ( .A(n5071), .Z(n5072) );
  XOR2_X1 U6223 ( .A(n5073), .B(n5072), .Z(n5090) );
  INV_X1 U6224 ( .A(n5693), .ZN(n6148) );
  AOI22_X1 U6225 ( .A1(n5075), .A2(n6148), .B1(n5074), .B2(n5688), .ZN(n6141)
         );
  OAI21_X1 U6226 ( .B1(n6151), .B2(n6130), .A(n6141), .ZN(n6121) );
  NOR2_X1 U6227 ( .A1(n5077), .A2(n5076), .ZN(n6150) );
  NAND2_X1 U6228 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U6229 ( .B1(n6149), .B2(n6160), .A(n6187), .ZN(n6177) );
  NAND2_X1 U6230 ( .A1(n6150), .A2(n6177), .ZN(n6156) );
  NOR2_X1 U6231 ( .A1(n5078), .A2(n6156), .ZN(n6137) );
  NAND2_X1 U6232 ( .A1(n6130), .A2(n6137), .ZN(n6125) );
  AOI21_X1 U6233 ( .B1(n3554), .B2(n5079), .A(n6125), .ZN(n5081) );
  AOI22_X1 U6234 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6121), .B1(n5081), .B2(n5080), .ZN(n5085) );
  INV_X1 U6235 ( .A(n5082), .ZN(n5960) );
  INV_X1 U6236 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5083) );
  NOR2_X1 U6237 ( .A1(n6193), .A2(n5083), .ZN(n5087) );
  AOI21_X1 U6238 ( .B1(n6180), .B2(n5960), .A(n5087), .ZN(n5084) );
  OAI211_X1 U6239 ( .C1(n5090), .C2(n5881), .A(n5085), .B(n5084), .ZN(U3008)
         );
  AND2_X1 U6240 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5086)
         );
  AOI211_X1 U6241 ( .C1(n5622), .C2(n5965), .A(n5087), .B(n5086), .ZN(n5089)
         );
  NAND2_X1 U6242 ( .A1(n5966), .A2(n6105), .ZN(n5088) );
  OAI211_X1 U6243 ( .C1(n5090), .C2(n5924), .A(n5089), .B(n5088), .ZN(U2976)
         );
  NOR2_X1 U6244 ( .A1(n5068), .A2(n5092), .ZN(n5093) );
  OR2_X1 U6245 ( .A1(n5091), .A2(n5093), .ZN(n5615) );
  XOR2_X1 U6246 ( .A(n5095), .B(n5094), .Z(n5872) );
  AOI22_X1 U6247 ( .A1(n5872), .A2(n5512), .B1(EBX_REG_17__SCAN_IN), .B2(n5511), .ZN(n5096) );
  OAI21_X1 U6248 ( .B1(n5615), .B2(n5228), .A(n5096), .ZN(U2842) );
  NOR2_X2 U6249 ( .A1(n6019), .A2(n5097), .ZN(n6016) );
  AOI22_X1 U6250 ( .A1(n6016), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6019), .ZN(n5102) );
  AND2_X1 U6251 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6252 ( .A1(n6020), .A2(DATAI_1_), .ZN(n5101) );
  OAI211_X1 U6253 ( .C1(n5615), .C2(n5831), .A(n5102), .B(n5101), .ZN(U2874)
         );
  NAND2_X1 U6254 ( .A1(n5104), .A2(n5103), .ZN(n5106) );
  XNOR2_X1 U6255 ( .A(n3558), .B(n6117), .ZN(n5105) );
  XNOR2_X1 U6256 ( .A(n5106), .B(n5105), .ZN(n6114) );
  INV_X1 U6257 ( .A(n6114), .ZN(n5111) );
  INV_X1 U6258 ( .A(n5151), .ZN(n5109) );
  AOI22_X1 U6259 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5580), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5107) );
  OAI21_X1 U6260 ( .B1(n6110), .B2(n5140), .A(n5107), .ZN(n5108) );
  AOI21_X1 U6261 ( .B1(n5109), .B2(n6105), .A(n5108), .ZN(n5110) );
  OAI21_X1 U6262 ( .B1(n5111), .B2(n5924), .A(n5110), .ZN(U2975) );
  INV_X1 U6263 ( .A(n6679), .ZN(n6572) );
  NOR3_X1 U6264 ( .A1(n6972), .A2(n6942), .A3(n6572), .ZN(n6562) );
  NAND2_X1 U6265 ( .A1(n5112), .A2(n4299), .ZN(n6570) );
  INV_X1 U6266 ( .A(n6570), .ZN(n5113) );
  OR2_X1 U6267 ( .A1(n6178), .A2(n5113), .ZN(n5114) );
  OR2_X1 U6268 ( .A1(n6562), .A2(n5114), .ZN(n5115) );
  AND2_X2 U6269 ( .A1(n6011), .A2(n5118), .ZN(n6687) );
  INV_X1 U6270 ( .A(n5119), .ZN(n5137) );
  INV_X1 U6271 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5135) );
  NOR2_X1 U6272 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5125) );
  INV_X1 U6273 ( .A(n5125), .ZN(n5127) );
  NAND2_X1 U6274 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5127), .ZN(n5120) );
  NOR2_X1 U6275 ( .A1(n3673), .A2(n5120), .ZN(n5121) );
  AND3_X1 U6276 ( .A1(n5123), .A2(n5122), .A3(n5125), .ZN(n5124) );
  INV_X1 U6277 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6704) );
  NAND3_X1 U6278 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5460) );
  INV_X1 U6279 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6602) );
  NOR3_X1 U6280 ( .A1(n6704), .A2(n5460), .A3(n6602), .ZN(n5152) );
  NAND4_X1 U6281 ( .A1(n5152), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(REIP_REG_8__SCAN_IN), .ZN(n5132) );
  INV_X1 U6282 ( .A(n5132), .ZN(n5141) );
  OAI21_X1 U6283 ( .B1(n5962), .B2(n5141), .A(n6011), .ZN(n5967) );
  AOI22_X1 U6284 ( .A1(n6000), .A2(n6120), .B1(REIP_REG_9__SCAN_IN), .B2(n5967), .ZN(n5134) );
  NAND2_X1 U6285 ( .A1(n5126), .A2(n5125), .ZN(n6554) );
  INV_X1 U6286 ( .A(n6554), .ZN(n5130) );
  INV_X1 U6287 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6288 ( .A1(n5128), .A2(n5127), .ZN(n5129) );
  OAI22_X1 U6289 ( .A1(n3395), .A2(n5130), .B1(n3290), .B2(n5129), .ZN(n5131)
         );
  INV_X1 U6290 ( .A(n6011), .ZN(n5459) );
  NOR3_X1 U6291 ( .A1(n6401), .A2(STATE2_REG_1__SCAN_IN), .A3(n5459), .ZN(
        n5964) );
  NOR3_X1 U6292 ( .A1(n5962), .A2(REIP_REG_9__SCAN_IN), .A3(n5132), .ZN(n5968)
         );
  AOI211_X1 U6293 ( .C1(n6686), .C2(EBX_REG_9__SCAN_IN), .A(n5964), .B(n5968), 
        .ZN(n5133) );
  OAI211_X1 U6294 ( .C1(n5135), .C2(n5977), .A(n5134), .B(n5133), .ZN(n5136)
         );
  AOI21_X1 U6295 ( .B1(n6687), .B2(n5137), .A(n5136), .ZN(n5138) );
  OAI21_X1 U6296 ( .B1(n5802), .B2(n5139), .A(n5138), .ZN(U2818) );
  INV_X1 U6297 ( .A(n5140), .ZN(n5149) );
  INV_X1 U6298 ( .A(n5962), .ZN(n5461) );
  NAND2_X1 U6299 ( .A1(n5141), .A2(REIP_REG_9__SCAN_IN), .ZN(n5961) );
  INV_X1 U6300 ( .A(n5961), .ZN(n5142) );
  NAND2_X1 U6301 ( .A1(n5142), .A2(REIP_REG_10__SCAN_IN), .ZN(n5146) );
  INV_X1 U6302 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U6303 ( .A1(n5146), .A2(n6610), .ZN(n5230) );
  INV_X1 U6304 ( .A(n5230), .ZN(n5143) );
  NAND2_X1 U6305 ( .A1(n5461), .A2(n5143), .ZN(n5145) );
  AND2_X1 U6306 ( .A1(n5145), .A2(n6011), .ZN(n5950) );
  OAI22_X1 U6307 ( .A1(n5950), .A2(n6610), .B1(n6692), .B2(n6112), .ZN(n5148)
         );
  AOI22_X1 U6308 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6686), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6685), .ZN(n5144) );
  INV_X1 U6309 ( .A(n5964), .ZN(n5982) );
  OAI211_X1 U6310 ( .C1(n5146), .C2(n5145), .A(n5144), .B(n5982), .ZN(n5147)
         );
  AOI211_X1 U6311 ( .C1(n6687), .C2(n5149), .A(n5148), .B(n5147), .ZN(n5150)
         );
  OAI21_X1 U6312 ( .B1(n5151), .B2(n5802), .A(n5150), .ZN(U2816) );
  OAI21_X1 U6313 ( .B1(n5962), .B2(n5152), .A(n6011), .ZN(n5985) );
  AOI22_X1 U6314 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6686), .B1(
        REIP_REG_6__SCAN_IN), .B2(n5985), .ZN(n5153) );
  OAI211_X1 U6315 ( .C1(n5977), .C2(n5154), .A(n5153), .B(n5982), .ZN(n5157)
         );
  INV_X1 U6316 ( .A(n5460), .ZN(n5155) );
  NAND2_X1 U6317 ( .A1(n5461), .A2(n5155), .ZN(n5462) );
  NOR2_X1 U6318 ( .A1(n5462), .A2(n6704), .ZN(n5986) );
  NAND2_X1 U6319 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5986), .ZN(n5973) );
  OAI22_X1 U6320 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5973), .B1(n6692), .B2(n6142), .ZN(n5156) );
  AOI211_X1 U6321 ( .C1(n6687), .C2(n5158), .A(n5157), .B(n5156), .ZN(n5159)
         );
  OAI21_X1 U6322 ( .B1(n5802), .B2(n5160), .A(n5159), .ZN(U2821) );
  OR2_X1 U6323 ( .A1(n5091), .A2(n5162), .ZN(n5163) );
  AND2_X1 U6324 ( .A1(n5206), .A2(n5163), .ZN(n6012) );
  INV_X1 U6325 ( .A(n6012), .ZN(n5170) );
  XNOR2_X1 U6326 ( .A(n5165), .B(n5164), .ZN(n5166) );
  OR2_X1 U6327 ( .A1(n5167), .A2(n5166), .ZN(n5207) );
  NAND2_X1 U6328 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  AND2_X1 U6329 ( .A1(n5207), .A2(n5168), .ZN(n5946) );
  AOI22_X1 U6330 ( .A1(n5946), .A2(n5512), .B1(EBX_REG_18__SCAN_IN), .B2(n5511), .ZN(n5169) );
  OAI21_X1 U6331 ( .B1(n5170), .B2(n5228), .A(n5169), .ZN(U2841) );
  NAND2_X1 U6332 ( .A1(n5320), .A2(n5171), .ZN(n5172) );
  NOR2_X1 U6333 ( .A1(n5962), .A2(REIP_REG_1__SCAN_IN), .ZN(n5999) );
  INV_X1 U6334 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6598) );
  NOR3_X1 U6335 ( .A1(n5999), .A2(n5459), .A3(n6598), .ZN(n5995) );
  INV_X1 U6336 ( .A(n5995), .ZN(n5174) );
  INV_X1 U6337 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U6338 ( .B1(n5962), .B2(n6664), .A(n6598), .ZN(n5173) );
  NAND2_X1 U6339 ( .A1(n5174), .A2(n5173), .ZN(n5182) );
  INV_X1 U6340 ( .A(n6109), .ZN(n5175) );
  AOI22_X1 U6341 ( .A1(n6685), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6687), 
        .B2(n5175), .ZN(n5181) );
  AOI22_X1 U6342 ( .A1(n6000), .A2(n6192), .B1(n6686), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5180) );
  INV_X1 U6343 ( .A(n5176), .ZN(n5177) );
  AND2_X1 U6344 ( .A1(n5320), .A2(n5177), .ZN(n6005) );
  NAND2_X1 U6345 ( .A1(n6005), .A2(n5178), .ZN(n5179) );
  AND4_X1 U6346 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n5183)
         );
  OAI21_X1 U6347 ( .B1(n5981), .B2(n6100), .A(n5183), .ZN(U2825) );
  CLKBUF_X1 U6348 ( .A(n5184), .Z(n5185) );
  INV_X1 U6349 ( .A(n5186), .ZN(n5187) );
  NOR2_X1 U6350 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  XNOR2_X1 U6351 ( .A(n5185), .B(n5189), .ZN(n5202) );
  NOR2_X1 U6352 ( .A1(n6193), .A2(n6613), .ZN(n5199) );
  AND2_X1 U6353 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5190)
         );
  AOI211_X1 U6354 ( .C1(n5622), .C2(n5954), .A(n5199), .B(n5190), .ZN(n5192)
         );
  NAND2_X1 U6355 ( .A1(n5955), .A2(n6105), .ZN(n5191) );
  OAI211_X1 U6356 ( .C1(n5202), .C2(n5924), .A(n5192), .B(n5191), .ZN(U2974)
         );
  INV_X1 U6357 ( .A(n5688), .ZN(n5193) );
  OAI22_X1 U6358 ( .A1(n5195), .A2(n5693), .B1(n5194), .B2(n5193), .ZN(n6111)
         );
  INV_X1 U6359 ( .A(n5196), .ZN(n6118) );
  AOI211_X1 U6360 ( .C1(n5197), .C2(n6117), .A(n5252), .B(n6118), .ZN(n5198)
         );
  AOI21_X1 U6361 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6111), .A(n5198), 
        .ZN(n5201) );
  AOI21_X1 U6362 ( .B1(n6180), .B2(n5952), .A(n5199), .ZN(n5200) );
  OAI211_X1 U6363 ( .C1(n5202), .C2(n5881), .A(n5201), .B(n5200), .ZN(U3006)
         );
  AOI21_X1 U6364 ( .B1(n5206), .B2(n5205), .A(n5204), .ZN(n5597) );
  INV_X1 U6365 ( .A(n5597), .ZN(n5244) );
  XOR2_X1 U6366 ( .A(n5208), .B(n5207), .Z(n5857) );
  AOI22_X1 U6367 ( .A1(n5857), .A2(n5512), .B1(n5511), .B2(EBX_REG_19__SCAN_IN), .ZN(n5209) );
  OAI21_X1 U6368 ( .B1(n5244), .B2(n5228), .A(n5209), .ZN(U2840) );
  AOI22_X1 U6369 ( .A1(n6016), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6019), .ZN(n5211) );
  NAND2_X1 U6370 ( .A1(n6020), .A2(DATAI_3_), .ZN(n5210) );
  OAI211_X1 U6371 ( .C1(n5244), .C2(n5831), .A(n5211), .B(n5210), .ZN(U2872)
         );
  NAND2_X1 U6372 ( .A1(n5962), .A2(n6011), .ZN(n5392) );
  OAI22_X1 U6373 ( .A1(n5212), .A2(n5811), .B1(n6692), .B2(n5706), .ZN(n5213)
         );
  AOI21_X1 U6374 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5392), .A(n5213), .ZN(n5216)
         );
  NAND2_X1 U6375 ( .A1(n5977), .A2(n5998), .ZN(n5214) );
  AOI22_X1 U6376 ( .A1(n5214), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6005), 
        .B2(n6528), .ZN(n5215) );
  OAI211_X1 U6377 ( .C1(n5981), .C2(n5217), .A(n5216), .B(n5215), .ZN(U2827)
         );
  NAND2_X1 U6378 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NAND2_X1 U6379 ( .A1(n5284), .A2(n5221), .ZN(n5823) );
  MUX2_X1 U6380 ( .A(n5224), .B(n5223), .S(n5222), .Z(n5226) );
  XNOR2_X1 U6381 ( .A(n5226), .B(n5225), .ZN(n5826) );
  AOI22_X1 U6382 ( .A1(n5826), .A2(n5512), .B1(EBX_REG_20__SCAN_IN), .B2(n5511), .ZN(n5227) );
  OAI21_X1 U6383 ( .B1(n5823), .B2(n5228), .A(n5227), .ZN(U2839) );
  NAND2_X1 U6384 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5229) );
  NAND2_X1 U6385 ( .A1(n5461), .A2(n5230), .ZN(n5444) );
  INV_X1 U6386 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6989) );
  OAI21_X1 U6387 ( .B1(n5229), .B2(n5444), .A(n6989), .ZN(n5235) );
  NAND4_X1 U6388 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5230), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5239) );
  INV_X1 U6389 ( .A(n5239), .ZN(n5418) );
  OAI21_X1 U6390 ( .B1(n5962), .B2(n5418), .A(n6011), .ZN(n5427) );
  AOI21_X1 U6391 ( .B1(n6687), .B2(n5270), .A(n5964), .ZN(n5231) );
  OAI21_X1 U6392 ( .B1(n6692), .B2(n5897), .A(n5231), .ZN(n5234) );
  OAI22_X1 U6393 ( .A1(n6803), .A2(n5811), .B1(n5232), .B2(n5977), .ZN(n5233)
         );
  AOI211_X1 U6394 ( .C1(n5235), .C2(n5427), .A(n5234), .B(n5233), .ZN(n5236)
         );
  OAI21_X1 U6395 ( .B1(n5273), .B2(n5802), .A(n5236), .ZN(U2813) );
  OAI21_X1 U6396 ( .B1(n5977), .B2(n6804), .A(n5982), .ZN(n5237) );
  AOI21_X1 U6397 ( .B1(n6687), .B2(n5594), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6398 ( .B1(n5811), .B2(n3733), .A(n5238), .ZN(n5242) );
  INV_X1 U6399 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6623) );
  INV_X1 U6400 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6620) );
  NOR2_X1 U6401 ( .A1(n6623), .A2(n6620), .ZN(n5821) );
  INV_X1 U6402 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6617) );
  NOR2_X1 U6403 ( .A1(n5239), .A2(n6617), .ZN(n5411) );
  NAND3_X1 U6404 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        n5411), .ZN(n5315) );
  OAI21_X1 U6405 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5942), .ZN(n5240) );
  OAI21_X1 U6406 ( .B1(n5459), .B2(n5315), .A(n5392), .ZN(n5944) );
  OAI22_X1 U6407 ( .A1(n5821), .A2(n5240), .B1(n5944), .B2(n6623), .ZN(n5241)
         );
  AOI211_X1 U6408 ( .C1(n5857), .C2(n6000), .A(n5242), .B(n5241), .ZN(n5243)
         );
  OAI21_X1 U6409 ( .B1(n5244), .B2(n5802), .A(n5243), .ZN(U2808) );
  XOR2_X1 U6410 ( .A(n5247), .B(n5246), .Z(n5262) );
  INV_X1 U6411 ( .A(n5248), .ZN(n5436) );
  AND2_X1 U6412 ( .A1(n5580), .A2(REIP_REG_13__SCAN_IN), .ZN(n5259) );
  AOI21_X1 U6413 ( .B1(n6099), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5259), 
        .ZN(n5249) );
  OAI21_X1 U6414 ( .B1(n6110), .B2(n5441), .A(n5249), .ZN(n5250) );
  AOI21_X1 U6415 ( .B1(n5436), .B2(n6105), .A(n5250), .ZN(n5251) );
  OAI21_X1 U6416 ( .B1(n5262), .B2(n5924), .A(n5251), .ZN(U2973) );
  INV_X1 U6417 ( .A(n5437), .ZN(n5260) );
  NAND2_X1 U6418 ( .A1(n5252), .A2(n3559), .ZN(n5902) );
  NOR2_X1 U6419 ( .A1(n5254), .A2(n5253), .ZN(n5255) );
  AOI211_X1 U6420 ( .C1(n5257), .C2(n5256), .A(n5255), .B(n6111), .ZN(n5901)
         );
  OAI22_X1 U6421 ( .A1(n6118), .A2(n5902), .B1(n5901), .B2(n3559), .ZN(n5258)
         );
  AOI211_X1 U6422 ( .C1(n6180), .C2(n5260), .A(n5259), .B(n5258), .ZN(n5261)
         );
  OAI21_X1 U6423 ( .B1(n5262), .B2(n5881), .A(n5261), .ZN(U3005) );
  INV_X1 U6424 ( .A(n5265), .ZN(n5267) );
  NOR2_X1 U6425 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6426 ( .A(n5264), .B(n5268), .ZN(n5905) );
  NAND2_X1 U6427 ( .A1(n5905), .A2(n3824), .ZN(n5272) );
  NAND2_X1 U6428 ( .A1(n6178), .A2(REIP_REG_14__SCAN_IN), .ZN(n5898) );
  OAI21_X1 U6429 ( .B1(n5610), .B2(n5232), .A(n5898), .ZN(n5269) );
  AOI21_X1 U6430 ( .B1(n5622), .B2(n5270), .A(n5269), .ZN(n5271) );
  OAI211_X1 U6431 ( .C1(n5590), .C2(n5273), .A(n5272), .B(n5271), .ZN(U2972)
         );
  OAI21_X1 U6432 ( .B1(n5275), .B2(n5277), .A(n5388), .ZN(n5816) );
  INV_X1 U6433 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U6434 ( .A1(n5278), .A2(n5279), .ZN(n5280) );
  NAND2_X1 U6435 ( .A1(n5394), .A2(n5280), .ZN(n5820) );
  OAI222_X1 U6436 ( .A1(n5514), .A2(n5816), .B1(n5505), .B2(n5812), .C1(n5820), 
        .C2(n5507), .ZN(U2837) );
  OR2_X1 U6437 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U6438 ( .A1(n5278), .A2(n5283), .ZN(n5680) );
  AOI21_X1 U6439 ( .B1(n5285), .B2(n5284), .A(n5275), .ZN(n5843) );
  INV_X1 U6440 ( .A(n5843), .ZN(n5409) );
  OAI222_X1 U6441 ( .A1(n5402), .A2(n5505), .B1(n5507), .B2(n5680), .C1(n5409), 
        .C2(n5514), .ZN(U2838) );
  XNOR2_X1 U6442 ( .A(n3558), .B(n6760), .ZN(n5287) );
  XNOR2_X1 U6443 ( .A(n5288), .B(n5287), .ZN(n5893) );
  NAND2_X1 U6444 ( .A1(n5893), .A2(n3824), .ZN(n5291) );
  NOR2_X1 U6445 ( .A1(n6193), .A2(n6617), .ZN(n5890) );
  NOR2_X1 U6446 ( .A1(n6110), .A2(n5430), .ZN(n5289) );
  AOI211_X1 U6447 ( .C1(n6099), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5890), 
        .B(n5289), .ZN(n5290) );
  OAI211_X1 U6448 ( .C1(n5590), .C2(n5435), .A(n5291), .B(n5290), .ZN(U2971)
         );
  XNOR2_X1 U6449 ( .A(n3558), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5592)
         );
  NAND2_X1 U6450 ( .A1(n5593), .A2(n5592), .ZN(n5591) );
  INV_X1 U6451 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U6452 ( .A1(n5591), .A2(n5292), .ZN(n5584) );
  NAND2_X1 U6453 ( .A1(n5584), .A2(n3136), .ZN(n5294) );
  INV_X1 U6454 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5703) );
  XNOR2_X1 U6455 ( .A(n5296), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5578)
         );
  NOR2_X1 U6456 ( .A1(n5577), .A2(n5578), .ZN(n5576) );
  NOR2_X1 U6457 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5569)
         );
  NAND2_X1 U6458 ( .A1(n5576), .A2(n5569), .ZN(n5559) );
  INV_X1 U6459 ( .A(n5576), .ZN(n5295) );
  OAI21_X1 U6460 ( .B1(n5296), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5295), 
        .ZN(n5571) );
  NAND3_X1 U6461 ( .A1(n5603), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6462 ( .A(n5298), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5314)
         );
  NOR2_X1 U6463 ( .A1(n5393), .A2(n5299), .ZN(n5300) );
  OR2_X1 U6464 ( .A1(n5502), .A2(n5300), .ZN(n6693) );
  INV_X1 U6465 ( .A(n6693), .ZN(n5301) );
  AND2_X1 U6466 ( .A1(n6178), .A2(REIP_REG_24__SCAN_IN), .ZN(n5308) );
  AOI21_X1 U6467 ( .B1(n5301), .B2(n6180), .A(n5308), .ZN(n5305) );
  INV_X1 U6468 ( .A(n5302), .ZN(n5303) );
  OAI211_X1 U6469 ( .C1(INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n5664), .A(n5661), .B(n5303), .ZN(n5304) );
  OAI211_X1 U6470 ( .C1(n5314), .C2(n5881), .A(n5305), .B(n5304), .ZN(U2994)
         );
  NOR2_X1 U6471 ( .A1(n5610), .A2(n5306), .ZN(n5307) );
  AOI211_X1 U6472 ( .C1(n5622), .C2(n6688), .A(n5308), .B(n5307), .ZN(n5313)
         );
  INV_X1 U6473 ( .A(n5309), .ZN(n5310) );
  XOR2_X1 U6474 ( .A(n5311), .B(n5310), .Z(n6697) );
  NAND2_X1 U6475 ( .A1(n6697), .A2(n6105), .ZN(n5312) );
  OAI211_X1 U6476 ( .C1(n5314), .C2(n5924), .A(n5313), .B(n5312), .ZN(U2962)
         );
  INV_X1 U6477 ( .A(n5517), .ZN(n5327) );
  INV_X1 U6478 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6632) );
  INV_X1 U6479 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6903) );
  INV_X1 U6480 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6625) );
  NAND4_X1 U6481 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5942), .ZN(n5808) );
  NOR2_X1 U6482 ( .A1(n6625), .A2(n5808), .ZN(n5815) );
  NAND2_X1 U6483 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5815), .ZN(n5390) );
  NOR2_X1 U6484 ( .A1(n6903), .A2(n5390), .ZN(n5800) );
  NAND2_X1 U6485 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5800), .ZN(n5797) );
  NOR2_X1 U6486 ( .A1(n6632), .A2(n5797), .ZN(n5791) );
  NAND2_X1 U6487 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5791), .ZN(n5787) );
  NAND2_X1 U6488 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5318) );
  NOR2_X1 U6489 ( .A1(n5787), .A2(n5318), .ZN(n5378) );
  INV_X1 U6490 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U6491 ( .A1(n5378), .A2(n6637), .ZN(n5375) );
  INV_X1 U6492 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6925) );
  NAND3_X1 U6493 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5316) );
  NOR3_X1 U6494 ( .A1(n5459), .A2(n5316), .A3(n5315), .ZN(n5809) );
  NAND4_X1 U6495 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5809), .ZN(n5391) );
  NOR3_X1 U6496 ( .A1(n6925), .A2(n6632), .A3(n5391), .ZN(n5317) );
  INV_X1 U6497 ( .A(n5392), .ZN(n5810) );
  AOI21_X1 U6498 ( .B1(n5317), .B2(REIP_REG_26__SCAN_IN), .A(n5810), .ZN(n5792) );
  AOI21_X1 U6499 ( .B1(n5461), .B2(n5318), .A(n5792), .ZN(n5772) );
  NAND2_X1 U6500 ( .A1(n5375), .A2(n5772), .ZN(n5385) );
  AND4_X1 U6501 ( .A1(n5320), .A2(n5319), .A3(EBX_REG_31__SCAN_IN), .A4(n6554), 
        .ZN(n5321) );
  AOI21_X1 U6502 ( .B1(n6685), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5321), 
        .ZN(n5324) );
  OAI21_X1 U6503 ( .B1(n6637), .B2(REIP_REG_31__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5322) );
  OAI211_X1 U6504 ( .C1(REIP_REG_31__SCAN_IN), .C2(REIP_REG_30__SCAN_IN), .A(
        n5378), .B(n5322), .ZN(n5323) );
  OAI211_X1 U6505 ( .C1(n5328), .C2(n6692), .A(n5324), .B(n5323), .ZN(n5325)
         );
  AOI21_X1 U6506 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5385), .A(n5325), .ZN(n5326) );
  OAI21_X1 U6507 ( .B1(n5327), .B2(n5802), .A(n5326), .ZN(U2796) );
  OAI22_X1 U6508 ( .A1(n5328), .A2(n5507), .B1(n5128), .B2(n5505), .ZN(U2828)
         );
  OR2_X1 U6509 ( .A1(n5603), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5544)
         );
  INV_X1 U6510 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U6511 ( .A1(n6738), .A2(n5533), .ZN(n5637) );
  OR2_X1 U6512 ( .A1(n5544), .A2(n5637), .ZN(n5357) );
  NOR3_X1 U6513 ( .A1(n5547), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5357), 
        .ZN(n5330) );
  NOR2_X1 U6514 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  INV_X1 U6515 ( .A(n5333), .ZN(n5347) );
  NAND2_X1 U6516 ( .A1(n5339), .A2(n5478), .ZN(n5334) );
  NAND2_X1 U6517 ( .A1(n5334), .A2(n5337), .ZN(n5335) );
  INV_X1 U6518 ( .A(n5337), .ZN(n5338) );
  OAI211_X1 U6519 ( .C1(n5478), .C2(n5340), .A(n5339), .B(n5338), .ZN(n5341)
         );
  NAND2_X1 U6520 ( .A1(n5580), .A2(REIP_REG_30__SCAN_IN), .ZN(n5351) );
  INV_X1 U6521 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5343) );
  NAND3_X1 U6522 ( .A1(n5644), .A2(n5344), .A3(n5343), .ZN(n5345) );
  OAI211_X1 U6523 ( .C1(n5471), .C2(n6195), .A(n5351), .B(n5345), .ZN(n5346)
         );
  AOI21_X1 U6524 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5347), .A(n5346), 
        .ZN(n5348) );
  OAI21_X1 U6525 ( .B1(n3122), .B2(n5881), .A(n5348), .ZN(U2988) );
  AOI21_X1 U6526 ( .B1(n5350), .B2(n5362), .A(n5349), .ZN(n5377) );
  INV_X1 U6527 ( .A(n5351), .ZN(n5352) );
  AOI21_X1 U6528 ( .B1(n6099), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5352), 
        .ZN(n5353) );
  OAI21_X1 U6529 ( .B1(n6110), .B2(n5379), .A(n5353), .ZN(n5354) );
  AOI21_X1 U6530 ( .B1(n5377), .B2(n6105), .A(n5354), .ZN(n5355) );
  OAI21_X1 U6531 ( .B1(n3122), .B2(n5924), .A(n5355), .ZN(U2956) );
  INV_X1 U6532 ( .A(n5628), .ZN(n5638) );
  OAI22_X1 U6533 ( .A1(n5539), .A2(n5638), .B1(n5547), .B2(n5357), .ZN(n5358)
         );
  XNOR2_X1 U6534 ( .A(n5358), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5635)
         );
  INV_X1 U6535 ( .A(n5370), .ZN(n5363) );
  NAND2_X1 U6536 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5359)
         );
  NAND2_X1 U6537 ( .A1(n5580), .A2(REIP_REG_29__SCAN_IN), .ZN(n5630) );
  OAI211_X1 U6538 ( .C1(n6110), .C2(n5363), .A(n3137), .B(n3123), .ZN(n5364)
         );
  INV_X1 U6539 ( .A(n5364), .ZN(n5365) );
  OAI21_X1 U6540 ( .B1(n5635), .B2(n5924), .A(n5365), .ZN(U2957) );
  AOI22_X1 U6541 ( .A1(n6016), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6019), .ZN(n5368) );
  NAND2_X1 U6542 ( .A1(n6020), .A2(DATAI_13_), .ZN(n5367) );
  OAI211_X1 U6543 ( .C1(n5366), .C2(n5831), .A(n5368), .B(n5367), .ZN(U2862)
         );
  XOR2_X1 U6544 ( .A(n5369), .B(n5478), .Z(n5631) );
  INV_X1 U6545 ( .A(n5631), .ZN(n5374) );
  AOI22_X1 U6546 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6685), .B1(n6687), 
        .B2(n5370), .ZN(n5372) );
  NAND2_X1 U6547 ( .A1(n6686), .A2(EBX_REG_29__SCAN_IN), .ZN(n5371) );
  OAI211_X1 U6548 ( .C1(n5772), .C2(n6637), .A(n5372), .B(n5371), .ZN(n5373)
         );
  AOI21_X1 U6549 ( .B1(n5374), .B2(n6000), .A(n5373), .ZN(n5376) );
  OAI211_X1 U6550 ( .C1(n5366), .C2(n5802), .A(n5376), .B(n5375), .ZN(U2798)
         );
  OAI222_X1 U6551 ( .A1(n6895), .A2(n5505), .B1(n5507), .B2(n5631), .C1(n5514), 
        .C2(n5366), .ZN(U2830) );
  INV_X1 U6552 ( .A(n5377), .ZN(n5522) );
  INV_X1 U6553 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6644) );
  AND3_X1 U6554 ( .A1(n5378), .A2(REIP_REG_29__SCAN_IN), .A3(n6644), .ZN(n5384) );
  INV_X1 U6555 ( .A(n5379), .ZN(n5380) );
  AOI22_X1 U6556 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6685), .B1(n6687), 
        .B2(n5380), .ZN(n5382) );
  NAND2_X1 U6557 ( .A1(n6686), .A2(EBX_REG_30__SCAN_IN), .ZN(n5381) );
  OAI211_X1 U6558 ( .C1(n5471), .C2(n6692), .A(n5382), .B(n5381), .ZN(n5383)
         );
  OAI21_X1 U6559 ( .B1(n5522), .B2(n5802), .A(n5386), .ZN(U2797) );
  INV_X1 U6560 ( .A(n5310), .ZN(n5387) );
  AOI21_X1 U6561 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n5567) );
  INV_X1 U6562 ( .A(n5567), .ZN(n5529) );
  NAND2_X1 U6563 ( .A1(n6903), .A2(n5390), .ZN(n5400) );
  AND2_X1 U6564 ( .A1(n5392), .A2(n5391), .ZN(n6689) );
  AOI21_X1 U6565 ( .B1(n5395), .B2(n5394), .A(n5393), .ZN(n5665) );
  INV_X1 U6566 ( .A(n5665), .ZN(n5398) );
  OAI22_X1 U6567 ( .A1(n6956), .A2(n5811), .B1(n5565), .B2(n5977), .ZN(n5396)
         );
  AOI21_X1 U6568 ( .B1(n6687), .B2(n5563), .A(n5396), .ZN(n5397) );
  OAI21_X1 U6569 ( .B1(n5398), .B2(n6692), .A(n5397), .ZN(n5399) );
  AOI21_X1 U6570 ( .B1(n5400), .B2(n6689), .A(n5399), .ZN(n5401) );
  OAI21_X1 U6571 ( .B1(n5529), .B2(n5802), .A(n5401), .ZN(U2804) );
  NOR2_X1 U6572 ( .A1(n5810), .A2(n5809), .ZN(n5822) );
  NOR2_X1 U6573 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5808), .ZN(n5404) );
  OAI22_X1 U6574 ( .A1(n5402), .A2(n5811), .B1(n6790), .B2(n5977), .ZN(n5403)
         );
  AOI211_X1 U6575 ( .C1(n5822), .C2(REIP_REG_21__SCAN_IN), .A(n5404), .B(n5403), .ZN(n5408) );
  INV_X1 U6576 ( .A(n5579), .ZN(n5405) );
  OAI22_X1 U6577 ( .A1(n5680), .A2(n6692), .B1(n5405), .B2(n5998), .ZN(n5406)
         );
  INV_X1 U6578 ( .A(n5406), .ZN(n5407) );
  OAI211_X1 U6579 ( .C1(n5409), .C2(n5802), .A(n5408), .B(n5407), .ZN(U2806)
         );
  NAND2_X1 U6580 ( .A1(n6686), .A2(EBX_REG_17__SCAN_IN), .ZN(n5410) );
  OAI211_X1 U6581 ( .C1(n5998), .C2(n5607), .A(n5410), .B(n5982), .ZN(n5414)
         );
  AND2_X1 U6582 ( .A1(n5461), .A2(n5411), .ZN(n5420) );
  AOI21_X1 U6583 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5420), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5412) );
  OAI22_X1 U6584 ( .A1(n5944), .A2(n5412), .B1(n5609), .B2(n5977), .ZN(n5413)
         );
  AOI211_X1 U6585 ( .C1(n6000), .C2(n5872), .A(n5414), .B(n5413), .ZN(n5415)
         );
  OAI21_X1 U6586 ( .B1(n5615), .B2(n5802), .A(n5415), .ZN(U2810) );
  INV_X1 U6587 ( .A(n5880), .ZN(n5425) );
  INV_X1 U6588 ( .A(n5621), .ZN(n5416) );
  OAI22_X1 U6589 ( .A1(n5811), .A2(n5417), .B1(n5416), .B2(n5998), .ZN(n5424)
         );
  INV_X1 U6591 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U6592 ( .A1(n6617), .A2(n5418), .ZN(n5419) );
  NOR2_X1 U6593 ( .A1(n5962), .A2(n5419), .ZN(n5432) );
  OAI33_X1 U6594 ( .A1(1'b0), .A2(n5420), .A3(REIP_REG_16__SCAN_IN), .B1(n6912), .B2(n5427), .B3(n5432), .ZN(n5422) );
  OAI211_X1 U6595 ( .C1(n5977), .C2(n6733), .A(n5422), .B(n5982), .ZN(n5423)
         );
  AOI211_X1 U6596 ( .C1(n5425), .C2(n6000), .A(n5424), .B(n5423), .ZN(n5426)
         );
  OAI21_X1 U6597 ( .B1(n6015), .B2(n5802), .A(n5426), .ZN(U2811) );
  AOI22_X1 U6598 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6686), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5427), .ZN(n5428) );
  OAI211_X1 U6599 ( .C1(n5977), .C2(n5429), .A(n5428), .B(n5982), .ZN(n5433)
         );
  OAI22_X1 U6600 ( .A1(n6692), .A2(n5889), .B1(n5430), .B2(n5998), .ZN(n5431)
         );
  NOR3_X1 U6601 ( .A1(n5433), .A2(n5432), .A3(n5431), .ZN(n5434) );
  OAI21_X1 U6602 ( .B1(n5435), .B2(n5802), .A(n5434), .ZN(U2812) );
  NAND2_X1 U6603 ( .A1(n5436), .A2(n6696), .ZN(n5448) );
  OAI22_X1 U6604 ( .A1(n5438), .A2(n5811), .B1(n6692), .B2(n5437), .ZN(n5439)
         );
  AOI211_X1 U6605 ( .C1(n6685), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5439), 
        .B(n5964), .ZN(n5447) );
  NOR2_X1 U6606 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5444), .ZN(n5953) );
  INV_X1 U6607 ( .A(n5953), .ZN(n5440) );
  NAND2_X1 U6608 ( .A1(n5950), .A2(n5440), .ZN(n5443) );
  INV_X1 U6609 ( .A(n5441), .ZN(n5442) );
  AOI22_X1 U6610 ( .A1(n5443), .A2(REIP_REG_13__SCAN_IN), .B1(n5442), .B2(
        n6687), .ZN(n5446) );
  INV_X1 U6611 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6613) );
  OR3_X1 U6612 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6613), .A3(n5444), .ZN(n5445)
         );
  NAND4_X1 U6613 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(U2814)
         );
  NAND2_X1 U6614 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5974) );
  NOR3_X1 U6615 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5974), .A3(n5973), .ZN(n5455)
         );
  AOI22_X1 U6616 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6685), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5967), .ZN(n5449) );
  OAI211_X1 U6617 ( .C1(n5811), .C2(n5450), .A(n5449), .B(n5982), .ZN(n5454)
         );
  OAI22_X1 U6618 ( .A1(n6692), .A2(n5452), .B1(n5998), .B2(n5451), .ZN(n5453)
         );
  NOR3_X1 U6619 ( .A1(n5455), .A2(n5454), .A3(n5453), .ZN(n5456) );
  OAI21_X1 U6620 ( .B1(n5802), .B2(n5457), .A(n5456), .ZN(U2819) );
  INV_X1 U6621 ( .A(n5458), .ZN(n5465) );
  AOI21_X1 U6622 ( .B1(n5461), .B2(n5460), .A(n5459), .ZN(n5993) );
  OAI221_X1 U6623 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5462), .C1(n6704), .C2(
        n5993), .A(n5982), .ZN(n5463) );
  AOI21_X1 U6624 ( .B1(n6685), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5463), 
        .ZN(n5464) );
  OAI21_X1 U6625 ( .B1(n5998), .B2(n5465), .A(n5464), .ZN(n5468) );
  INV_X1 U6626 ( .A(n6005), .ZN(n5466) );
  OAI22_X1 U6627 ( .A1(n5811), .A2(n3684), .B1(n5466), .B2(n5909), .ZN(n5467)
         );
  AOI211_X1 U6628 ( .C1(n6000), .C2(n6170), .A(n5468), .B(n5467), .ZN(n5469)
         );
  OAI21_X1 U6629 ( .B1(n5981), .B2(n5470), .A(n5469), .ZN(U2823) );
  INV_X1 U6630 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5472) );
  OAI222_X1 U6631 ( .A1(n5514), .A2(n5522), .B1(n5505), .B2(n5472), .C1(n5471), 
        .C2(n5507), .ZN(U2829) );
  NOR2_X1 U6632 ( .A1(n5485), .A2(n5473), .ZN(n5474) );
  OR2_X1 U6633 ( .A1(n5475), .A2(n5474), .ZN(n5535) );
  NOR2_X1 U6634 ( .A1(n5482), .A2(n5476), .ZN(n5477) );
  OR2_X1 U6635 ( .A1(n5478), .A2(n5477), .ZN(n5776) );
  OAI22_X1 U6636 ( .A1(n5776), .A2(n5507), .B1(n6748), .B2(n5505), .ZN(n5479)
         );
  INV_X1 U6637 ( .A(n5479), .ZN(n5480) );
  OAI21_X1 U6638 ( .B1(n5535), .B2(n5514), .A(n5480), .ZN(U2831) );
  INV_X1 U6639 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5487) );
  AND2_X1 U6640 ( .A1(n5494), .A2(n5481), .ZN(n5483) );
  OR2_X1 U6641 ( .A1(n5483), .A2(n5482), .ZN(n5777) );
  AND2_X1 U6642 ( .A1(n5490), .A2(n5484), .ZN(n5486) );
  OAI222_X1 U6643 ( .A1(n5487), .A2(n5505), .B1(n5507), .B2(n5777), .C1(n5783), 
        .C2(n5514), .ZN(U2832) );
  INV_X1 U6644 ( .A(n5490), .ZN(n5491) );
  AOI21_X1 U6645 ( .B1(n5492), .B2(n5489), .A(n5491), .ZN(n5835) );
  INV_X1 U6646 ( .A(n5835), .ZN(n5789) );
  INV_X1 U6647 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5497) );
  INV_X1 U6648 ( .A(n5500), .ZN(n5496) );
  INV_X1 U6649 ( .A(n5493), .ZN(n5495) );
  OAI21_X1 U6650 ( .B1(n5496), .B2(n5495), .A(n5494), .ZN(n5788) );
  OAI222_X1 U6651 ( .A1(n5514), .A2(n5789), .B1(n5505), .B2(n5497), .C1(n5788), 
        .C2(n5507), .ZN(U2833) );
  OAI21_X1 U6652 ( .B1(n5499), .B2(n5498), .A(n5489), .ZN(n5803) );
  OAI21_X1 U6653 ( .B1(n5502), .B2(n5501), .A(n5500), .ZN(n5801) );
  INV_X1 U6654 ( .A(n5801), .ZN(n5503) );
  AOI22_X1 U6655 ( .A1(n5503), .A2(n5512), .B1(n5511), .B2(EBX_REG_25__SCAN_IN), .ZN(n5504) );
  OAI21_X1 U6656 ( .B1(n5803), .B2(n5514), .A(n5504), .ZN(U2834) );
  OAI22_X1 U6657 ( .A1(n6693), .A2(n5507), .B1(n5506), .B2(n5505), .ZN(n5508)
         );
  AOI21_X1 U6658 ( .B1(n6697), .B2(n5509), .A(n5508), .ZN(n5510) );
  INV_X1 U6659 ( .A(n5510), .ZN(U2835) );
  AOI22_X1 U6660 ( .A1(n5665), .A2(n5512), .B1(n5511), .B2(EBX_REG_23__SCAN_IN), .ZN(n5513) );
  OAI21_X1 U6661 ( .B1(n5529), .B2(n5514), .A(n5513), .ZN(U2836) );
  NAND3_X1 U6662 ( .A1(n5517), .A2(n5516), .A3(n5515), .ZN(n5519) );
  AOI22_X1 U6663 ( .A1(n6016), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6019), .ZN(n5518) );
  NAND2_X1 U6664 ( .A1(n5519), .A2(n5518), .ZN(U2860) );
  AOI22_X1 U6665 ( .A1(n6016), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6019), .ZN(n5521) );
  NAND2_X1 U6666 ( .A1(n6020), .A2(DATAI_14_), .ZN(n5520) );
  OAI211_X1 U6667 ( .C1(n5522), .C2(n5831), .A(n5521), .B(n5520), .ZN(U2861)
         );
  AOI22_X1 U6668 ( .A1(n6020), .A2(DATAI_11_), .B1(n6019), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6669 ( .A1(n6016), .A2(DATAI_27_), .ZN(n5523) );
  OAI211_X1 U6670 ( .C1(n5783), .C2(n5831), .A(n5524), .B(n5523), .ZN(U2864)
         );
  AOI22_X1 U6671 ( .A1(n6020), .A2(DATAI_9_), .B1(n6019), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6672 ( .A1(n6016), .A2(DATAI_25_), .ZN(n5525) );
  OAI211_X1 U6673 ( .C1(n5803), .C2(n5831), .A(n5526), .B(n5525), .ZN(U2866)
         );
  AOI22_X1 U6674 ( .A1(n6016), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6019), .ZN(n5528) );
  NAND2_X1 U6675 ( .A1(n6020), .A2(DATAI_7_), .ZN(n5527) );
  OAI211_X1 U6676 ( .C1(n5529), .C2(n5831), .A(n5528), .B(n5527), .ZN(U2868)
         );
  INV_X1 U6677 ( .A(n5539), .ZN(n5532) );
  OAI22_X1 U6678 ( .A1(n5532), .A2(n5531), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5530), .ZN(n5534) );
  XNOR2_X1 U6679 ( .A(n5534), .B(n5533), .ZN(n5643) );
  NAND2_X1 U6680 ( .A1(n6178), .A2(REIP_REG_28__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U6681 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5536)
         );
  OAI211_X1 U6682 ( .C1(n6110), .C2(n5769), .A(n5640), .B(n5536), .ZN(n5537)
         );
  AOI21_X1 U6683 ( .B1(n5832), .B2(n6105), .A(n5537), .ZN(n5538) );
  OAI21_X1 U6684 ( .B1(n5643), .B2(n5924), .A(n5538), .ZN(U2958) );
  INV_X1 U6685 ( .A(n3577), .ZN(n5552) );
  OAI21_X1 U6686 ( .B1(n5552), .B2(n5544), .A(n5539), .ZN(n5540) );
  XNOR2_X1 U6687 ( .A(n5540), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5650)
         );
  NAND2_X1 U6688 ( .A1(n5580), .A2(REIP_REG_27__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U6689 ( .B1(n5610), .B2(n6762), .A(n5646), .ZN(n5542) );
  NOR2_X1 U6690 ( .A1(n5783), .A2(n5590), .ZN(n5541) );
  AOI211_X1 U6691 ( .C1(n5622), .C2(n5778), .A(n5542), .B(n5541), .ZN(n5543)
         );
  OAI21_X1 U6692 ( .B1(n5650), .B2(n5924), .A(n5543), .ZN(U2959) );
  INV_X1 U6693 ( .A(n5544), .ZN(n5545) );
  NOR2_X1 U6694 ( .A1(n5546), .A2(n5545), .ZN(n5548) );
  XOR2_X1 U6695 ( .A(n5548), .B(n5547), .Z(n5656) );
  NAND2_X1 U6696 ( .A1(n6178), .A2(REIP_REG_26__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6697 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5549)
         );
  OAI211_X1 U6698 ( .C1(n6110), .C2(n5795), .A(n5653), .B(n5549), .ZN(n5550)
         );
  AOI21_X1 U6699 ( .B1(n5835), .B2(n6105), .A(n5550), .ZN(n5551) );
  OAI21_X1 U6700 ( .B1(n5656), .B2(n5924), .A(n5551), .ZN(U2960) );
  OAI21_X1 U6701 ( .B1(n5554), .B2(n5553), .A(n5552), .ZN(n5555) );
  INV_X1 U6702 ( .A(n5555), .ZN(n5663) );
  NAND2_X1 U6703 ( .A1(n5580), .A2(REIP_REG_25__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U6704 ( .B1(n5610), .B2(n5796), .A(n5659), .ZN(n5557) );
  NOR2_X1 U6705 ( .A1(n5803), .A2(n5590), .ZN(n5556) );
  AOI211_X1 U6706 ( .C1(n5622), .C2(n5799), .A(n5557), .B(n5556), .ZN(n5558)
         );
  OAI21_X1 U6707 ( .B1(n5663), .B2(n5924), .A(n5558), .ZN(U2961) );
  NAND3_X1 U6708 ( .A1(n5603), .A2(n5697), .A3(n5674), .ZN(n5560) );
  OAI21_X1 U6709 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5562) );
  XNOR2_X1 U6710 ( .A(n5562), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5672)
         );
  NAND2_X1 U6711 ( .A1(n5622), .A2(n5563), .ZN(n5564) );
  NAND2_X1 U6712 ( .A1(n6178), .A2(REIP_REG_23__SCAN_IN), .ZN(n5666) );
  OAI211_X1 U6713 ( .C1(n5610), .C2(n5565), .A(n5564), .B(n5666), .ZN(n5566)
         );
  AOI21_X1 U6714 ( .B1(n5567), .B2(n6105), .A(n5566), .ZN(n5568) );
  OAI21_X1 U6715 ( .B1(n5672), .B2(n5924), .A(n5568), .ZN(U2963) );
  AOI21_X1 U6716 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5617), .A(n5569), 
        .ZN(n5570) );
  XNOR2_X1 U6717 ( .A(n5571), .B(n5570), .ZN(n5679) );
  INV_X1 U6718 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6719 ( .A1(n5580), .A2(REIP_REG_22__SCAN_IN), .ZN(n5676) );
  OAI21_X1 U6720 ( .B1(n5610), .B2(n5572), .A(n5676), .ZN(n5574) );
  NOR2_X1 U6721 ( .A1(n5816), .A2(n5590), .ZN(n5573) );
  AOI211_X1 U6722 ( .C1(n5622), .C2(n5817), .A(n5574), .B(n5573), .ZN(n5575)
         );
  OAI21_X1 U6723 ( .B1(n5679), .B2(n5924), .A(n5575), .ZN(U2964) );
  AOI21_X1 U6724 ( .B1(n5578), .B2(n5577), .A(n5576), .ZN(n5687) );
  NAND2_X1 U6725 ( .A1(n5622), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U6726 ( .A1(n5580), .A2(REIP_REG_21__SCAN_IN), .ZN(n5681) );
  OAI211_X1 U6727 ( .C1(n5610), .C2(n6790), .A(n5581), .B(n5681), .ZN(n5582)
         );
  AOI21_X1 U6728 ( .B1(n5843), .B2(n6105), .A(n5582), .ZN(n5583) );
  OAI21_X1 U6729 ( .B1(n5687), .B2(n5924), .A(n5583), .ZN(U2965) );
  XNOR2_X1 U6730 ( .A(n5296), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5585)
         );
  XNOR2_X1 U6731 ( .A(n5584), .B(n5585), .ZN(n5696) );
  NAND2_X1 U6732 ( .A1(n5696), .A2(n3824), .ZN(n5589) );
  INV_X1 U6733 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5586) );
  NOR2_X1 U6734 ( .A1(n6193), .A2(n5586), .ZN(n5700) );
  NOR2_X1 U6735 ( .A1(n6110), .A2(n5824), .ZN(n5587) );
  AOI211_X1 U6736 ( .C1(n6099), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5700), 
        .B(n5587), .ZN(n5588) );
  OAI211_X1 U6737 ( .C1(n5590), .C2(n5823), .A(n5589), .B(n5588), .ZN(U2966)
         );
  OAI21_X1 U6738 ( .B1(n5593), .B2(n5592), .A(n5591), .ZN(n5859) );
  NAND2_X1 U6739 ( .A1(n5622), .A2(n5594), .ZN(n5595) );
  NAND2_X1 U6740 ( .A1(n6178), .A2(REIP_REG_19__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U6741 ( .C1(n5610), .C2(n6804), .A(n5595), .B(n5855), .ZN(n5596)
         );
  AOI21_X1 U6742 ( .B1(n5597), .B2(n6105), .A(n5596), .ZN(n5598) );
  OAI21_X1 U6743 ( .B1(n5859), .B2(n5924), .A(n5598), .ZN(U2967) );
  NAND2_X1 U6744 ( .A1(n5599), .A2(n5600), .ZN(n5616) );
  OR3_X1 U6745 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5850) );
  INV_X1 U6746 ( .A(n5850), .ZN(n5601) );
  AOI22_X1 U6747 ( .A1(n5616), .A2(n5601), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n3558), .ZN(n5849) );
  INV_X1 U6748 ( .A(n5851), .ZN(n5606) );
  NOR2_X1 U6749 ( .A1(n5603), .A2(n3569), .ZN(n5620) );
  XNOR2_X1 U6750 ( .A(n3558), .B(n5690), .ZN(n5604) );
  OAI21_X1 U6751 ( .B1(n5606), .B2(n5620), .A(n5604), .ZN(n5605) );
  OAI21_X1 U6752 ( .B1(n5849), .B2(n5606), .A(n5605), .ZN(n5873) );
  NAND2_X1 U6753 ( .A1(n5873), .A2(n3824), .ZN(n5614) );
  INV_X1 U6754 ( .A(n5607), .ZN(n5612) );
  INV_X1 U6755 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5608) );
  OAI22_X1 U6756 ( .A1(n5610), .A2(n5609), .B1(n6193), .B2(n5608), .ZN(n5611)
         );
  AOI21_X1 U6757 ( .B1(n5612), .B2(n5622), .A(n5611), .ZN(n5613) );
  OAI211_X1 U6758 ( .C1(n5590), .C2(n5615), .A(n5614), .B(n5613), .ZN(U2969)
         );
  INV_X1 U6759 ( .A(n5616), .ZN(n5619) );
  AOI21_X1 U6760 ( .B1(n3569), .B2(n5617), .A(n5620), .ZN(n5618) );
  OAI22_X1 U6761 ( .A1(n5620), .A2(n5851), .B1(n5619), .B2(n5618), .ZN(n5882)
         );
  AOI22_X1 U6762 ( .A1(n6099), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6178), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U6763 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  OAI211_X1 U6764 ( .C1(n6015), .C2(n5590), .A(n5624), .B(n5623), .ZN(n5625)
         );
  INV_X1 U6765 ( .A(n5625), .ZN(n5626) );
  OAI21_X1 U6766 ( .B1(n5882), .B2(n5924), .A(n5626), .ZN(U2970) );
  NAND3_X1 U6767 ( .A1(n5644), .A2(n5628), .A3(n5627), .ZN(n5629) );
  OAI211_X1 U6768 ( .C1(n5631), .C2(n6195), .A(n5630), .B(n5629), .ZN(n5632)
         );
  AOI21_X1 U6769 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5633), .A(n5632), 
        .ZN(n5634) );
  OAI21_X1 U6770 ( .B1(n5635), .B2(n5881), .A(n5634), .ZN(U2989) );
  INV_X1 U6771 ( .A(n5636), .ZN(n5648) );
  NAND3_X1 U6772 ( .A1(n5644), .A2(n5638), .A3(n5637), .ZN(n5639) );
  OAI211_X1 U6773 ( .C1(n5776), .C2(n6195), .A(n5640), .B(n5639), .ZN(n5641)
         );
  AOI21_X1 U6774 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5648), .A(n5641), 
        .ZN(n5642) );
  OAI21_X1 U6775 ( .B1(n5643), .B2(n5881), .A(n5642), .ZN(U2990) );
  NAND2_X1 U6776 ( .A1(n5644), .A2(n6738), .ZN(n5645) );
  OAI211_X1 U6777 ( .C1(n5777), .C2(n6195), .A(n5646), .B(n5645), .ZN(n5647)
         );
  AOI21_X1 U6778 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5648), .A(n5647), 
        .ZN(n5649) );
  OAI21_X1 U6779 ( .B1(n5650), .B2(n5881), .A(n5649), .ZN(U2991) );
  OAI211_X1 U6780 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5657), .B(n5651), .ZN(n5652) );
  OAI211_X1 U6781 ( .C1(n5788), .C2(n6195), .A(n5653), .B(n5652), .ZN(n5654)
         );
  AOI21_X1 U6782 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5661), .A(n5654), 
        .ZN(n5655) );
  OAI21_X1 U6783 ( .B1(n5656), .B2(n5881), .A(n5655), .ZN(U2992) );
  NAND2_X1 U6784 ( .A1(n5657), .A2(n6913), .ZN(n5658) );
  OAI211_X1 U6785 ( .C1(n5801), .C2(n6195), .A(n5659), .B(n5658), .ZN(n5660)
         );
  AOI21_X1 U6786 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5661), .A(n5660), 
        .ZN(n5662) );
  OAI21_X1 U6787 ( .B1(n5663), .B2(n5881), .A(n5662), .ZN(U2993) );
  INV_X1 U6788 ( .A(n5664), .ZN(n5668) );
  NAND2_X1 U6789 ( .A1(n5665), .A2(n6180), .ZN(n5667) );
  OAI211_X1 U6790 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5668), .A(n5667), .B(n5666), .ZN(n5669) );
  AOI21_X1 U6791 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5670), .A(n5669), 
        .ZN(n5671) );
  OAI21_X1 U6792 ( .B1(n5672), .B2(n5881), .A(n5671), .ZN(U2995) );
  OR3_X1 U6793 ( .A1(n5682), .A2(n5674), .A3(n5673), .ZN(n5675) );
  OAI211_X1 U6794 ( .C1(n5820), .C2(n6195), .A(n5676), .B(n5675), .ZN(n5677)
         );
  AOI21_X1 U6795 ( .B1(n5685), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5677), 
        .ZN(n5678) );
  OAI21_X1 U6796 ( .B1(n5679), .B2(n5881), .A(n5678), .ZN(U2996) );
  NOR2_X1 U6797 ( .A1(n5680), .A2(n6195), .ZN(n5684) );
  OAI21_X1 U6798 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5682), .A(n5681), 
        .ZN(n5683) );
  AOI211_X1 U6799 ( .C1(n5685), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5684), .B(n5683), .ZN(n5686) );
  OAI21_X1 U6800 ( .B1(n5687), .B2(n5881), .A(n5686), .ZN(U2997) );
  OAI21_X1 U6801 ( .B1(n5690), .B2(n5689), .A(n5688), .ZN(n5691) );
  OAI21_X1 U6802 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n5871) );
  NOR2_X1 U6803 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6160), .ZN(n5694)
         );
  NOR2_X1 U6804 ( .A1(n5871), .A2(n5694), .ZN(n5864) );
  NAND2_X1 U6805 ( .A1(n5878), .A2(n5865), .ZN(n5695) );
  AND2_X1 U6806 ( .A1(n5864), .A2(n5695), .ZN(n5858) );
  NAND2_X1 U6807 ( .A1(n5696), .A2(n6190), .ZN(n5702) );
  NOR3_X1 U6808 ( .A1(n5863), .A2(n5698), .A3(n5697), .ZN(n5699) );
  AOI211_X1 U6809 ( .C1(n5826), .C2(n6180), .A(n5700), .B(n5699), .ZN(n5701)
         );
  OAI211_X1 U6810 ( .C1(n5858), .C2(n5703), .A(n5702), .B(n5701), .ZN(U2998)
         );
  INV_X1 U6811 ( .A(n5704), .ZN(n5713) );
  OAI21_X1 U6812 ( .B1(n6195), .B2(n5706), .A(n5705), .ZN(n5707) );
  AOI21_X1 U6813 ( .B1(n6190), .B2(n5708), .A(n5707), .ZN(n5712) );
  OAI21_X1 U6814 ( .B1(n5710), .B2(n5709), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5711) );
  NAND3_X1 U6815 ( .A1(n5713), .A2(n5712), .A3(n5711), .ZN(U3018) );
  OAI211_X1 U6816 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4585), .A(n6203), .B(
        n6447), .ZN(n5714) );
  OAI21_X1 U6817 ( .B1(n5716), .B2(n5715), .A(n5714), .ZN(n5718) );
  MUX2_X1 U6818 ( .A(n5718), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n5717), 
        .Z(U3464) );
  INV_X1 U6819 ( .A(n5719), .ZN(n5722) );
  INV_X1 U6820 ( .A(n5720), .ZN(n5721) );
  OAI22_X1 U6821 ( .A1(n5722), .A2(n6661), .B1(n5721), .B2(n6558), .ZN(n5723)
         );
  MUX2_X1 U6822 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5723), .S(n6659), 
        .Z(U3456) );
  NOR3_X1 U6823 ( .A1(n6289), .A2(n4585), .A3(n6353), .ZN(n5724) );
  NOR2_X1 U6824 ( .A1(n5724), .A2(n6401), .ZN(n6247) );
  OR2_X1 U6825 ( .A1(n6454), .A2(n5725), .ZN(n6246) );
  INV_X1 U6826 ( .A(n6246), .ZN(n5726) );
  NAND3_X1 U6827 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6397), .A3(n6534), .ZN(n6243) );
  NOR2_X1 U6828 ( .A1(n6355), .A2(n6243), .ZN(n5759) );
  AOI21_X1 U6829 ( .B1(n5726), .B2(n6528), .A(n5759), .ZN(n5729) );
  INV_X1 U6830 ( .A(n6243), .ZN(n5727) );
  OAI21_X1 U6831 ( .B1(n6447), .B2(n5727), .A(n6406), .ZN(n5728) );
  AOI21_X1 U6832 ( .B1(n6247), .B2(n5729), .A(n5728), .ZN(n5765) );
  INV_X1 U6833 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5734) );
  INV_X1 U6834 ( .A(n6247), .ZN(n5730) );
  OAI22_X1 U6835 ( .A1(n5730), .A2(n5729), .B1(n6243), .B2(n6568), .ZN(n5762)
         );
  AOI22_X1 U6836 ( .A1(n6456), .A2(n5759), .B1(n6267), .B2(n6399), .ZN(n5731)
         );
  OAI21_X1 U6837 ( .B1(n6460), .B2(n6275), .A(n5731), .ZN(n5732) );
  AOI21_X1 U6838 ( .B1(n5762), .B2(n6457), .A(n5732), .ZN(n5733) );
  OAI21_X1 U6839 ( .B1(n5765), .B2(n5734), .A(n5733), .ZN(U3060) );
  INV_X1 U6840 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5738) );
  AOI22_X1 U6841 ( .A1(n6464), .A2(n5759), .B1(n6267), .B2(n6367), .ZN(n5735)
         );
  OAI21_X1 U6842 ( .B1(n6468), .B2(n6275), .A(n5735), .ZN(n5736) );
  AOI21_X1 U6843 ( .B1(n5762), .B2(n6465), .A(n5736), .ZN(n5737) );
  OAI21_X1 U6844 ( .B1(n5765), .B2(n5738), .A(n5737), .ZN(U3061) );
  INV_X1 U6845 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5742) );
  AOI22_X1 U6846 ( .A1(n6472), .A2(n5759), .B1(n6267), .B2(n6370), .ZN(n5739)
         );
  OAI21_X1 U6847 ( .B1(n6474), .B2(n6275), .A(n5739), .ZN(n5740) );
  AOI21_X1 U6848 ( .B1(n5762), .B2(n6473), .A(n5740), .ZN(n5741) );
  OAI21_X1 U6849 ( .B1(n5765), .B2(n5742), .A(n5741), .ZN(U3062) );
  INV_X1 U6850 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5746) );
  AOI22_X1 U6851 ( .A1(n6480), .A2(n5759), .B1(n6267), .B2(n6420), .ZN(n5743)
         );
  OAI21_X1 U6852 ( .B1(n6482), .B2(n6275), .A(n5743), .ZN(n5744) );
  AOI21_X1 U6853 ( .B1(n5762), .B2(n6481), .A(n5744), .ZN(n5745) );
  OAI21_X1 U6854 ( .B1(n5765), .B2(n5746), .A(n5745), .ZN(U3063) );
  INV_X1 U6855 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5750) );
  AOI22_X1 U6856 ( .A1(n6488), .A2(n5759), .B1(n6267), .B2(n6377), .ZN(n5747)
         );
  OAI21_X1 U6857 ( .B1(n6490), .B2(n6275), .A(n5747), .ZN(n5748) );
  AOI21_X1 U6858 ( .B1(n5762), .B2(n6489), .A(n5748), .ZN(n5749) );
  OAI21_X1 U6859 ( .B1(n5765), .B2(n5750), .A(n5749), .ZN(U3064) );
  INV_X1 U6860 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5754) );
  AOI22_X1 U6861 ( .A1(n6496), .A2(n5759), .B1(n6267), .B2(n6380), .ZN(n5751)
         );
  OAI21_X1 U6862 ( .B1(n6498), .B2(n6275), .A(n5751), .ZN(n5752) );
  AOI21_X1 U6863 ( .B1(n5762), .B2(n6497), .A(n5752), .ZN(n5753) );
  OAI21_X1 U6864 ( .B1(n5765), .B2(n5754), .A(n5753), .ZN(U3065) );
  INV_X1 U6865 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5758) );
  AOI22_X1 U6866 ( .A1(n6504), .A2(n5759), .B1(n6267), .B2(n6383), .ZN(n5755)
         );
  OAI21_X1 U6867 ( .B1(n6506), .B2(n6275), .A(n5755), .ZN(n5756) );
  AOI21_X1 U6868 ( .B1(n5762), .B2(n6505), .A(n5756), .ZN(n5757) );
  OAI21_X1 U6869 ( .B1(n5765), .B2(n5758), .A(n5757), .ZN(U3066) );
  INV_X1 U6870 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5764) );
  AOI22_X1 U6871 ( .A1(n6513), .A2(n5759), .B1(n6267), .B2(n6388), .ZN(n5760)
         );
  OAI21_X1 U6872 ( .B1(n6517), .B2(n6275), .A(n5760), .ZN(n5761) );
  AOI21_X1 U6873 ( .B1(n5762), .B2(n6515), .A(n5761), .ZN(n5763) );
  OAI21_X1 U6874 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(U3067) );
  AND2_X1 U6875 ( .A1(n6039), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6876 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5767), .A(n5766), .ZN(
        n5768) );
  INV_X1 U6877 ( .A(n5768), .ZN(U2788) );
  INV_X1 U6878 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6778) );
  OAI22_X1 U6879 ( .A1(n4276), .A2(n5977), .B1(n5998), .B2(n5769), .ZN(n5770)
         );
  AOI21_X1 U6880 ( .B1(n6686), .B2(EBX_REG_28__SCAN_IN), .A(n5770), .ZN(n5771)
         );
  OAI21_X1 U6881 ( .B1(n5772), .B2(n6778), .A(n5771), .ZN(n5773) );
  AOI21_X1 U6882 ( .B1(n5832), .B2(n6696), .A(n5773), .ZN(n5775) );
  INV_X1 U6883 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6634) );
  OR3_X1 U6884 ( .A1(n6634), .A2(n5787), .A3(REIP_REG_28__SCAN_IN), .ZN(n5774)
         );
  OAI211_X1 U6885 ( .C1(n6692), .C2(n5776), .A(n5775), .B(n5774), .ZN(U2799)
         );
  INV_X1 U6886 ( .A(n5777), .ZN(n5785) );
  INV_X1 U6887 ( .A(n5778), .ZN(n5779) );
  OAI22_X1 U6888 ( .A1(n6762), .A2(n5977), .B1(n5998), .B2(n5779), .ZN(n5780)
         );
  AOI21_X1 U6889 ( .B1(n6686), .B2(EBX_REG_27__SCAN_IN), .A(n5780), .ZN(n5782)
         );
  NAND2_X1 U6890 ( .A1(n5792), .A2(REIP_REG_27__SCAN_IN), .ZN(n5781) );
  OAI211_X1 U6891 ( .C1(n5783), .C2(n5802), .A(n5782), .B(n5781), .ZN(n5784)
         );
  AOI21_X1 U6892 ( .B1(n5785), .B2(n6000), .A(n5784), .ZN(n5786) );
  OAI21_X1 U6893 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5787), .A(n5786), .ZN(U2800) );
  AOI22_X1 U6894 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6686), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6685), .ZN(n5794) );
  OAI22_X1 U6895 ( .A1(n5789), .A2(n5802), .B1(n5788), .B2(n6692), .ZN(n5790)
         );
  AOI221_X1 U6896 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5792), .C1(n5791), .C2(
        n5792), .A(n5790), .ZN(n5793) );
  OAI211_X1 U6897 ( .C1(n5795), .C2(n5998), .A(n5794), .B(n5793), .ZN(U2801)
         );
  OAI22_X1 U6898 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5797), .B1(n5796), .B2(
        n5977), .ZN(n5798) );
  AOI21_X1 U6899 ( .B1(n5799), .B2(n6687), .A(n5798), .ZN(n5806) );
  AND2_X1 U6900 ( .A1(n5800), .A2(n6925), .ZN(n6695) );
  OAI22_X1 U6901 ( .A1(n5803), .A2(n5802), .B1(n5801), .B2(n6692), .ZN(n5804)
         );
  AOI221_X1 U6902 ( .B1(n6695), .B2(REIP_REG_25__SCAN_IN), .C1(n6689), .C2(
        REIP_REG_25__SCAN_IN), .A(n5804), .ZN(n5805) );
  OAI211_X1 U6903 ( .C1(n5807), .C2(n5811), .A(n5806), .B(n5805), .ZN(U2802)
         );
  INV_X1 U6904 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6628) );
  OAI22_X1 U6905 ( .A1(n5810), .A2(n5809), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5808), .ZN(n5814) );
  OAI22_X1 U6906 ( .A1(n5812), .A2(n5811), .B1(n5572), .B2(n5977), .ZN(n5813)
         );
  AOI221_X1 U6907 ( .B1(n5815), .B2(n6628), .C1(n5814), .C2(
        REIP_REG_22__SCAN_IN), .A(n5813), .ZN(n5819) );
  INV_X1 U6908 ( .A(n5816), .ZN(n5840) );
  AOI22_X1 U6909 ( .A1(n5840), .A2(n6696), .B1(n5817), .B2(n6687), .ZN(n5818)
         );
  OAI211_X1 U6910 ( .C1(n5820), .C2(n6692), .A(n5819), .B(n5818), .ZN(U2805)
         );
  AOI21_X1 U6911 ( .B1(n5821), .B2(n5942), .A(REIP_REG_20__SCAN_IN), .ZN(n5830) );
  INV_X1 U6912 ( .A(n5822), .ZN(n5829) );
  AOI22_X1 U6913 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6686), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6685), .ZN(n5828) );
  INV_X1 U6914 ( .A(n5823), .ZN(n5846) );
  INV_X1 U6915 ( .A(n5824), .ZN(n5825) );
  AOI222_X1 U6916 ( .A1(n5826), .A2(n6000), .B1(n5846), .B2(n6696), .C1(n5825), 
        .C2(n6687), .ZN(n5827) );
  OAI211_X1 U6917 ( .C1(n5830), .C2(n5829), .A(n5828), .B(n5827), .ZN(U2807)
         );
  INV_X1 U6918 ( .A(n5831), .ZN(n6017) );
  AOI22_X1 U6919 ( .A1(n5832), .A2(n6017), .B1(n6016), .B2(DATAI_28_), .ZN(
        n5834) );
  AOI22_X1 U6920 ( .A1(n6020), .A2(DATAI_12_), .B1(n6019), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6921 ( .A1(n5834), .A2(n5833), .ZN(U2863) );
  AOI22_X1 U6922 ( .A1(n5835), .A2(n6017), .B1(n6016), .B2(DATAI_26_), .ZN(
        n5837) );
  AOI22_X1 U6923 ( .A1(n6020), .A2(DATAI_10_), .B1(n6019), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6924 ( .A1(n5837), .A2(n5836), .ZN(U2865) );
  AOI22_X1 U6925 ( .A1(n6697), .A2(n6017), .B1(DATAI_24_), .B2(n6016), .ZN(
        n5839) );
  AOI22_X1 U6926 ( .A1(n6020), .A2(DATAI_8_), .B1(n6019), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U6927 ( .A1(n5839), .A2(n5838), .ZN(U2867) );
  AOI22_X1 U6928 ( .A1(n5840), .A2(n6017), .B1(n6016), .B2(DATAI_22_), .ZN(
        n5842) );
  AOI22_X1 U6929 ( .A1(n6020), .A2(DATAI_6_), .B1(n6019), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U6930 ( .A1(n5842), .A2(n5841), .ZN(U2869) );
  AOI22_X1 U6931 ( .A1(n5843), .A2(n6017), .B1(n6016), .B2(DATAI_21_), .ZN(
        n5845) );
  AOI22_X1 U6932 ( .A1(n6020), .A2(DATAI_5_), .B1(n6019), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U6933 ( .A1(n5845), .A2(n5844), .ZN(U2870) );
  AOI22_X1 U6934 ( .A1(n5846), .A2(n6017), .B1(n6016), .B2(DATAI_20_), .ZN(
        n5848) );
  AOI22_X1 U6935 ( .A1(n6020), .A2(DATAI_4_), .B1(n6019), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6936 ( .A1(n5848), .A2(n5847), .ZN(U2871) );
  AOI22_X1 U6937 ( .A1(n6178), .A2(REIP_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6099), .ZN(n5854) );
  AOI21_X1 U6938 ( .B1(n5851), .B2(n5850), .A(n5849), .ZN(n5852) );
  XNOR2_X1 U6939 ( .A(n5852), .B(n5865), .ZN(n5867) );
  AOI22_X1 U6940 ( .A1(n5867), .A2(n3824), .B1(n6105), .B2(n6012), .ZN(n5853)
         );
  OAI211_X1 U6941 ( .C1(n6110), .C2(n5949), .A(n5854), .B(n5853), .ZN(U2968)
         );
  INV_X1 U6942 ( .A(n5855), .ZN(n5856) );
  AOI21_X1 U6943 ( .B1(n5857), .B2(n6180), .A(n5856), .ZN(n5862) );
  OAI22_X1 U6944 ( .A1(n5859), .A2(n5881), .B1(n5858), .B2(n6702), .ZN(n5860)
         );
  INV_X1 U6945 ( .A(n5860), .ZN(n5861) );
  OAI211_X1 U6946 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5863), .A(n5862), .B(n5861), .ZN(U2999) );
  NAND2_X1 U6947 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5865), .ZN(n5870) );
  OAI22_X1 U6948 ( .A1(n5865), .A2(n5864), .B1(n6193), .B2(n6620), .ZN(n5866)
         );
  INV_X1 U6949 ( .A(n5866), .ZN(n5869) );
  AOI22_X1 U6950 ( .A1(n5867), .A2(n6190), .B1(n6180), .B2(n5946), .ZN(n5868)
         );
  OAI211_X1 U6951 ( .C1(n5876), .C2(n5870), .A(n5869), .B(n5868), .ZN(U3000)
         );
  AOI22_X1 U6952 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5871), .B1(n6178), .B2(REIP_REG_17__SCAN_IN), .ZN(n5875) );
  AOI22_X1 U6953 ( .A1(n5873), .A2(n6190), .B1(n6180), .B2(n5872), .ZN(n5874)
         );
  OAI211_X1 U6954 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5876), .A(n5875), .B(n5874), .ZN(U3001) );
  AND2_X1 U6955 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  OR2_X1 U6956 ( .A1(n6111), .A2(n5879), .ZN(n5888) );
  OAI22_X1 U6957 ( .A1(n5880), .A2(n6195), .B1(n6912), .B2(n6193), .ZN(n5884)
         );
  NOR2_X1 U6958 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  AOI211_X1 U6959 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5888), .A(n5884), .B(n5883), .ZN(n5887) );
  OAI211_X1 U6960 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5892), .B(n5885), .ZN(n5886) );
  NAND2_X1 U6961 ( .A1(n5887), .A2(n5886), .ZN(U3002) );
  INV_X1 U6962 ( .A(n5888), .ZN(n5896) );
  INV_X1 U6963 ( .A(n5889), .ZN(n5891) );
  AOI21_X1 U6964 ( .B1(n5891), .B2(n6180), .A(n5890), .ZN(n5895) );
  AOI22_X1 U6965 ( .A1(n5893), .A2(n6190), .B1(n5892), .B2(n6760), .ZN(n5894)
         );
  OAI211_X1 U6966 ( .C1(n5896), .C2(n6760), .A(n5895), .B(n5894), .ZN(U3003)
         );
  INV_X1 U6967 ( .A(n5897), .ZN(n5900) );
  INV_X1 U6968 ( .A(n5898), .ZN(n5899) );
  AOI21_X1 U6969 ( .B1(n5900), .B2(n6180), .A(n5899), .ZN(n5907) );
  OAI21_X1 U6970 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(n5904) );
  AOI22_X1 U6971 ( .A1(n5905), .A2(n6190), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5904), .ZN(n5906) );
  OAI211_X1 U6972 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n5908), .A(n5907), .B(n5906), .ZN(U3004) );
  INV_X1 U6973 ( .A(n5909), .ZN(n5913) );
  INV_X1 U6974 ( .A(n5910), .ZN(n5911) );
  NAND3_X1 U6975 ( .A1(n5913), .A2(n5912), .A3(n5911), .ZN(n5914) );
  OAI22_X1 U6976 ( .A1(n5915), .A2(n5914), .B1(n4577), .B2(n6659), .ZN(U3455)
         );
  AOI21_X1 U6977 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6595), .A(n6588), .ZN(n5922) );
  INV_X1 U6978 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5916) );
  NAND2_X1 U6979 ( .A1(n6588), .A2(STATE_REG_1__SCAN_IN), .ZN(n6684) );
  INV_X1 U6980 ( .A(n6684), .ZN(n6594) );
  AOI21_X1 U6981 ( .B1(n5922), .B2(n5916), .A(n6594), .ZN(U2789) );
  NAND2_X1 U6982 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6679), .ZN(n5920) );
  OAI21_X1 U6983 ( .B1(n5918), .B2(n5917), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5919) );
  OAI21_X1 U6984 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5920), .A(n5919), .ZN(
        U2790) );
  INV_X1 U6985 ( .A(n6594), .ZN(n6674) );
  NOR2_X1 U6986 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5923) );
  OAI21_X1 U6987 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5923), .A(n6684), .ZN(n5921)
         );
  OAI21_X1 U6988 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6674), .A(n5921), .ZN(
        U2791) );
  NOR2_X1 U6989 ( .A1(n6594), .A2(n5922), .ZN(n6650) );
  OAI21_X1 U6990 ( .B1(n5923), .B2(BS16_N), .A(n6650), .ZN(n6648) );
  OAI21_X1 U6991 ( .B1(n6650), .B2(n6353), .A(n6648), .ZN(U2792) );
  OAI21_X1 U6992 ( .B1(n5926), .B2(n5925), .A(n5924), .ZN(U2793) );
  NOR4_X1 U6993 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5936) );
  NOR4_X1 U6994 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5935) );
  INV_X1 U6995 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6649) );
  INV_X1 U6996 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6668) );
  NOR4_X1 U6997 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6998 ( .B1(n6649), .B2(n6668), .A(n5927), .ZN(n5933) );
  NOR4_X1 U6999 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5931) );
  NOR4_X1 U7000 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5930) );
  NOR4_X1 U7001 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5929) );
  NOR4_X1 U7002 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5928) );
  NAND4_X1 U7003 ( .A1(n5931), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n5932)
         );
  NOR4_X1 U7004 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_22__SCAN_IN), .A3(n5933), .A4(n5932), .ZN(n5934) );
  NAND3_X1 U7005 ( .A1(n5936), .A2(n5935), .A3(n5934), .ZN(n5938) );
  NOR2_X1 U7006 ( .A1(REIP_REG_1__SCAN_IN), .A2(n5938), .ZN(n5939) );
  INV_X1 U7007 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5937) );
  NOR2_X1 U7008 ( .A1(REIP_REG_0__SCAN_IN), .A2(n5938), .ZN(n6663) );
  NAND3_X1 U7009 ( .A1(n6663), .A2(n6649), .A3(n6668), .ZN(n5940) );
  OAI221_X1 U7010 ( .B1(n5939), .B2(n5937), .C1(n5939), .C2(n5938), .A(n5940), 
        .ZN(U2794) );
  INV_X1 U7011 ( .A(n5938), .ZN(n6671) );
  INV_X1 U7012 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7013 ( .A1(n5939), .A2(n6649), .ZN(n6669) );
  OAI211_X1 U7014 ( .C1(n6671), .C2(n5941), .A(n5940), .B(n6669), .ZN(U2795)
         );
  AOI22_X1 U7015 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6686), .B1(n5942), .B2(n6620), .ZN(n5943) );
  OAI21_X1 U7016 ( .B1(n5944), .B2(n6620), .A(n5943), .ZN(n5945) );
  AOI211_X1 U7017 ( .C1(n6685), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5964), 
        .B(n5945), .ZN(n5948) );
  AOI22_X1 U7018 ( .A1(n6012), .A2(n6696), .B1(n5946), .B2(n6000), .ZN(n5947)
         );
  OAI211_X1 U7019 ( .C1(n5949), .C2(n5998), .A(n5948), .B(n5947), .ZN(U2809)
         );
  INV_X1 U7020 ( .A(n5950), .ZN(n5951) );
  AOI22_X1 U7021 ( .A1(n6000), .A2(n5952), .B1(REIP_REG_12__SCAN_IN), .B2(
        n5951), .ZN(n5959) );
  AOI211_X1 U7022 ( .C1(n6685), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5964), 
        .B(n5953), .ZN(n5958) );
  AOI22_X1 U7023 ( .A1(n5955), .A2(n6696), .B1(n6687), .B2(n5954), .ZN(n5957)
         );
  NAND2_X1 U7024 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6686), .ZN(n5956) );
  NAND4_X1 U7025 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(U2815)
         );
  AOI22_X1 U7026 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6686), .B1(n6000), .B2(n5960), .ZN(n5972) );
  NOR3_X1 U7027 ( .A1(n5962), .A2(REIP_REG_10__SCAN_IN), .A3(n5961), .ZN(n5963) );
  AOI211_X1 U7028 ( .C1(n6685), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5964), 
        .B(n5963), .ZN(n5971) );
  AOI22_X1 U7029 ( .A1(n5966), .A2(n6696), .B1(n6687), .B2(n5965), .ZN(n5970)
         );
  OAI21_X1 U7030 ( .B1(n5968), .B2(n5967), .A(REIP_REG_10__SCAN_IN), .ZN(n5969) );
  NAND4_X1 U7031 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(U2817)
         );
  INV_X1 U7032 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6606) );
  INV_X1 U7033 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6604) );
  AOI21_X1 U7034 ( .B1(n6606), .B2(n6604), .A(n5973), .ZN(n5975) );
  AOI22_X1 U7035 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5985), .B1(n5975), .B2(n5974), .ZN(n5980) );
  AOI22_X1 U7036 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6686), .B1(n6000), .B2(n6136), 
        .ZN(n5976) );
  OAI211_X1 U7037 ( .C1(n5977), .C2(n3828), .A(n5976), .B(n5982), .ZN(n5978)
         );
  AOI21_X1 U7038 ( .B1(n6079), .B2(n6696), .A(n5978), .ZN(n5979) );
  OAI211_X1 U7039 ( .C1(n6082), .C2(n5998), .A(n5980), .B(n5979), .ZN(U2820)
         );
  AOI22_X1 U7040 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6686), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6685), .ZN(n5983) );
  OAI211_X1 U7041 ( .C1(n6692), .C2(n6159), .A(n5983), .B(n5982), .ZN(n5984)
         );
  AOI21_X1 U7042 ( .B1(n6087), .B2(n6002), .A(n5984), .ZN(n5988) );
  OAI21_X1 U7043 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5986), .A(n5985), .ZN(n5987)
         );
  OAI211_X1 U7044 ( .C1(n5998), .C2(n6090), .A(n5988), .B(n5987), .ZN(U2822)
         );
  AOI22_X1 U7045 ( .A1(n6179), .A2(n6000), .B1(n6686), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5992) );
  NAND2_X1 U7046 ( .A1(n6002), .A2(n6095), .ZN(n5991) );
  AOI22_X1 U7047 ( .A1(n6005), .A2(n5989), .B1(n6685), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5990) );
  AND3_X1 U7048 ( .A1(n5992), .A2(n5991), .A3(n5990), .ZN(n5997) );
  INV_X1 U7049 ( .A(n5993), .ZN(n5994) );
  OAI21_X1 U7050 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5995), .A(n5994), .ZN(n5996)
         );
  OAI211_X1 U7051 ( .C1(n5998), .C2(n6098), .A(n5997), .B(n5996), .ZN(U2824)
         );
  AOI21_X1 U7052 ( .B1(n6685), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5999), 
        .ZN(n6010) );
  AOI22_X1 U7053 ( .A1(n6000), .A2(n4427), .B1(n6686), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6008) );
  NAND2_X1 U7054 ( .A1(n6002), .A2(n6001), .ZN(n6007) );
  INV_X1 U7055 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6003) );
  AOI22_X1 U7056 ( .A1(n6005), .A2(n6004), .B1(n6687), .B2(n6003), .ZN(n6006)
         );
  AND3_X1 U7057 ( .A1(n6008), .A2(n6007), .A3(n6006), .ZN(n6009) );
  OAI211_X1 U7058 ( .C1(n6011), .C2(n6664), .A(n6010), .B(n6009), .ZN(U2826)
         );
  AOI22_X1 U7059 ( .A1(n6012), .A2(n6017), .B1(n6016), .B2(DATAI_18_), .ZN(
        n6014) );
  AOI22_X1 U7060 ( .A1(n6020), .A2(DATAI_2_), .B1(n6019), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7061 ( .A1(n6014), .A2(n6013), .ZN(U2873) );
  INV_X1 U7062 ( .A(n6015), .ZN(n6018) );
  AOI22_X1 U7063 ( .A1(n6018), .A2(n6017), .B1(n6016), .B2(DATAI_16_), .ZN(
        n6022) );
  AOI22_X1 U7064 ( .A1(n6020), .A2(DATAI_0_), .B1(n6019), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7065 ( .A1(n6022), .A2(n6021), .ZN(U2875) );
  AOI22_X1 U7066 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7067 ( .B1(n4550), .B2(n6051), .A(n6024), .ZN(U2908) );
  AOI22_X1 U7068 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7069 ( .B1(n6026), .B2(n6051), .A(n6025), .ZN(U2909) );
  INV_X1 U7070 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6028) );
  AOI22_X1 U7071 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7072 ( .B1(n6028), .B2(n6051), .A(n6027), .ZN(U2910) );
  INV_X1 U7073 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6030) );
  AOI22_X1 U7074 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7075 ( .B1(n6030), .B2(n6051), .A(n6029), .ZN(U2911) );
  INV_X1 U7076 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U7077 ( .A1(DATAO_REG_11__SCAN_IN), .A2(n6049), .B1(
        LWORD_REG_11__SCAN_IN), .B2(n6677), .ZN(n6031) );
  OAI21_X1 U7078 ( .B1(n6032), .B2(n6051), .A(n6031), .ZN(U2912) );
  AOI22_X1 U7079 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U7080 ( .B1(n4442), .B2(n6051), .A(n6033), .ZN(U2913) );
  INV_X1 U7081 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6035) );
  AOI22_X1 U7082 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7083 ( .B1(n6035), .B2(n6051), .A(n6034), .ZN(U2914) );
  INV_X1 U7084 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6037) );
  AOI22_X1 U7085 ( .A1(DATAO_REG_8__SCAN_IN), .A2(n6049), .B1(
        LWORD_REG_8__SCAN_IN), .B2(n6677), .ZN(n6036) );
  OAI21_X1 U7086 ( .B1(n6037), .B2(n6051), .A(n6036), .ZN(U2915) );
  AOI22_X1 U7087 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7088 ( .B1(n3829), .B2(n6051), .A(n6038), .ZN(U2916) );
  AOI22_X1 U7089 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6677), .B1(n6039), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U7090 ( .B1(n3954), .B2(n6051), .A(n6040), .ZN(U2917) );
  AOI22_X1 U7091 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7092 ( .B1(n3948), .B2(n6051), .A(n6041), .ZN(U2918) );
  AOI22_X1 U7093 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U7094 ( .B1(n6043), .B2(n6051), .A(n6042), .ZN(U2919) );
  AOI22_X1 U7095 ( .A1(DATAO_REG_3__SCAN_IN), .A2(n6049), .B1(
        LWORD_REG_3__SCAN_IN), .B2(n6677), .ZN(n6044) );
  OAI21_X1 U7096 ( .B1(n6045), .B2(n6051), .A(n6044), .ZN(U2920) );
  AOI22_X1 U7097 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6046) );
  OAI21_X1 U7098 ( .B1(n4454), .B2(n6051), .A(n6046), .ZN(U2921) );
  AOI22_X1 U7099 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6047) );
  OAI21_X1 U7100 ( .B1(n6048), .B2(n6051), .A(n6047), .ZN(U2922) );
  AOI22_X1 U7101 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6677), .B1(n6049), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6050) );
  OAI21_X1 U7102 ( .B1(n4444), .B2(n6051), .A(n6050), .ZN(U2923) );
  INV_X1 U7103 ( .A(n6052), .ZN(n6061) );
  NAND2_X1 U7104 ( .A1(n6061), .A2(DATAI_8_), .ZN(n6063) );
  INV_X1 U7105 ( .A(n6063), .ZN(n6053) );
  AOI21_X1 U7106 ( .B1(n6071), .B2(UWORD_REG_8__SCAN_IN), .A(n6053), .ZN(n6054) );
  OAI21_X1 U7107 ( .B1(n7002), .B2(n6060), .A(n6054), .ZN(U2932) );
  NAND2_X1 U7108 ( .A1(n6061), .A2(DATAI_9_), .ZN(n6065) );
  INV_X1 U7109 ( .A(n6065), .ZN(n6055) );
  AOI21_X1 U7110 ( .B1(n6071), .B2(UWORD_REG_9__SCAN_IN), .A(n6055), .ZN(n6056) );
  OAI21_X1 U7111 ( .B1(n6707), .B2(n6060), .A(n6056), .ZN(U2933) );
  AOI22_X1 U7112 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6072), .B1(
        UWORD_REG_11__SCAN_IN), .B2(n6071), .ZN(n6057) );
  NAND2_X1 U7113 ( .A1(n6061), .A2(DATAI_11_), .ZN(n6067) );
  NAND2_X1 U7114 ( .A1(n6057), .A2(n6067), .ZN(U2935) );
  NAND2_X1 U7115 ( .A1(n6061), .A2(DATAI_12_), .ZN(n6069) );
  INV_X1 U7116 ( .A(n6069), .ZN(n6058) );
  AOI21_X1 U7117 ( .B1(n6071), .B2(UWORD_REG_12__SCAN_IN), .A(n6058), .ZN(
        n6059) );
  OAI21_X1 U7118 ( .B1(n6780), .B2(n6060), .A(n6059), .ZN(U2936) );
  AOI22_X1 U7119 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6072), .B1(n6071), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7120 ( .A1(n6061), .A2(DATAI_13_), .ZN(n6073) );
  NAND2_X1 U7121 ( .A1(n6062), .A2(n6073), .ZN(U2937) );
  AOI22_X1 U7122 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6072), .B1(n6071), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7123 ( .A1(n6064), .A2(n6063), .ZN(U2947) );
  AOI22_X1 U7124 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6072), .B1(
        LWORD_REG_9__SCAN_IN), .B2(n6071), .ZN(n6066) );
  NAND2_X1 U7125 ( .A1(n6066), .A2(n6065), .ZN(U2948) );
  AOI22_X1 U7126 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6072), .B1(n6071), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7127 ( .A1(n6068), .A2(n6067), .ZN(U2950) );
  AOI22_X1 U7128 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6072), .B1(n6071), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7129 ( .A1(n6070), .A2(n6069), .ZN(U2951) );
  AOI22_X1 U7130 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6072), .B1(n6071), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7131 ( .A1(n6074), .A2(n6073), .ZN(U2952) );
  AOI22_X1 U7132 ( .A1(n6178), .A2(REIP_REG_7__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n6099), .ZN(n6081) );
  OAI21_X1 U7133 ( .B1(n6075), .B2(n6077), .A(n6076), .ZN(n6078) );
  INV_X1 U7134 ( .A(n6078), .ZN(n6138) );
  AOI22_X1 U7135 ( .A1(n6138), .A2(n3824), .B1(n6105), .B2(n6079), .ZN(n6080)
         );
  OAI211_X1 U7136 ( .C1(n6110), .C2(n6082), .A(n6081), .B(n6080), .ZN(U2979)
         );
  AOI22_X1 U7137 ( .A1(n6178), .A2(REIP_REG_5__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6099), .ZN(n6089) );
  OAI21_X1 U7138 ( .B1(n6083), .B2(n6085), .A(n6084), .ZN(n6086) );
  INV_X1 U7139 ( .A(n6086), .ZN(n6164) );
  AOI22_X1 U7140 ( .A1(n6164), .A2(n3824), .B1(n6105), .B2(n6087), .ZN(n6088)
         );
  OAI211_X1 U7141 ( .C1(n6110), .C2(n6090), .A(n6089), .B(n6088), .ZN(U2981)
         );
  AOI22_X1 U7142 ( .A1(n6178), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6099), .ZN(n6097) );
  OAI21_X1 U7143 ( .B1(n6091), .B2(n6093), .A(n6092), .ZN(n6094) );
  INV_X1 U7144 ( .A(n6094), .ZN(n6181) );
  AOI22_X1 U7145 ( .A1(n6181), .A2(n3824), .B1(n6105), .B2(n6095), .ZN(n6096)
         );
  OAI211_X1 U7146 ( .C1(n6110), .C2(n6098), .A(n6097), .B(n6096), .ZN(U2983)
         );
  AOI22_X1 U7147 ( .A1(n6178), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6099), .ZN(n6108) );
  INV_X1 U7148 ( .A(n6100), .ZN(n6106) );
  CLKBUF_X1 U7149 ( .A(n6101), .Z(n6102) );
  XNOR2_X1 U7150 ( .A(n6102), .B(n3422), .ZN(n6103) );
  XNOR2_X1 U7151 ( .A(n6104), .B(n6103), .ZN(n6191) );
  AOI22_X1 U7152 ( .A1(n6106), .A2(n6105), .B1(n6191), .B2(n3824), .ZN(n6107)
         );
  OAI211_X1 U7153 ( .C1(n6110), .C2(n6109), .A(n6108), .B(n6107), .ZN(U2984)
         );
  INV_X1 U7154 ( .A(n6111), .ZN(n6116) );
  OAI22_X1 U7155 ( .A1(n6195), .A2(n6112), .B1(n6610), .B2(n6193), .ZN(n6113)
         );
  AOI21_X1 U7156 ( .B1(n6114), .B2(n6190), .A(n6113), .ZN(n6115) );
  OAI221_X1 U7157 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6118), .C1(
        n6117), .C2(n6116), .A(n6115), .ZN(U3007) );
  AOI21_X1 U7158 ( .B1(n6180), .B2(n6120), .A(n6119), .ZN(n6124) );
  AOI22_X1 U7159 ( .A1(n6122), .A2(n6190), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6121), .ZN(n6123) );
  OAI211_X1 U7160 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6125), .A(n6124), 
        .B(n6123), .ZN(U3009) );
  INV_X1 U7161 ( .A(n6126), .ZN(n6127) );
  AOI21_X1 U7162 ( .B1(n6180), .B2(n6128), .A(n6127), .ZN(n6134) );
  INV_X1 U7163 ( .A(n6129), .ZN(n6132) );
  AOI21_X1 U7164 ( .B1(n6135), .B2(n6723), .A(n6130), .ZN(n6131) );
  AOI22_X1 U7165 ( .A1(n6132), .A2(n6190), .B1(n6137), .B2(n6131), .ZN(n6133)
         );
  OAI211_X1 U7166 ( .C1(n6141), .C2(n6135), .A(n6134), .B(n6133), .ZN(U3010)
         );
  AOI22_X1 U7167 ( .A1(n6180), .A2(n6136), .B1(n6178), .B2(REIP_REG_7__SCAN_IN), .ZN(n6140) );
  AOI22_X1 U7168 ( .A1(n6138), .A2(n6190), .B1(n6137), .B2(n6723), .ZN(n6139)
         );
  OAI211_X1 U7169 ( .C1(n6141), .C2(n6723), .A(n6140), .B(n6139), .ZN(U3011)
         );
  INV_X1 U7170 ( .A(n6142), .ZN(n6145) );
  INV_X1 U7171 ( .A(n6143), .ZN(n6144) );
  AOI21_X1 U7172 ( .B1(n6180), .B2(n6145), .A(n6144), .ZN(n6155) );
  INV_X1 U7173 ( .A(n6146), .ZN(n6147) );
  AOI22_X1 U7174 ( .A1(n6149), .A2(n6148), .B1(n6187), .B2(n6147), .ZN(n6200)
         );
  OAI21_X1 U7175 ( .B1(n6151), .B2(n6150), .A(n6200), .ZN(n6157) );
  INV_X1 U7176 ( .A(n6152), .ZN(n6153) );
  AOI22_X1 U7177 ( .A1(n6157), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n6153), 
        .B2(n6190), .ZN(n6154) );
  OAI211_X1 U7178 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6156), .A(n6155), 
        .B(n6154), .ZN(U3012) );
  OAI21_X1 U7179 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6158), .A(n6157), 
        .ZN(n6166) );
  OAI22_X1 U7180 ( .A1(n6195), .A2(n6159), .B1(n6602), .B2(n6193), .ZN(n6163)
         );
  NOR3_X1 U7181 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6161), .A3(n6160), 
        .ZN(n6162) );
  AOI211_X1 U7182 ( .C1(n6164), .C2(n6190), .A(n6163), .B(n6162), .ZN(n6165)
         );
  NAND2_X1 U7183 ( .A1(n6166), .A2(n6165), .ZN(U3013) );
  NOR2_X1 U7184 ( .A1(n6757), .A2(n6167), .ZN(n6176) );
  OAI211_X1 U7185 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6177), .B(n6189), .ZN(n6175) );
  INV_X1 U7186 ( .A(n6168), .ZN(n6169) );
  AOI21_X1 U7187 ( .B1(n6180), .B2(n6170), .A(n6169), .ZN(n6174) );
  OAI21_X1 U7188 ( .B1(n6187), .B2(n6189), .A(n6200), .ZN(n6182) );
  INV_X1 U7189 ( .A(n6171), .ZN(n6172) );
  AOI22_X1 U7190 ( .A1(n6182), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6190), 
        .B2(n6172), .ZN(n6173) );
  OAI211_X1 U7191 ( .C1(n6176), .C2(n6175), .A(n6174), .B(n6173), .ZN(U3014)
         );
  NAND2_X1 U7192 ( .A1(n6189), .A2(n6177), .ZN(n6185) );
  AOI22_X1 U7193 ( .A1(n6180), .A2(n6179), .B1(n6178), .B2(REIP_REG_3__SCAN_IN), .ZN(n6184) );
  AOI22_X1 U7194 ( .A1(n6182), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6190), 
        .B2(n6181), .ZN(n6183) );
  OAI211_X1 U7195 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6185), .A(n6184), 
        .B(n6183), .ZN(U3015) );
  NAND2_X1 U7196 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6186), .ZN(n6201)
         );
  AOI221_X1 U7197 ( .B1(n3422), .B2(n6189), .C1(n6188), .C2(n6189), .A(n6187), 
        .ZN(n6198) );
  AND2_X1 U7198 ( .A1(n6191), .A2(n6190), .ZN(n6197) );
  INV_X1 U7199 ( .A(n6192), .ZN(n6194) );
  OAI22_X1 U7200 ( .A1(n6195), .A2(n6194), .B1(n6598), .B2(n6193), .ZN(n6196)
         );
  NOR3_X1 U7201 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n6199) );
  OAI221_X1 U7202 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6201), .C1(n3422), .C2(n6200), .A(n6199), .ZN(U3016) );
  NOR2_X1 U7203 ( .A1(n6983), .A2(n6202), .ZN(U3019) );
  INV_X1 U7204 ( .A(n6203), .ZN(n6402) );
  AOI21_X1 U7205 ( .B1(n6204), .B2(n6402), .A(n6401), .ZN(n6205) );
  NOR2_X1 U7206 ( .A1(n6206), .A2(n6205), .ZN(n6213) );
  NOR2_X1 U7207 ( .A1(n6398), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6234)
         );
  AOI21_X1 U7208 ( .B1(n6207), .B2(n6528), .A(n6234), .ZN(n6212) );
  INV_X1 U7209 ( .A(n6212), .ZN(n6208) );
  OAI21_X1 U7210 ( .B1(n6213), .B2(n6208), .A(n6406), .ZN(n6209) );
  AOI21_X1 U7211 ( .B1(n6401), .B2(n6211), .A(n6209), .ZN(n6239) );
  INV_X1 U7212 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6922) );
  AOI22_X1 U7213 ( .A1(n6456), .A2(n6234), .B1(n6399), .B2(n6233), .ZN(n6215)
         );
  OR3_X1 U7214 ( .A1(n3934), .A2(n6210), .A3(n6396), .ZN(n6271) );
  INV_X1 U7215 ( .A(n6271), .ZN(n6236) );
  OAI22_X1 U7216 ( .A1(n6213), .A2(n6212), .B1(n6211), .B2(n6568), .ZN(n6235)
         );
  AOI22_X1 U7217 ( .A1(n6364), .A2(n6236), .B1(n6457), .B2(n6235), .ZN(n6214)
         );
  OAI211_X1 U7218 ( .C1(n6239), .C2(n6922), .A(n6215), .B(n6214), .ZN(U3044)
         );
  INV_X1 U7219 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U7220 ( .A1(n6464), .A2(n6234), .B1(n6367), .B2(n6233), .ZN(n6217)
         );
  AOI22_X1 U7221 ( .A1(n6414), .A2(n6236), .B1(n6465), .B2(n6235), .ZN(n6216)
         );
  OAI211_X1 U7222 ( .C1(n6239), .C2(n6218), .A(n6217), .B(n6216), .ZN(U3045)
         );
  INV_X1 U7223 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6221) );
  AOI22_X1 U7224 ( .A1(n6472), .A2(n6234), .B1(n6370), .B2(n6233), .ZN(n6220)
         );
  AOI22_X1 U7225 ( .A1(n6417), .A2(n6236), .B1(n6473), .B2(n6235), .ZN(n6219)
         );
  OAI211_X1 U7226 ( .C1(n6239), .C2(n6221), .A(n6220), .B(n6219), .ZN(U3046)
         );
  INV_X1 U7227 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6224) );
  AOI22_X1 U7228 ( .A1(n6480), .A2(n6234), .B1(n6420), .B2(n6233), .ZN(n6223)
         );
  AOI22_X1 U7229 ( .A1(n6373), .A2(n6236), .B1(n6481), .B2(n6235), .ZN(n6222)
         );
  OAI211_X1 U7230 ( .C1(n6239), .C2(n6224), .A(n6223), .B(n6222), .ZN(U3047)
         );
  INV_X1 U7231 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6227) );
  AOI22_X1 U7232 ( .A1(n6488), .A2(n6234), .B1(n6377), .B2(n6233), .ZN(n6226)
         );
  AOI22_X1 U7233 ( .A1(n6424), .A2(n6236), .B1(n6489), .B2(n6235), .ZN(n6225)
         );
  OAI211_X1 U7234 ( .C1(n6239), .C2(n6227), .A(n6226), .B(n6225), .ZN(U3048)
         );
  INV_X1 U7235 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6230) );
  AOI22_X1 U7236 ( .A1(n6496), .A2(n6234), .B1(n6380), .B2(n6233), .ZN(n6229)
         );
  AOI22_X1 U7237 ( .A1(n6427), .A2(n6236), .B1(n6497), .B2(n6235), .ZN(n6228)
         );
  OAI211_X1 U7238 ( .C1(n6239), .C2(n6230), .A(n6229), .B(n6228), .ZN(U3049)
         );
  INV_X1 U7239 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U7240 ( .A1(n6504), .A2(n6234), .B1(n6383), .B2(n6233), .ZN(n6232)
         );
  AOI22_X1 U7241 ( .A1(n6430), .A2(n6236), .B1(n6505), .B2(n6235), .ZN(n6231)
         );
  OAI211_X1 U7242 ( .C1(n6239), .C2(n6807), .A(n6232), .B(n6231), .ZN(U3050)
         );
  INV_X1 U7243 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6811) );
  AOI22_X1 U7244 ( .A1(n6513), .A2(n6234), .B1(n6388), .B2(n6233), .ZN(n6238)
         );
  AOI22_X1 U7245 ( .A1(n6433), .A2(n6236), .B1(n6515), .B2(n6235), .ZN(n6237)
         );
  OAI211_X1 U7246 ( .C1(n6239), .C2(n6811), .A(n6238), .B(n6237), .ZN(U3051)
         );
  INV_X1 U7247 ( .A(n6240), .ZN(n6241) );
  OAI22_X1 U7248 ( .A1(n6242), .A2(n6454), .B1(n6453), .B2(n6241), .ZN(n6266)
         );
  NOR2_X1 U7249 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6243), .ZN(n6265)
         );
  AOI22_X1 U7250 ( .A1(n6457), .A2(n6266), .B1(n6456), .B2(n6265), .ZN(n6252)
         );
  INV_X1 U7251 ( .A(n6265), .ZN(n6245) );
  AOI211_X1 U7252 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6245), .A(n6442), .B(
        n6244), .ZN(n6250) );
  OAI211_X1 U7253 ( .C1(n6248), .C2(n6271), .A(n6247), .B(n6246), .ZN(n6249)
         );
  NAND2_X1 U7254 ( .A1(n6250), .A2(n6249), .ZN(n6268) );
  AOI22_X1 U7255 ( .A1(n6268), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6364), 
        .B2(n6267), .ZN(n6251) );
  OAI211_X1 U7256 ( .C1(n6458), .C2(n6271), .A(n6252), .B(n6251), .ZN(U3052)
         );
  AOI22_X1 U7257 ( .A1(n6465), .A2(n6266), .B1(n6464), .B2(n6265), .ZN(n6254)
         );
  AOI22_X1 U7258 ( .A1(n6268), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6414), 
        .B2(n6267), .ZN(n6253) );
  OAI211_X1 U7259 ( .C1(n6466), .C2(n6271), .A(n6254), .B(n6253), .ZN(U3053)
         );
  AOI22_X1 U7260 ( .A1(n6473), .A2(n6266), .B1(n6472), .B2(n6265), .ZN(n6256)
         );
  AOI22_X1 U7261 ( .A1(n6268), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6417), 
        .B2(n6267), .ZN(n6255) );
  OAI211_X1 U7262 ( .C1(n6479), .C2(n6271), .A(n6256), .B(n6255), .ZN(U3054)
         );
  AOI22_X1 U7263 ( .A1(n6481), .A2(n6266), .B1(n6480), .B2(n6265), .ZN(n6258)
         );
  AOI22_X1 U7264 ( .A1(n6268), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6373), 
        .B2(n6267), .ZN(n6257) );
  OAI211_X1 U7265 ( .C1(n6487), .C2(n6271), .A(n6258), .B(n6257), .ZN(U3055)
         );
  AOI22_X1 U7266 ( .A1(n6489), .A2(n6266), .B1(n6488), .B2(n6265), .ZN(n6260)
         );
  AOI22_X1 U7267 ( .A1(n6268), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6424), 
        .B2(n6267), .ZN(n6259) );
  OAI211_X1 U7268 ( .C1(n6495), .C2(n6271), .A(n6260), .B(n6259), .ZN(U3056)
         );
  AOI22_X1 U7269 ( .A1(n6497), .A2(n6266), .B1(n6496), .B2(n6265), .ZN(n6262)
         );
  AOI22_X1 U7270 ( .A1(n6268), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6427), 
        .B2(n6267), .ZN(n6261) );
  OAI211_X1 U7271 ( .C1(n6503), .C2(n6271), .A(n6262), .B(n6261), .ZN(U3057)
         );
  AOI22_X1 U7272 ( .A1(n6505), .A2(n6266), .B1(n6504), .B2(n6265), .ZN(n6264)
         );
  AOI22_X1 U7273 ( .A1(n6268), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6430), 
        .B2(n6267), .ZN(n6263) );
  OAI211_X1 U7274 ( .C1(n6511), .C2(n6271), .A(n6264), .B(n6263), .ZN(U3058)
         );
  AOI22_X1 U7275 ( .A1(n6515), .A2(n6266), .B1(n6513), .B2(n6265), .ZN(n6270)
         );
  AOI22_X1 U7276 ( .A1(n6268), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6433), 
        .B2(n6267), .ZN(n6269) );
  OAI211_X1 U7277 ( .C1(n6524), .C2(n6271), .A(n6270), .B(n6269), .ZN(U3059)
         );
  AOI22_X1 U7278 ( .A1(n6457), .A2(n6273), .B1(n6456), .B2(n6272), .ZN(n6279)
         );
  INV_X1 U7279 ( .A(n6274), .ZN(n6277) );
  INV_X1 U7280 ( .A(n6275), .ZN(n6276) );
  AOI22_X1 U7281 ( .A1(n6277), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6399), 
        .B2(n6276), .ZN(n6278) );
  OAI211_X1 U7282 ( .C1(n6460), .C2(n6280), .A(n6279), .B(n6278), .ZN(U3068)
         );
  AND2_X1 U7283 ( .A1(n6281), .A2(n6324), .ZN(n6286) );
  INV_X1 U7284 ( .A(n6282), .ZN(n6312) );
  AOI21_X1 U7285 ( .B1(n6283), .B2(n6528), .A(n6312), .ZN(n6285) );
  INV_X1 U7286 ( .A(n6285), .ZN(n6284) );
  AOI22_X1 U7287 ( .A1(n6286), .A2(n6284), .B1(n6288), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n6318) );
  AOI22_X1 U7288 ( .A1(n6456), .A2(n6312), .B1(n6399), .B2(n6313), .ZN(n6291)
         );
  NAND2_X1 U7289 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  OAI211_X1 U7290 ( .C1(n6288), .C2(n6447), .A(n6406), .B(n6287), .ZN(n6314)
         );
  AOI22_X1 U7291 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6314), .B1(n6364), 
        .B2(n6311), .ZN(n6290) );
  OAI211_X1 U7292 ( .C1(n6318), .C2(n6292), .A(n6291), .B(n6290), .ZN(U3076)
         );
  AOI22_X1 U7293 ( .A1(n6464), .A2(n6312), .B1(n6414), .B2(n6311), .ZN(n6294)
         );
  AOI22_X1 U7294 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6314), .B1(n6367), 
        .B2(n6313), .ZN(n6293) );
  OAI211_X1 U7295 ( .C1(n6318), .C2(n6295), .A(n6294), .B(n6293), .ZN(U3077)
         );
  AOI22_X1 U7296 ( .A1(n6472), .A2(n6312), .B1(n6417), .B2(n6311), .ZN(n6297)
         );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6314), .B1(n6370), 
        .B2(n6313), .ZN(n6296) );
  OAI211_X1 U7298 ( .C1(n6318), .C2(n6298), .A(n6297), .B(n6296), .ZN(U3078)
         );
  AOI22_X1 U7299 ( .A1(n6480), .A2(n6312), .B1(n6420), .B2(n6313), .ZN(n6300)
         );
  AOI22_X1 U7300 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6314), .B1(n6373), 
        .B2(n6311), .ZN(n6299) );
  OAI211_X1 U7301 ( .C1(n6318), .C2(n6301), .A(n6300), .B(n6299), .ZN(U3079)
         );
  AOI22_X1 U7302 ( .A1(n6488), .A2(n6312), .B1(n6377), .B2(n6313), .ZN(n6303)
         );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6314), .B1(n6424), 
        .B2(n6311), .ZN(n6302) );
  OAI211_X1 U7304 ( .C1(n6318), .C2(n6304), .A(n6303), .B(n6302), .ZN(U3080)
         );
  AOI22_X1 U7305 ( .A1(n6496), .A2(n6312), .B1(n6380), .B2(n6313), .ZN(n6306)
         );
  AOI22_X1 U7306 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6314), .B1(n6427), 
        .B2(n6311), .ZN(n6305) );
  OAI211_X1 U7307 ( .C1(n6318), .C2(n6307), .A(n6306), .B(n6305), .ZN(U3081)
         );
  AOI22_X1 U7308 ( .A1(n6504), .A2(n6312), .B1(n6430), .B2(n6311), .ZN(n6309)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6314), .B1(n6383), 
        .B2(n6313), .ZN(n6308) );
  OAI211_X1 U7310 ( .C1(n6318), .C2(n6310), .A(n6309), .B(n6308), .ZN(U3082)
         );
  AOI22_X1 U7311 ( .A1(n6513), .A2(n6312), .B1(n6433), .B2(n6311), .ZN(n6316)
         );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6314), .B1(n6388), 
        .B2(n6313), .ZN(n6315) );
  OAI211_X1 U7313 ( .C1(n6318), .C2(n6317), .A(n6316), .B(n6315), .ZN(U3083)
         );
  INV_X1 U7314 ( .A(n6319), .ZN(n6455) );
  NAND2_X1 U7315 ( .A1(n6321), .A2(n6320), .ZN(n6452) );
  OAI22_X1 U7316 ( .A1(n6455), .A2(n6357), .B1(n6322), .B2(n6452), .ZN(n6348)
         );
  NAND3_X1 U7317 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6539), .A3(n6534), .ZN(n6361) );
  NOR2_X1 U7318 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6361), .ZN(n6347)
         );
  AOI22_X1 U7319 ( .A1(n6457), .A2(n6348), .B1(n6456), .B2(n6347), .ZN(n6334)
         );
  AOI21_X1 U7320 ( .B1(n6332), .B2(n6352), .A(n6353), .ZN(n6331) );
  OAI21_X1 U7321 ( .B1(n6325), .B2(n6357), .A(n6324), .ZN(n6330) );
  AOI21_X1 U7322 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6452), .A(n6326), .ZN(
        n6445) );
  INV_X1 U7323 ( .A(n6347), .ZN(n6328) );
  AOI21_X1 U7324 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6328), .A(n6327), .ZN(
        n6329) );
  OAI211_X1 U7325 ( .C1(n6331), .C2(n6330), .A(n6445), .B(n6329), .ZN(n6349)
         );
  AOI22_X1 U7326 ( .A1(n6349), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6364), 
        .B2(n6389), .ZN(n6333) );
  OAI211_X1 U7327 ( .C1(n6458), .C2(n6352), .A(n6334), .B(n6333), .ZN(U3084)
         );
  AOI22_X1 U7328 ( .A1(n6465), .A2(n6348), .B1(n6464), .B2(n6347), .ZN(n6336)
         );
  AOI22_X1 U7329 ( .A1(n6349), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6414), 
        .B2(n6389), .ZN(n6335) );
  OAI211_X1 U7330 ( .C1(n6466), .C2(n6352), .A(n6336), .B(n6335), .ZN(U3085)
         );
  AOI22_X1 U7331 ( .A1(n6473), .A2(n6348), .B1(n6472), .B2(n6347), .ZN(n6338)
         );
  AOI22_X1 U7332 ( .A1(n6349), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6417), 
        .B2(n6389), .ZN(n6337) );
  OAI211_X1 U7333 ( .C1(n6479), .C2(n6352), .A(n6338), .B(n6337), .ZN(U3086)
         );
  AOI22_X1 U7334 ( .A1(n6481), .A2(n6348), .B1(n6480), .B2(n6347), .ZN(n6340)
         );
  AOI22_X1 U7335 ( .A1(n6349), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6373), 
        .B2(n6389), .ZN(n6339) );
  OAI211_X1 U7336 ( .C1(n6487), .C2(n6352), .A(n6340), .B(n6339), .ZN(U3087)
         );
  AOI22_X1 U7337 ( .A1(n6489), .A2(n6348), .B1(n6488), .B2(n6347), .ZN(n6342)
         );
  AOI22_X1 U7338 ( .A1(n6349), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6424), 
        .B2(n6389), .ZN(n6341) );
  OAI211_X1 U7339 ( .C1(n6495), .C2(n6352), .A(n6342), .B(n6341), .ZN(U3088)
         );
  AOI22_X1 U7340 ( .A1(n6497), .A2(n6348), .B1(n6496), .B2(n6347), .ZN(n6344)
         );
  AOI22_X1 U7341 ( .A1(n6349), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6427), 
        .B2(n6389), .ZN(n6343) );
  OAI211_X1 U7342 ( .C1(n6503), .C2(n6352), .A(n6344), .B(n6343), .ZN(U3089)
         );
  AOI22_X1 U7343 ( .A1(n6505), .A2(n6348), .B1(n6504), .B2(n6347), .ZN(n6346)
         );
  AOI22_X1 U7344 ( .A1(n6349), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6430), 
        .B2(n6389), .ZN(n6345) );
  OAI211_X1 U7345 ( .C1(n6511), .C2(n6352), .A(n6346), .B(n6345), .ZN(U3090)
         );
  AOI22_X1 U7346 ( .A1(n6515), .A2(n6348), .B1(n6513), .B2(n6347), .ZN(n6351)
         );
  AOI22_X1 U7347 ( .A1(n6349), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6433), 
        .B2(n6389), .ZN(n6350) );
  OAI211_X1 U7348 ( .C1(n6524), .C2(n6352), .A(n6351), .B(n6350), .ZN(U3091)
         );
  OAI21_X1 U7349 ( .B1(n6354), .B2(n6353), .A(n6447), .ZN(n6363) );
  NOR2_X1 U7350 ( .A1(n6355), .A2(n6361), .ZN(n6387) );
  INV_X1 U7351 ( .A(n6387), .ZN(n6356) );
  OAI21_X1 U7352 ( .B1(n6358), .B2(n6357), .A(n6356), .ZN(n6360) );
  OAI21_X1 U7353 ( .B1(n6363), .B2(n6360), .A(n6406), .ZN(n6359) );
  AOI21_X1 U7354 ( .B1(n6401), .B2(n6361), .A(n6359), .ZN(n6395) );
  INV_X1 U7355 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7356 ( .A1(n6389), .A2(n6399), .B1(n6456), .B2(n6387), .ZN(n6366)
         );
  INV_X1 U7357 ( .A(n6360), .ZN(n6362) );
  OAI22_X1 U7358 ( .A1(n6363), .A2(n6362), .B1(n6361), .B2(n6568), .ZN(n6391)
         );
  AOI22_X1 U7359 ( .A1(n6391), .A2(n6457), .B1(n6390), .B2(n6364), .ZN(n6365)
         );
  OAI211_X1 U7360 ( .C1(n6395), .C2(n6904), .A(n6366), .B(n6365), .ZN(U3092)
         );
  INV_X1 U7361 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6977) );
  AOI22_X1 U7362 ( .A1(n6389), .A2(n6367), .B1(n6464), .B2(n6387), .ZN(n6369)
         );
  AOI22_X1 U7363 ( .A1(n6391), .A2(n6465), .B1(n6390), .B2(n6414), .ZN(n6368)
         );
  OAI211_X1 U7364 ( .C1(n6395), .C2(n6977), .A(n6369), .B(n6368), .ZN(U3093)
         );
  INV_X1 U7365 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7366 ( .A1(n6390), .A2(n6417), .B1(n6472), .B2(n6387), .ZN(n6372)
         );
  AOI22_X1 U7367 ( .A1(n6391), .A2(n6473), .B1(n6370), .B2(n6389), .ZN(n6371)
         );
  OAI211_X1 U7368 ( .C1(n6395), .C2(n6772), .A(n6372), .B(n6371), .ZN(U3094)
         );
  INV_X1 U7369 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6376) );
  AOI22_X1 U7370 ( .A1(n6390), .A2(n6373), .B1(n6480), .B2(n6387), .ZN(n6375)
         );
  AOI22_X1 U7371 ( .A1(n6391), .A2(n6481), .B1(n6420), .B2(n6389), .ZN(n6374)
         );
  OAI211_X1 U7372 ( .C1(n6395), .C2(n6376), .A(n6375), .B(n6374), .ZN(U3095)
         );
  INV_X1 U7373 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7374 ( .A1(n6390), .A2(n6424), .B1(n6488), .B2(n6387), .ZN(n6379)
         );
  AOI22_X1 U7375 ( .A1(n6391), .A2(n6489), .B1(n6377), .B2(n6389), .ZN(n6378)
         );
  OAI211_X1 U7376 ( .C1(n6395), .C2(n6732), .A(n6379), .B(n6378), .ZN(U3096)
         );
  INV_X1 U7377 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U7378 ( .A1(n6390), .A2(n6427), .B1(n6496), .B2(n6387), .ZN(n6382)
         );
  AOI22_X1 U7379 ( .A1(n6391), .A2(n6497), .B1(n6380), .B2(n6389), .ZN(n6381)
         );
  OAI211_X1 U7380 ( .C1(n6395), .C2(n6954), .A(n6382), .B(n6381), .ZN(U3097)
         );
  INV_X1 U7381 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U7382 ( .A1(n6390), .A2(n6430), .B1(n6504), .B2(n6387), .ZN(n6385)
         );
  AOI22_X1 U7383 ( .A1(n6391), .A2(n6505), .B1(n6383), .B2(n6389), .ZN(n6384)
         );
  OAI211_X1 U7384 ( .C1(n6395), .C2(n6386), .A(n6385), .B(n6384), .ZN(U3098)
         );
  INV_X1 U7385 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6394) );
  AOI22_X1 U7386 ( .A1(n6389), .A2(n6388), .B1(n6513), .B2(n6387), .ZN(n6393)
         );
  AOI22_X1 U7387 ( .A1(n6391), .A2(n6515), .B1(n6390), .B2(n6433), .ZN(n6392)
         );
  OAI211_X1 U7388 ( .C1(n6395), .C2(n6394), .A(n6393), .B(n6392), .ZN(U3099)
         );
  NOR2_X1 U7389 ( .A1(n6398), .A2(n6397), .ZN(n6435) );
  INV_X1 U7390 ( .A(n6440), .ZN(n6421) );
  AOI22_X1 U7391 ( .A1(n6456), .A2(n6435), .B1(n6421), .B2(n6399), .ZN(n6413)
         );
  INV_X1 U7392 ( .A(n6409), .ZN(n6407) );
  INV_X1 U7393 ( .A(n6400), .ZN(n6403) );
  AOI21_X1 U7394 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6408) );
  AOI21_X1 U7395 ( .B1(n6404), .B2(n6528), .A(n6435), .ZN(n6410) );
  NAND2_X1 U7396 ( .A1(n6408), .A2(n6410), .ZN(n6405) );
  OAI211_X1 U7397 ( .C1(n6447), .C2(n6407), .A(n6406), .B(n6405), .ZN(n6437)
         );
  INV_X1 U7398 ( .A(n6408), .ZN(n6411) );
  OAI22_X1 U7399 ( .A1(n6411), .A2(n6410), .B1(n6409), .B2(n6568), .ZN(n6436)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6437), .B1(n6457), 
        .B2(n6436), .ZN(n6412) );
  OAI211_X1 U7401 ( .C1(n6460), .C2(n6523), .A(n6413), .B(n6412), .ZN(U3108)
         );
  INV_X1 U7402 ( .A(n6523), .ZN(n6434) );
  AOI22_X1 U7403 ( .A1(n6464), .A2(n6435), .B1(n6434), .B2(n6414), .ZN(n6416)
         );
  AOI22_X1 U7404 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6437), .B1(n6465), 
        .B2(n6436), .ZN(n6415) );
  OAI211_X1 U7405 ( .C1(n6466), .C2(n6440), .A(n6416), .B(n6415), .ZN(U3109)
         );
  AOI22_X1 U7406 ( .A1(n6472), .A2(n6435), .B1(n6434), .B2(n6417), .ZN(n6419)
         );
  AOI22_X1 U7407 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6437), .B1(n6473), 
        .B2(n6436), .ZN(n6418) );
  OAI211_X1 U7408 ( .C1(n6479), .C2(n6440), .A(n6419), .B(n6418), .ZN(U3110)
         );
  AOI22_X1 U7409 ( .A1(n6480), .A2(n6435), .B1(n6421), .B2(n6420), .ZN(n6423)
         );
  AOI22_X1 U7410 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6437), .B1(n6481), 
        .B2(n6436), .ZN(n6422) );
  OAI211_X1 U7411 ( .C1(n6482), .C2(n6523), .A(n6423), .B(n6422), .ZN(U3111)
         );
  AOI22_X1 U7412 ( .A1(n6488), .A2(n6435), .B1(n6434), .B2(n6424), .ZN(n6426)
         );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6437), .B1(n6489), 
        .B2(n6436), .ZN(n6425) );
  OAI211_X1 U7414 ( .C1(n6495), .C2(n6440), .A(n6426), .B(n6425), .ZN(U3112)
         );
  AOI22_X1 U7415 ( .A1(n6496), .A2(n6435), .B1(n6434), .B2(n6427), .ZN(n6429)
         );
  AOI22_X1 U7416 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6437), .B1(n6497), 
        .B2(n6436), .ZN(n6428) );
  OAI211_X1 U7417 ( .C1(n6503), .C2(n6440), .A(n6429), .B(n6428), .ZN(U3113)
         );
  AOI22_X1 U7418 ( .A1(n6504), .A2(n6435), .B1(n6434), .B2(n6430), .ZN(n6432)
         );
  AOI22_X1 U7419 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6437), .B1(n6505), 
        .B2(n6436), .ZN(n6431) );
  OAI211_X1 U7420 ( .C1(n6511), .C2(n6440), .A(n6432), .B(n6431), .ZN(U3114)
         );
  AOI22_X1 U7421 ( .A1(n6513), .A2(n6435), .B1(n6434), .B2(n6433), .ZN(n6439)
         );
  AOI22_X1 U7422 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6437), .B1(n6515), 
        .B2(n6436), .ZN(n6438) );
  OAI211_X1 U7423 ( .C1(n6524), .C2(n6440), .A(n6439), .B(n6438), .ZN(U3115)
         );
  NOR2_X1 U7424 ( .A1(n6441), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6512)
         );
  INV_X1 U7425 ( .A(n6512), .ZN(n6443) );
  AOI21_X1 U7426 ( .B1(n6443), .B2(STATE2_REG_3__SCAN_IN), .A(n6442), .ZN(
        n6444) );
  AND2_X1 U7427 ( .A1(n6445), .A2(n6444), .ZN(n6451) );
  NAND2_X1 U7428 ( .A1(n6516), .A2(n6523), .ZN(n6446) );
  NAND2_X1 U7429 ( .A1(n6446), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6448) );
  OAI211_X1 U7430 ( .C1(n6449), .C2(n6454), .A(n6448), .B(n6447), .ZN(n6450)
         );
  INV_X1 U7431 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6940) );
  OAI22_X1 U7432 ( .A1(n6455), .A2(n6454), .B1(n6453), .B2(n6452), .ZN(n6514)
         );
  AOI22_X1 U7433 ( .A1(n6457), .A2(n6514), .B1(n6456), .B2(n6512), .ZN(n6463)
         );
  OR2_X1 U7434 ( .A1(n6523), .A2(n6458), .ZN(n6459) );
  OAI21_X1 U7435 ( .B1(n6516), .B2(n6460), .A(n6459), .ZN(n6461) );
  INV_X1 U7436 ( .A(n6461), .ZN(n6462) );
  OAI211_X1 U7437 ( .C1(n6519), .C2(n6940), .A(n6463), .B(n6462), .ZN(U3116)
         );
  INV_X1 U7438 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7439 ( .A1(n6465), .A2(n6514), .B1(n6464), .B2(n6512), .ZN(n6471)
         );
  OR2_X1 U7440 ( .A1(n6523), .A2(n6466), .ZN(n6467) );
  OAI21_X1 U7441 ( .B1(n6516), .B2(n6468), .A(n6467), .ZN(n6469) );
  INV_X1 U7442 ( .A(n6469), .ZN(n6470) );
  OAI211_X1 U7443 ( .C1(n6519), .C2(n6960), .A(n6471), .B(n6470), .ZN(U3117)
         );
  AOI22_X1 U7444 ( .A1(n6473), .A2(n6514), .B1(n6472), .B2(n6512), .ZN(n6478)
         );
  INV_X1 U7445 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6475) );
  OAI22_X1 U7446 ( .A1(n6519), .A2(n6475), .B1(n6474), .B2(n6516), .ZN(n6476)
         );
  INV_X1 U7447 ( .A(n6476), .ZN(n6477) );
  OAI211_X1 U7448 ( .C1(n6479), .C2(n6523), .A(n6478), .B(n6477), .ZN(U3118)
         );
  AOI22_X1 U7449 ( .A1(n6481), .A2(n6514), .B1(n6480), .B2(n6512), .ZN(n6486)
         );
  INV_X1 U7450 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6483) );
  OAI22_X1 U7451 ( .A1(n6519), .A2(n6483), .B1(n6482), .B2(n6516), .ZN(n6484)
         );
  INV_X1 U7452 ( .A(n6484), .ZN(n6485) );
  OAI211_X1 U7453 ( .C1(n6487), .C2(n6523), .A(n6486), .B(n6485), .ZN(U3119)
         );
  AOI22_X1 U7454 ( .A1(n6489), .A2(n6514), .B1(n6488), .B2(n6512), .ZN(n6494)
         );
  INV_X1 U7455 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6491) );
  OAI22_X1 U7456 ( .A1(n6519), .A2(n6491), .B1(n6490), .B2(n6516), .ZN(n6492)
         );
  INV_X1 U7457 ( .A(n6492), .ZN(n6493) );
  OAI211_X1 U7458 ( .C1(n6495), .C2(n6523), .A(n6494), .B(n6493), .ZN(U3120)
         );
  AOI22_X1 U7459 ( .A1(n6497), .A2(n6514), .B1(n6496), .B2(n6512), .ZN(n6502)
         );
  INV_X1 U7460 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6499) );
  OAI22_X1 U7461 ( .A1(n6519), .A2(n6499), .B1(n6498), .B2(n6516), .ZN(n6500)
         );
  INV_X1 U7462 ( .A(n6500), .ZN(n6501) );
  OAI211_X1 U7463 ( .C1(n6503), .C2(n6523), .A(n6502), .B(n6501), .ZN(U3121)
         );
  AOI22_X1 U7464 ( .A1(n6505), .A2(n6514), .B1(n6504), .B2(n6512), .ZN(n6510)
         );
  INV_X1 U7465 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6507) );
  OAI22_X1 U7466 ( .A1(n6519), .A2(n6507), .B1(n6506), .B2(n6516), .ZN(n6508)
         );
  INV_X1 U7467 ( .A(n6508), .ZN(n6509) );
  OAI211_X1 U7468 ( .C1(n6511), .C2(n6523), .A(n6510), .B(n6509), .ZN(U3122)
         );
  AOI22_X1 U7469 ( .A1(n6515), .A2(n6514), .B1(n6513), .B2(n6512), .ZN(n6522)
         );
  INV_X1 U7470 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6518) );
  OAI22_X1 U7471 ( .A1(n6519), .A2(n6518), .B1(n6517), .B2(n6516), .ZN(n6520)
         );
  INV_X1 U7472 ( .A(n6520), .ZN(n6521) );
  OAI211_X1 U7473 ( .C1(n6524), .C2(n6523), .A(n6522), .B(n6521), .ZN(U3123)
         );
  NOR2_X1 U7474 ( .A1(n6525), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6526)
         );
  AOI21_X1 U7475 ( .B1(n6528), .B2(n6527), .A(n6526), .ZN(n6657) );
  NAND2_X1 U7476 ( .A1(n6529), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6662) );
  AND2_X1 U7477 ( .A1(n6662), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6530)
         );
  NAND2_X1 U7478 ( .A1(n6657), .A2(n6530), .ZN(n6533) );
  INV_X1 U7479 ( .A(n6533), .ZN(n6536) );
  OAI211_X1 U7480 ( .C1(n6534), .C2(n6533), .A(n6532), .B(n6531), .ZN(n6535)
         );
  OAI21_X1 U7481 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6536), .A(n6535), 
        .ZN(n6537) );
  AOI222_X1 U7482 ( .A1(n6539), .A2(n6538), .B1(n6539), .B2(n6537), .C1(n6538), 
        .C2(n6537), .ZN(n6542) );
  INV_X1 U7483 ( .A(n6540), .ZN(n6541) );
  AOI222_X1 U7484 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6542), .B1(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6541), .C1(n6542), .C2(n6541), 
        .ZN(n6550) );
  OAI21_X1 U7485 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6543), 
        .ZN(n6544) );
  NAND4_X1 U7486 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(n6548)
         );
  AOI211_X1 U7487 ( .C1(n6550), .C2(n6983), .A(n6549), .B(n6548), .ZN(n6551)
         );
  INV_X1 U7488 ( .A(n6551), .ZN(n6563) );
  NOR2_X1 U7489 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6892), .ZN(n6576) );
  NOR3_X1 U7490 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6568), .A3(n6892), .ZN(
        n6552) );
  OAI22_X1 U7491 ( .A1(n6555), .A2(n6554), .B1(n6553), .B2(n6552), .ZN(n6556)
         );
  AOI221_X1 U7492 ( .B1(n6972), .B2(n6557), .C1(n6563), .C2(n6557), .A(n6556), 
        .ZN(n6651) );
  NOR2_X1 U7493 ( .A1(n6576), .A2(n6651), .ZN(n6560) );
  OAI21_X1 U7494 ( .B1(n6572), .B2(n6558), .A(n6972), .ZN(n6559) );
  OAI22_X1 U7495 ( .A1(n6972), .A2(n6560), .B1(n6651), .B2(n6559), .ZN(n6561)
         );
  AOI211_X1 U7496 ( .C1(n6566), .C2(n6563), .A(n6562), .B(n6561), .ZN(n6564)
         );
  OAI21_X1 U7497 ( .B1(n6972), .B2(n6565), .A(n6564), .ZN(U3148) );
  AOI21_X1 U7498 ( .B1(n6567), .B2(n6892), .A(n6566), .ZN(n6571) );
  NAND2_X1 U7499 ( .A1(n6972), .A2(n6568), .ZN(n6573) );
  OAI211_X1 U7500 ( .C1(n6651), .C2(n6576), .A(STATE2_REG_1__SCAN_IN), .B(
        n6573), .ZN(n6569) );
  OAI211_X1 U7501 ( .C1(n6651), .C2(n6571), .A(n6570), .B(n6569), .ZN(U3149)
         );
  NAND3_X1 U7502 ( .A1(n6573), .A2(n6572), .A3(n6652), .ZN(n6575) );
  OAI21_X1 U7503 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(U3150) );
  INV_X1 U7504 ( .A(n6650), .ZN(n6577) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6577), .ZN(U3151) );
  AND2_X1 U7506 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6577), .ZN(U3152) );
  AND2_X1 U7507 ( .A1(n6577), .A2(DATAWIDTH_REG_29__SCAN_IN), .ZN(U3153) );
  AND2_X1 U7508 ( .A1(n6577), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6577), .ZN(U3155) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6577), .ZN(U3156) );
  AND2_X1 U7511 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6577), .ZN(U3157) );
  AND2_X1 U7512 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6577), .ZN(U3158) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6577), .ZN(U3159) );
  AND2_X1 U7514 ( .A1(n6577), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U7515 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6577), .ZN(U3161) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6577), .ZN(U3162) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6577), .ZN(U3163) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6577), .ZN(U3164) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6577), .ZN(U3165) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6577), .ZN(U3166) );
  AND2_X1 U7521 ( .A1(n6577), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6577), .ZN(U3168) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6577), .ZN(U3169) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6577), .ZN(U3170) );
  AND2_X1 U7525 ( .A1(n6577), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6577), .ZN(U3172) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6577), .ZN(U3173) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6577), .ZN(U3174) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6577), .ZN(U3175) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6577), .ZN(U3176) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6577), .ZN(U3177) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6577), .ZN(U3178) );
  AND2_X1 U7533 ( .A1(n6577), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6577), .ZN(U3180) );
  AOI22_X1 U7535 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6593) );
  AND2_X1 U7536 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6581) );
  INV_X1 U7537 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6579) );
  INV_X1 U7538 ( .A(NA_N), .ZN(n6586) );
  AOI221_X1 U7539 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6586), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6590) );
  AOI221_X1 U7540 ( .B1(n6581), .B2(n6684), .C1(n6579), .C2(n6674), .A(n6590), 
        .ZN(n6578) );
  OAI21_X1 U7541 ( .B1(n6585), .B2(n6593), .A(n6578), .ZN(U3181) );
  NOR2_X1 U7542 ( .A1(n6588), .A2(n6579), .ZN(n6587) );
  NAND2_X1 U7543 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6580) );
  OAI21_X1 U7544 ( .B1(n6587), .B2(n6581), .A(n6580), .ZN(n6582) );
  OAI211_X1 U7545 ( .C1(n6584), .C2(n6892), .A(n6583), .B(n6582), .ZN(U3182)
         );
  AOI21_X1 U7546 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6592) );
  AOI221_X1 U7547 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6892), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6589) );
  AOI221_X1 U7548 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6589), .C2(HOLD), .A(n6588), .ZN(n6591) );
  OAI22_X1 U7549 ( .A1(n6593), .A2(n6592), .B1(n6591), .B2(n6590), .ZN(U3183)
         );
  INV_X1 U7550 ( .A(n6638), .ZN(n6643) );
  NAND2_X1 U7551 ( .A1(n6595), .A2(n6594), .ZN(n6640) );
  INV_X1 U7552 ( .A(n6640), .ZN(n6641) );
  AOI22_X1 U7553 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6674), .ZN(n6596) );
  OAI21_X1 U7554 ( .B1(n6664), .B2(n6643), .A(n6596), .ZN(U3184) );
  AOI22_X1 U7555 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6674), .ZN(n6597) );
  OAI21_X1 U7556 ( .B1(n6598), .B2(n6643), .A(n6597), .ZN(U3185) );
  INV_X1 U7557 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U7558 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6674), .ZN(n6599) );
  OAI21_X1 U7559 ( .B1(n6810), .B2(n6643), .A(n6599), .ZN(U3186) );
  AOI22_X1 U7560 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6674), .ZN(n6600) );
  OAI21_X1 U7561 ( .B1(n6704), .B2(n6643), .A(n6600), .ZN(U3187) );
  AOI22_X1 U7562 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6674), .ZN(n6601) );
  OAI21_X1 U7563 ( .B1(n6602), .B2(n6643), .A(n6601), .ZN(U3188) );
  AOI22_X1 U7564 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6674), .ZN(n6603) );
  OAI21_X1 U7565 ( .B1(n6604), .B2(n6643), .A(n6603), .ZN(U3189) );
  AOI22_X1 U7566 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6674), .ZN(n6605) );
  OAI21_X1 U7567 ( .B1(n6606), .B2(n6643), .A(n6605), .ZN(U3190) );
  AOI22_X1 U7568 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6674), .ZN(n6607) );
  OAI21_X1 U7569 ( .B1(n5057), .B2(n6640), .A(n6607), .ZN(U3191) );
  AOI22_X1 U7570 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6674), .ZN(n6608) );
  OAI21_X1 U7571 ( .B1(n5057), .B2(n6643), .A(n6608), .ZN(U3192) );
  AOI22_X1 U7572 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6674), .ZN(n6609) );
  OAI21_X1 U7573 ( .B1(n6610), .B2(n6640), .A(n6609), .ZN(U3193) );
  AOI222_X1 U7574 ( .A1(n6641), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6674), .C1(REIP_REG_11__SCAN_IN), .C2(
        n6638), .ZN(n6611) );
  INV_X1 U7575 ( .A(n6611), .ZN(U3194) );
  AOI22_X1 U7576 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6674), .ZN(n6612) );
  OAI21_X1 U7577 ( .B1(n6613), .B2(n6643), .A(n6612), .ZN(U3195) );
  AOI22_X1 U7578 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6684), .ZN(n6614) );
  OAI21_X1 U7579 ( .B1(n6989), .B2(n6640), .A(n6614), .ZN(U3196) );
  AOI22_X1 U7580 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6674), .ZN(n6615) );
  OAI21_X1 U7581 ( .B1(n6989), .B2(n6643), .A(n6615), .ZN(U3197) );
  AOI22_X1 U7582 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6674), .ZN(n6616) );
  OAI21_X1 U7583 ( .B1(n6617), .B2(n6643), .A(n6616), .ZN(U3198) );
  AOI22_X1 U7584 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6674), .ZN(n6618) );
  OAI21_X1 U7585 ( .B1(n6912), .B2(n6643), .A(n6618), .ZN(U3199) );
  AOI22_X1 U7586 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6684), .ZN(n6619) );
  OAI21_X1 U7587 ( .B1(n6620), .B2(n6640), .A(n6619), .ZN(U3200) );
  AOI22_X1 U7588 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6674), .ZN(n6621) );
  OAI21_X1 U7589 ( .B1(n6623), .B2(n6640), .A(n6621), .ZN(U3201) );
  AOI22_X1 U7590 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6684), .ZN(n6622) );
  OAI21_X1 U7591 ( .B1(n6623), .B2(n6643), .A(n6622), .ZN(U3202) );
  AOI22_X1 U7592 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6674), .ZN(n6624) );
  OAI21_X1 U7593 ( .B1(n6625), .B2(n6640), .A(n6624), .ZN(U3203) );
  AOI22_X1 U7594 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6684), .ZN(n6626) );
  OAI21_X1 U7595 ( .B1(n6628), .B2(n6640), .A(n6626), .ZN(U3204) );
  AOI22_X1 U7596 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6674), .ZN(n6627) );
  OAI21_X1 U7597 ( .B1(n6628), .B2(n6643), .A(n6627), .ZN(U3205) );
  AOI22_X1 U7598 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6674), .ZN(n6629) );
  OAI21_X1 U7599 ( .B1(n6903), .B2(n6643), .A(n6629), .ZN(U3206) );
  AOI22_X1 U7600 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6684), .ZN(n6630) );
  OAI21_X1 U7601 ( .B1(n6925), .B2(n6643), .A(n6630), .ZN(U3207) );
  AOI22_X1 U7602 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6674), .ZN(n6631) );
  OAI21_X1 U7603 ( .B1(n6632), .B2(n6643), .A(n6631), .ZN(U3208) );
  AOI22_X1 U7604 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6684), .ZN(n6633) );
  OAI21_X1 U7605 ( .B1(n6634), .B2(n6640), .A(n6633), .ZN(U3209) );
  AOI22_X1 U7606 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6684), .ZN(n6635) );
  OAI21_X1 U7607 ( .B1(n6778), .B2(n6640), .A(n6635), .ZN(U3210) );
  AOI22_X1 U7608 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6684), .ZN(n6636) );
  OAI21_X1 U7609 ( .B1(n6637), .B2(n6640), .A(n6636), .ZN(U3211) );
  AOI22_X1 U7610 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6638), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6684), .ZN(n6639) );
  OAI21_X1 U7611 ( .B1(n6644), .B2(n6640), .A(n6639), .ZN(U3212) );
  AOI22_X1 U7612 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6641), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6684), .ZN(n6642) );
  OAI21_X1 U7613 ( .B1(n6644), .B2(n6643), .A(n6642), .ZN(U3213) );
  MUX2_X1 U7614 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6684), .Z(U3445) );
  OAI22_X1 U7615 ( .A1(n6684), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n6594), .ZN(n6645) );
  INV_X1 U7616 ( .A(n6645), .ZN(U3446) );
  OAI22_X1 U7617 ( .A1(n6684), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n6594), .ZN(n6646) );
  INV_X1 U7618 ( .A(n6646), .ZN(U3447) );
  MUX2_X1 U7619 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6684), .Z(U3448) );
  OAI21_X1 U7620 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6650), .A(n6648), .ZN(
        n6647) );
  INV_X1 U7621 ( .A(n6647), .ZN(U3451) );
  OAI21_X1 U7622 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(U3452) );
  INV_X1 U7623 ( .A(n6651), .ZN(n6654) );
  OAI211_X1 U7624 ( .C1(n6942), .C2(n6654), .A(n6653), .B(n6652), .ZN(U3453)
         );
  AOI21_X1 U7625 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n4406), .A(n6655), .ZN(
        n6656) );
  OAI211_X1 U7626 ( .C1(n6657), .C2(n6661), .A(n6659), .B(n6656), .ZN(n6658)
         );
  OAI21_X1 U7627 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6659), .A(n6658), 
        .ZN(n6660) );
  OAI21_X1 U7628 ( .B1(n6662), .B2(n6661), .A(n6660), .ZN(U3461) );
  NAND2_X1 U7629 ( .A1(n6663), .A2(n6664), .ZN(n6670) );
  INV_X1 U7630 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6665) );
  OAI21_X1 U7631 ( .B1(n6665), .B2(n6664), .A(n6671), .ZN(n6666) );
  OAI21_X1 U7632 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6671), .A(n6666), .ZN(
        n6667) );
  OAI221_X1 U7633 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6669), .C1(n6668), 
        .C2(n6670), .A(n6667), .ZN(U3468) );
  OAI21_X1 U7634 ( .B1(n6671), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6670), .ZN(
        n6672) );
  INV_X1 U7635 ( .A(n6672), .ZN(U3469) );
  NAND2_X1 U7636 ( .A1(n6674), .A2(W_R_N_REG_SCAN_IN), .ZN(n6673) );
  OAI21_X1 U7637 ( .B1(n6674), .B2(READREQUEST_REG_SCAN_IN), .A(n6673), .ZN(
        U3470) );
  AOI211_X1 U7638 ( .C1(n6677), .C2(n6892), .A(n6676), .B(n6675), .ZN(n6683)
         );
  OAI211_X1 U7639 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3395), .A(n6678), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6680) );
  AOI21_X1 U7640 ( .B1(n6680), .B2(STATE2_REG_0__SCAN_IN), .A(n6679), .ZN(
        n6682) );
  NAND2_X1 U7641 ( .A1(n6683), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6681) );
  OAI21_X1 U7642 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(U3472) );
  MUX2_X1 U7643 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6684), .Z(U3473) );
  AOI22_X1 U7644 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6686), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6685), .ZN(n6691) );
  AOI22_X1 U7645 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6689), .B1(n6688), .B2(
        n6687), .ZN(n6690) );
  OAI211_X1 U7646 ( .C1(n6693), .C2(n6692), .A(n6691), .B(n6690), .ZN(n6694)
         );
  AOI211_X1 U7647 ( .C1(n6697), .C2(n6696), .A(n6695), .B(n6694), .ZN(n7025)
         );
  INV_X1 U7648 ( .A(keyinput75), .ZN(n6699) );
  AOI22_X1 U7649 ( .A1(n4442), .A2(keyinput16), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(n6699), .ZN(n6698) );
  OAI221_X1 U7650 ( .B1(n4442), .B2(keyinput16), .C1(n6699), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6698), .ZN(n6711) );
  INV_X1 U7651 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U7652 ( .A1(n6702), .A2(keyinput35), .B1(n6701), .B2(keyinput13), 
        .ZN(n6700) );
  OAI221_X1 U7653 ( .B1(n6702), .B2(keyinput35), .C1(n6701), .C2(keyinput13), 
        .A(n6700), .ZN(n6710) );
  AOI22_X1 U7654 ( .A1(n4848), .A2(keyinput77), .B1(keyinput32), .B2(n6704), 
        .ZN(n6703) );
  OAI221_X1 U7655 ( .B1(n4848), .B2(keyinput77), .C1(n6704), .C2(keyinput32), 
        .A(n6703), .ZN(n6709) );
  AOI22_X1 U7656 ( .A1(n6707), .A2(keyinput69), .B1(n6706), .B2(keyinput89), 
        .ZN(n6705) );
  OAI221_X1 U7657 ( .B1(n6707), .B2(keyinput69), .C1(n6706), .C2(keyinput89), 
        .A(n6705), .ZN(n6708) );
  NOR4_X1 U7658 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n7023)
         );
  INV_X1 U7659 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6714) );
  AOI22_X1 U7660 ( .A1(keyinput12), .A2(n6712), .B1(keyinput15), .B2(n6714), 
        .ZN(n6713) );
  OAI21_X1 U7661 ( .B1(keyinput15), .B2(n6714), .A(n6713), .ZN(n6727) );
  INV_X1 U7662 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6717) );
  INV_X1 U7663 ( .A(keyinput85), .ZN(n6716) );
  AOI22_X1 U7664 ( .A1(n6717), .A2(keyinput84), .B1(ADDRESS_REG_10__SCAN_IN), 
        .B2(n6716), .ZN(n6715) );
  OAI221_X1 U7665 ( .B1(n6717), .B2(keyinput84), .C1(n6716), .C2(
        ADDRESS_REG_10__SCAN_IN), .A(n6715), .ZN(n6726) );
  INV_X1 U7666 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6720) );
  INV_X1 U7667 ( .A(keyinput79), .ZN(n6719) );
  AOI22_X1 U7668 ( .A1(n6720), .A2(keyinput53), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n6719), .ZN(n6718) );
  OAI221_X1 U7669 ( .B1(n6720), .B2(keyinput53), .C1(n6719), .C2(
        DATAO_REG_16__SCAN_IN), .A(n6718), .ZN(n6725) );
  INV_X1 U7670 ( .A(keyinput97), .ZN(n6722) );
  AOI22_X1 U7671 ( .A1(n6723), .A2(keyinput88), .B1(DATAWIDTH_REG_15__SCAN_IN), 
        .B2(n6722), .ZN(n6721) );
  OAI221_X1 U7672 ( .B1(n6723), .B2(keyinput88), .C1(n6722), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6721), .ZN(n6724) );
  NOR4_X1 U7673 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n7022)
         );
  INV_X1 U7674 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6730) );
  INV_X1 U7675 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6729) );
  AOI22_X1 U7676 ( .A1(n6730), .A2(keyinput109), .B1(keyinput56), .B2(n6729), 
        .ZN(n6728) );
  OAI221_X1 U7677 ( .B1(n6730), .B2(keyinput109), .C1(n6729), .C2(keyinput56), 
        .A(n6728), .ZN(n6825) );
  AOI22_X1 U7678 ( .A1(n6733), .A2(keyinput66), .B1(n6732), .B2(keyinput28), 
        .ZN(n6731) );
  OAI221_X1 U7679 ( .B1(n6733), .B2(keyinput66), .C1(n6732), .C2(keyinput28), 
        .A(n6731), .ZN(n6824) );
  INV_X1 U7680 ( .A(keyinput34), .ZN(n6735) );
  OAI22_X1 U7681 ( .A1(keyinput68), .A2(n6736), .B1(n6735), .B2(DATAI_17_), 
        .ZN(n6734) );
  AOI221_X1 U7682 ( .B1(n6736), .B2(keyinput68), .C1(n6735), .C2(DATAI_17_), 
        .A(n6734), .ZN(n6755) );
  OAI22_X1 U7683 ( .A1(n5487), .A2(keyinput80), .B1(n6738), .B2(keyinput8), 
        .ZN(n6737) );
  AOI221_X1 U7684 ( .B1(n5487), .B2(keyinput80), .C1(keyinput8), .C2(n6738), 
        .A(n6737), .ZN(n6754) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7686 ( .A1(n5212), .A2(keyinput91), .B1(n6740), .B2(keyinput61), 
        .ZN(n6739) );
  OAI221_X1 U7687 ( .B1(n5212), .B2(keyinput91), .C1(n6740), .C2(keyinput61), 
        .A(n6739), .ZN(n6752) );
  INV_X1 U7688 ( .A(keyinput45), .ZN(n6742) );
  AOI22_X1 U7689 ( .A1(n6743), .A2(keyinput122), .B1(DATAO_REG_8__SCAN_IN), 
        .B2(n6742), .ZN(n6741) );
  OAI221_X1 U7690 ( .B1(n6743), .B2(keyinput122), .C1(n6742), .C2(
        DATAO_REG_8__SCAN_IN), .A(n6741), .ZN(n6751) );
  INV_X1 U7691 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7692 ( .A1(n6745), .A2(keyinput92), .B1(n4852), .B2(keyinput87), 
        .ZN(n6744) );
  OAI221_X1 U7693 ( .B1(n6745), .B2(keyinput92), .C1(n4852), .C2(keyinput87), 
        .A(n6744), .ZN(n6750) );
  INV_X1 U7694 ( .A(keyinput90), .ZN(n6747) );
  AOI22_X1 U7695 ( .A1(n6748), .A2(keyinput37), .B1(BE_N_REG_0__SCAN_IN), .B2(
        n6747), .ZN(n6746) );
  OAI221_X1 U7696 ( .B1(n6748), .B2(keyinput37), .C1(n6747), .C2(
        BE_N_REG_0__SCAN_IN), .A(n6746), .ZN(n6749) );
  NOR4_X1 U7697 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6753)
         );
  NAND3_X1 U7698 ( .A1(n6755), .A2(n6754), .A3(n6753), .ZN(n6823) );
  AOI22_X1 U7699 ( .A1(n6757), .A2(keyinput7), .B1(n3520), .B2(keyinput111), 
        .ZN(n6756) );
  OAI221_X1 U7700 ( .B1(n6757), .B2(keyinput7), .C1(n3520), .C2(keyinput111), 
        .A(n6756), .ZN(n6769) );
  INV_X1 U7701 ( .A(keyinput55), .ZN(n6759) );
  AOI22_X1 U7702 ( .A1(n6760), .A2(keyinput46), .B1(DATAWIDTH_REG_28__SCAN_IN), 
        .B2(n6759), .ZN(n6758) );
  OAI221_X1 U7703 ( .B1(n6760), .B2(keyinput46), .C1(n6759), .C2(
        DATAWIDTH_REG_28__SCAN_IN), .A(n6758), .ZN(n6768) );
  INV_X1 U7704 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7705 ( .A1(n6763), .A2(keyinput114), .B1(keyinput123), .B2(n6762), 
        .ZN(n6761) );
  OAI221_X1 U7706 ( .B1(n6763), .B2(keyinput114), .C1(n6762), .C2(keyinput123), 
        .A(n6761), .ZN(n6767) );
  XOR2_X1 U7707 ( .A(n4276), .B(keyinput40), .Z(n6765) );
  XNOR2_X1 U7708 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput70), .ZN(
        n6764) );
  NAND2_X1 U7709 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  NOR4_X1 U7710 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6821)
         );
  INV_X1 U7711 ( .A(keyinput65), .ZN(n6771) );
  AOI22_X1 U7712 ( .A1(n6772), .A2(keyinput30), .B1(DATAI_19_), .B2(n6771), 
        .ZN(n6770) );
  OAI221_X1 U7713 ( .B1(n6772), .B2(keyinput30), .C1(n6771), .C2(DATAI_19_), 
        .A(n6770), .ZN(n6785) );
  INV_X1 U7714 ( .A(keyinput71), .ZN(n6774) );
  AOI22_X1 U7715 ( .A1(n6775), .A2(keyinput98), .B1(UWORD_REG_3__SCAN_IN), 
        .B2(n6774), .ZN(n6773) );
  OAI221_X1 U7716 ( .B1(n6775), .B2(keyinput98), .C1(n6774), .C2(
        UWORD_REG_3__SCAN_IN), .A(n6773), .ZN(n6784) );
  INV_X1 U7717 ( .A(keyinput102), .ZN(n6777) );
  AOI22_X1 U7718 ( .A1(n6778), .A2(keyinput127), .B1(DATAWIDTH_REG_1__SCAN_IN), 
        .B2(n6777), .ZN(n6776) );
  OAI221_X1 U7719 ( .B1(n6778), .B2(keyinput127), .C1(n6777), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(n6776), .ZN(n6783) );
  AOI22_X1 U7720 ( .A1(n6781), .A2(keyinput126), .B1(n6780), .B2(keyinput50), 
        .ZN(n6779) );
  OAI221_X1 U7721 ( .B1(n6781), .B2(keyinput126), .C1(n6780), .C2(keyinput50), 
        .A(n6779), .ZN(n6782) );
  NOR4_X1 U7722 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6820)
         );
  INV_X1 U7723 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6788) );
  INV_X1 U7724 ( .A(keyinput31), .ZN(n6787) );
  AOI22_X1 U7725 ( .A1(n6788), .A2(keyinput110), .B1(DATAI_4_), .B2(n6787), 
        .ZN(n6786) );
  OAI221_X1 U7726 ( .B1(n6788), .B2(keyinput110), .C1(n6787), .C2(DATAI_4_), 
        .A(n6786), .ZN(n6801) );
  AOI22_X1 U7727 ( .A1(n6791), .A2(keyinput19), .B1(keyinput39), .B2(n6790), 
        .ZN(n6789) );
  OAI221_X1 U7728 ( .B1(n6791), .B2(keyinput19), .C1(n6790), .C2(keyinput39), 
        .A(n6789), .ZN(n6800) );
  INV_X1 U7729 ( .A(keyinput25), .ZN(n6793) );
  AOI22_X1 U7730 ( .A1(n6794), .A2(keyinput72), .B1(MEMORYFETCH_REG_SCAN_IN), 
        .B2(n6793), .ZN(n6792) );
  OAI221_X1 U7731 ( .B1(n6794), .B2(keyinput72), .C1(n6793), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6792), .ZN(n6799) );
  INV_X1 U7732 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6797) );
  INV_X1 U7733 ( .A(keyinput120), .ZN(n6796) );
  AOI22_X1 U7734 ( .A1(n6797), .A2(keyinput67), .B1(ADDRESS_REG_6__SCAN_IN), 
        .B2(n6796), .ZN(n6795) );
  OAI221_X1 U7735 ( .B1(n6797), .B2(keyinput67), .C1(n6796), .C2(
        ADDRESS_REG_6__SCAN_IN), .A(n6795), .ZN(n6798) );
  NOR4_X1 U7736 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6819)
         );
  AOI22_X1 U7737 ( .A1(n6804), .A2(keyinput2), .B1(n6803), .B2(keyinput104), 
        .ZN(n6802) );
  OAI221_X1 U7738 ( .B1(n6804), .B2(keyinput2), .C1(n6803), .C2(keyinput104), 
        .A(n6802), .ZN(n6817) );
  INV_X1 U7739 ( .A(keyinput3), .ZN(n6806) );
  AOI22_X1 U7740 ( .A1(n6807), .A2(keyinput96), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n6806), .ZN(n6805) );
  OAI221_X1 U7741 ( .B1(n6807), .B2(keyinput96), .C1(n6806), .C2(
        DATAO_REG_25__SCAN_IN), .A(n6805), .ZN(n6816) );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6809) );
  AOI22_X1 U7743 ( .A1(n6810), .A2(keyinput6), .B1(n6809), .B2(keyinput29), 
        .ZN(n6808) );
  OAI221_X1 U7744 ( .B1(n6810), .B2(keyinput6), .C1(n6809), .C2(keyinput29), 
        .A(n6808), .ZN(n6815) );
  XOR2_X1 U7745 ( .A(n6811), .B(keyinput27), .Z(n6813) );
  XNOR2_X1 U7746 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput36), .ZN(
        n6812) );
  NAND2_X1 U7747 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NOR4_X1 U7748 ( .A1(n6817), .A2(n6816), .A3(n6815), .A4(n6814), .ZN(n6818)
         );
  NAND4_X1 U7749 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6822)
         );
  NOR4_X1 U7750 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .ZN(n7021)
         );
  INV_X1 U7751 ( .A(keyinput77), .ZN(n6826) );
  NAND4_X1 U7752 ( .A1(keyinput69), .A2(keyinput75), .A3(keyinput89), .A4(
        n6826), .ZN(n6827) );
  NOR3_X1 U7753 ( .A1(keyinput79), .A2(keyinput35), .A3(n6827), .ZN(n6839) );
  NAND2_X1 U7754 ( .A1(keyinput126), .A2(keyinput71), .ZN(n6828) );
  NOR3_X1 U7755 ( .A1(keyinput30), .A2(keyinput65), .A3(n6828), .ZN(n6829) );
  NAND3_X1 U7756 ( .A1(keyinput32), .A2(keyinput98), .A3(n6829), .ZN(n6837) );
  INV_X1 U7757 ( .A(keyinput88), .ZN(n6830) );
  NAND4_X1 U7758 ( .A1(keyinput84), .A2(keyinput85), .A3(keyinput53), .A4(
        n6830), .ZN(n6831) );
  NOR4_X1 U7759 ( .A1(keyinput101), .A2(keyinput15), .A3(keyinput97), .A4(
        n6831), .ZN(n6835) );
  NOR2_X1 U7760 ( .A1(keyinput102), .A2(keyinput114), .ZN(n6832) );
  NAND3_X1 U7761 ( .A1(keyinput55), .A2(keyinput111), .A3(n6832), .ZN(n6833)
         );
  NOR3_X1 U7762 ( .A1(keyinput46), .A2(keyinput70), .A3(n6833), .ZN(n6834) );
  NAND4_X1 U7763 ( .A1(n6835), .A2(keyinput40), .A3(keyinput7), .A4(n6834), 
        .ZN(n6836) );
  NOR4_X1 U7764 ( .A1(keyinput50), .A2(keyinput127), .A3(n6837), .A4(n6836), 
        .ZN(n6838) );
  NAND4_X1 U7765 ( .A1(keyinput13), .A2(keyinput16), .A3(n6839), .A4(n6838), 
        .ZN(n6887) );
  NAND2_X1 U7766 ( .A1(keyinput108), .A2(keyinput81), .ZN(n6840) );
  NOR3_X1 U7767 ( .A1(keyinput124), .A2(keyinput23), .A3(n6840), .ZN(n6885) );
  NOR4_X1 U7768 ( .A1(keyinput112), .A2(keyinput63), .A3(keyinput59), .A4(
        keyinput1), .ZN(n6884) );
  NAND2_X1 U7769 ( .A1(keyinput10), .A2(keyinput25), .ZN(n6841) );
  NOR3_X1 U7770 ( .A1(keyinput83), .A2(keyinput86), .A3(n6841), .ZN(n6842) );
  NAND3_X1 U7771 ( .A1(keyinput43), .A2(keyinput18), .A3(n6842), .ZN(n6851) );
  INV_X1 U7772 ( .A(keyinput0), .ZN(n6920) );
  NOR4_X1 U7773 ( .A1(keyinput107), .A2(keyinput64), .A3(keyinput76), .A4(
        n6920), .ZN(n6849) );
  NAND2_X1 U7774 ( .A1(keyinput58), .A2(keyinput95), .ZN(n6843) );
  NOR3_X1 U7775 ( .A1(keyinput78), .A2(keyinput4), .A3(n6843), .ZN(n6848) );
  NAND2_X1 U7776 ( .A1(keyinput33), .A2(keyinput103), .ZN(n6844) );
  NOR3_X1 U7777 ( .A1(keyinput118), .A2(keyinput74), .A3(n6844), .ZN(n6847) );
  NAND2_X1 U7778 ( .A1(keyinput41), .A2(keyinput5), .ZN(n6845) );
  NOR3_X1 U7779 ( .A1(keyinput17), .A2(keyinput24), .A3(n6845), .ZN(n6846) );
  NAND4_X1 U7780 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6850)
         );
  NOR4_X1 U7781 ( .A1(keyinput49), .A2(keyinput105), .A3(n6851), .A4(n6850), 
        .ZN(n6883) );
  NAND4_X1 U7782 ( .A1(keyinput68), .A2(keyinput34), .A3(keyinput8), .A4(
        keyinput66), .ZN(n6881) );
  NOR2_X1 U7783 ( .A1(keyinput123), .A2(keyinput28), .ZN(n6852) );
  NAND3_X1 U7784 ( .A1(keyinput80), .A2(keyinput109), .A3(n6852), .ZN(n6880)
         );
  NOR4_X1 U7785 ( .A1(keyinput3), .A2(keyinput36), .A3(keyinput27), .A4(
        keyinput6), .ZN(n6863) );
  NAND2_X1 U7786 ( .A1(keyinput2), .A2(keyinput96), .ZN(n6853) );
  NOR3_X1 U7787 ( .A1(keyinput87), .A2(keyinput29), .A3(n6853), .ZN(n6862) );
  NAND4_X1 U7788 ( .A1(keyinput61), .A2(keyinput37), .A3(keyinput90), .A4(
        keyinput92), .ZN(n6860) );
  NOR2_X1 U7789 ( .A1(keyinput56), .A2(keyinput122), .ZN(n6854) );
  NAND3_X1 U7790 ( .A1(keyinput45), .A2(keyinput91), .A3(n6854), .ZN(n6859) );
  NOR2_X1 U7791 ( .A1(keyinput67), .A2(keyinput120), .ZN(n6855) );
  NAND3_X1 U7792 ( .A1(keyinput31), .A2(keyinput72), .A3(n6855), .ZN(n6858) );
  NOR2_X1 U7793 ( .A1(keyinput19), .A2(keyinput110), .ZN(n6856) );
  NAND3_X1 U7794 ( .A1(keyinput104), .A2(keyinput39), .A3(n6856), .ZN(n6857)
         );
  NOR4_X1 U7795 ( .A1(n6860), .A2(n6859), .A3(n6858), .A4(n6857), .ZN(n6861)
         );
  NAND3_X1 U7796 ( .A1(n6863), .A2(n6862), .A3(n6861), .ZN(n6879) );
  NOR2_X1 U7797 ( .A1(keyinput51), .A2(keyinput93), .ZN(n6864) );
  NAND3_X1 U7798 ( .A1(keyinput9), .A2(keyinput47), .A3(n6864), .ZN(n6865) );
  NOR3_X1 U7799 ( .A1(keyinput94), .A2(keyinput26), .A3(n6865), .ZN(n6877) );
  NAND4_X1 U7800 ( .A1(keyinput117), .A2(keyinput38), .A3(keyinput121), .A4(
        keyinput60), .ZN(n6875) );
  NOR2_X1 U7801 ( .A1(keyinput113), .A2(keyinput52), .ZN(n6866) );
  NAND3_X1 U7802 ( .A1(keyinput20), .A2(keyinput42), .A3(n6866), .ZN(n6874) );
  NAND2_X1 U7803 ( .A1(keyinput125), .A2(keyinput62), .ZN(n6867) );
  NOR3_X1 U7804 ( .A1(keyinput82), .A2(keyinput116), .A3(n6867), .ZN(n6872) );
  INV_X1 U7805 ( .A(keyinput22), .ZN(n6970) );
  NOR4_X1 U7806 ( .A1(keyinput106), .A2(keyinput73), .A3(keyinput11), .A4(
        n6970), .ZN(n6871) );
  NOR4_X1 U7807 ( .A1(keyinput54), .A2(keyinput119), .A3(keyinput14), .A4(
        keyinput100), .ZN(n6870) );
  NAND2_X1 U7808 ( .A1(keyinput57), .A2(keyinput21), .ZN(n6868) );
  NOR3_X1 U7809 ( .A1(keyinput44), .A2(keyinput115), .A3(n6868), .ZN(n6869) );
  NAND4_X1 U7810 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6873)
         );
  NOR3_X1 U7811 ( .A1(n6875), .A2(n6874), .A3(n6873), .ZN(n6876) );
  NAND4_X1 U7812 ( .A1(keyinput48), .A2(keyinput99), .A3(n6877), .A4(n6876), 
        .ZN(n6878) );
  NOR4_X1 U7813 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6882)
         );
  NAND4_X1 U7814 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6886)
         );
  OAI21_X1 U7815 ( .B1(n6887), .B2(n6886), .A(keyinput12), .ZN(n7019) );
  INV_X1 U7816 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6889) );
  AOI22_X1 U7817 ( .A1(n6889), .A2(keyinput86), .B1(keyinput49), .B2(n4550), 
        .ZN(n6888) );
  OAI221_X1 U7818 ( .B1(n6889), .B2(keyinput86), .C1(n4550), .C2(keyinput49), 
        .A(n6888), .ZN(n6901) );
  INV_X1 U7819 ( .A(keyinput83), .ZN(n6891) );
  AOI22_X1 U7820 ( .A1(n6892), .A2(keyinput105), .B1(ADDRESS_REG_25__SCAN_IN), 
        .B2(n6891), .ZN(n6890) );
  OAI221_X1 U7821 ( .B1(n6892), .B2(keyinput105), .C1(n6891), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n6890), .ZN(n6900) );
  INV_X1 U7822 ( .A(keyinput10), .ZN(n6894) );
  AOI22_X1 U7823 ( .A1(n6895), .A2(keyinput43), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n6894), .ZN(n6893) );
  OAI221_X1 U7824 ( .B1(n6895), .B2(keyinput43), .C1(n6894), .C2(
        DATAO_REG_23__SCAN_IN), .A(n6893), .ZN(n6899) );
  INV_X1 U7825 ( .A(keyinput112), .ZN(n6897) );
  AOI22_X1 U7826 ( .A1(n4828), .A2(keyinput18), .B1(DATAI_20_), .B2(n6897), 
        .ZN(n6896) );
  OAI221_X1 U7827 ( .B1(n4828), .B2(keyinput18), .C1(n6897), .C2(DATAI_20_), 
        .A(n6896), .ZN(n6898) );
  NOR4_X1 U7828 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6951)
         );
  AOI22_X1 U7829 ( .A1(n6904), .A2(keyinput63), .B1(keyinput59), .B2(n6903), 
        .ZN(n6902) );
  OAI221_X1 U7830 ( .B1(n6904), .B2(keyinput63), .C1(n6903), .C2(keyinput59), 
        .A(n6902), .ZN(n6917) );
  INV_X1 U7831 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6907) );
  INV_X1 U7832 ( .A(keyinput124), .ZN(n6906) );
  AOI22_X1 U7833 ( .A1(n6907), .A2(keyinput1), .B1(BYTEENABLE_REG_1__SCAN_IN), 
        .B2(n6906), .ZN(n6905) );
  OAI221_X1 U7834 ( .B1(n6907), .B2(keyinput1), .C1(n6906), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6905), .ZN(n6916) );
  INV_X1 U7835 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n6910) );
  INV_X1 U7836 ( .A(keyinput81), .ZN(n6909) );
  AOI22_X1 U7837 ( .A1(n6910), .A2(keyinput108), .B1(DATAWIDTH_REG_3__SCAN_IN), 
        .B2(n6909), .ZN(n6908) );
  OAI221_X1 U7838 ( .B1(n6910), .B2(keyinput108), .C1(n6909), .C2(
        DATAWIDTH_REG_3__SCAN_IN), .A(n6908), .ZN(n6915) );
  AOI22_X1 U7839 ( .A1(n6913), .A2(keyinput23), .B1(keyinput95), .B2(n6912), 
        .ZN(n6911) );
  OAI221_X1 U7840 ( .B1(n6913), .B2(keyinput23), .C1(n6912), .C2(keyinput95), 
        .A(n6911), .ZN(n6914) );
  NOR4_X1 U7841 ( .A1(n6917), .A2(n6916), .A3(n6915), .A4(n6914), .ZN(n6950)
         );
  INV_X1 U7842 ( .A(keyinput17), .ZN(n6919) );
  AOI22_X1 U7843 ( .A1(n6920), .A2(LWORD_REG_9__SCAN_IN), .B1(
        DATAWIDTH_REG_22__SCAN_IN), .B2(n6919), .ZN(n6918) );
  OAI221_X1 U7844 ( .B1(n6920), .B2(LWORD_REG_9__SCAN_IN), .C1(n6919), .C2(
        DATAWIDTH_REG_22__SCAN_IN), .A(n6918), .ZN(n6932) );
  AOI22_X1 U7845 ( .A1(n6922), .A2(keyinput64), .B1(keyinput76), .B2(n6499), 
        .ZN(n6921) );
  OAI221_X1 U7846 ( .B1(n6922), .B2(keyinput64), .C1(n6499), .C2(keyinput76), 
        .A(n6921), .ZN(n6931) );
  INV_X1 U7847 ( .A(keyinput78), .ZN(n6924) );
  AOI22_X1 U7848 ( .A1(n6925), .A2(keyinput58), .B1(DATAI_6_), .B2(n6924), 
        .ZN(n6923) );
  OAI221_X1 U7849 ( .B1(n6925), .B2(keyinput58), .C1(n6924), .C2(DATAI_6_), 
        .A(n6923), .ZN(n6930) );
  INV_X1 U7850 ( .A(keyinput107), .ZN(n6926) );
  XOR2_X1 U7851 ( .A(ADDRESS_REG_2__SCAN_IN), .B(n6926), .Z(n6928) );
  XNOR2_X1 U7852 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput4), .ZN(
        n6927) );
  NAND2_X1 U7853 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  NOR4_X1 U7854 ( .A1(n6932), .A2(n6931), .A3(n6930), .A4(n6929), .ZN(n6949)
         );
  INV_X1 U7855 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U7856 ( .A1(n6934), .A2(keyinput5), .B1(keyinput41), .B2(n5608), 
        .ZN(n6933) );
  OAI221_X1 U7857 ( .B1(n6934), .B2(keyinput5), .C1(n5608), .C2(keyinput41), 
        .A(n6933), .ZN(n6947) );
  INV_X1 U7858 ( .A(keyinput24), .ZN(n6936) );
  AOI22_X1 U7859 ( .A1(n6937), .A2(keyinput118), .B1(UWORD_REG_14__SCAN_IN), 
        .B2(n6936), .ZN(n6935) );
  OAI221_X1 U7860 ( .B1(n6937), .B2(keyinput118), .C1(n6936), .C2(
        UWORD_REG_14__SCAN_IN), .A(n6935), .ZN(n6946) );
  INV_X1 U7861 ( .A(keyinput103), .ZN(n6939) );
  AOI22_X1 U7862 ( .A1(n6940), .A2(keyinput74), .B1(DATAI_15_), .B2(n6939), 
        .ZN(n6938) );
  OAI221_X1 U7863 ( .B1(n6940), .B2(keyinput74), .C1(n6939), .C2(DATAI_15_), 
        .A(n6938), .ZN(n6945) );
  AOI22_X1 U7864 ( .A1(n6943), .A2(keyinput33), .B1(n6942), .B2(keyinput113), 
        .ZN(n6941) );
  OAI221_X1 U7865 ( .B1(n6943), .B2(keyinput33), .C1(n6942), .C2(keyinput113), 
        .A(n6941), .ZN(n6944) );
  NOR4_X1 U7866 ( .A1(n6947), .A2(n6946), .A3(n6945), .A4(n6944), .ZN(n6948)
         );
  NAND4_X1 U7867 ( .A1(n6951), .A2(n6950), .A3(n6949), .A4(n6948), .ZN(n7018)
         );
  INV_X1 U7868 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7869 ( .A1(n6954), .A2(keyinput20), .B1(keyinput117), .B2(n6953), 
        .ZN(n6952) );
  OAI221_X1 U7870 ( .B1(n6954), .B2(keyinput20), .C1(n6953), .C2(keyinput117), 
        .A(n6952), .ZN(n6967) );
  AOI22_X1 U7871 ( .A1(n6957), .A2(keyinput38), .B1(keyinput52), .B2(n6956), 
        .ZN(n6955) );
  OAI221_X1 U7872 ( .B1(n6957), .B2(keyinput38), .C1(n6956), .C2(keyinput52), 
        .A(n6955), .ZN(n6966) );
  INV_X1 U7873 ( .A(keyinput121), .ZN(n6959) );
  AOI22_X1 U7874 ( .A1(n6960), .A2(keyinput42), .B1(ADDRESS_REG_3__SCAN_IN), 
        .B2(n6959), .ZN(n6958) );
  OAI221_X1 U7875 ( .B1(n6960), .B2(keyinput42), .C1(n6959), .C2(
        ADDRESS_REG_3__SCAN_IN), .A(n6958), .ZN(n6965) );
  INV_X1 U7876 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6963) );
  INV_X1 U7877 ( .A(keyinput106), .ZN(n6962) );
  AOI22_X1 U7878 ( .A1(n6963), .A2(keyinput60), .B1(UWORD_REG_11__SCAN_IN), 
        .B2(n6962), .ZN(n6961) );
  OAI221_X1 U7879 ( .B1(n6963), .B2(keyinput60), .C1(n6962), .C2(
        UWORD_REG_11__SCAN_IN), .A(n6961), .ZN(n6964) );
  NOR4_X1 U7880 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n7016)
         );
  INV_X1 U7881 ( .A(keyinput73), .ZN(n6969) );
  AOI22_X1 U7882 ( .A1(n6970), .A2(UWORD_REG_6__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n6969), .ZN(n6968) );
  OAI221_X1 U7883 ( .B1(n6970), .B2(UWORD_REG_6__SCAN_IN), .C1(n6969), .C2(
        BE_N_REG_1__SCAN_IN), .A(n6968), .ZN(n6981) );
  AOI22_X1 U7884 ( .A1(n6973), .A2(keyinput11), .B1(n6972), .B2(keyinput62), 
        .ZN(n6971) );
  OAI221_X1 U7885 ( .B1(n6973), .B2(keyinput11), .C1(n6972), .C2(keyinput62), 
        .A(n6971), .ZN(n6980) );
  AOI22_X1 U7886 ( .A1(n5572), .A2(keyinput82), .B1(n5738), .B2(keyinput125), 
        .ZN(n6974) );
  OAI221_X1 U7887 ( .B1(n5572), .B2(keyinput82), .C1(n5738), .C2(keyinput125), 
        .A(n6974), .ZN(n6979) );
  INV_X1 U7888 ( .A(keyinput9), .ZN(n6976) );
  AOI22_X1 U7889 ( .A1(n6977), .A2(keyinput116), .B1(UWORD_REG_7__SCAN_IN), 
        .B2(n6976), .ZN(n6975) );
  OAI221_X1 U7890 ( .B1(n6977), .B2(keyinput116), .C1(n6976), .C2(
        UWORD_REG_7__SCAN_IN), .A(n6975), .ZN(n6978) );
  NOR4_X1 U7891 ( .A1(n6981), .A2(n6980), .A3(n6979), .A4(n6978), .ZN(n7015)
         );
  AOI22_X1 U7892 ( .A1(n4233), .A2(keyinput99), .B1(n6983), .B2(keyinput21), 
        .ZN(n6982) );
  OAI221_X1 U7893 ( .B1(n4233), .B2(keyinput99), .C1(n6983), .C2(keyinput21), 
        .A(n6982), .ZN(n6996) );
  INV_X1 U7894 ( .A(keyinput47), .ZN(n6985) );
  AOI22_X1 U7895 ( .A1(n6986), .A2(keyinput26), .B1(DATAO_REG_11__SCAN_IN), 
        .B2(n6985), .ZN(n6984) );
  OAI221_X1 U7896 ( .B1(n6986), .B2(keyinput26), .C1(n6985), .C2(
        DATAO_REG_11__SCAN_IN), .A(n6984), .ZN(n6995) );
  INV_X1 U7897 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7898 ( .A1(n6989), .A2(keyinput51), .B1(n6988), .B2(keyinput94), 
        .ZN(n6987) );
  OAI221_X1 U7899 ( .B1(n6989), .B2(keyinput51), .C1(n6988), .C2(keyinput94), 
        .A(n6987), .ZN(n6994) );
  INV_X1 U7900 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6990) );
  XOR2_X1 U7901 ( .A(n6990), .B(keyinput93), .Z(n6992) );
  XNOR2_X1 U7902 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput48), .ZN(n6991)
         );
  NAND2_X1 U7903 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  NOR4_X1 U7904 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n7014)
         );
  INV_X1 U7905 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6999) );
  INV_X1 U7906 ( .A(keyinput44), .ZN(n6998) );
  AOI22_X1 U7907 ( .A1(n6999), .A2(keyinput57), .B1(ADDRESS_REG_9__SCAN_IN), 
        .B2(n6998), .ZN(n6997) );
  OAI221_X1 U7908 ( .B1(n6999), .B2(keyinput57), .C1(n6998), .C2(
        ADDRESS_REG_9__SCAN_IN), .A(n6997), .ZN(n7012) );
  INV_X1 U7909 ( .A(keyinput54), .ZN(n7001) );
  AOI22_X1 U7910 ( .A1(n7002), .A2(keyinput115), .B1(DATAO_REG_3__SCAN_IN), 
        .B2(n7001), .ZN(n7000) );
  OAI221_X1 U7911 ( .B1(n7002), .B2(keyinput115), .C1(n7001), .C2(
        DATAO_REG_3__SCAN_IN), .A(n7000), .ZN(n7011) );
  INV_X1 U7912 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n7005) );
  INV_X1 U7913 ( .A(keyinput14), .ZN(n7004) );
  AOI22_X1 U7914 ( .A1(n7005), .A2(keyinput119), .B1(DATAWIDTH_REG_29__SCAN_IN), .B2(n7004), .ZN(n7003) );
  OAI221_X1 U7915 ( .B1(n7005), .B2(keyinput119), .C1(n7004), .C2(
        DATAWIDTH_REG_29__SCAN_IN), .A(n7003), .ZN(n7010) );
  INV_X1 U7916 ( .A(keyinput100), .ZN(n7007) );
  AOI22_X1 U7917 ( .A1(n7008), .A2(keyinput101), .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(n7007), .ZN(n7006) );
  OAI221_X1 U7918 ( .B1(n7008), .B2(keyinput101), .C1(n7007), .C2(
        DATAWIDTH_REG_11__SCAN_IN), .A(n7006), .ZN(n7009) );
  NOR4_X1 U7919 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), .ZN(n7013)
         );
  NAND4_X1 U7920 ( .A1(n7016), .A2(n7015), .A3(n7014), .A4(n7013), .ZN(n7017)
         );
  AOI211_X1 U7921 ( .C1(INSTQUEUE_REG_4__2__SCAN_IN), .C2(n7019), .A(n7018), 
        .B(n7017), .ZN(n7020) );
  NAND4_X1 U7922 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7024)
         );
  XOR2_X1 U7923 ( .A(n7025), .B(n7024), .Z(U2803) );
  CLKBUF_X1 U3570 ( .A(n3365), .Z(n4285) );
  OAI211_X1 U3586 ( .C1(n4038), .C2(n6943), .A(n3995), .B(n3994), .ZN(n3996)
         );
  CLKBUF_X1 U3591 ( .A(n3267), .Z(n4493) );
  NOR2_X2 U3620 ( .A1(n5362), .A2(n5350), .ZN(n5349) );
  CLKBUF_X1 U3649 ( .A(n5161), .Z(n5206) );
  CLKBUF_X1 U3657 ( .A(n5356), .Z(n5539) );
  CLKBUF_X1 U3733 ( .A(n3907), .Z(n4585) );
  CLKBUF_X1 U3763 ( .A(n3914), .Z(n6528) );
  NAND2_X1 U3804 ( .A1(n5475), .A2(n5360), .ZN(n5362) );
  CLKBUF_X1 U3926 ( .A(n6039), .Z(n6049) );
  AOI211_X1 U4162 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5385), .A(n5384), .B(n5383), .ZN(n5386) );
  INV_X2 U5281 ( .A(n6687), .ZN(n5998) );
endmodule

