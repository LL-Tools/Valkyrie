

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591;

  AOI21_X1 U7148 ( .B1(n14682), .B2(n15251), .A(n14681), .ZN(n14986) );
  NAND2_X1 U7150 ( .A1(n12439), .A2(n12438), .ZN(n12437) );
  OAI21_X1 U7151 ( .B1(n13806), .B2(n9223), .A(n9101), .ZN(n13628) );
  BUF_X1 U7152 ( .A(n12696), .Z(n6417) );
  AND2_X1 U7153 ( .A1(n8972), .A2(n8971), .ZN(n14025) );
  XNOR2_X1 U7154 ( .A(n14031), .B(n13884), .ZN(n13913) );
  AND2_X1 U7155 ( .A1(n8956), .A2(n8955), .ZN(n13912) );
  CLKBUF_X2 U7156 ( .A(n13377), .Z(n6404) );
  INV_X1 U7157 ( .A(n11355), .ZN(n11538) );
  NAND2_X1 U7158 ( .A1(n8466), .A2(n8465), .ZN(n11776) );
  CLKBUF_X2 U7159 ( .A(n8772), .Z(n13926) );
  BUF_X1 U7160 ( .A(n12298), .Z(n6402) );
  INV_X1 U7161 ( .A(n6401), .ZN(n11352) );
  INV_X1 U7162 ( .A(n7116), .ZN(n9574) );
  BUF_X4 U7164 ( .A(n10800), .Z(n12203) );
  INV_X2 U7165 ( .A(n8389), .ZN(n8437) );
  INV_X1 U7166 ( .A(n13218), .ZN(n11426) );
  CLKBUF_X2 U7167 ( .A(n13366), .Z(n6408) );
  CLKBUF_X2 U7169 ( .A(n13215), .Z(n6407) );
  INV_X1 U7170 ( .A(n13369), .ZN(n9091) );
  XNOR2_X1 U7171 ( .A(n10106), .B(n10071), .ZN(n10105) );
  AND2_X1 U7172 ( .A1(n13024), .A2(n12055), .ZN(n8051) );
  INV_X2 U7173 ( .A(n6406), .ZN(n9350) );
  NAND2_X1 U7174 ( .A1(n9347), .A2(n10065), .ZN(n9637) );
  INV_X1 U7175 ( .A(n13198), .ZN(n13452) );
  NAND2_X1 U7176 ( .A1(n8697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8699) );
  INV_X1 U7177 ( .A(n13377), .ZN(n13215) );
  AND2_X1 U7178 ( .A1(n7780), .A2(n9758), .ZN(n7779) );
  NAND2_X2 U7179 ( .A1(n14248), .A2(n10758), .ZN(n12273) );
  INV_X1 U7180 ( .A(n11341), .ZN(n6415) );
  CLKBUF_X2 U7181 ( .A(n14253), .Z(n14427) );
  NAND2_X1 U7182 ( .A1(n7204), .A2(n7203), .ZN(n7202) );
  NOR2_X1 U7183 ( .A1(n7975), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U7184 ( .A1(n8456), .A2(n6872), .ZN(n10987) );
  BUF_X1 U7185 ( .A(n9109), .Z(n9282) );
  INV_X1 U7186 ( .A(n9162), .ZN(n9218) );
  AND2_X1 U7187 ( .A1(n7549), .A2(n13872), .ZN(n13803) );
  INV_X1 U7188 ( .A(n12273), .ZN(n12316) );
  NAND2_X1 U7189 ( .A1(n14720), .A2(n14700), .ZN(n14697) );
  OR2_X1 U7190 ( .A1(n14710), .A2(n14750), .ZN(n14751) );
  INV_X1 U7191 ( .A(n14970), .ZN(n14260) );
  OAI21_X1 U7192 ( .B1(n12437), .B2(n7573), .A(n7570), .ZN(n12199) );
  INV_X1 U7193 ( .A(n10431), .ZN(n6875) );
  INV_X1 U7194 ( .A(n10193), .ZN(n9092) );
  INV_X1 U7195 ( .A(n13584), .ZN(n13633) );
  AND2_X1 U7196 ( .A1(n8913), .A2(n8912), .ZN(n13609) );
  INV_X1 U7197 ( .A(n13235), .ZN(n11637) );
  OAI211_X1 U7199 ( .C1(n9160), .C2(n10086), .A(n8783), .B(n8782), .ZN(n15368)
         );
  XNOR2_X1 U7200 ( .A(n8711), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13197) );
  INV_X1 U7201 ( .A(n9376), .ZN(n9786) );
  INV_X2 U7202 ( .A(n11538), .ZN(n12313) );
  NAND2_X1 U7203 ( .A1(n7026), .A2(n11871), .ZN(n12014) );
  NAND2_X1 U7204 ( .A1(n8363), .A2(n8362), .ZN(n12770) );
  XNOR2_X1 U7205 ( .A(n7924), .B(n7923), .ZN(n10880) );
  INV_X1 U7206 ( .A(n11577), .ZN(n14046) );
  OAI21_X1 U7207 ( .B1(n11530), .B2(n9160), .A(n9161), .ZN(n13972) );
  AND2_X1 U7208 ( .A1(n9229), .A2(n9228), .ZN(n13640) );
  BUF_X1 U7209 ( .A(n9970), .Z(n6405) );
  INV_X1 U7210 ( .A(n9384), .ZN(n9844) );
  CLKBUF_X3 U7211 ( .A(n10880), .Z(n13031) );
  AND2_X1 U7213 ( .A1(n9001), .A2(n9000), .ZN(n13878) );
  INV_X1 U7214 ( .A(n15222), .ZN(n15237) );
  AND3_X1 U7215 ( .A1(n6540), .A2(n7912), .A3(n8556), .ZN(n6400) );
  NAND2_X1 U7217 ( .A1(n10741), .A2(n10758), .ZN(n12298) );
  OR2_X2 U7218 ( .A1(n8110), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8124) );
  AND2_X2 U7219 ( .A1(n9328), .A2(n9396), .ZN(n9546) );
  INV_X4 U7220 ( .A(n8784), .ZN(n9079) );
  NAND4_X4 U7221 ( .A1(n8771), .A2(n8770), .A3(n8769), .A4(n8768), .ZN(n13448)
         );
  INV_X2 U7222 ( .A(n8784), .ZN(n8742) );
  NAND3_X2 U7223 ( .A1(n7722), .A2(n7721), .A3(n7719), .ZN(n11829) );
  NAND2_X2 U7224 ( .A1(n10409), .A2(n10408), .ZN(n10716) );
  INV_X4 U7225 ( .A(n8714), .ZN(n10065) );
  NAND2_X1 U7226 ( .A1(n10193), .A2(n6409), .ZN(n9160) );
  OAI211_X2 U7227 ( .C1(n9160), .C2(n10088), .A(n8741), .B(n8740), .ZN(n15361)
         );
  AOI21_X2 U7229 ( .B1(n12842), .B2(n6486), .A(n7488), .ZN(n12795) );
  NAND2_X2 U7230 ( .A1(n8476), .A2(n8475), .ZN(n12842) );
  XNOR2_X2 U7231 ( .A(n10872), .B(n10877), .ZN(n10870) );
  NAND2_X2 U7232 ( .A1(n6982), .A2(n10630), .ZN(n10872) );
  XNOR2_X1 U7233 ( .A(n8161), .B(n8160), .ZN(n11722) );
  XNOR2_X2 U7234 ( .A(n10406), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n10179) );
  NAND2_X2 U7235 ( .A1(n10178), .A2(n10177), .ZN(n10406) );
  AND2_X1 U7236 ( .A1(n13197), .A2(n13196), .ZN(n13377) );
  NAND2_X2 U7237 ( .A1(n10039), .A2(n10038), .ZN(n10051) );
  NAND2_X4 U7238 ( .A1(n10199), .A2(n10205), .ZN(n10193) );
  XNOR2_X2 U7239 ( .A(n8699), .B(n8698), .ZN(n10199) );
  XNOR2_X2 U7240 ( .A(n12525), .B(n11732), .ZN(n12524) );
  NAND2_X2 U7241 ( .A1(n11720), .A2(n11719), .ZN(n12525) );
  OAI211_X2 U7242 ( .C1(n9160), .C2(n10084), .A(n8766), .B(n8765), .ZN(n13218)
         );
  NAND2_X1 U7243 ( .A1(n9333), .A2(n9334), .ZN(n9970) );
  XNOR2_X2 U7244 ( .A(n8600), .B(n14082), .ZN(n8602) );
  OAI21_X2 U7245 ( .B1(n13125), .B2(n9188), .A(n13093), .ZN(n13168) );
  AND2_X2 U7246 ( .A1(n7448), .A2(n7447), .ZN(n13125) );
  NOR2_X2 U7247 ( .A1(n9571), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9691) );
  INV_X1 U7249 ( .A(n9160), .ZN(n13366) );
  INV_X2 U7250 ( .A(n10065), .ZN(n6409) );
  INV_X2 U7251 ( .A(n10065), .ZN(n6410) );
  INV_X2 U7252 ( .A(n10065), .ZN(n10093) );
  AND2_X2 U7253 ( .A1(n7243), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U7254 ( .A1(n10053), .A2(n10052), .ZN(n10076) );
  XNOR2_X2 U7255 ( .A(n10068), .B(n10058), .ZN(n10067) );
  NAND2_X2 U7256 ( .A1(n7244), .A2(n10057), .ZN(n10068) );
  NOR3_X2 U7257 ( .A1(n12555), .A2(n12554), .A3(n12553), .ZN(n12582) );
  XOR2_X1 U7258 ( .A(n12140), .B(n12137), .Z(n6458) );
  NAND2_X1 U7259 ( .A1(n13718), .A2(n7836), .ZN(n13710) );
  NAND2_X1 U7260 ( .A1(n8704), .A2(n8703), .ZN(n13978) );
  NAND2_X1 U7261 ( .A1(n14368), .A2(n14800), .ZN(n14815) );
  INV_X2 U7262 ( .A(n13701), .ZN(n13741) );
  NAND2_X1 U7263 ( .A1(n9584), .A2(n9583), .ZN(n15022) );
  OR2_X2 U7264 ( .A1(n11824), .A2(n14447), .ZN(n11823) );
  CLKBUF_X1 U7265 ( .A(n8533), .Z(n12882) );
  XNOR2_X2 U7266 ( .A(n15419), .B(n12518), .ZN(n11454) );
  INV_X1 U7267 ( .A(n12519), .ZN(n11472) );
  INV_X1 U7268 ( .A(n14490), .ZN(n14306) );
  CLKBUF_X2 U7270 ( .A(n8050), .Z(n8347) );
  INV_X1 U7271 ( .A(n11343), .ZN(n14497) );
  CLKBUF_X2 U7272 ( .A(n14513), .Z(P1_U4016) );
  BUF_X2 U7273 ( .A(n8050), .Z(n8442) );
  INV_X2 U7274 ( .A(n15170), .ZN(n11342) );
  INV_X1 U7275 ( .A(n13449), .ZN(n10482) );
  NAND4_X2 U7276 ( .A1(n9354), .A2(n9356), .A3(n9355), .A4(n9357), .ZN(n14498)
         );
  NOR2_X1 U7277 ( .A1(n11840), .A2(n11574), .ZN(n9715) );
  INV_X2 U7278 ( .A(n8743), .ZN(n9042) );
  NAND2_X4 U7279 ( .A1(n7198), .A2(n7197), .ZN(n8714) );
  NAND2_X1 U7280 ( .A1(n8052), .A2(n7930), .ZN(n8074) );
  NAND3_X1 U7281 ( .A1(n9361), .A2(n7769), .A3(n9342), .ZN(n9370) );
  CLKBUF_X2 U7282 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n10501) );
  NOR2_X1 U7283 ( .A1(n12137), .A2(n8506), .ZN(n8524) );
  NAND2_X1 U7284 ( .A1(n13666), .A2(n13905), .ZN(n6773) );
  NAND2_X1 U7285 ( .A1(n13665), .A2(n13664), .ZN(n13666) );
  NAND2_X1 U7286 ( .A1(n13665), .A2(n7713), .ZN(n13650) );
  NAND2_X1 U7287 ( .A1(n8493), .A2(n8492), .ZN(n12756) );
  NAND2_X1 U7288 ( .A1(n7665), .A2(n6513), .ZN(n14651) );
  AOI211_X1 U7289 ( .C1(n13938), .C2(n13949), .A(n13660), .B(n13659), .ZN(
        n13661) );
  NAND2_X1 U7290 ( .A1(n12363), .A2(n12185), .ZN(n12439) );
  NAND2_X1 U7291 ( .A1(n7564), .A2(n7562), .ZN(n12363) );
  NAND2_X1 U7292 ( .A1(n14765), .A2(n7191), .ZN(n14749) );
  NAND2_X1 U7293 ( .A1(n7177), .A2(n7176), .ZN(n14675) );
  NAND2_X1 U7294 ( .A1(n6925), .A2(n7075), .ZN(n15144) );
  OAI21_X2 U7295 ( .B1(n14779), .B2(n14780), .A(n9603), .ZN(n14764) );
  NOR2_X1 U7296 ( .A1(n7600), .A2(n13415), .ZN(n7599) );
  OR2_X1 U7297 ( .A1(n13516), .A2(n13532), .ZN(n13536) );
  XNOR2_X1 U7298 ( .A(n12623), .B(n12630), .ZN(n12615) );
  CLKBUF_X1 U7299 ( .A(n14918), .Z(n6642) );
  NAND2_X1 U7300 ( .A1(n7741), .A2(n7740), .ZN(n12831) );
  NOR2_X1 U7301 ( .A1(n12240), .A2(n12239), .ZN(n12244) );
  NAND2_X1 U7302 ( .A1(n11979), .A2(n15308), .ZN(n7305) );
  NAND2_X1 U7303 ( .A1(n7025), .A2(n7587), .ZN(n12448) );
  NAND2_X1 U7304 ( .A1(n12744), .A2(n9903), .ZN(n8499) );
  CLKBUF_X1 U7305 ( .A(n7202), .Z(n7201) );
  OR2_X1 U7306 ( .A1(n7824), .A2(n7822), .ZN(n6457) );
  NAND2_X1 U7307 ( .A1(n12014), .A2(n7242), .ZN(n7025) );
  NAND2_X1 U7308 ( .A1(n7306), .A2(n11939), .ZN(n11979) );
  NAND2_X1 U7309 ( .A1(n11599), .A2(n15549), .ZN(n11939) );
  AOI21_X1 U7310 ( .B1(n6419), .B2(n7150), .A(n6434), .ZN(n7145) );
  INV_X1 U7311 ( .A(n14815), .ZN(n6411) );
  OAI21_X1 U7312 ( .B1(n13607), .B2(n7790), .A(n7788), .ZN(n13914) );
  AND2_X1 U7313 ( .A1(n9206), .A2(n9205), .ZN(n13667) );
  NAND2_X1 U7314 ( .A1(n11323), .A2(n9430), .ZN(n11705) );
  AND2_X1 U7315 ( .A1(n13622), .A2(n7812), .ZN(n7808) );
  AND2_X1 U7316 ( .A1(n6429), .A2(n7552), .ZN(n7551) );
  NAND2_X1 U7317 ( .A1(n9108), .A2(n9107), .ZN(n13988) );
  NAND2_X1 U7318 ( .A1(n9562), .A2(n9561), .ZN(n15034) );
  NAND2_X1 U7319 ( .A1(n8008), .A2(n8007), .ZN(n12788) );
  OAI21_X1 U7320 ( .B1(n7037), .B2(n11020), .A(n7033), .ZN(n11288) );
  AND2_X1 U7321 ( .A1(n8280), .A2(n8279), .ZN(n12473) );
  INV_X1 U7322 ( .A(n13912), .ZN(n14031) );
  AND2_X1 U7323 ( .A1(n10704), .A2(n10667), .ZN(n10672) );
  NAND2_X1 U7324 ( .A1(n9007), .A2(n9006), .ZN(n14013) );
  NAND2_X1 U7325 ( .A1(n6552), .A2(n7588), .ZN(n7587) );
  OR2_X1 U7326 ( .A1(n9052), .A2(n10819), .ZN(n9086) );
  OAI21_X2 U7327 ( .B1(n11199), .B2(n9748), .A(n9747), .ZN(n11296) );
  NAND2_X1 U7328 ( .A1(n9534), .A2(n9533), .ZN(n15046) );
  OR2_X1 U7329 ( .A1(n14303), .A2(n14489), .ZN(n14938) );
  NAND2_X1 U7330 ( .A1(n7062), .A2(n8934), .ZN(n14036) );
  NAND2_X1 U7331 ( .A1(n9472), .A2(n9471), .ZN(n14303) );
  INV_X2 U7332 ( .A(n13554), .ZN(n13938) );
  NAND2_X1 U7333 ( .A1(n7131), .A2(n15543), .ZN(n8329) );
  NAND3_X1 U7334 ( .A1(n7546), .A2(n7547), .A3(n7545), .ZN(n11793) );
  NAND2_X2 U7335 ( .A1(n13880), .A2(n10015), .ZN(n13931) );
  INV_X2 U7336 ( .A(n13880), .ZN(n13940) );
  NAND2_X1 U7337 ( .A1(n9460), .A2(n9459), .ZN(n15079) );
  NAND2_X1 U7338 ( .A1(n8876), .A2(n8875), .ZN(n14051) );
  NOR2_X1 U7339 ( .A1(n12012), .A2(n12516), .ZN(n12013) );
  OR2_X1 U7340 ( .A1(n9059), .A2(n13160), .ZN(n9095) );
  NAND2_X1 U7341 ( .A1(n8176), .A2(n8175), .ZN(n12469) );
  NAND2_X1 U7342 ( .A1(n9794), .A2(n15237), .ZN(n15215) );
  INV_X2 U7343 ( .A(n15220), .ZN(n6412) );
  NAND2_X1 U7344 ( .A1(n7223), .A2(n11005), .ZN(n8047) );
  NAND2_X1 U7345 ( .A1(n7160), .A2(n9432), .ZN(n14956) );
  XNOR2_X1 U7346 ( .A(n13235), .B(n13445), .ZN(n13401) );
  NAND2_X1 U7347 ( .A1(n7938), .A2(n7937), .ZN(n8253) );
  AND2_X1 U7348 ( .A1(n14277), .A2(n14278), .ZN(n14439) );
  NAND4_X2 U7349 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n12878)
         );
  AND3_X1 U7350 ( .A1(n8024), .A2(n8023), .A3(n6498), .ZN(n11005) );
  NOR2_X1 U7351 ( .A1(n8986), .A2(n11502), .ZN(n8985) );
  OR2_X2 U7352 ( .A1(n8211), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8237) );
  AOI22_X1 U7353 ( .A1(n7158), .A2(n7056), .B1(n8833), .B2(n8644), .ZN(n7054)
         );
  BUF_X4 U7354 ( .A(n11352), .Z(n12315) );
  AND4_X1 U7355 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n11866)
         );
  NAND2_X1 U7356 ( .A1(n7302), .A2(n10104), .ZN(n10176) );
  NAND4_X2 U7357 ( .A1(n9395), .A2(n9394), .A3(n9393), .A4(n9392), .ZN(n14495)
         );
  NAND2_X1 U7358 ( .A1(n8029), .A2(n7400), .ZN(n8063) );
  NAND2_X1 U7359 ( .A1(n8029), .A2(n10065), .ZN(n8062) );
  INV_X2 U7360 ( .A(n11341), .ZN(n10744) );
  NAND2_X2 U7361 ( .A1(n7796), .A2(n7794), .ZN(n13450) );
  BUF_X2 U7362 ( .A(n8051), .Z(n8441) );
  INV_X2 U7363 ( .A(n9585), .ZN(n9785) );
  AND2_X2 U7364 ( .A1(n7951), .A2(n13024), .ZN(n8091) );
  OAI211_X1 U7365 ( .C1(n9637), .C2(n10086), .A(n9386), .B(n9385), .ZN(n15222)
         );
  AND3_X2 U7366 ( .A1(n9365), .A2(n9364), .A3(n9363), .ZN(n14268) );
  AND3_X1 U7367 ( .A1(n8724), .A2(n7344), .A3(n8723), .ZN(n13198) );
  NAND4_X1 U7368 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(n13449)
         );
  INV_X1 U7369 ( .A(n15361), .ZN(n11266) );
  OR2_X1 U7370 ( .A1(n13197), .A2(n8712), .ZN(n10909) );
  NAND2_X1 U7371 ( .A1(n9343), .A2(n7397), .ZN(n14970) );
  INV_X2 U7372 ( .A(n9637), .ZN(n9845) );
  NOR2_X1 U7373 ( .A1(n7057), .A2(n7058), .ZN(n7056) );
  CLKBUF_X1 U7374 ( .A(n9347), .Z(n7116) );
  INV_X1 U7375 ( .A(n8710), .ZN(n8711) );
  INV_X1 U7376 ( .A(n8745), .ZN(n8960) );
  NAND2_X1 U7377 ( .A1(n7853), .A2(n7539), .ZN(n10017) );
  NAND2_X1 U7378 ( .A1(n9334), .A2(n9335), .ZN(n9539) );
  CLKBUF_X1 U7379 ( .A(n8745), .Z(n9223) );
  NAND2_X2 U7380 ( .A1(n9332), .A2(n9335), .ZN(n9376) );
  AND3_X1 U7381 ( .A1(n8656), .A2(n8951), .A3(n8907), .ZN(n8657) );
  OR2_X1 U7382 ( .A1(n13369), .A2(n10089), .ZN(n8741) );
  XNOR2_X1 U7383 ( .A(n8125), .B(n8139), .ZN(n11144) );
  NAND2_X1 U7384 ( .A1(n8662), .A2(n8929), .ZN(n6738) );
  INV_X2 U7385 ( .A(n7728), .ZN(n9289) );
  NAND2_X2 U7386 ( .A1(n15106), .A2(n9784), .ZN(n9347) );
  AND2_X1 U7387 ( .A1(n8648), .A2(n7275), .ZN(n7274) );
  INV_X1 U7388 ( .A(n9334), .ZN(n9332) );
  NAND2_X1 U7389 ( .A1(n7102), .A2(n7099), .ZN(n11840) );
  NAND2_X1 U7390 ( .A1(n8619), .A2(n8615), .ZN(n13195) );
  NAND2_X1 U7391 ( .A1(n9709), .A2(n9708), .ZN(n11531) );
  NAND2_X1 U7392 ( .A1(n9714), .A2(n9713), .ZN(n11574) );
  XNOR2_X1 U7393 ( .A(n9573), .B(P1_IR_REG_19__SCAN_IN), .ZN(n14246) );
  XNOR2_X1 U7394 ( .A(n7189), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9334) );
  OAI21_X1 U7395 ( .B1(n13018), .B2(P3_IR_REG_30__SCAN_IN), .A(n6528), .ZN(
        n7157) );
  NAND2_X1 U7396 ( .A1(n9340), .A2(n7683), .ZN(n15106) );
  OR2_X1 U7397 ( .A1(n8124), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U7398 ( .A1(n9700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7004) );
  MUX2_X1 U7399 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9339), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9340) );
  NAND2_X1 U7400 ( .A1(n9713), .A2(n7082), .ZN(n7102) );
  NOR2_X1 U7401 ( .A1(n7101), .A2(n7100), .ZN(n7099) );
  XNOR2_X1 U7402 ( .A(n10051), .B(n10049), .ZN(n10047) );
  NAND2_X1 U7403 ( .A1(n7118), .A2(n7121), .ZN(n14089) );
  INV_X1 U7404 ( .A(n13373), .ZN(n6414) );
  NAND2_X1 U7405 ( .A1(n6471), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7121) );
  NOR2_X1 U7406 ( .A1(n8555), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7297) );
  BUF_X1 U7407 ( .A(n7946), .Z(n7949) );
  OR2_X1 U7408 ( .A1(n9711), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U7409 ( .A1(n7105), .A2(n7104), .ZN(n8114) );
  INV_X1 U7410 ( .A(n10065), .ZN(n7400) );
  AND2_X1 U7411 ( .A1(n7982), .A2(n7589), .ZN(n8270) );
  AND2_X1 U7412 ( .A1(n8706), .A2(n8705), .ZN(n8997) );
  AND2_X1 U7413 ( .A1(n7343), .A2(n7342), .ZN(n8599) );
  XNOR2_X1 U7414 ( .A(n6836), .B(n7459), .ZN(n10727) );
  NOR2_X1 U7415 ( .A1(n9705), .A2(n9318), .ZN(n9329) );
  INV_X1 U7416 ( .A(n8185), .ZN(n7982) );
  INV_X1 U7417 ( .A(n9705), .ZN(n7715) );
  INV_X1 U7418 ( .A(n8092), .ZN(n7105) );
  AND2_X1 U7419 ( .A1(n7736), .A2(n7461), .ZN(n7217) );
  OR2_X1 U7420 ( .A1(n8080), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U7421 ( .A1(n10045), .A2(n10044), .ZN(n10055) );
  NAND2_X1 U7422 ( .A1(n7932), .A2(n7931), .ZN(n8092) );
  AND2_X1 U7423 ( .A1(n8695), .A2(n8592), .ZN(n7843) );
  NAND2_X1 U7424 ( .A1(n7255), .A2(n7927), .ZN(n7198) );
  INV_X1 U7425 ( .A(n8074), .ZN(n7932) );
  AND2_X1 U7426 ( .A1(n7923), .A2(n7920), .ZN(n7461) );
  NOR2_X1 U7427 ( .A1(n9316), .A2(n9336), .ZN(n7082) );
  AND3_X1 U7428 ( .A1(n8591), .A2(n8590), .A3(n9236), .ZN(n8695) );
  NOR2_X1 U7429 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7913) );
  NOR2_X1 U7430 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7915) );
  INV_X1 U7431 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8557) );
  INV_X1 U7432 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9361) );
  NOR2_X1 U7433 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7914) );
  INV_X1 U7434 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7104) );
  NOR2_X1 U7435 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8558) );
  INV_X1 U7436 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8556) );
  NOR2_X1 U7437 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7909) );
  NOR3_X1 U7438 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n8589) );
  INV_X4 U7439 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7440 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8081) );
  NOR2_X1 U7441 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n9693) );
  INV_X4 U7442 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7443 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9694) );
  NOR2_X1 U7444 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n9313) );
  NOR2_X1 U7445 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8594) );
  NOR2_X2 U7446 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8041) );
  INV_X1 U7447 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7979) );
  INV_X1 U7448 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8780) );
  INV_X1 U7449 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8812) );
  NOR2_X1 U7450 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8593) );
  INV_X1 U7451 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9409) );
  INV_X4 U7452 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7453 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9321) );
  INV_X1 U7454 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8014) );
  INV_X1 U7455 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7931) );
  INV_X1 U7456 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8778) );
  INV_X1 U7457 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7910) );
  NOR2_X1 U7458 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8595) );
  NOR3_X2 U7459 ( .A1(n8553), .A2(n8552), .A3(n7133), .ZN(n7132) );
  NOR2_X2 U7460 ( .A1(n13653), .A2(n13947), .ZN(n13601) );
  XNOR2_X2 U7461 ( .A(n8739), .B(n8738), .ZN(n13458) );
  INV_X2 U7462 ( .A(n6415), .ZN(n6416) );
  AOI21_X2 U7463 ( .B1(n13710), .B2(n13638), .A(n7042), .ZN(n13694) );
  OR2_X2 U7464 ( .A1(n12993), .A2(n12473), .ZN(n12813) );
  XNOR2_X2 U7465 ( .A(n14019), .B(n13620), .ZN(n13622) );
  NOR2_X2 U7466 ( .A1(n13705), .A2(n13962), .ZN(n13689) );
  NAND3_X2 U7467 ( .A1(n13768), .A2(n6431), .A3(n13708), .ZN(n13705) );
  AOI21_X2 U7468 ( .B1(n10744), .B2(n14499), .A(n10743), .ZN(n10855) );
  XNOR2_X1 U7469 ( .A(n8306), .B(n8305), .ZN(n12696) );
  OAI211_X1 U7470 ( .C1(n13369), .C2(n10083), .A(n8815), .B(n8814), .ZN(n8816)
         );
  OAI22_X2 U7471 ( .A1(n14109), .A2(n7009), .B1(n7010), .B2(n7008), .ZN(n12240) );
  NAND2_X2 U7472 ( .A1(n14187), .A2(n12104), .ZN(n14109) );
  NOR2_X2 U7473 ( .A1(n11265), .A2(n15361), .ZN(n11264) );
  OR2_X1 U7474 ( .A1(n10017), .A2(n13200), .ZN(n11265) );
  NAND2_X1 U7475 ( .A1(n8120), .A2(n11456), .ZN(n7294) );
  NAND2_X1 U7476 ( .A1(n6738), .A2(n8951), .ZN(n6737) );
  NAND2_X1 U7477 ( .A1(n13319), .A2(n6714), .ZN(n13322) );
  OAI21_X1 U7478 ( .B1(n13313), .B2(n7639), .A(n6715), .ZN(n6714) );
  NOR2_X1 U7479 ( .A1(n13318), .A2(n6716), .ZN(n6715) );
  INV_X1 U7480 ( .A(n12055), .ZN(n7951) );
  NAND2_X1 U7481 ( .A1(n9898), .A2(n9897), .ZN(n7761) );
  NAND2_X1 U7482 ( .A1(n7469), .A2(n7470), .ZN(n8498) );
  INV_X1 U7483 ( .A(n7471), .ZN(n7470) );
  OAI21_X1 U7484 ( .B1(n8494), .B2(n7472), .A(n8496), .ZN(n7471) );
  NOR2_X1 U7485 ( .A1(n9900), .A2(n7142), .ZN(n7141) );
  AOI21_X1 U7486 ( .B1(n7518), .B2(n7871), .A(n6545), .ZN(n7517) );
  OR2_X1 U7487 ( .A1(n9274), .A2(n15559), .ZN(n9288) );
  NAND2_X1 U7488 ( .A1(n13818), .A2(n13627), .ZN(n13793) );
  INV_X1 U7489 ( .A(n13618), .ZN(n7812) );
  OR2_X1 U7490 ( .A1(n7554), .A2(n13741), .ZN(n7836) );
  NAND2_X1 U7491 ( .A1(n7047), .A2(n7343), .ZN(n7046) );
  AND2_X1 U7492 ( .A1(n8610), .A2(n7043), .ZN(n7047) );
  AND2_X1 U7493 ( .A1(n8695), .A2(n7044), .ZN(n7043) );
  AND2_X1 U7494 ( .A1(n8592), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7044) );
  AND2_X1 U7495 ( .A1(n7458), .A2(n7456), .ZN(n7453) );
  INV_X1 U7496 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7456) );
  NOR3_X1 U7497 ( .A1(n14408), .A2(n14697), .A3(n14983), .ZN(n9974) );
  OR2_X1 U7498 ( .A1(n9644), .A2(n9629), .ZN(n9631) );
  OR2_X1 U7499 ( .A1(n9775), .A2(n6573), .ZN(n7182) );
  INV_X1 U7500 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9326) );
  INV_X1 U7501 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9325) );
  INV_X1 U7502 ( .A(n8441), .ZN(n8409) );
  NOR2_X1 U7503 ( .A1(n14136), .A2(n7685), .ZN(n7684) );
  INV_X1 U7504 ( .A(n12255), .ZN(n7685) );
  NOR2_X1 U7505 ( .A1(n14408), .A2(n7726), .ZN(n7725) );
  NAND2_X1 U7506 ( .A1(n14421), .A2(n7727), .ZN(n7726) );
  OAI21_X1 U7507 ( .B1(n14226), .B2(n14983), .A(n9780), .ZN(n14689) );
  NAND2_X1 U7508 ( .A1(n7112), .A2(SI_23_), .ZN(n9152) );
  AND2_X1 U7509 ( .A1(n11938), .A2(n7307), .ZN(n7306) );
  INV_X1 U7510 ( .A(n11946), .ZN(n7307) );
  NAND2_X1 U7511 ( .A1(n11947), .A2(n11946), .ZN(n11980) );
  NAND2_X1 U7512 ( .A1(n8136), .A2(n11443), .ZN(n7293) );
  AND2_X1 U7513 ( .A1(n8322), .A2(n8321), .ZN(n6674) );
  AOI21_X1 U7514 ( .B1(n6432), .B2(n6721), .A(n6423), .ZN(n6718) );
  AND2_X1 U7515 ( .A1(n13318), .A2(n7636), .ZN(n7635) );
  NAND2_X1 U7516 ( .A1(n7639), .A2(n7638), .ZN(n7636) );
  AND2_X1 U7517 ( .A1(n6737), .A2(n8663), .ZN(n8664) );
  INV_X1 U7518 ( .A(n11728), .ZN(n7374) );
  AND2_X1 U7519 ( .A1(n13341), .A2(n13327), .ZN(n13332) );
  INV_X1 U7520 ( .A(n14409), .ZN(n7281) );
  INV_X1 U7521 ( .A(n9757), .ZN(n7781) );
  OR2_X1 U7522 ( .A1(n7782), .A2(n7781), .ZN(n7780) );
  NOR2_X1 U7523 ( .A1(n9191), .A2(n6752), .ZN(n6751) );
  INV_X1 U7524 ( .A(n9174), .ZN(n6752) );
  INV_X1 U7525 ( .A(n12205), .ZN(n7585) );
  OAI21_X1 U7526 ( .B1(n12592), .B2(P3_REG2_REG_13__SCAN_IN), .A(n12591), .ZN(
        n6828) );
  INV_X1 U7527 ( .A(n7743), .ZN(n7742) );
  OAI21_X1 U7528 ( .B1(n12857), .B2(n7744), .A(n9889), .ZN(n7743) );
  OR2_X1 U7529 ( .A1(n12520), .A2(n9872), .ZN(n8457) );
  NAND2_X1 U7530 ( .A1(n7496), .A2(n8412), .ZN(n8525) );
  OR2_X1 U7531 ( .A1(n12715), .A2(n12511), .ZN(n8504) );
  NOR2_X1 U7532 ( .A1(n7766), .A2(n12725), .ZN(n7765) );
  OR2_X1 U7533 ( .A1(n12980), .A2(n12798), .ZN(n9895) );
  OR2_X1 U7534 ( .A1(n12974), .A2(n12375), .ZN(n8488) );
  NAND2_X1 U7535 ( .A1(n7153), .A2(n6509), .ZN(n12031) );
  AND2_X1 U7536 ( .A1(n6430), .A2(n8246), .ZN(n7589) );
  AND2_X1 U7537 ( .A1(n7910), .A2(n7591), .ZN(n7590) );
  NAND2_X1 U7538 ( .A1(n7602), .A2(n6493), .ZN(n7093) );
  NOR2_X1 U7539 ( .A1(n13711), .A2(n13719), .ZN(n7602) );
  AOI21_X1 U7540 ( .B1(n13322), .B2(n13321), .A(n13320), .ZN(n13324) );
  INV_X1 U7541 ( .A(n14089), .ZN(n8603) );
  INV_X1 U7542 ( .A(n9221), .ZN(n9219) );
  INV_X1 U7543 ( .A(n7837), .ZN(n7825) );
  INV_X1 U7544 ( .A(n13572), .ZN(n7316) );
  NAND2_X1 U7545 ( .A1(n14025), .A2(n13568), .ZN(n13570) );
  NAND2_X1 U7546 ( .A1(n11413), .A2(n13235), .ZN(n7340) );
  AND2_X1 U7547 ( .A1(n13682), .A2(n13967), .ZN(n7042) );
  NAND2_X1 U7548 ( .A1(n13428), .A2(n13195), .ZN(n13423) );
  NOR2_X1 U7549 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8587) );
  NOR2_X1 U7550 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8586) );
  INV_X1 U7551 ( .A(n9768), .ZN(n6963) );
  OR2_X1 U7552 ( .A1(n15028), .A2(n14827), .ZN(n14368) );
  AND2_X1 U7553 ( .A1(n9568), .A2(n7172), .ZN(n7171) );
  OR2_X1 U7554 ( .A1(n7174), .A2(n7173), .ZN(n7172) );
  AND2_X1 U7555 ( .A1(n9767), .A2(n9765), .ZN(n7772) );
  INV_X1 U7556 ( .A(n14895), .ZN(n7681) );
  NAND2_X1 U7557 ( .A1(n14920), .A2(n14919), .ZN(n14918) );
  INV_X1 U7558 ( .A(n7723), .ZN(n7722) );
  NAND2_X1 U7559 ( .A1(n11357), .A2(n11377), .ZN(n7723) );
  NAND2_X1 U7560 ( .A1(n9741), .A2(n14268), .ZN(n14267) );
  AND2_X1 U7561 ( .A1(n7183), .A2(n7178), .ZN(n14701) );
  OR2_X1 U7562 ( .A1(n9826), .A2(n9825), .ZN(n9830) );
  NOR2_X1 U7563 ( .A1(n6614), .A2(n7284), .ZN(n7283) );
  INV_X1 U7564 ( .A(n8691), .ZN(n7284) );
  NAND2_X1 U7565 ( .A1(n6742), .A2(n8681), .ZN(n9072) );
  OAI21_X1 U7566 ( .B1(n9002), .B2(n7613), .A(n6740), .ZN(n6742) );
  NOR2_X1 U7567 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7699) );
  AND2_X1 U7568 ( .A1(n8663), .A2(n8655), .ZN(n8951) );
  OAI21_X1 U7569 ( .B1(n7158), .B2(n8833), .A(n7055), .ZN(n8852) );
  NAND2_X1 U7570 ( .A1(n11597), .A2(n11596), .ZN(n11941) );
  OR2_X1 U7571 ( .A1(n11594), .A2(n11593), .ZN(n11597) );
  AND2_X1 U7572 ( .A1(n12336), .A2(n7584), .ZN(n7583) );
  OR2_X1 U7573 ( .A1(n12484), .A2(n7585), .ZN(n7584) );
  AND2_X1 U7574 ( .A1(n7221), .A2(n9919), .ZN(n7220) );
  OR2_X1 U7575 ( .A1(n10586), .A2(n10607), .ZN(n7433) );
  NAND2_X1 U7576 ( .A1(n10586), .A2(n10607), .ZN(n10729) );
  NAND2_X1 U7577 ( .A1(n7364), .A2(n10634), .ZN(n7363) );
  INV_X1 U7578 ( .A(n10646), .ZN(n7364) );
  NAND2_X1 U7579 ( .A1(n12639), .A2(n6822), .ZN(n12610) );
  AND2_X1 U7580 ( .A1(n12608), .A2(n12630), .ZN(n6825) );
  NAND2_X1 U7581 ( .A1(n7423), .A2(n6996), .ZN(n7422) );
  NAND2_X1 U7582 ( .A1(n12649), .A2(n12666), .ZN(n12672) );
  OR2_X1 U7583 ( .A1(n8390), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12065) );
  NAND2_X1 U7584 ( .A1(n6708), .A2(n6524), .ZN(n7142) );
  NAND2_X1 U7585 ( .A1(n7760), .A2(n7758), .ZN(n6708) );
  INV_X1 U7586 ( .A(n9897), .ZN(n7758) );
  INV_X1 U7587 ( .A(n12831), .ZN(n7147) );
  NOR2_X1 U7588 ( .A1(n7478), .A2(n7476), .ZN(n7475) );
  INV_X1 U7589 ( .A(n8470), .ZN(n7476) );
  NOR2_X1 U7590 ( .A1(n6468), .A2(n7480), .ZN(n7479) );
  INV_X1 U7591 ( .A(n8463), .ZN(n7480) );
  AND2_X1 U7593 ( .A1(n9951), .A2(n11134), .ZN(n12889) );
  NAND2_X1 U7594 ( .A1(n8498), .A2(n6435), .ZN(n7485) );
  INV_X1 U7595 ( .A(n12144), .ZN(n12880) );
  NAND2_X1 U7596 ( .A1(n9956), .A2(n9909), .ZN(n12883) );
  NOR2_X1 U7597 ( .A1(n10508), .A2(n10571), .ZN(n10807) );
  OR2_X1 U7598 ( .A1(n9936), .A2(n10806), .ZN(n12048) );
  OAI21_X1 U7599 ( .B1(n9920), .B2(P3_D_REG_1__SCAN_IN), .A(n9921), .ZN(n10690) );
  NAND2_X1 U7600 ( .A1(n13018), .A2(n7229), .ZN(n7227) );
  NOR2_X1 U7601 ( .A1(n13017), .A2(n7230), .ZN(n7229) );
  OAI211_X1 U7602 ( .C1(n7949), .C2(n7947), .A(n7226), .B(n7228), .ZN(n7952)
         );
  NAND2_X1 U7603 ( .A1(n13017), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U7604 ( .A1(n7949), .A2(n6511), .ZN(n7226) );
  NAND2_X1 U7605 ( .A1(n7901), .A2(n7900), .ZN(n7523) );
  OAI21_X1 U7606 ( .B1(n8449), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8450) );
  AOI21_X1 U7607 ( .B1(n8281), .B2(n7502), .A(n7501), .ZN(n7500) );
  INV_X1 U7608 ( .A(n7890), .ZN(n7501) );
  INV_X1 U7609 ( .A(n7887), .ZN(n7502) );
  AOI21_X1 U7610 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6723) );
  INV_X1 U7611 ( .A(n7884), .ZN(n6724) );
  INV_X1 U7612 ( .A(n7535), .ZN(n6725) );
  OR2_X1 U7613 ( .A1(n8184), .A2(n8183), .ZN(n7877) );
  AOI21_X1 U7614 ( .B1(n6547), .B2(n7514), .A(n6444), .ZN(n7511) );
  NAND2_X1 U7615 ( .A1(n6681), .A2(n6683), .ZN(n6680) );
  INV_X1 U7616 ( .A(n6683), .ZN(n6682) );
  NOR2_X1 U7617 ( .A1(n8015), .A2(n6684), .ZN(n6683) );
  XNOR2_X1 U7618 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n7857) );
  NAND2_X1 U7619 ( .A1(n9163), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U7620 ( .A1(n13168), .A2(n9208), .ZN(n13167) );
  INV_X1 U7621 ( .A(n9289), .ZN(n13365) );
  INV_X1 U7622 ( .A(n9223), .ZN(n9294) );
  NAND2_X1 U7623 ( .A1(n8602), .A2(n8603), .ZN(n8784) );
  AND2_X1 U7624 ( .A1(n8601), .A2(n14089), .ZN(n8743) );
  NAND2_X1 U7625 ( .A1(n8601), .A2(n8603), .ZN(n8745) );
  OAI21_X1 U7626 ( .B1(n10661), .B2(n10660), .A(n6790), .ZN(n10707) );
  OR2_X1 U7627 ( .A1(n10663), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6790) );
  OR2_X1 U7628 ( .A1(n10707), .A2(n10708), .ZN(n6789) );
  NOR2_X1 U7629 ( .A1(n11499), .A2(n6793), .ZN(n15309) );
  AND2_X1 U7630 ( .A1(n11504), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U7631 ( .A1(n7051), .A2(n7050), .ZN(n13720) );
  NAND2_X1 U7632 ( .A1(n13632), .A2(n7053), .ZN(n7050) );
  NAND2_X1 U7633 ( .A1(n13765), .A2(n13580), .ZN(n7708) );
  NAND2_X1 U7634 ( .A1(n13776), .A2(n13579), .ZN(n13765) );
  INV_X1 U7635 ( .A(n6759), .ZN(n6758) );
  OAI21_X1 U7636 ( .B1(n7806), .B2(n6761), .A(n13835), .ZN(n6759) );
  AOI21_X1 U7637 ( .B1(n13563), .B2(n6754), .A(n6522), .ZN(n6753) );
  INV_X1 U7638 ( .A(n11746), .ZN(n6754) );
  NOR2_X1 U7639 ( .A1(n6414), .A2(n13421), .ZN(n10905) );
  INV_X1 U7640 ( .A(n6777), .ZN(n6776) );
  OAI22_X1 U7641 ( .A1(n13668), .A2(n13871), .B1(n13869), .B2(n13667), .ZN(
        n6777) );
  INV_X1 U7642 ( .A(n13604), .ZN(n13947) );
  OR2_X1 U7643 ( .A1(n15384), .A2(n9226), .ZN(n6774) );
  AND2_X2 U7644 ( .A1(n13423), .A2(n10905), .ZN(n15377) );
  AND3_X1 U7645 ( .A1(n8737), .A2(n8593), .A3(n8738), .ZN(n6764) );
  INV_X1 U7646 ( .A(n14085), .ZN(n7120) );
  AND2_X2 U7647 ( .A1(n8594), .A2(n8595), .ZN(n8596) );
  NAND2_X1 U7648 ( .A1(n9606), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9642) );
  INV_X1 U7649 ( .A(n9607), .ZN(n9606) );
  OR2_X1 U7650 ( .A1(n9642), .A2(n9641), .ZN(n9644) );
  AOI21_X1 U7651 ( .B1(n7015), .B2(n7017), .A(n7014), .ZN(n7013) );
  INV_X1 U7652 ( .A(n14195), .ZN(n7014) );
  NOR2_X1 U7653 ( .A1(n14152), .A2(n7690), .ZN(n7022) );
  AND2_X1 U7654 ( .A1(n9626), .A2(n9625), .ZN(n14225) );
  OR2_X1 U7655 ( .A1(n14722), .A2(n9785), .ZN(n9626) );
  XNOR2_X1 U7656 ( .A(n14626), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14636) );
  OR2_X1 U7657 ( .A1(n14408), .A2(n14478), .ZN(n9687) );
  AND2_X1 U7658 ( .A1(n9792), .A2(n9791), .ZN(n14420) );
  OR3_X1 U7659 ( .A1(n14663), .A2(n9785), .A3(n14662), .ZN(n9792) );
  AND2_X1 U7660 ( .A1(n6887), .A2(n9677), .ZN(n14226) );
  OR2_X1 U7661 ( .A1(n14684), .A2(n9785), .ZN(n6887) );
  NOR2_X1 U7662 ( .A1(n14675), .A2(n14689), .ZN(n14676) );
  AND2_X1 U7663 ( .A1(n9663), .A2(n9662), .ZN(n14679) );
  NAND2_X1 U7664 ( .A1(n9655), .A2(n9654), .ZN(n14395) );
  XNOR2_X1 U7665 ( .A(n9615), .B(n14784), .ZN(n14768) );
  XNOR2_X1 U7666 ( .A(n15017), .B(n14484), .ZN(n14780) );
  NAND2_X1 U7667 ( .A1(n15028), .A2(n14827), .ZN(n14800) );
  AND4_X1 U7668 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n14861)
         );
  OR2_X1 U7669 ( .A1(n15053), .A2(n14862), .ZN(n14342) );
  NAND2_X1 U7670 ( .A1(n14876), .A2(n14877), .ZN(n9764) );
  OR2_X1 U7671 ( .A1(n14432), .A2(n14511), .ZN(n14933) );
  AND2_X1 U7672 ( .A1(n9836), .A2(n9835), .ZN(n14981) );
  AND2_X1 U7673 ( .A1(n14750), .A2(n9616), .ZN(n7191) );
  NAND2_X1 U7674 ( .A1(n9783), .A2(n9782), .ZN(n15251) );
  NAND2_X1 U7675 ( .A1(n12313), .A2(n9737), .ZN(n15247) );
  OR2_X1 U7676 ( .A1(n14248), .A2(n9803), .ZN(n9737) );
  INV_X1 U7677 ( .A(n15247), .ZN(n15263) );
  INV_X1 U7678 ( .A(n15255), .ZN(n15259) );
  NAND2_X1 U7679 ( .A1(n7190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7189) );
  AND2_X1 U7680 ( .A1(n9329), .A2(n7787), .ZN(n7083) );
  NAND2_X1 U7681 ( .A1(n11160), .A2(n11159), .ZN(n7071) );
  NOR2_X1 U7682 ( .A1(n15140), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6926) );
  NAND2_X1 U7683 ( .A1(n15140), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U7684 ( .A1(n15144), .A2(n6921), .ZN(n15151) );
  INV_X1 U7685 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6922) );
  AND2_X1 U7686 ( .A1(n7998), .A2(n7997), .ZN(n12357) );
  NAND2_X1 U7687 ( .A1(n7990), .A2(n7989), .ZN(n12909) );
  INV_X1 U7688 ( .A(n12432), .ZN(n12752) );
  INV_X1 U7689 ( .A(n12706), .ZN(n7109) );
  NAND2_X1 U7690 ( .A1(n7110), .A2(n12707), .ZN(n6908) );
  NAND2_X1 U7691 ( .A1(n6670), .A2(n6669), .ZN(n13600) );
  INV_X1 U7692 ( .A(n6770), .ZN(n6769) );
  NAND2_X1 U7693 ( .A1(n6774), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U7694 ( .A1(n12160), .A2(n9845), .ZN(n6886) );
  OR2_X1 U7695 ( .A1(n11335), .A2(n9637), .ZN(n9640) );
  OR2_X1 U7696 ( .A1(n14432), .A2(n9784), .ZN(n14935) );
  NAND2_X1 U7697 ( .A1(n9636), .A2(n9635), .ZN(n14712) );
  AOI22_X1 U7698 ( .A1(n14087), .A2(n9845), .B1(n9844), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U7699 ( .A1(n6947), .A2(n7249), .ZN(n15122) );
  OR2_X1 U7700 ( .A1(n15120), .A2(n7252), .ZN(n7249) );
  NOR2_X1 U7701 ( .A1(n15120), .A2(n7251), .ZN(n7250) );
  AND2_X2 U7702 ( .A1(n7304), .A2(n7303), .ZN(n15140) );
  NOR2_X1 U7703 ( .A1(n11007), .A2(n8035), .ZN(n6655) );
  NAND2_X1 U7704 ( .A1(n14259), .A2(n14970), .ZN(n14263) );
  INV_X1 U7705 ( .A(n7291), .ZN(n7290) );
  INV_X1 U7706 ( .A(n13231), .ZN(n6687) );
  NOR2_X1 U7707 ( .A1(n13234), .A2(n13231), .ZN(n6688) );
  OAI22_X1 U7708 ( .A1(n13228), .A2(n7651), .B1(n13229), .B2(n7650), .ZN(
        n13232) );
  NOR2_X1 U7709 ( .A1(n13239), .A2(n13236), .ZN(n7644) );
  NAND2_X1 U7710 ( .A1(n13239), .A2(n13236), .ZN(n7643) );
  NOR2_X1 U7711 ( .A1(n14284), .A2(n14281), .ZN(n7385) );
  NAND2_X1 U7712 ( .A1(n14284), .A2(n14281), .ZN(n7384) );
  INV_X1 U7713 ( .A(n13255), .ZN(n7629) );
  NAND2_X1 U7714 ( .A1(n7632), .A2(n7631), .ZN(n7630) );
  OAI21_X1 U7715 ( .B1(n6929), .B2(n6927), .A(n7380), .ZN(n14299) );
  OR2_X1 U7716 ( .A1(n14294), .A2(n7381), .ZN(n7380) );
  OAI21_X1 U7717 ( .B1(n14291), .B2(n14292), .A(n6445), .ZN(n6929) );
  AOI21_X1 U7718 ( .B1(n14291), .B2(n14292), .A(n6928), .ZN(n6927) );
  NAND2_X1 U7719 ( .A1(n14368), .A2(n14427), .ZN(n7261) );
  NAND2_X1 U7720 ( .A1(n14800), .A2(n14414), .ZN(n7260) );
  NOR2_X1 U7721 ( .A1(n13297), .A2(n7649), .ZN(n7648) );
  NOR2_X1 U7722 ( .A1(n6647), .A2(n6646), .ZN(n6645) );
  INV_X1 U7723 ( .A(n12787), .ZN(n6646) );
  NAND2_X1 U7724 ( .A1(n6939), .A2(n7390), .ZN(n6937) );
  INV_X1 U7725 ( .A(n6936), .ZN(n6935) );
  OAI21_X1 U7726 ( .B1(n6938), .B2(n7390), .A(n14384), .ZN(n6936) );
  NOR2_X1 U7727 ( .A1(n6808), .A2(n11692), .ZN(n6807) );
  OAI21_X1 U7728 ( .B1(n14391), .B2(n7395), .A(n7084), .ZN(n14398) );
  OR2_X1 U7729 ( .A1(n14393), .A2(n7396), .ZN(n7084) );
  OAI21_X1 U7730 ( .B1(n14390), .B2(n14389), .A(n6537), .ZN(n7395) );
  INV_X1 U7731 ( .A(n13521), .ZN(n6802) );
  INV_X1 U7732 ( .A(n6807), .ZN(n6803) );
  OAI21_X1 U7733 ( .B1(n7122), .B2(n6799), .A(n6797), .ZN(n6801) );
  OR2_X1 U7734 ( .A1(n6454), .A2(n6798), .ZN(n6797) );
  OR2_X1 U7735 ( .A1(n6454), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6799) );
  INV_X1 U7736 ( .A(n11690), .ZN(n6798) );
  AND2_X1 U7737 ( .A1(n14249), .A2(n14248), .ZN(n14411) );
  XNOR2_X1 U7738 ( .A(n14246), .B(n14245), .ZN(n14415) );
  INV_X1 U7739 ( .A(n6841), .ZN(n6840) );
  OAI21_X1 U7740 ( .B1(n11933), .B2(n6842), .A(n14613), .ZN(n6841) );
  INV_X1 U7741 ( .A(n6624), .ZN(n6842) );
  NAND2_X1 U7742 ( .A1(n8851), .A2(n8647), .ZN(n7275) );
  OAI21_X1 U7743 ( .B1(n6409), .B2(n8621), .A(n8620), .ZN(n8643) );
  NAND2_X1 U7744 ( .A1(n10093), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8620) );
  INV_X1 U7745 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U7746 ( .A1(n7561), .A2(n7558), .ZN(n7557) );
  INV_X1 U7747 ( .A(n11470), .ZN(n7558) );
  INV_X1 U7748 ( .A(n11679), .ZN(n7561) );
  INV_X1 U7749 ( .A(n11677), .ZN(n7560) );
  NOR2_X1 U7750 ( .A1(n12372), .A2(n7575), .ZN(n7574) );
  INV_X1 U7751 ( .A(n12188), .ZN(n7575) );
  AND2_X1 U7752 ( .A1(n11284), .A2(n11289), .ZN(n7240) );
  AND2_X1 U7753 ( .A1(n10649), .A2(n10615), .ZN(n10616) );
  OR2_X1 U7754 ( .A1(n10614), .A2(n10625), .ZN(n10615) );
  NOR2_X1 U7755 ( .A1(n10650), .A2(n6832), .ZN(n6831) );
  OAI21_X1 U7756 ( .B1(n10649), .B2(n10650), .A(n7429), .ZN(n7428) );
  NAND2_X1 U7757 ( .A1(n10655), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7429) );
  OAI21_X1 U7758 ( .B1(n10651), .B2(n7426), .A(n7425), .ZN(n10881) );
  NAND2_X1 U7759 ( .A1(n7430), .A2(n10871), .ZN(n7426) );
  NAND2_X1 U7760 ( .A1(n7428), .A2(n10871), .ZN(n7425) );
  OR2_X1 U7761 ( .A1(n11721), .A2(n6821), .ZN(n6820) );
  AND2_X1 U7762 ( .A1(n6403), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6821) );
  INV_X1 U7763 ( .A(n6820), .ZN(n11723) );
  NAND2_X1 U7764 ( .A1(n7373), .A2(n7374), .ZN(n7370) );
  OR2_X1 U7765 ( .A1(n11396), .A2(n7371), .ZN(n7368) );
  NAND2_X1 U7766 ( .A1(n7374), .A2(n7375), .ZN(n7371) );
  NAND2_X1 U7767 ( .A1(n12560), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7203) );
  OR2_X1 U7768 ( .A1(n12657), .A2(n12606), .ZN(n6918) );
  NAND2_X1 U7769 ( .A1(n6632), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U7770 ( .A1(n12666), .A2(n12627), .ZN(n6985) );
  OR2_X1 U7771 ( .A1(n6991), .A2(n12677), .ZN(n6987) );
  INV_X1 U7772 ( .A(n12627), .ZN(n6993) );
  NAND2_X1 U7773 ( .A1(n7106), .A2(n12779), .ZN(n8492) );
  INV_X1 U7774 ( .A(n12968), .ZN(n7106) );
  NOR2_X1 U7775 ( .A1(n8253), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8252) );
  NOR2_X2 U7776 ( .A1(n8237), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7938) );
  INV_X1 U7777 ( .A(n8456), .ZN(n7465) );
  NAND2_X1 U7778 ( .A1(n8104), .A2(n8457), .ZN(n9871) );
  NAND2_X1 U7779 ( .A1(n11023), .A2(n10998), .ZN(n8455) );
  INV_X1 U7780 ( .A(n9902), .ZN(n7763) );
  OR2_X1 U7781 ( .A1(n12986), .A2(n8336), .ZN(n8486) );
  OR2_X1 U7782 ( .A1(n12868), .A2(n12513), .ZN(n8471) );
  OR2_X1 U7783 ( .A1(n6459), .A2(n7749), .ZN(n7748) );
  AND2_X1 U7784 ( .A1(n6448), .A2(n6588), .ZN(n7136) );
  INV_X1 U7785 ( .A(n11442), .ZN(n7138) );
  INV_X1 U7786 ( .A(n9878), .ZN(n7137) );
  NOR2_X1 U7787 ( .A1(n6459), .A2(n7752), .ZN(n7751) );
  INV_X1 U7788 ( .A(n9879), .ZN(n7752) );
  AOI21_X1 U7789 ( .B1(n11565), .B2(n9879), .A(n7754), .ZN(n7753) );
  NOR2_X1 U7790 ( .A1(n6882), .A2(n9877), .ZN(n6878) );
  INV_X1 U7791 ( .A(n6883), .ZN(n6882) );
  NOR2_X1 U7792 ( .A1(n7460), .A2(n6884), .ZN(n6883) );
  INV_X1 U7793 ( .A(n8464), .ZN(n6884) );
  INV_X1 U7794 ( .A(n8465), .ZN(n7460) );
  INV_X1 U7795 ( .A(n8466), .ZN(n6880) );
  NAND2_X1 U7796 ( .A1(n11445), .A2(n9878), .ZN(n11566) );
  NAND2_X1 U7797 ( .A1(n10931), .A2(n10930), .ZN(n10929) );
  NAND2_X1 U7798 ( .A1(n9918), .A2(n6436), .ZN(n7222) );
  INV_X1 U7799 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U7800 ( .A1(n7525), .A2(n7522), .ZN(n7521) );
  INV_X1 U7801 ( .A(n6623), .ZN(n7522) );
  INV_X1 U7802 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8559) );
  AOI21_X1 U7803 ( .B1(n7500), .B2(n7503), .A(n7498), .ZN(n7497) );
  INV_X1 U7804 ( .A(n8265), .ZN(n7498) );
  NOR2_X1 U7805 ( .A1(n8098), .A2(n7509), .ZN(n7508) );
  INV_X1 U7806 ( .A(n7866), .ZN(n7509) );
  INV_X1 U7807 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U7808 ( .A1(n10060), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7864) );
  INV_X1 U7809 ( .A(n7435), .ZN(n7434) );
  OAI21_X1 U7810 ( .B1(n6469), .B2(n7436), .A(n9018), .ZN(n7435) );
  INV_X1 U7811 ( .A(n8984), .ZN(n7436) );
  AND2_X1 U7812 ( .A1(n8985), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9008) );
  OR4_X1 U7813 ( .A1(n13410), .A2(n13835), .A3(n13859), .A4(n13622), .ZN(
        n13411) );
  OAI211_X1 U7814 ( .C1(n13360), .C2(n13359), .A(n13358), .B(n13357), .ZN(
        n13361) );
  AND2_X1 U7815 ( .A1(n13389), .A2(n13383), .ZN(n7655) );
  INV_X1 U7816 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U7817 ( .A1(n13674), .A2(n6463), .ZN(n7800) );
  NAND2_X1 U7818 ( .A1(n9199), .A2(n9198), .ZN(n9221) );
  AOI21_X1 U7819 ( .B1(n7326), .B2(n7328), .A(n7323), .ZN(n7322) );
  INV_X1 U7820 ( .A(n13588), .ZN(n7323) );
  AND2_X1 U7821 ( .A1(n7053), .A2(n7815), .ZN(n7052) );
  NOR2_X1 U7822 ( .A1(n9095), .A2(n13075), .ZN(n6653) );
  OAI21_X1 U7823 ( .B1(n13866), .B2(n7320), .A(n7319), .ZN(n7318) );
  INV_X1 U7824 ( .A(n13859), .ZN(n7319) );
  INV_X1 U7825 ( .A(n14013), .ZN(n7553) );
  OR2_X1 U7826 ( .A1(n13373), .A2(n11129), .ZN(n10195) );
  AND2_X1 U7827 ( .A1(n13888), .A2(n14025), .ZN(n13872) );
  NOR2_X1 U7828 ( .A1(n14036), .A2(n14041), .ZN(n7543) );
  INV_X1 U7829 ( .A(n10905), .ZN(n9302) );
  NAND2_X1 U7830 ( .A1(n10004), .A2(n9999), .ZN(n10481) );
  NAND2_X1 U7831 ( .A1(n10905), .A2(n13195), .ZN(n8772) );
  OR2_X1 U7832 ( .A1(n13962), .A2(n13667), .ZN(n13392) );
  INV_X1 U7833 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9231) );
  AND2_X1 U7834 ( .A1(n8696), .A2(n8611), .ZN(n9232) );
  AND2_X1 U7835 ( .A1(n8763), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6870) );
  AND2_X1 U7836 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6871), .ZN(n6868) );
  INV_X1 U7837 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U7838 ( .A1(n7006), .A2(n7005), .ZN(n10856) );
  OR2_X1 U7839 ( .A1(n6405), .A2(n10249), .ZN(n9367) );
  OR2_X1 U7840 ( .A1(n9376), .A2(n10262), .ZN(n7195) );
  NAND2_X1 U7841 ( .A1(n9966), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U7842 ( .A1(n11616), .A2(n6843), .ZN(n11928) );
  OR2_X1 U7843 ( .A1(n11617), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U7844 ( .A1(n9780), .A2(n14689), .ZN(n7785) );
  NOR2_X1 U7845 ( .A1(n9772), .A2(n6573), .ZN(n7179) );
  INV_X1 U7846 ( .A(n14702), .ZN(n7181) );
  NOR2_X1 U7847 ( .A1(n14877), .A2(n7678), .ZN(n7677) );
  INV_X1 U7848 ( .A(n9519), .ZN(n7678) );
  NOR2_X1 U7849 ( .A1(n14303), .A2(n15079), .ZN(n7733) );
  OR2_X1 U7850 ( .A1(n7657), .A2(n7855), .ZN(n7162) );
  AND2_X1 U7851 ( .A1(n9478), .A2(n7658), .ZN(n7657) );
  AND2_X1 U7852 ( .A1(n11863), .A2(n9756), .ZN(n7782) );
  INV_X1 U7853 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9422) );
  INV_X1 U7854 ( .A(n11317), .ZN(n6973) );
  NAND2_X1 U7855 ( .A1(n9416), .A2(n14440), .ZN(n11301) );
  AND2_X1 U7856 ( .A1(n6748), .A2(n6451), .ZN(n6743) );
  XNOR2_X1 U7857 ( .A(n9823), .B(n9818), .ZN(n9267) );
  AND2_X1 U7858 ( .A1(n9156), .A2(n6617), .ZN(n7108) );
  NOR2_X1 U7859 ( .A1(n9696), .A2(n9702), .ZN(n7081) );
  NAND2_X1 U7860 ( .A1(n8672), .A2(n10546), .ZN(n8675) );
  INV_X1 U7861 ( .A(n8671), .ZN(n7606) );
  INV_X1 U7862 ( .A(n8927), .ZN(n8659) );
  INV_X1 U7863 ( .A(n8796), .ZN(n7593) );
  NAND2_X1 U7864 ( .A1(n7926), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7197) );
  INV_X1 U7865 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7927) );
  NAND3_X1 U7866 ( .A1(n6730), .A2(n6729), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7255) );
  INV_X1 U7867 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6729) );
  NAND2_X1 U7868 ( .A1(n10108), .A2(n10107), .ZN(n10168) );
  XNOR2_X1 U7869 ( .A(n10168), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n10167) );
  AOI21_X1 U7870 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n10720) );
  AOI21_X1 U7871 ( .B1(n7567), .B2(n7566), .A(n6476), .ZN(n7565) );
  INV_X1 U7872 ( .A(n12182), .ZN(n7566) );
  NAND2_X1 U7873 ( .A1(n7028), .A2(n7567), .ZN(n7564) );
  AOI21_X1 U7874 ( .B1(n7583), .B2(n7585), .A(n6551), .ZN(n7581) );
  NAND2_X1 U7875 ( .A1(n11182), .A2(n8017), .ZN(n7039) );
  INV_X1 U7876 ( .A(n12168), .ZN(n7588) );
  OAI211_X1 U7877 ( .C1(n10590), .C2(n10431), .A(n8045), .B(n8044), .ZN(n12888) );
  INV_X1 U7878 ( .A(n12878), .ZN(n11023) );
  OR2_X1 U7879 ( .A1(n11285), .A2(n7240), .ZN(n7035) );
  NAND2_X1 U7880 ( .A1(n7039), .A2(n7038), .ZN(n7036) );
  OR2_X1 U7881 ( .A1(n8551), .A2(n8550), .ZN(n7133) );
  AND3_X1 U7882 ( .A1(n8519), .A2(n8518), .A3(n8517), .ZN(n8530) );
  AND2_X1 U7883 ( .A1(n8447), .A2(n8446), .ZN(n12062) );
  AND2_X1 U7884 ( .A1(n7377), .A2(n7376), .ZN(n10527) );
  OR2_X1 U7885 ( .A1(n13031), .A2(n11013), .ZN(n7377) );
  NAND2_X1 U7886 ( .A1(n13031), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7376) );
  NAND2_X1 U7887 ( .A1(n6638), .A2(n10729), .ZN(n10731) );
  NAND2_X1 U7888 ( .A1(n10612), .A2(n10728), .ZN(n10733) );
  NAND2_X1 U7889 ( .A1(n7432), .A2(n7431), .ZN(n10612) );
  NAND2_X1 U7890 ( .A1(n10607), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7431) );
  NAND2_X1 U7891 ( .A1(n7088), .A2(n7087), .ZN(n10631) );
  NAND2_X1 U7892 ( .A1(n13031), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7087) );
  OR2_X1 U7893 ( .A1(n13031), .A2(n6832), .ZN(n7088) );
  NAND2_X1 U7894 ( .A1(n10616), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10651) );
  AOI21_X1 U7895 ( .B1(n10884), .B2(n10882), .A(n10883), .ZN(n11138) );
  NAND2_X1 U7896 ( .A1(n7361), .A2(n7366), .ZN(n7356) );
  NAND2_X1 U7897 ( .A1(n7355), .A2(n7366), .ZN(n7354) );
  AOI21_X1 U7898 ( .B1(n7361), .B2(n7363), .A(n7360), .ZN(n7359) );
  INV_X1 U7899 ( .A(n10878), .ZN(n7360) );
  NAND2_X1 U7900 ( .A1(n11152), .A2(n11153), .ZN(n11396) );
  NAND2_X1 U7901 ( .A1(n6978), .A2(n11137), .ZN(n11380) );
  XNOR2_X1 U7902 ( .A(n6820), .B(n11732), .ZN(n11724) );
  NOR2_X1 U7903 ( .A1(n12605), .A2(n12604), .ZN(n12631) );
  NAND3_X1 U7904 ( .A1(n6824), .A2(n12624), .A3(n6823), .ZN(n12639) );
  NAND2_X1 U7905 ( .A1(n6828), .A2(n12608), .ZN(n6824) );
  NAND2_X1 U7906 ( .A1(n6835), .A2(n12673), .ZN(n12674) );
  NAND2_X1 U7907 ( .A1(n7421), .A2(n12672), .ZN(n6835) );
  NAND2_X1 U7908 ( .A1(n8504), .A2(n8502), .ZN(n12207) );
  NAND2_X1 U7909 ( .A1(n7943), .A2(n7942), .ZN(n7975) );
  INV_X1 U7910 ( .A(n7992), .ZN(n7943) );
  AOI21_X1 U7911 ( .B1(n7151), .B2(n7149), .A(n6521), .ZN(n7148) );
  AOI21_X1 U7912 ( .B1(n7742), .B2(n7744), .A(n6484), .ZN(n7740) );
  INV_X1 U7913 ( .A(n7938), .ZN(n8239) );
  AND3_X1 U7914 ( .A1(n8229), .A2(n8228), .A3(n8227), .ZN(n12405) );
  NOR2_X1 U7915 ( .A1(n12046), .A2(n7756), .ZN(n7755) );
  INV_X1 U7916 ( .A(n9886), .ZN(n7756) );
  NOR2_X1 U7917 ( .A1(n6890), .A2(n6889), .ZN(n6888) );
  INV_X1 U7918 ( .A(n8472), .ZN(n6889) );
  NAND2_X1 U7919 ( .A1(n8191), .A2(n7936), .ZN(n8211) );
  INV_X1 U7920 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7936) );
  OR2_X2 U7921 ( .A1(n8164), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8177) );
  NAND2_X1 U7922 ( .A1(n11441), .A2(n11443), .ZN(n7481) );
  NAND2_X1 U7923 ( .A1(n7138), .A2(n9877), .ZN(n11445) );
  INV_X1 U7924 ( .A(n9871), .ZN(n11094) );
  CLKBUF_X1 U7925 ( .A(n10980), .Z(n10981) );
  NAND2_X1 U7926 ( .A1(n9950), .A2(n9949), .ZN(n11777) );
  OR2_X1 U7927 ( .A1(n8063), .A2(n10094), .ZN(n8024) );
  NAND2_X1 U7928 ( .A1(n10694), .A2(n10693), .ZN(n10696) );
  NAND2_X1 U7929 ( .A1(n8423), .A2(n8422), .ZN(n8526) );
  AOI21_X1 U7930 ( .B1(n12714), .B2(n8395), .A(n8394), .ZN(n12511) );
  AND2_X1 U7931 ( .A1(n6679), .A2(n6597), .ZN(n7140) );
  NAND2_X1 U7932 ( .A1(n7141), .A2(n7759), .ZN(n6679) );
  NAND2_X1 U7933 ( .A1(n7140), .A2(n6678), .ZN(n12741) );
  AND2_X1 U7934 ( .A1(n7139), .A2(n12742), .ZN(n6678) );
  NAND2_X1 U7935 ( .A1(n8373), .A2(n8497), .ZN(n12742) );
  NAND2_X1 U7936 ( .A1(n7473), .A2(n8494), .ZN(n12754) );
  INV_X1 U7937 ( .A(n12756), .ZN(n7473) );
  AND2_X1 U7938 ( .A1(n6700), .A2(n6701), .ZN(n6697) );
  AOI21_X1 U7939 ( .B1(n12774), .B2(n8491), .A(n8490), .ZN(n12764) );
  AND2_X1 U7940 ( .A1(n9891), .A2(n6488), .ZN(n7151) );
  NAND2_X1 U7941 ( .A1(n12831), .A2(n9890), .ZN(n7152) );
  AND2_X1 U7942 ( .A1(n12813), .A2(n8479), .ZN(n12822) );
  OR2_X1 U7943 ( .A1(n12387), .A2(n12514), .ZN(n8470) );
  NAND2_X1 U7944 ( .A1(n11911), .A2(n11913), .ZN(n7477) );
  AND2_X1 U7945 ( .A1(n8471), .A2(n8472), .ZN(n12034) );
  AND4_X1 U7946 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n12344)
         );
  AND2_X1 U7947 ( .A1(n8470), .A2(n8469), .ZN(n11913) );
  AOI21_X1 U7948 ( .B1(n7531), .B2(n7957), .A(n8380), .ZN(n7530) );
  AND2_X1 U7949 ( .A1(n7041), .A2(n6591), .ZN(n7040) );
  NAND2_X1 U7950 ( .A1(n6705), .A2(n7899), .ZN(n8359) );
  INV_X1 U7951 ( .A(n7899), .ZN(n6704) );
  AND2_X1 U7952 ( .A1(n7898), .A2(n7897), .ZN(n8338) );
  XNOR2_X1 U7953 ( .A(n8448), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U7954 ( .A1(n8555), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8448) );
  AND2_X1 U7955 ( .A1(n7894), .A2(n7893), .ZN(n8301) );
  INV_X1 U7956 ( .A(n6693), .ZN(n6692) );
  OAI21_X1 U7957 ( .B1(n7497), .B2(n6694), .A(n8301), .ZN(n6693) );
  INV_X1 U7958 ( .A(n7892), .ZN(n6694) );
  AND2_X1 U7959 ( .A1(n7890), .A2(n7889), .ZN(n8281) );
  INV_X1 U7960 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8221) );
  INV_X1 U7961 ( .A(n7880), .ZN(n7537) );
  AOI21_X1 U7962 ( .B1(n6550), .B2(n7880), .A(n7536), .ZN(n7535) );
  INV_X1 U7963 ( .A(n7882), .ZN(n7536) );
  AND2_X1 U7964 ( .A1(n10235), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7881) );
  AND2_X1 U7965 ( .A1(n10187), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7872) );
  INV_X1 U7966 ( .A(n7980), .ZN(n7981) );
  AND2_X1 U7967 ( .A1(n7738), .A2(n6540), .ZN(n6656) );
  AOI21_X1 U7968 ( .B1(n7517), .B2(n7515), .A(n6544), .ZN(n7514) );
  INV_X1 U7969 ( .A(n7871), .ZN(n7515) );
  INV_X1 U7970 ( .A(n7517), .ZN(n7516) );
  NAND2_X1 U7971 ( .A1(n8621), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7871) );
  INV_X1 U7972 ( .A(n8108), .ZN(n7518) );
  NAND2_X1 U7973 ( .A1(n7869), .A2(n7868), .ZN(n8109) );
  NAND2_X1 U7974 ( .A1(n10063), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U7975 ( .A1(n8086), .A2(n8087), .ZN(n7510) );
  NAND2_X1 U7976 ( .A1(n6553), .A2(n7860), .ZN(n6681) );
  NAND2_X1 U7977 ( .A1(n8058), .A2(n8014), .ZN(n8080) );
  AND2_X1 U7978 ( .A1(n8041), .A2(n7979), .ZN(n8058) );
  NAND2_X1 U7979 ( .A1(n7857), .A2(n7856), .ZN(n8020) );
  XNOR2_X1 U7980 ( .A(n8022), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10528) );
  AND2_X1 U7981 ( .A1(n10917), .A2(n10920), .ZN(n7441) );
  NAND2_X1 U7982 ( .A1(n10681), .A2(n6856), .ZN(n8791) );
  INV_X1 U7983 ( .A(n8773), .ZN(n6856) );
  NOR2_X1 U7984 ( .A1(n10110), .A2(n10065), .ZN(n7540) );
  XNOR2_X1 U7985 ( .A(n9109), .B(n6418), .ZN(n10825) );
  OR2_X1 U7986 ( .A1(n9139), .A2(n13065), .ZN(n9164) );
  OAI21_X1 U7987 ( .B1(n13149), .B2(n7450), .A(n6852), .ZN(n7448) );
  NAND2_X1 U7988 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  INV_X1 U7989 ( .A(n13058), .ZN(n7451) );
  INV_X1 U7990 ( .A(n13126), .ZN(n7447) );
  NAND2_X1 U7991 ( .A1(n11106), .A2(n8865), .ZN(n11063) );
  NAND2_X1 U7992 ( .A1(n13198), .A2(n13200), .ZN(n10908) );
  NAND2_X1 U7993 ( .A1(n8584), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9139) );
  INV_X1 U7994 ( .A(n9137), .ZN(n8584) );
  XNOR2_X1 U7995 ( .A(n6855), .B(n9146), .ZN(n13149) );
  INV_X1 U7996 ( .A(n13631), .ZN(n13740) );
  AND2_X1 U7997 ( .A1(n9281), .A2(n9280), .ZN(n13668) );
  AND2_X1 U7998 ( .A1(n9183), .A2(n9182), .ZN(n13637) );
  AND4_X1 U7999 ( .A1(n8920), .A2(n8919), .A3(n8918), .A4(n8917), .ZN(n13608)
         );
  NAND2_X1 U8000 ( .A1(n6819), .A2(n6815), .ZN(n6814) );
  INV_X1 U8001 ( .A(n6817), .ZN(n6815) );
  AOI21_X1 U8002 ( .B1(n15276), .B2(n15277), .A(n6818), .ZN(n6817) );
  INV_X1 U8003 ( .A(n13494), .ZN(n6818) );
  NAND2_X1 U8004 ( .A1(n10665), .A2(n10664), .ZN(n10702) );
  NAND2_X1 U8005 ( .A1(n6792), .A2(n6628), .ZN(n11668) );
  OR2_X1 U8006 ( .A1(n15309), .A2(n15310), .ZN(n6792) );
  NOR2_X1 U8007 ( .A1(n7122), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6796) );
  INV_X1 U8008 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U8009 ( .A1(n13346), .A2(n13345), .ZN(n13386) );
  NAND2_X1 U8010 ( .A1(n13371), .A2(n13370), .ZN(n13544) );
  INV_X1 U8011 ( .A(n13650), .ZN(n6670) );
  NOR2_X1 U8012 ( .A1(n7327), .A2(n13711), .ZN(n7326) );
  AND2_X1 U8013 ( .A1(n7710), .A2(n13587), .ZN(n7327) );
  INV_X1 U8014 ( .A(n13587), .ZN(n7328) );
  NAND2_X1 U8015 ( .A1(n7325), .A2(n13587), .ZN(n13699) );
  NAND2_X1 U8016 ( .A1(n7711), .A2(n7709), .ZN(n7325) );
  NAND2_X1 U8017 ( .A1(n7708), .A2(n7706), .ZN(n13758) );
  NOR2_X1 U8018 ( .A1(n13755), .A2(n7707), .ZN(n7706) );
  INV_X1 U8019 ( .A(n13581), .ZN(n7707) );
  INV_X1 U8020 ( .A(n6653), .ZN(n9111) );
  AND2_X1 U8021 ( .A1(n7832), .A2(n6473), .ZN(n7823) );
  INV_X1 U8022 ( .A(n13779), .ZN(n13578) );
  NAND2_X1 U8023 ( .A1(n13794), .A2(n13796), .ZN(n7712) );
  XNOR2_X1 U8024 ( .A(n13997), .B(n13628), .ZN(n13796) );
  NAND2_X1 U8025 ( .A1(n13834), .A2(n6504), .ZN(n13818) );
  NAND2_X1 U8026 ( .A1(n6640), .A2(n6437), .ZN(n7310) );
  INV_X1 U8027 ( .A(n13864), .ZN(n6640) );
  NAND2_X1 U8028 ( .A1(n7318), .A2(n7315), .ZN(n7309) );
  NOR2_X1 U8029 ( .A1(n7808), .A2(n13621), .ZN(n7805) );
  NAND2_X1 U8030 ( .A1(n7811), .A2(n13859), .ZN(n7807) );
  CLKBUF_X1 U8031 ( .A(n13864), .Z(n13865) );
  OR2_X1 U8032 ( .A1(n13569), .A2(n13568), .ZN(n13618) );
  NOR2_X1 U8033 ( .A1(n13619), .A2(n7814), .ZN(n7813) );
  INV_X1 U8034 ( .A(n13615), .ZN(n7814) );
  OAI21_X1 U8035 ( .B1(n13567), .B2(n13900), .A(n13903), .ZN(n7060) );
  OR2_X1 U8036 ( .A1(n14036), .A2(n13611), .ZN(n13903) );
  AND2_X1 U8037 ( .A1(n8894), .A2(n8893), .ZN(n11577) );
  NAND2_X1 U8038 ( .A1(n7339), .A2(n7337), .ZN(n7335) );
  NOR2_X1 U8039 ( .A1(n11035), .A2(n7704), .ZN(n7703) );
  INV_X1 U8040 ( .A(n11035), .ZN(n7701) );
  OR2_X1 U8041 ( .A1(n13374), .A2(n9302), .ZN(n10371) );
  INV_X1 U8042 ( .A(n13871), .ZN(n13885) );
  BUF_X1 U8043 ( .A(n13662), .Z(n13680) );
  INV_X1 U8044 ( .A(n15377), .ZN(n14024) );
  NAND2_X1 U8045 ( .A1(n8839), .A2(n8838), .ZN(n15376) );
  NAND2_X1 U8046 ( .A1(n8700), .A2(n8701), .ZN(n10205) );
  NAND2_X1 U8047 ( .A1(n7046), .A2(n7045), .ZN(n8700) );
  NOR2_X1 U8048 ( .A1(n6481), .A2(n7048), .ZN(n7045) );
  INV_X1 U8049 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8698) );
  INV_X1 U8050 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9236) );
  INV_X1 U8051 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7458) );
  AND3_X1 U8052 ( .A1(n6764), .A2(n8596), .A3(n6765), .ZN(n7343) );
  OR2_X1 U8053 ( .A1(n8891), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8910) );
  INV_X1 U8054 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8725) );
  INV_X1 U8055 ( .A(n7689), .ZN(n7688) );
  OAI21_X1 U8056 ( .B1(n14152), .B2(n7690), .A(n14224), .ZN(n7689) );
  OR2_X1 U8057 ( .A1(n9423), .A2(n9422), .ZN(n9448) );
  NOR2_X1 U8058 ( .A1(n14142), .A2(n7698), .ZN(n7697) );
  INV_X1 U8059 ( .A(n12090), .ZN(n7698) );
  INV_X1 U8060 ( .A(n14243), .ZN(n10761) );
  AOI21_X1 U8061 ( .B1(n7684), .B2(n7016), .A(n6542), .ZN(n7015) );
  INV_X1 U8062 ( .A(n14179), .ZN(n7016) );
  INV_X1 U8063 ( .A(n7684), .ZN(n7017) );
  NAND2_X1 U8064 ( .A1(n12085), .A2(n12084), .ZN(n14202) );
  NAND2_X1 U8065 ( .A1(n11352), .A2(n14499), .ZN(n7006) );
  XNOR2_X1 U8066 ( .A(n6893), .B(n14246), .ZN(n6892) );
  NAND2_X1 U8067 ( .A1(n14457), .A2(n6422), .ZN(n6893) );
  INV_X1 U8068 ( .A(n14468), .ZN(n6891) );
  NAND2_X1 U8069 ( .A1(n14425), .A2(n14424), .ZN(n6953) );
  NAND2_X1 U8070 ( .A1(n6949), .A2(n6950), .ZN(n6948) );
  AND2_X1 U8071 ( .A1(n9650), .A2(n9649), .ZN(n14171) );
  OR2_X1 U8072 ( .A1(n14757), .A2(n9785), .ZN(n9650) );
  INV_X1 U8073 ( .A(n7194), .ZN(n9741) );
  OR2_X1 U8074 ( .A1(n6405), .A2(n10246), .ZN(n9356) );
  NAND2_X1 U8075 ( .A1(n9350), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8076 ( .A1(n10248), .A2(n10247), .ZN(n14536) );
  NAND2_X1 U8077 ( .A1(n11932), .A2(n11933), .ZN(n14599) );
  NAND2_X1 U8078 ( .A1(n9828), .A2(n9827), .ZN(n14668) );
  NAND2_X1 U8079 ( .A1(n9619), .A2(n6452), .ZN(n14663) );
  NOR2_X1 U8080 ( .A1(n14732), .A2(n6977), .ZN(n6976) );
  INV_X1 U8081 ( .A(n14711), .ZN(n6977) );
  NAND2_X1 U8082 ( .A1(n14785), .A2(n6428), .ZN(n14771) );
  NAND2_X1 U8083 ( .A1(n7774), .A2(n7775), .ZN(n14769) );
  OAI21_X1 U8084 ( .B1(n6427), .B2(n7776), .A(n6474), .ZN(n7775) );
  INV_X1 U8085 ( .A(n14780), .ZN(n7776) );
  INV_X1 U8086 ( .A(n14768), .ZN(n14766) );
  AND2_X1 U8087 ( .A1(n9614), .A2(n9613), .ZN(n14784) );
  OR2_X1 U8088 ( .A1(n14197), .A2(n9785), .ZN(n9614) );
  AND2_X1 U8089 ( .A1(n6491), .A2(n9769), .ZN(n7778) );
  OAI21_X1 U8090 ( .B1(n7773), .B2(n6963), .A(n6961), .ZN(n9770) );
  AND2_X1 U8091 ( .A1(n7666), .A2(n7166), .ZN(n7165) );
  NAND2_X1 U8092 ( .A1(n7167), .A2(n7173), .ZN(n7166) );
  NOR2_X1 U8093 ( .A1(n6411), .A2(n7673), .ZN(n7672) );
  INV_X1 U8094 ( .A(n9569), .ZN(n7673) );
  NAND2_X1 U8095 ( .A1(n7169), .A2(n7171), .ZN(n9570) );
  OR2_X1 U8096 ( .A1(n14854), .A2(n7173), .ZN(n7169) );
  AND3_X1 U8097 ( .A1(n9581), .A2(n9580), .A3(n9579), .ZN(n14827) );
  NOR2_X1 U8098 ( .A1(n9559), .A2(n7175), .ZN(n7174) );
  INV_X1 U8099 ( .A(n9544), .ZN(n7175) );
  AND2_X1 U8100 ( .A1(n14900), .A2(n6569), .ZN(n14828) );
  NAND2_X1 U8101 ( .A1(n7773), .A2(n7772), .ZN(n14840) );
  AND2_X1 U8102 ( .A1(n14342), .A2(n14343), .ZN(n14877) );
  NAND2_X1 U8103 ( .A1(n9763), .A2(n14341), .ZN(n14876) );
  NAND2_X1 U8104 ( .A1(n9512), .A2(n9511), .ZN(n14901) );
  NAND2_X1 U8105 ( .A1(n6642), .A2(n7679), .ZN(n14893) );
  INV_X1 U8106 ( .A(n6967), .ZN(n6968) );
  INV_X1 U8107 ( .A(n14450), .ZN(n14919) );
  NAND2_X1 U8108 ( .A1(n11823), .A2(n7782), .ZN(n11862) );
  NOR2_X1 U8109 ( .A1(n14289), .A2(n14956), .ZN(n7721) );
  INV_X1 U8110 ( .A(n15215), .ZN(n7719) );
  NAND2_X1 U8111 ( .A1(n11705), .A2(n14443), .ZN(n11704) );
  NAND2_X1 U8112 ( .A1(n10093), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7401) );
  NAND2_X1 U8113 ( .A1(n14651), .A2(n6500), .ZN(n9983) );
  NAND2_X1 U8114 ( .A1(n9618), .A2(n9617), .ZN(n14995) );
  NAND2_X1 U8115 ( .A1(n11113), .A2(n9845), .ZN(n7262) );
  NAND2_X1 U8116 ( .A1(n9495), .A2(n9494), .ZN(n15065) );
  AND2_X1 U8117 ( .A1(n11574), .A2(P1_B_REG_SCAN_IN), .ZN(n9721) );
  NAND2_X1 U8118 ( .A1(n9833), .A2(n9832), .ZN(n9840) );
  XNOR2_X1 U8119 ( .A(n9830), .B(n9829), .ZN(n13342) );
  NAND2_X1 U8120 ( .A1(n6747), .A2(n6745), .ZN(n9823) );
  AOI21_X1 U8121 ( .B1(n6748), .B2(n6608), .A(n6746), .ZN(n6745) );
  NAND2_X1 U8122 ( .A1(n9157), .A2(n6743), .ZN(n6747) );
  NOR2_X1 U8123 ( .A1(n9213), .A2(n13037), .ZN(n6746) );
  INV_X1 U8124 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U8125 ( .A(n9215), .B(n9193), .ZN(n11783) );
  NAND2_X1 U8126 ( .A1(n6744), .A2(n6748), .ZN(n9215) );
  OR2_X1 U8127 ( .A1(n9157), .A2(n6750), .ZN(n6744) );
  NAND2_X1 U8128 ( .A1(n9546), .A2(n7715), .ZN(n9711) );
  INV_X1 U8129 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9703) );
  INV_X1 U8130 ( .A(n9711), .ZN(n9707) );
  NOR2_X1 U8131 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9706) );
  NAND2_X1 U8132 ( .A1(n7081), .A2(n7080), .ZN(n9719) );
  INV_X1 U8133 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U8134 ( .A1(n8692), .A2(n9150), .ZN(n8693) );
  OR2_X1 U8135 ( .A1(n9153), .A2(n9158), .ZN(n8692) );
  NOR2_X1 U8136 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6933) );
  INV_X1 U8137 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9692) );
  INV_X1 U8138 ( .A(n7597), .ZN(n7595) );
  OR2_X1 U8139 ( .A1(n9072), .A2(n15447), .ZN(n9104) );
  XNOR2_X1 U8140 ( .A(n7063), .B(n8931), .ZN(n10236) );
  OAI21_X1 U8141 ( .B1(n8950), .B2(n8928), .A(n8927), .ZN(n7063) );
  XNOR2_X1 U8142 ( .A(n8852), .B(n7276), .ZN(n10111) );
  INV_X1 U8143 ( .A(n8645), .ZN(n7276) );
  INV_X1 U8144 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9319) );
  OR2_X1 U8145 ( .A1(n11250), .A2(n11249), .ZN(n11252) );
  NAND2_X1 U8146 ( .A1(n11984), .A2(n11983), .ZN(n15115) );
  OR2_X1 U8147 ( .A1(n11982), .A2(n11981), .ZN(n11984) );
  NAND2_X1 U8148 ( .A1(n11468), .A2(n11467), .ZN(n11471) );
  NAND2_X1 U8149 ( .A1(n7582), .A2(n12205), .ZN(n12335) );
  INV_X1 U8150 ( .A(n12336), .ZN(n6673) );
  INV_X1 U8151 ( .A(n12744), .ZN(n12397) );
  NAND2_X1 U8152 ( .A1(n11020), .A2(n11019), .ZN(n11183) );
  INV_X1 U8153 ( .A(n12860), .ZN(n12417) );
  NAND2_X1 U8154 ( .A1(n8051), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7493) );
  NAND2_X1 U8155 ( .A1(n8091), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U8156 ( .A1(n8050), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U8157 ( .A1(n7027), .A2(n10805), .ZN(n7239) );
  INV_X1 U8158 ( .A(n12888), .ZN(n10812) );
  NAND2_X1 U8159 ( .A1(n11288), .A2(n11287), .ZN(n11468) );
  INV_X1 U8160 ( .A(n12497), .ZN(n12488) );
  NAND2_X1 U8161 ( .A1(n7225), .A2(n12176), .ZN(n12495) );
  NAND2_X1 U8162 ( .A1(n10564), .A2(n10563), .ZN(n12502) );
  NAND2_X1 U8163 ( .A1(n10575), .A2(n12891), .ZN(n12503) );
  INV_X1 U8164 ( .A(n12357), .ZN(n12767) );
  NAND2_X1 U8165 ( .A1(n8335), .A2(n8334), .ZN(n12805) );
  INV_X1 U8166 ( .A(n12473), .ZN(n12832) );
  NAND2_X1 U8167 ( .A1(n8299), .A2(n8298), .ZN(n12846) );
  INV_X1 U8168 ( .A(n12344), .ZN(n12513) );
  INV_X1 U8169 ( .A(n12450), .ZN(n12514) );
  NAND4_X1 U8170 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n12520)
         );
  CLKBUF_X1 U8171 ( .A(n8046), .Z(n12522) );
  XNOR2_X1 U8172 ( .A(n10527), .B(n7211), .ZN(n10530) );
  OAI21_X1 U8173 ( .B1(n10723), .B2(n10724), .A(n6479), .ZN(n10635) );
  XNOR2_X1 U8174 ( .A(n11380), .B(n11150), .ZN(n11378) );
  INV_X1 U8175 ( .A(n12660), .ZN(n7215) );
  AOI21_X1 U8176 ( .B1(n12661), .B2(n6996), .A(n7214), .ZN(n7213) );
  OAI21_X1 U8177 ( .B1(n12655), .B2(n15497), .A(n12654), .ZN(n7214) );
  INV_X1 U8178 ( .A(n7421), .ZN(n7420) );
  NAND2_X1 U8179 ( .A1(n7422), .A2(n12672), .ZN(n12650) );
  XNOR2_X1 U8180 ( .A(n12678), .B(n12677), .ZN(n7216) );
  NAND2_X1 U8181 ( .A1(n6988), .A2(n6989), .ZN(n12678) );
  AOI21_X1 U8182 ( .B1(n12628), .B2(n6991), .A(n6990), .ZN(n6989) );
  OR2_X1 U8183 ( .A1(n12628), .A2(n6995), .ZN(n6988) );
  AND2_X1 U8184 ( .A1(n10440), .A2(n10436), .ZN(n12688) );
  INV_X1 U8185 ( .A(n12704), .ZN(n7345) );
  NOR2_X1 U8186 ( .A1(n12701), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U8187 ( .A1(n7929), .A2(n7928), .ZN(n9906) );
  NAND2_X1 U8188 ( .A1(n6896), .A2(n7487), .ZN(n6895) );
  AOI21_X1 U8189 ( .B1(n12724), .B2(n12883), .A(n12723), .ZN(n12901) );
  NAND2_X1 U8190 ( .A1(n12722), .A2(n12721), .ZN(n12723) );
  NAND2_X1 U8191 ( .A1(n12744), .A2(n12880), .ZN(n12721) );
  INV_X1 U8192 ( .A(n7142), .ZN(n7757) );
  AOI21_X1 U8193 ( .B1(n12159), .B2(n8437), .A(n8307), .ZN(n12811) );
  NAND2_X1 U8194 ( .A1(n8290), .A2(n8289), .ZN(n12935) );
  OR2_X1 U8195 ( .A1(n8389), .A2(n7845), .ZN(n8103) );
  NAND2_X1 U8196 ( .A1(n6875), .A2(n6874), .ZN(n6873) );
  NAND2_X1 U8197 ( .A1(n8288), .A2(SI_4_), .ZN(n6876) );
  NAND2_X1 U8198 ( .A1(n8147), .A2(n8146), .ZN(n11882) );
  NAND2_X1 U8199 ( .A1(n8225), .A2(n8224), .ZN(n13006) );
  NAND2_X1 U8200 ( .A1(n8163), .A2(n8162), .ZN(n12022) );
  CLKBUF_X1 U8201 ( .A(n8571), .Z(n13027) );
  INV_X1 U8202 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8305) );
  OAI21_X1 U8203 ( .B1(n6425), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8306) );
  INV_X1 U8204 ( .A(n10528), .ZN(n7211) );
  AND3_X1 U8205 ( .A1(n8990), .A2(n8989), .A3(n8988), .ZN(n13620) );
  OR2_X1 U8206 ( .A1(n11335), .A2(n9160), .ZN(n8704) );
  AOI21_X1 U8207 ( .B1(n13167), .B2(n6859), .A(n9266), .ZN(n9285) );
  NOR2_X1 U8208 ( .A1(n6860), .A2(n13165), .ZN(n6859) );
  INV_X1 U8209 ( .A(n6860), .ZN(n6858) );
  AND4_X1 U8210 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n13256)
         );
  INV_X1 U8211 ( .A(n13692), .ZN(n13962) );
  INV_X1 U8212 ( .A(n13623), .ZN(n13870) );
  INV_X1 U8213 ( .A(n13667), .ZN(n13702) );
  INV_X1 U8214 ( .A(n13637), .ZN(n13682) );
  OR2_X1 U8215 ( .A1(n13722), .A2(n9223), .ZN(n9171) );
  NAND2_X1 U8216 ( .A1(n9118), .A2(n9117), .ZN(n13630) );
  NAND2_X1 U8217 ( .A1(n9066), .A2(n9065), .ZN(n13797) );
  INV_X1 U8218 ( .A(n13620), .ZN(n13886) );
  INV_X1 U8219 ( .A(n7797), .ZN(n7796) );
  AND2_X1 U8220 ( .A1(n7795), .A2(n8720), .ZN(n7794) );
  OAI21_X1 U8221 ( .B1(n8745), .B2(n8719), .A(n7729), .ZN(n7797) );
  NAND2_X1 U8222 ( .A1(n6791), .A2(n6517), .ZN(n10661) );
  OR2_X1 U8223 ( .A1(n10299), .A2(n10298), .ZN(n6791) );
  NAND2_X1 U8224 ( .A1(n10714), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8225 ( .A1(n13540), .A2(n15315), .ZN(n6784) );
  INV_X1 U8226 ( .A(n6783), .ZN(n6782) );
  CLKBUF_X1 U8227 ( .A(n13197), .Z(n13541) );
  OAI21_X1 U8228 ( .B1(n13540), .B2(n15300), .A(n6787), .ZN(n6786) );
  NAND2_X1 U8229 ( .A1(n13539), .A2(n15318), .ZN(n6787) );
  NOR2_X1 U8230 ( .A1(n15322), .A2(n6730), .ZN(n6779) );
  AND2_X1 U8231 ( .A1(n9273), .A2(n9272), .ZN(n13656) );
  NAND2_X1 U8232 ( .A1(n7802), .A2(n6463), .ZN(n6762) );
  NAND2_X1 U8233 ( .A1(n9078), .A2(n9077), .ZN(n13993) );
  OR2_X1 U8234 ( .A1(n11130), .A2(n9160), .ZN(n9078) );
  NAND2_X1 U8235 ( .A1(n13947), .A2(n15377), .ZN(n7542) );
  NOR2_X1 U8236 ( .A1(n6518), .A2(n6769), .ZN(n6767) );
  INV_X1 U8237 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14082) );
  AND4_X1 U8238 ( .A1(n6764), .A2(n7341), .A3(n6765), .A4(n8596), .ZN(n6763)
         );
  AND2_X1 U8239 ( .A1(n8598), .A2(n7049), .ZN(n7341) );
  INV_X1 U8240 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8598) );
  INV_X1 U8241 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U8242 ( .A1(n9681), .A2(n9680), .ZN(n14408) );
  NAND2_X1 U8243 ( .A1(n9593), .A2(n9592), .ZN(n15017) );
  OR2_X1 U8244 ( .A1(n11230), .A2(n9637), .ZN(n9593) );
  INV_X1 U8245 ( .A(n14152), .ZN(n7096) );
  AND4_X1 U8246 ( .A1(n9531), .A2(n9530), .A3(n9529), .A4(n9528), .ZN(n14862)
         );
  INV_X1 U8247 ( .A(n15000), .ZN(n14739) );
  OR2_X1 U8248 ( .A1(n11130), .A2(n9637), .ZN(n9584) );
  NAND2_X1 U8249 ( .A1(n10760), .A2(n10761), .ZN(n14198) );
  NAND2_X1 U8250 ( .A1(n11371), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15182) );
  NOR2_X2 U8251 ( .A1(n14231), .A2(n15259), .ZN(n14221) );
  NAND2_X1 U8252 ( .A1(n12289), .A2(n12288), .ZN(n14151) );
  OR2_X1 U8253 ( .A1(n12287), .A2(n12286), .ZN(n12288) );
  NAND2_X1 U8254 ( .A1(n7024), .A2(n12297), .ZN(n7023) );
  INV_X1 U8255 ( .A(n14224), .ZN(n7024) );
  AND4_X1 U8256 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n14345)
         );
  NAND2_X1 U8257 ( .A1(n9602), .A2(n9601), .ZN(n14484) );
  NAND2_X1 U8258 ( .A1(n9591), .A2(n9590), .ZN(n14816) );
  INV_X1 U8259 ( .A(n14827), .ZN(n14485) );
  NOR2_X1 U8260 ( .A1(n10312), .A2(n6472), .ZN(n14552) );
  NAND2_X1 U8261 ( .A1(n14561), .A2(n6837), .ZN(n10451) );
  AND2_X1 U8262 ( .A1(n10337), .A2(n10338), .ZN(n6837) );
  NAND2_X1 U8263 ( .A1(n14562), .A2(n14563), .ZN(n14561) );
  NOR2_X1 U8264 ( .A1(n10455), .A2(n10454), .ZN(n10769) );
  OAI21_X1 U8265 ( .B1(n14636), .B2(n14635), .A(n6848), .ZN(n6847) );
  OR2_X1 U8266 ( .A1(n14638), .A2(n14637), .ZN(n6848) );
  NAND2_X1 U8267 ( .A1(n14636), .A2(n15188), .ZN(n14634) );
  AND2_X1 U8268 ( .A1(n10161), .A2(n10159), .ZN(n15199) );
  XNOR2_X1 U8269 ( .A(n9847), .B(n9846), .ZN(n14640) );
  NOR2_X1 U8270 ( .A1(n9976), .A2(n14648), .ZN(n9847) );
  AOI21_X1 U8271 ( .B1(n7192), .B2(n15251), .A(n9793), .ZN(n9811) );
  OAI21_X1 U8272 ( .B1(n14676), .B2(n9781), .A(n14655), .ZN(n7192) );
  AND2_X1 U8273 ( .A1(n14683), .A2(n6480), .ZN(n14982) );
  INV_X1 U8274 ( .A(n14395), .ZN(n14700) );
  OAI21_X1 U8275 ( .B1(n14695), .B2(n14694), .A(n14693), .ZN(n14696) );
  NAND2_X1 U8276 ( .A1(n15220), .A2(n15263), .ZN(n14910) );
  OR2_X1 U8277 ( .A1(n9384), .A2(n10059), .ZN(n9364) );
  NAND2_X1 U8278 ( .A1(n7185), .A2(n6501), .ZN(n7187) );
  INV_X1 U8279 ( .A(n14737), .ZN(n7184) );
  OR2_X1 U8280 ( .A1(n14735), .A2(n14734), .ZN(n14736) );
  INV_X1 U8281 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15446) );
  AND2_X1 U8282 ( .A1(n7787), .A2(n9331), .ZN(n7786) );
  INV_X1 U8283 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U8284 ( .A1(n7071), .A2(n6490), .ZN(n11248) );
  NAND2_X1 U8285 ( .A1(n6663), .A2(n7086), .ZN(n7304) );
  NAND2_X1 U8286 ( .A1(n15121), .A2(n15120), .ZN(n7303) );
  AND2_X1 U8287 ( .A1(n6666), .A2(n7252), .ZN(n15121) );
  AND2_X1 U8288 ( .A1(n7077), .A2(n15141), .ZN(n7075) );
  NAND2_X1 U8289 ( .A1(n7622), .A2(n13216), .ZN(n7621) );
  INV_X1 U8290 ( .A(n13217), .ZN(n7622) );
  NOR2_X1 U8291 ( .A1(n13230), .A2(n13227), .ZN(n7651) );
  INV_X1 U8292 ( .A(n13227), .ZN(n7650) );
  NAND2_X1 U8293 ( .A1(n7378), .A2(n14264), .ZN(n14274) );
  NAND2_X1 U8294 ( .A1(n14263), .A2(n14262), .ZN(n14264) );
  OAI21_X1 U8295 ( .B1(n14261), .B2(n14414), .A(n14260), .ZN(n14262) );
  OAI21_X1 U8296 ( .B1(n14253), .B2(n14265), .A(n14269), .ZN(n14270) );
  AOI21_X1 U8297 ( .B1(n6657), .B2(n8170), .A(n11776), .ZN(n8200) );
  AOI21_X1 U8298 ( .B1(n7644), .B2(n7643), .A(n7641), .ZN(n7640) );
  INV_X1 U8299 ( .A(n13243), .ZN(n7641) );
  NAND2_X1 U8300 ( .A1(n6956), .A2(n14285), .ZN(n6955) );
  NAND2_X1 U8301 ( .A1(n7385), .A2(n7384), .ZN(n7382) );
  OAI21_X1 U8302 ( .B1(n14282), .B2(n7385), .A(n7384), .ZN(n6958) );
  NAND2_X1 U8303 ( .A1(n6555), .A2(n7630), .ZN(n7627) );
  NAND2_X1 U8304 ( .A1(n7630), .A2(n6507), .ZN(n7628) );
  INV_X1 U8305 ( .A(n14290), .ZN(n6928) );
  AND2_X1 U8306 ( .A1(n14309), .A2(n14350), .ZN(n6945) );
  NOR2_X1 U8307 ( .A1(n6946), .A2(n14340), .ZN(n6941) );
  AOI21_X1 U8308 ( .B1(n14364), .B2(n14365), .A(n6514), .ZN(n7389) );
  INV_X1 U8309 ( .A(n14364), .ZN(n7388) );
  NAND2_X1 U8310 ( .A1(n7261), .A2(n7260), .ZN(n14369) );
  INV_X1 U8311 ( .A(n8337), .ZN(n6660) );
  INV_X1 U8312 ( .A(n8354), .ZN(n6647) );
  NAND2_X1 U8313 ( .A1(n13297), .A2(n7649), .ZN(n7646) );
  OR2_X1 U8314 ( .A1(n13295), .A2(n7647), .ZN(n7645) );
  OR2_X1 U8315 ( .A1(n7648), .A2(n13294), .ZN(n7647) );
  NAND2_X1 U8316 ( .A1(n13300), .A2(n6720), .ZN(n6719) );
  AND2_X1 U8317 ( .A1(n13298), .A2(n6722), .ZN(n6721) );
  INV_X1 U8318 ( .A(n13300), .ZN(n6722) );
  INV_X1 U8319 ( .A(n14380), .ZN(n6938) );
  NAND2_X1 U8320 ( .A1(n7259), .A2(n7386), .ZN(n7256) );
  NAND2_X1 U8321 ( .A1(n7387), .A2(n6411), .ZN(n7386) );
  NAND2_X1 U8322 ( .A1(n7389), .A2(n7388), .ZN(n7387) );
  NOR2_X1 U8323 ( .A1(n7300), .A2(n12757), .ZN(n7299) );
  INV_X1 U8324 ( .A(n8372), .ZN(n7300) );
  NAND2_X1 U8325 ( .A1(n13315), .A2(n13312), .ZN(n7638) );
  NAND2_X1 U8326 ( .A1(n7282), .A2(n7124), .ZN(n14390) );
  NAND2_X1 U8327 ( .A1(n14386), .A2(n14385), .ZN(n7282) );
  INV_X1 U8328 ( .A(n14392), .ZN(n7396) );
  INV_X1 U8329 ( .A(n7638), .ZN(n6716) );
  NOR2_X1 U8330 ( .A1(n13315), .A2(n13312), .ZN(n7639) );
  AOI21_X1 U8331 ( .B1(n7616), .B2(n8677), .A(n7615), .ZN(n7614) );
  NAND2_X1 U8332 ( .A1(n8675), .A2(SI_17_), .ZN(n7616) );
  NOR2_X1 U8333 ( .A1(n8675), .A2(SI_17_), .ZN(n7615) );
  NOR3_X1 U8334 ( .A1(n13400), .A2(n13399), .A3(n13398), .ZN(n13403) );
  NOR2_X1 U8335 ( .A1(n8938), .A2(n8937), .ZN(n8936) );
  NOR2_X1 U8336 ( .A1(n8878), .A2(n8877), .ZN(n6654) );
  OR2_X1 U8337 ( .A1(n14447), .A2(n7659), .ZN(n7658) );
  INV_X1 U8338 ( .A(n7848), .ZN(n6741) );
  AOI21_X1 U8339 ( .B1(n7612), .B2(n7617), .A(n6519), .ZN(n7611) );
  OAI21_X1 U8340 ( .B1(n8676), .B2(n7617), .A(n7614), .ZN(n9052) );
  AOI21_X1 U8341 ( .B1(n8664), .B2(n7609), .A(n6543), .ZN(n7608) );
  NOR2_X1 U8342 ( .A1(n8657), .A2(n8670), .ZN(n7609) );
  NAND2_X1 U8343 ( .A1(n6737), .A2(n6736), .ZN(n7610) );
  NOR2_X1 U8344 ( .A1(n8670), .A2(n6739), .ZN(n6736) );
  INV_X1 U8345 ( .A(n8641), .ZN(n7058) );
  NAND2_X1 U8346 ( .A1(n10070), .A2(n10069), .ZN(n10106) );
  INV_X1 U8347 ( .A(n8550), .ZN(n8512) );
  NOR2_X1 U8348 ( .A1(n12140), .A2(n6644), .ZN(n6643) );
  INV_X1 U8349 ( .A(n8413), .ZN(n6644) );
  NAND2_X1 U8350 ( .A1(n7207), .A2(n10513), .ZN(n10437) );
  NAND2_X1 U8351 ( .A1(n10528), .A2(n6516), .ZN(n7207) );
  NAND2_X1 U8352 ( .A1(n10528), .A2(n6510), .ZN(n10441) );
  NAND2_X1 U8353 ( .A1(n7354), .A2(n7353), .ZN(n7352) );
  INV_X1 U8354 ( .A(n11146), .ZN(n7353) );
  OAI21_X1 U8355 ( .B1(n7352), .B2(n7350), .A(n7365), .ZN(n7349) );
  OR2_X1 U8356 ( .A1(n11144), .A2(n11145), .ZN(n7365) );
  INV_X1 U8357 ( .A(n7356), .ZN(n7350) );
  OR2_X1 U8358 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  NOR2_X2 U8359 ( .A1(n8293), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7131) );
  INV_X1 U8360 ( .A(n9888), .ZN(n7744) );
  NAND2_X1 U8361 ( .A1(n10809), .A2(n11005), .ZN(n10802) );
  OR2_X1 U8362 ( .A1(n12935), .A2(n12846), .ZN(n12812) );
  INV_X1 U8363 ( .A(n11454), .ZN(n11456) );
  AND2_X1 U8364 ( .A1(n7983), .A2(n7590), .ZN(n7041) );
  NAND2_X1 U8365 ( .A1(n7535), .A2(n8183), .ZN(n6728) );
  AOI21_X1 U8366 ( .B1(n7535), .B2(n7537), .A(n8219), .ZN(n7534) );
  INV_X1 U8367 ( .A(n7876), .ZN(n7538) );
  NAND2_X1 U8368 ( .A1(n7877), .A2(n7876), .ZN(n8204) );
  INV_X1 U8369 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7286) );
  INV_X1 U8370 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7459) );
  INV_X1 U8371 ( .A(n7862), .ZN(n6684) );
  NAND2_X1 U8372 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7412) );
  INV_X1 U8373 ( .A(n13052), .ZN(n7437) );
  OAI21_X1 U8374 ( .B1(n13059), .B2(n6854), .A(n7449), .ZN(n6853) );
  NAND2_X1 U8375 ( .A1(n9147), .A2(n9148), .ZN(n7449) );
  AND2_X1 U8376 ( .A1(n13060), .A2(n13062), .ZN(n6854) );
  NAND2_X1 U8377 ( .A1(n13060), .A2(n13633), .ZN(n7452) );
  NAND2_X1 U8378 ( .A1(n13087), .A2(n9130), .ZN(n6855) );
  NAND2_X1 U8379 ( .A1(n11208), .A2(n6865), .ZN(n6864) );
  INV_X1 U8380 ( .A(n8868), .ZN(n6865) );
  OAI21_X1 U8381 ( .B1(n6795), .B2(n7122), .A(n6800), .ZN(n13530) );
  OR2_X1 U8382 ( .A1(n11666), .A2(n6454), .ZN(n6795) );
  NOR2_X1 U8383 ( .A1(n6801), .A2(n6629), .ZN(n6800) );
  NAND2_X1 U8384 ( .A1(n13586), .A2(n13585), .ZN(n7710) );
  NOR2_X1 U8385 ( .A1(n13982), .A2(n13978), .ZN(n7555) );
  OAI211_X1 U8386 ( .C1(n7819), .C2(n7824), .A(n7818), .B(n7816), .ZN(n7815)
         );
  NAND2_X1 U8387 ( .A1(n6426), .A2(n7832), .ZN(n7819) );
  NAND2_X1 U8388 ( .A1(n7823), .A2(n6426), .ZN(n7818) );
  AND2_X1 U8389 ( .A1(n7803), .A2(n13624), .ZN(n6755) );
  INV_X1 U8390 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8973) );
  INV_X1 U8391 ( .A(n13610), .ZN(n7792) );
  INV_X1 U8392 ( .A(n13606), .ZN(n7789) );
  NAND2_X1 U8393 ( .A1(n8936), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8974) );
  AND2_X1 U8394 ( .A1(n7090), .A2(n13903), .ZN(n6641) );
  INV_X1 U8395 ( .A(n7091), .ZN(n7090) );
  OAI21_X1 U8396 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n7091) );
  NAND2_X1 U8397 ( .A1(n6654), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8915) );
  INV_X1 U8398 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8914) );
  OR2_X1 U8399 ( .A1(n8915), .A2(n8914), .ZN(n8938) );
  INV_X1 U8400 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8877) );
  INV_X1 U8401 ( .A(n6654), .ZN(n8896) );
  AND2_X1 U8402 ( .A1(n7544), .A2(n11491), .ZN(n7547) );
  INV_X1 U8403 ( .A(n7548), .ZN(n7544) );
  NAND2_X1 U8404 ( .A1(n11409), .A2(n11637), .ZN(n7548) );
  AND2_X1 U8405 ( .A1(n11034), .A2(n15368), .ZN(n11035) );
  NAND2_X1 U8406 ( .A1(n7705), .A2(n11033), .ZN(n11647) );
  NOR2_X1 U8407 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7049), .ZN(n7048) );
  NOR2_X1 U8408 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n8590) );
  INV_X1 U8409 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8705) );
  NOR2_X1 U8410 ( .A1(n11242), .A2(n9498), .ZN(n6903) );
  INV_X1 U8411 ( .A(n9499), .ZN(n9497) );
  INV_X1 U8412 ( .A(n14404), .ZN(n7379) );
  NAND2_X1 U8413 ( .A1(n7278), .A2(n6952), .ZN(n6949) );
  NAND2_X1 U8414 ( .A1(n14422), .A2(n14423), .ZN(n6952) );
  OR2_X1 U8415 ( .A1(n6842), .A2(n6625), .ZN(n6839) );
  OR2_X1 U8416 ( .A1(n6840), .A2(n6625), .ZN(n6838) );
  NOR2_X1 U8417 ( .A1(n14227), .A2(n14153), .ZN(n6897) );
  AND3_X1 U8418 ( .A1(n9653), .A2(n9651), .A3(n14733), .ZN(n9652) );
  AND2_X1 U8419 ( .A1(n7778), .A2(n6474), .ZN(n7777) );
  NAND2_X1 U8420 ( .A1(n6961), .A2(n6963), .ZN(n6959) );
  NOR2_X1 U8421 ( .A1(n9577), .A2(n9576), .ZN(n6906) );
  NOR2_X1 U8422 ( .A1(n7670), .A2(n7168), .ZN(n7167) );
  INV_X1 U8423 ( .A(n7171), .ZN(n7168) );
  AOI21_X1 U8424 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n7666) );
  INV_X1 U8425 ( .A(n14371), .ZN(n7667) );
  INV_X1 U8426 ( .A(n7672), .ZN(n7668) );
  INV_X1 U8427 ( .A(n9558), .ZN(n7173) );
  INV_X1 U8428 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9536) );
  NOR2_X1 U8429 ( .A1(n15053), .A2(n15046), .ZN(n7718) );
  NAND2_X1 U8430 ( .A1(n15053), .A2(n14862), .ZN(n14343) );
  AOI21_X1 U8431 ( .B1(n7779), .B2(n7781), .A(n6520), .ZN(n6967) );
  NAND2_X1 U8432 ( .A1(n6967), .A2(n6966), .ZN(n6965) );
  INV_X1 U8433 ( .A(n9390), .ZN(n6902) );
  NAND2_X1 U8434 ( .A1(n14267), .A2(n7852), .ZN(n14436) );
  NAND2_X1 U8435 ( .A1(n14258), .A2(n14260), .ZN(n10840) );
  AND2_X1 U8436 ( .A1(n14652), .A2(n15263), .ZN(n7663) );
  AND2_X1 U8437 ( .A1(n6428), .A2(n7731), .ZN(n7730) );
  INV_X1 U8438 ( .A(n14247), .ZN(n14416) );
  AND2_X1 U8439 ( .A1(n11131), .A2(n14917), .ZN(n9804) );
  NOR3_X1 U8440 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n9314) );
  INV_X1 U8441 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9317) );
  INV_X1 U8442 ( .A(n9318), .ZN(n7716) );
  INV_X1 U8443 ( .A(n6751), .ZN(n6750) );
  AOI21_X1 U8444 ( .B1(n6749), .B2(n6751), .A(n6612), .ZN(n6748) );
  INV_X1 U8445 ( .A(n7108), .ZN(n6749) );
  NAND2_X1 U8446 ( .A1(n8683), .A2(SI_21_), .ZN(n8686) );
  NAND2_X1 U8447 ( .A1(n8658), .A2(n10158), .ZN(n8927) );
  OR2_X1 U8448 ( .A1(n9469), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9479) );
  AOI21_X1 U8449 ( .B1(n7274), .B2(n7277), .A(n6533), .ZN(n7272) );
  INV_X1 U8450 ( .A(n8647), .ZN(n7277) );
  XNOR2_X1 U8451 ( .A(n8649), .B(SI_9_), .ZN(n8869) );
  OR2_X1 U8452 ( .A1(n9521), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9440) );
  XNOR2_X1 U8453 ( .A(n8640), .B(SI_6_), .ZN(n8796) );
  INV_X1 U8454 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U8455 ( .A1(n11169), .A2(n11168), .ZN(n11250) );
  NAND2_X1 U8456 ( .A1(n6999), .A2(n6997), .ZN(n12623) );
  AOI21_X1 U8457 ( .B1(n7201), .B2(n6998), .A(n12602), .ZN(n6997) );
  NOR2_X1 U8458 ( .A1(n12579), .A2(n12567), .ZN(n6998) );
  NOR2_X1 U8459 ( .A1(n7241), .A2(n12013), .ZN(n12018) );
  INV_X1 U8460 ( .A(n12014), .ZN(n7241) );
  INV_X1 U8461 ( .A(n10943), .ZN(n7231) );
  NAND2_X1 U8462 ( .A1(n7237), .A2(n7239), .ZN(n7238) );
  AND2_X1 U8463 ( .A1(n12192), .A2(n7571), .ZN(n7570) );
  NAND2_X1 U8464 ( .A1(n7572), .A2(n12191), .ZN(n7571) );
  INV_X1 U8465 ( .A(n7574), .ZN(n7572) );
  INV_X1 U8466 ( .A(n12191), .ZN(n7573) );
  NAND2_X1 U8467 ( .A1(n7224), .A2(n12494), .ZN(n12401) );
  NAND2_X1 U8468 ( .A1(n12456), .A2(n12375), .ZN(n12424) );
  NAND2_X1 U8469 ( .A1(n7556), .A2(n7559), .ZN(n11873) );
  AOI21_X1 U8470 ( .B1(n11679), .B2(n7560), .A(n6495), .ZN(n7559) );
  NAND2_X1 U8471 ( .A1(n11471), .A2(n7557), .ZN(n7556) );
  NAND2_X1 U8472 ( .A1(n8053), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7492) );
  NOR2_X1 U8473 ( .A1(n6534), .A2(n12013), .ZN(n7242) );
  AND2_X1 U8474 ( .A1(n12165), .A2(n12164), .ZN(n12381) );
  INV_X1 U8475 ( .A(n15413), .ZN(n11290) );
  NAND2_X1 U8476 ( .A1(n13013), .A2(n10557), .ZN(n10571) );
  NAND2_X1 U8477 ( .A1(n8405), .A2(n7495), .ZN(n8505) );
  AND2_X1 U8478 ( .A1(n12510), .A2(n8404), .ZN(n7495) );
  NAND4_X1 U8479 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(n8046)
         );
  NAND2_X1 U8480 ( .A1(n10521), .A2(n10520), .ZN(n10592) );
  NAND2_X1 U8481 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U8482 ( .A1(n13031), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6911) );
  OR2_X1 U8483 ( .A1(n13031), .A2(n10583), .ZN(n6912) );
  XNOR2_X1 U8484 ( .A(n6910), .B(n6909), .ZN(n10581) );
  XNOR2_X1 U8485 ( .A(n10608), .B(n10602), .ZN(n10606) );
  NAND2_X1 U8486 ( .A1(n10606), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6981) );
  INV_X1 U8487 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U8488 ( .A1(n10651), .A2(n10649), .ZN(n7427) );
  NAND2_X1 U8489 ( .A1(n10628), .A2(n10627), .ZN(n10648) );
  NOR2_X1 U8490 ( .A1(n10881), .A2(n6829), .ZN(n10637) );
  AND2_X1 U8491 ( .A1(n6830), .A2(n7424), .ZN(n6829) );
  AOI21_X1 U8492 ( .B1(n10616), .B2(n6831), .A(n10871), .ZN(n6830) );
  NAND2_X1 U8493 ( .A1(n10637), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U8494 ( .A1(n6914), .A2(n6913), .ZN(n11152) );
  NAND2_X1 U8495 ( .A1(n7351), .A2(n10635), .ZN(n6913) );
  INV_X1 U8496 ( .A(n7349), .ZN(n6914) );
  INV_X1 U8497 ( .A(n7352), .ZN(n7351) );
  AOI21_X1 U8498 ( .B1(n6833), .B2(n11385), .A(n11386), .ZN(n11721) );
  OR2_X1 U8499 ( .A1(n11396), .A2(n11394), .ZN(n7369) );
  OAI21_X1 U8500 ( .B1(n7405), .B2(n11724), .A(n7407), .ZN(n12545) );
  NAND2_X1 U8501 ( .A1(n12529), .A2(n12536), .ZN(n7406) );
  NAND2_X1 U8502 ( .A1(n7368), .A2(n7370), .ZN(n12532) );
  AND2_X1 U8503 ( .A1(n7368), .A2(n6585), .ZN(n12555) );
  XNOR2_X1 U8504 ( .A(n7202), .B(n12573), .ZN(n12569) );
  NAND2_X1 U8505 ( .A1(n6827), .A2(n6826), .ZN(n12609) );
  INV_X1 U8506 ( .A(n6828), .ZN(n6827) );
  INV_X1 U8507 ( .A(n12610), .ZN(n12611) );
  NAND2_X1 U8508 ( .A1(n12611), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12640) );
  OR2_X1 U8509 ( .A1(n12607), .A2(n12606), .ZN(n6920) );
  NAND2_X1 U8510 ( .A1(n6917), .A2(n6915), .ZN(n12658) );
  OR2_X1 U8511 ( .A1(n12607), .A2(n6918), .ZN(n6917) );
  OAI21_X1 U8512 ( .B1(n6919), .B2(n12657), .A(n12656), .ZN(n6916) );
  NAND2_X1 U8513 ( .A1(n7422), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7421) );
  AND2_X1 U8514 ( .A1(n12627), .A2(n12666), .ZN(n6991) );
  OAI211_X1 U8515 ( .C1(n12628), .C2(n6986), .A(n6630), .B(n6983), .ZN(n12692)
         );
  NAND2_X1 U8516 ( .A1(n6992), .A2(n6424), .ZN(n6986) );
  NOR2_X1 U8517 ( .A1(n7348), .A2(n12690), .ZN(n7347) );
  INV_X1 U8518 ( .A(n12703), .ZN(n7348) );
  NAND2_X1 U8519 ( .A1(n7130), .A2(n7944), .ZN(n8390) );
  AOI21_X1 U8520 ( .B1(n7486), .B2(n9904), .A(n7484), .ZN(n7483) );
  INV_X1 U8521 ( .A(n8501), .ZN(n7484) );
  NAND2_X1 U8522 ( .A1(n7767), .A2(n7765), .ZN(n12719) );
  INV_X1 U8523 ( .A(n7155), .ZN(n7154) );
  AOI21_X1 U8524 ( .B1(n7767), .B2(n9905), .A(n7487), .ZN(n7155) );
  INV_X1 U8525 ( .A(n7107), .ZN(n8344) );
  INV_X1 U8526 ( .A(n7131), .ZN(n8308) );
  NAND2_X1 U8527 ( .A1(n12841), .A2(n8478), .ZN(n12835) );
  INV_X1 U8528 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7937) );
  NOR2_X2 U8529 ( .A1(n8177), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U8530 ( .A1(n7935), .A2(n7934), .ZN(n8164) );
  INV_X1 U8531 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7934) );
  INV_X1 U8532 ( .A(n8148), .ZN(n7935) );
  NAND2_X1 U8533 ( .A1(n7103), .A2(n7933), .ZN(n8128) );
  INV_X1 U8534 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n7933) );
  INV_X1 U8535 ( .A(n8114), .ZN(n7103) );
  OR2_X2 U8536 ( .A1(n8128), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8148) );
  AND2_X1 U8537 ( .A1(n8457), .A2(n7464), .ZN(n7466) );
  INV_X1 U8538 ( .A(n12520), .ZN(n11289) );
  INV_X1 U8539 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U8540 ( .A1(n8455), .A2(n8454), .ZN(n10936) );
  INV_X1 U8541 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15542) );
  INV_X1 U8542 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15543) );
  NOR2_X1 U8543 ( .A1(n12062), .A2(n12142), .ZN(n12066) );
  INV_X1 U8544 ( .A(n12207), .ZN(n9907) );
  OAI211_X1 U8545 ( .C1(n12733), .C2(n7764), .A(n7762), .B(n9911), .ZN(n12139)
         );
  NAND2_X1 U8546 ( .A1(n7765), .A2(n7763), .ZN(n7762) );
  INV_X1 U8547 ( .A(n7765), .ZN(n7764) );
  INV_X1 U8548 ( .A(n9899), .ZN(n12765) );
  CLKBUF_X1 U8549 ( .A(n12776), .Z(n12778) );
  INV_X1 U8550 ( .A(n7489), .ZN(n7488) );
  AOI21_X1 U8551 ( .B1(n8483), .B2(n6503), .A(n7491), .ZN(n7489) );
  NAND2_X1 U8552 ( .A1(n12842), .A2(n12845), .ZN(n12841) );
  NAND2_X1 U8553 ( .A1(n12858), .A2(n12857), .ZN(n12856) );
  AND2_X1 U8554 ( .A1(n8241), .A2(n8240), .ZN(n12500) );
  INV_X1 U8555 ( .A(n7746), .ZN(n7745) );
  OAI21_X1 U8556 ( .B1(n7753), .B2(n7748), .A(n9881), .ZN(n7746) );
  NAND2_X1 U8557 ( .A1(n11566), .A2(n7751), .ZN(n7750) );
  AND2_X1 U8558 ( .A1(n8201), .A2(n8467), .ZN(n11800) );
  AOI21_X1 U8559 ( .B1(n6881), .B2(n6883), .A(n6880), .ZN(n6879) );
  INV_X1 U8560 ( .A(n7479), .ZN(n6881) );
  OR2_X1 U8561 ( .A1(n9944), .A2(n9936), .ZN(n10508) );
  NAND2_X1 U8562 ( .A1(n8420), .A2(n8419), .ZN(n8434) );
  NAND2_X1 U8563 ( .A1(n7920), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7918) );
  AOI21_X1 U8564 ( .B1(n7905), .B2(n7533), .A(n7532), .ZN(n7531) );
  INV_X1 U8565 ( .A(n7903), .ZN(n7533) );
  INV_X1 U8566 ( .A(n7906), .ZN(n7532) );
  NAND2_X1 U8567 ( .A1(n7922), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7924) );
  XNOR2_X1 U8568 ( .A(n8568), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U8569 ( .A1(n7524), .A2(n7526), .ZN(n7520) );
  NOR2_X1 U8570 ( .A1(n7999), .A2(n6707), .ZN(n6706) );
  INV_X1 U8571 ( .A(n7898), .ZN(n6707) );
  NAND2_X1 U8572 ( .A1(n7297), .A2(n7986), .ZN(n8449) );
  INV_X1 U8573 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7986) );
  AOI21_X1 U8574 ( .B1(n6692), .B2(n6694), .A(n6691), .ZN(n6690) );
  INV_X1 U8575 ( .A(n7894), .ZN(n6691) );
  AND2_X1 U8576 ( .A1(n7896), .A2(n7895), .ZN(n8323) );
  AND2_X1 U8577 ( .A1(n7892), .A2(n7891), .ZN(n8265) );
  INV_X1 U8578 ( .A(n8281), .ZN(n7503) );
  INV_X1 U8579 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U8580 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n6713), .ZN(n6712) );
  AND3_X2 U8581 ( .A1(n7413), .A2(n7411), .A3(n7410), .ZN(n10590) );
  OR2_X1 U8582 ( .A1(n8041), .A2(n7412), .ZN(n7411) );
  NAND2_X1 U8583 ( .A1(n13017), .A2(n7979), .ZN(n7410) );
  INV_X1 U8584 ( .A(n8058), .ZN(n7413) );
  NAND2_X1 U8585 ( .A1(n8967), .A2(n6469), .ZN(n13049) );
  NAND2_X1 U8586 ( .A1(n6855), .A2(n9146), .ZN(n13059) );
  NAND2_X1 U8587 ( .A1(n13926), .A2(n13448), .ZN(n8773) );
  OR2_X1 U8588 ( .A1(n13041), .A2(n6861), .ZN(n6860) );
  INV_X1 U8589 ( .A(n9212), .ZN(n6861) );
  NAND2_X1 U8590 ( .A1(n6652), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8858) );
  INV_X1 U8591 ( .A(n8841), .ZN(n6652) );
  INV_X1 U8592 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8857) );
  OR2_X1 U8593 ( .A1(n8858), .A2(n8857), .ZN(n8878) );
  NAND2_X1 U8594 ( .A1(n13114), .A2(n6505), .ZN(n7444) );
  NOR2_X1 U8595 ( .A1(n6527), .A2(n7445), .ZN(n7443) );
  NAND2_X1 U8596 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8818) );
  NAND2_X1 U8597 ( .A1(n6857), .A2(n9027), .ZN(n13115) );
  OAI21_X1 U8598 ( .B1(n8967), .B2(n7436), .A(n7434), .ZN(n6857) );
  AND2_X1 U8599 ( .A1(n7444), .A2(n9071), .ZN(n9102) );
  NAND2_X1 U8600 ( .A1(n8922), .A2(n11583), .ZN(n11608) );
  OAI21_X1 U8601 ( .B1(n11063), .B2(n6866), .A(n6863), .ZN(n11583) );
  INV_X1 U8602 ( .A(n11208), .ZN(n6866) );
  AND2_X1 U8603 ( .A1(n7442), .A2(n6864), .ZN(n6863) );
  AND2_X1 U8604 ( .A1(n8906), .A2(n8887), .ZN(n7442) );
  NAND2_X1 U8605 ( .A1(n9008), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U8606 ( .A1(n13115), .A2(n13116), .ZN(n13114) );
  NAND2_X1 U8607 ( .A1(n8582), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8841) );
  INV_X1 U8608 ( .A(n8820), .ZN(n8582) );
  OR2_X1 U8609 ( .A1(n8974), .A2(n8973), .ZN(n8986) );
  AND3_X1 U8610 ( .A1(n9295), .A2(n9262), .A3(n10382), .ZN(n9303) );
  NAND2_X1 U8611 ( .A1(n7603), .A2(n7601), .ZN(n7600) );
  AND2_X1 U8612 ( .A1(n6557), .A2(n7092), .ZN(n7601) );
  NOR2_X1 U8613 ( .A1(n7093), .A2(n13674), .ZN(n7092) );
  NAND2_X1 U8614 ( .A1(n13389), .A2(n6497), .ZN(n7652) );
  AND4_X1 U8615 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(n13611)
         );
  NAND2_X1 U8616 ( .A1(n8742), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7795) );
  OR2_X1 U8617 ( .A1(n8745), .A2(n8721), .ZN(n8723) );
  AND2_X1 U8618 ( .A1(n8722), .A2(n6576), .ZN(n7344) );
  NAND2_X1 U8619 ( .A1(n10215), .A2(n10214), .ZN(n13470) );
  NAND2_X1 U8620 ( .A1(n6816), .A2(n15276), .ZN(n15275) );
  OR2_X1 U8621 ( .A1(n15278), .A2(n15277), .ZN(n6816) );
  OR2_X1 U8622 ( .A1(n8853), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8871) );
  OR2_X1 U8623 ( .A1(n10702), .A2(n10703), .ZN(n10704) );
  NOR2_X1 U8624 ( .A1(n15298), .A2(n15299), .ZN(n15297) );
  NOR2_X1 U8625 ( .A1(n15297), .A2(n6794), .ZN(n11499) );
  OR2_X1 U8626 ( .A1(n10958), .A2(n10959), .ZN(n6794) );
  NAND2_X1 U8627 ( .A1(n6665), .A2(n6664), .ZN(n13537) );
  INV_X1 U8628 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13160) );
  INV_X1 U8629 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n13075) );
  NOR2_X1 U8630 ( .A1(n7603), .A2(n13920), .ZN(n6669) );
  OAI21_X1 U8631 ( .B1(n13694), .B2(n7800), .A(n7798), .ZN(n13658) );
  INV_X1 U8632 ( .A(n13639), .ZN(n7799) );
  NAND2_X1 U8633 ( .A1(n13658), .A2(n13657), .ZN(n6731) );
  AND2_X1 U8634 ( .A1(n9288), .A2(n9275), .ZN(n13654) );
  NOR2_X1 U8635 ( .A1(n13657), .A2(n7714), .ZN(n7713) );
  INV_X1 U8636 ( .A(n13591), .ZN(n7714) );
  NAND2_X1 U8637 ( .A1(n13694), .A2(n13639), .ZN(n7802) );
  AND2_X1 U8638 ( .A1(n9200), .A2(n9221), .ZN(n13690) );
  NAND2_X1 U8639 ( .A1(n13768), .A2(n6431), .ZN(n13724) );
  XNOR2_X1 U8640 ( .A(n13972), .B(n13741), .ZN(n13719) );
  NAND2_X1 U8641 ( .A1(n13768), .A2(n7555), .ZN(n13732) );
  AND2_X1 U8642 ( .A1(n13768), .A2(n13754), .ZN(n13749) );
  AND2_X1 U8643 ( .A1(n7817), .A2(n7815), .ZN(n13748) );
  NAND2_X1 U8644 ( .A1(n6653), .A2(n8583), .ZN(n9137) );
  NOR2_X1 U8645 ( .A1(n14004), .A2(n7550), .ZN(n7549) );
  CLKBUF_X1 U8646 ( .A(n13794), .Z(n13795) );
  NAND2_X1 U8647 ( .A1(n7317), .A2(n7312), .ZN(n7311) );
  INV_X1 U8648 ( .A(n7318), .ZN(n7317) );
  OR2_X1 U8649 ( .A1(n13865), .A2(n7320), .ZN(n7312) );
  AND2_X1 U8650 ( .A1(n9038), .A2(n9011), .ZN(n13854) );
  NAND2_X1 U8651 ( .A1(n13872), .A2(n6429), .ZN(n13851) );
  NAND2_X1 U8652 ( .A1(n13912), .A2(n13884), .ZN(n7059) );
  INV_X1 U8653 ( .A(n7791), .ZN(n7790) );
  AOI21_X1 U8654 ( .B1(n7791), .B2(n7789), .A(n6538), .ZN(n7788) );
  NOR2_X1 U8655 ( .A1(n13612), .A2(n7792), .ZN(n7791) );
  NAND2_X1 U8656 ( .A1(n11814), .A2(n7543), .ZN(n13924) );
  NAND2_X1 U8657 ( .A1(n11814), .A2(n13609), .ZN(n13927) );
  NOR2_X1 U8658 ( .A1(n11654), .A2(n6418), .ZN(n11085) );
  NAND2_X1 U8659 ( .A1(n11261), .A2(n10483), .ZN(n11031) );
  XNOR2_X1 U8660 ( .A(n13449), .B(n15361), .ZN(n13396) );
  NAND2_X1 U8661 ( .A1(n11260), .A2(n13396), .ZN(n11261) );
  INV_X1 U8662 ( .A(n13946), .ZN(n7270) );
  INV_X1 U8663 ( .A(n13656), .ZN(n13950) );
  AND2_X1 U8664 ( .A1(n15371), .A2(n10909), .ZN(n15381) );
  INV_X1 U8665 ( .A(n9235), .ZN(n9248) );
  NOR2_X1 U8666 ( .A1(n6868), .A2(n6870), .ZN(n6867) );
  OR2_X1 U8667 ( .A1(n8798), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U8668 ( .A1(n8714), .A2(n8627), .ZN(n8727) );
  NAND2_X1 U8669 ( .A1(n9497), .A2(n6903), .ZN(n9526) );
  OR2_X1 U8670 ( .A1(n14109), .A2(n14110), .ZN(n14107) );
  OR2_X2 U8671 ( .A1(n12273), .A2(n15216), .ZN(n11341) );
  OR2_X1 U8672 ( .A1(n9537), .A2(n9536), .ZN(n9552) );
  INV_X1 U8673 ( .A(n12111), .ZN(n7011) );
  INV_X1 U8674 ( .A(n12124), .ZN(n7692) );
  NAND2_X1 U8675 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9390) );
  INV_X1 U8676 ( .A(n10856), .ZN(n10783) );
  NAND2_X1 U8677 ( .A1(n9497), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U8678 ( .A1(n10745), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10747) );
  OR2_X1 U8679 ( .A1(n12273), .A2(n10837), .ZN(n10746) );
  OR2_X1 U8680 ( .A1(n9564), .A2(n9563), .ZN(n9577) );
  NAND2_X1 U8681 ( .A1(n9550), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9564) );
  INV_X1 U8682 ( .A(n9552), .ZN(n9550) );
  OR2_X1 U8683 ( .A1(n14432), .A2(n9804), .ZN(n11368) );
  AND4_X1 U8684 ( .A1(n9369), .A2(n9368), .A3(n9367), .A4(n9366), .ZN(n11343)
         );
  NAND2_X1 U8685 ( .A1(n14500), .A2(n14501), .ZN(n14517) );
  NAND2_X1 U8686 ( .A1(n9396), .A2(n9409), .ZN(n9411) );
  OAI21_X1 U8687 ( .B1(n9479), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9492) );
  NOR2_X1 U8688 ( .A1(n14580), .A2(n6845), .ZN(n14577) );
  OR2_X1 U8689 ( .A1(n14578), .A2(n14579), .ZN(n6845) );
  NOR2_X1 U8690 ( .A1(n14577), .A2(n6844), .ZN(n11239) );
  AND2_X1 U8691 ( .A1(n14586), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U8692 ( .A1(n11239), .A2(n11240), .ZN(n11616) );
  INV_X1 U8693 ( .A(n14652), .ZN(n14656) );
  NAND2_X1 U8694 ( .A1(n9975), .A2(n9976), .ZN(n14670) );
  NAND2_X1 U8695 ( .A1(n9669), .A2(n7661), .ZN(n7665) );
  NOR2_X1 U8696 ( .A1(n9679), .A2(n7662), .ZN(n7661) );
  INV_X1 U8697 ( .A(n9668), .ZN(n7662) );
  OR2_X1 U8698 ( .A1(n9778), .A2(n9777), .ZN(n7783) );
  AND2_X1 U8699 ( .A1(n9779), .A2(n7785), .ZN(n7784) );
  NAND2_X1 U8700 ( .A1(n7180), .A2(n9776), .ZN(n7176) );
  AND2_X1 U8701 ( .A1(n9672), .A2(n9657), .ZN(n14698) );
  AND2_X1 U8702 ( .A1(n9631), .A2(n9630), .ZN(n14743) );
  AND2_X1 U8703 ( .A1(n14785), .A2(n14790), .ZN(n14770) );
  NAND2_X1 U8704 ( .A1(n6906), .A2(n6905), .ZN(n9607) );
  NOR2_X1 U8705 ( .A1(n14182), .A2(n9594), .ZN(n6905) );
  INV_X1 U8706 ( .A(n6906), .ZN(n9595) );
  AOI21_X1 U8707 ( .B1(n7680), .B2(n7677), .A(n6443), .ZN(n7675) );
  INV_X1 U8708 ( .A(n7677), .ZN(n7676) );
  NAND2_X1 U8709 ( .A1(n14900), .A2(n7718), .ZN(n14859) );
  NOR2_X1 U8710 ( .A1(n14951), .A2(n15065), .ZN(n7732) );
  INV_X1 U8711 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U8712 ( .A1(n6899), .A2(n6898), .ZN(n9499) );
  NOR2_X1 U8713 ( .A1(n10456), .A2(n9482), .ZN(n6898) );
  INV_X1 U8714 ( .A(n9483), .ZN(n6899) );
  NAND2_X1 U8715 ( .A1(n6901), .A2(n6508), .ZN(n9463) );
  INV_X1 U8716 ( .A(n9448), .ZN(n6901) );
  NAND2_X1 U8717 ( .A1(n6900), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9483) );
  INV_X1 U8718 ( .A(n9463), .ZN(n6900) );
  NAND2_X1 U8719 ( .A1(n11827), .A2(n9454), .ZN(n11855) );
  NAND2_X1 U8720 ( .A1(n11704), .A2(n9439), .ZN(n11828) );
  NAND2_X1 U8721 ( .A1(n11828), .A2(n14447), .ZN(n11827) );
  NAND2_X1 U8722 ( .A1(n6613), .A2(n7770), .ZN(n11709) );
  NOR2_X1 U8723 ( .A1(n9751), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U8724 ( .A1(n9754), .A2(n9753), .ZN(n7200) );
  AND2_X1 U8725 ( .A1(n7770), .A2(n9750), .ZN(n11320) );
  NOR2_X1 U8726 ( .A1(n14289), .A2(n15215), .ZN(n7720) );
  NAND2_X1 U8727 ( .A1(n6902), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9403) );
  NOR2_X1 U8728 ( .A1(n7723), .A2(n15215), .ZN(n11326) );
  NOR2_X1 U8729 ( .A1(n15215), .A2(n15245), .ZN(n11307) );
  AND2_X1 U8730 ( .A1(n11298), .A2(n9401), .ZN(n14442) );
  NAND2_X1 U8731 ( .A1(n9374), .A2(n14272), .ZN(n11119) );
  OR2_X1 U8732 ( .A1(n9735), .A2(n10751), .ZN(n14658) );
  NAND2_X1 U8733 ( .A1(n10837), .A2(n14260), .ZN(n11045) );
  INV_X1 U8734 ( .A(n14935), .ZN(n14880) );
  INV_X1 U8735 ( .A(n14933), .ZN(n14897) );
  AND2_X1 U8736 ( .A1(n14652), .A2(n15251), .ZN(n9986) );
  AND2_X1 U8737 ( .A1(n14749), .A2(n14714), .ZN(n14735) );
  AND2_X1 U8738 ( .A1(n14756), .A2(n15216), .ZN(n15004) );
  NOR2_X1 U8739 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7787) );
  XNOR2_X1 U8740 ( .A(n9840), .B(n9834), .ZN(n13367) );
  XNOR2_X1 U8741 ( .A(n9267), .B(SI_27_), .ZN(n12160) );
  INV_X1 U8742 ( .A(n9710), .ZN(n7101) );
  NOR2_X1 U8743 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7100) );
  NAND2_X1 U8744 ( .A1(n9175), .A2(n9174), .ZN(n9192) );
  INV_X1 U8745 ( .A(n7081), .ZN(n9717) );
  NAND2_X1 U8746 ( .A1(n7264), .A2(n6515), .ZN(n9106) );
  OR2_X1 U8747 ( .A1(n8685), .A2(SI_20_), .ZN(n7263) );
  NAND2_X1 U8748 ( .A1(n9691), .A2(n9690), .ZN(n9698) );
  NAND2_X1 U8749 ( .A1(n8676), .A2(n8675), .ZN(n9030) );
  OAI21_X1 U8750 ( .B1(n8949), .B2(n8950), .A(n8948), .ZN(n8952) );
  INV_X1 U8751 ( .A(n6738), .ZN(n8948) );
  XNOR2_X1 U8752 ( .A(n8870), .B(n8869), .ZN(n10144) );
  NAND2_X1 U8753 ( .A1(n7273), .A2(n8647), .ZN(n8870) );
  NAND2_X1 U8754 ( .A1(n8852), .A2(n8645), .ZN(n7273) );
  OR2_X1 U8755 ( .A1(n9411), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U8756 ( .A(n8832), .B(n8833), .ZN(n10096) );
  OAI21_X1 U8757 ( .B1(n8714), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n7113), .ZN(
        n8760) );
  NAND2_X1 U8758 ( .A1(n8714), .A2(n10085), .ZN(n7113) );
  NAND2_X1 U8759 ( .A1(n9346), .A2(n8727), .ZN(n8713) );
  INV_X1 U8760 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7243) );
  XNOR2_X1 U8761 ( .A(n10033), .B(n10042), .ZN(n10037) );
  XNOR2_X1 U8762 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n10033) );
  NAND2_X1 U8763 ( .A1(n10170), .A2(n10169), .ZN(n10404) );
  OR2_X1 U8764 ( .A1(n10167), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10170) );
  INV_X1 U8765 ( .A(n11247), .ZN(n7070) );
  NOR2_X1 U8766 ( .A1(n7070), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7067) );
  OR2_X1 U8767 ( .A1(n11163), .A2(n11162), .ZN(n11164) );
  INV_X1 U8768 ( .A(n7254), .ZN(n7251) );
  NAND2_X1 U8769 ( .A1(n15110), .A2(n15111), .ZN(n7254) );
  INV_X1 U8770 ( .A(n15110), .ZN(n7253) );
  OR2_X1 U8771 ( .A1(n15127), .A2(n15126), .ZN(n15129) );
  NAND2_X1 U8772 ( .A1(n11471), .A2(n11470), .ZN(n11678) );
  NAND2_X1 U8773 ( .A1(n12018), .A2(n12017), .ZN(n12165) );
  NAND2_X1 U8774 ( .A1(n7238), .A2(n7235), .ZN(n10946) );
  NOR2_X1 U8775 ( .A1(n12361), .A2(n7563), .ZN(n7562) );
  INV_X1 U8776 ( .A(n7565), .ZN(n7563) );
  NAND2_X1 U8777 ( .A1(n7564), .A2(n7565), .ZN(n12362) );
  NOR2_X1 U8778 ( .A1(n7586), .A2(n7583), .ZN(n7579) );
  NAND2_X1 U8779 ( .A1(n7581), .A2(n12208), .ZN(n7580) );
  NAND2_X1 U8780 ( .A1(n11680), .A2(n11679), .ZN(n11870) );
  NAND2_X1 U8781 ( .A1(n11678), .A2(n11677), .ZN(n11680) );
  INV_X1 U8782 ( .A(n12788), .ZN(n12375) );
  NAND2_X1 U8783 ( .A1(n12437), .A2(n12188), .ZN(n12371) );
  AND4_X1 U8784 ( .A1(n8181), .A2(n8180), .A3(n8179), .A4(n8178), .ZN(n12386)
         );
  CLKBUF_X1 U8785 ( .A(n12401), .Z(n12402) );
  AOI21_X1 U8786 ( .B1(n12748), .B2(n8395), .A(n7978), .ZN(n12432) );
  AND4_X1 U8787 ( .A1(n8197), .A2(n8196), .A3(n8195), .A4(n8194), .ZN(n12450)
         );
  INV_X1 U8788 ( .A(n12779), .ZN(n12459) );
  AND2_X1 U8789 ( .A1(n7568), .A2(n7569), .ZN(n12476) );
  NAND2_X1 U8790 ( .A1(n12402), .A2(n12182), .ZN(n7568) );
  NAND2_X1 U8791 ( .A1(n7039), .A2(n7038), .ZN(n7037) );
  INV_X1 U8792 ( .A(n7034), .ZN(n7033) );
  OAI21_X1 U8793 ( .B1(n7036), .B2(n11019), .A(n7035), .ZN(n7034) );
  NOR2_X1 U8794 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  NOR2_X1 U8795 ( .A1(n11527), .A2(n9938), .ZN(n7504) );
  XNOR2_X1 U8796 ( .A(n7132), .B(n6417), .ZN(n8554) );
  OR2_X1 U8797 ( .A1(n8524), .A2(n7474), .ZN(n8578) );
  NAND2_X1 U8798 ( .A1(n8352), .A2(n8351), .ZN(n12798) );
  OAI211_X1 U8799 ( .C1(n8409), .C2(n12999), .A(n8256), .B(n8255), .ZN(n12860)
         );
  INV_X1 U8800 ( .A(n12405), .ZN(n12847) );
  INV_X1 U8801 ( .A(n12386), .ZN(n12515) );
  NAND4_X1 U8802 ( .A1(n8097), .A2(n8096), .A3(n8095), .A4(n8094), .ZN(n12519)
         );
  NAND2_X1 U8803 ( .A1(n8051), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8026) );
  XNOR2_X1 U8804 ( .A(n10590), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10516) );
  OAI22_X1 U8805 ( .A1(n10582), .A2(n10581), .B1(n6909), .B2(n6910), .ZN(
        n10604) );
  NAND2_X1 U8806 ( .A1(n7433), .A2(n10729), .ZN(n10587) );
  INV_X1 U8807 ( .A(n10631), .ZN(n10632) );
  INV_X1 U8808 ( .A(n7357), .ZN(n10879) );
  AOI21_X1 U8809 ( .B1(n10635), .B2(n7358), .A(n7089), .ZN(n7357) );
  INV_X1 U8810 ( .A(n7363), .ZN(n7358) );
  NAND2_X1 U8811 ( .A1(n6627), .A2(n7354), .ZN(n11147) );
  NOR2_X1 U8812 ( .A1(n11384), .A2(n7419), .ZN(n11139) );
  AOI21_X1 U8813 ( .B1(n11396), .B2(n11395), .A(n11394), .ZN(n11727) );
  NAND2_X1 U8814 ( .A1(n11382), .A2(n11381), .ZN(n11718) );
  NAND2_X1 U8815 ( .A1(n12527), .A2(n12526), .ZN(n12562) );
  NOR2_X1 U8816 ( .A1(n12549), .A2(n12550), .ZN(n12593) );
  NAND2_X1 U8817 ( .A1(n7001), .A2(n7000), .ZN(n12572) );
  NAND2_X1 U8818 ( .A1(n7201), .A2(n12573), .ZN(n7000) );
  OR2_X1 U8819 ( .A1(n12569), .A2(n12568), .ZN(n7001) );
  NAND2_X1 U8820 ( .A1(n12572), .A2(n12578), .ZN(n12613) );
  AOI21_X1 U8821 ( .B1(n12639), .B2(n7404), .A(n6635), .ZN(n7403) );
  XNOR2_X1 U8822 ( .A(n12703), .B(n12702), .ZN(n12668) );
  NOR2_X1 U8823 ( .A1(n12668), .A2(n12669), .ZN(n12701) );
  OAI21_X1 U8824 ( .B1(n13026), .B2(n8389), .A(n8388), .ZN(n12715) );
  NAND2_X1 U8825 ( .A1(n7146), .A2(n7148), .ZN(n12804) );
  NAND2_X1 U8826 ( .A1(n7147), .A2(n7151), .ZN(n7146) );
  NAND2_X1 U8827 ( .A1(n12032), .A2(n9886), .ZN(n12047) );
  NAND2_X1 U8828 ( .A1(n8236), .A2(n8235), .ZN(n12942) );
  NAND2_X1 U8829 ( .A1(n8473), .A2(n8472), .ZN(n12043) );
  NAND2_X1 U8830 ( .A1(n8210), .A2(n8209), .ZN(n12868) );
  NAND2_X1 U8831 ( .A1(n12896), .A2(n11003), .ZN(n12876) );
  NAND2_X1 U8832 ( .A1(n7481), .A2(n7479), .ZN(n6885) );
  NAND2_X1 U8833 ( .A1(n7481), .A2(n8463), .ZN(n11564) );
  INV_X1 U8834 ( .A(n11469), .ZN(n15419) );
  NAND2_X1 U8835 ( .A1(n7468), .A2(n8456), .ZN(n11092) );
  NAND2_X1 U8836 ( .A1(n10981), .A2(n10982), .ZN(n7468) );
  NAND2_X2 U8837 ( .A1(n10696), .A2(n12891), .ZN(n12896) );
  AND2_X1 U8838 ( .A1(n10698), .A2(n10697), .ZN(n12855) );
  AND2_X1 U8839 ( .A1(n15589), .A2(n15423), .ZN(n12939) );
  INV_X1 U8840 ( .A(n12939), .ZN(n12905) );
  AND2_X2 U8841 ( .A1(n10694), .A2(n9941), .ZN(n15589) );
  INV_X1 U8842 ( .A(n8508), .ZN(n12950) );
  INV_X1 U8843 ( .A(n8526), .ZN(n12068) );
  NAND2_X1 U8844 ( .A1(n8405), .A2(n8404), .ZN(n7496) );
  NAND2_X1 U8845 ( .A1(n9906), .A2(n15423), .ZN(n7134) );
  AOI21_X1 U8846 ( .B1(n6651), .B2(n12883), .A(n6649), .ZN(n12952) );
  INV_X1 U8847 ( .A(n6650), .ZN(n6649) );
  XNOR2_X1 U8848 ( .A(n12733), .B(n12734), .ZN(n6651) );
  AOI22_X1 U8849 ( .A1(n12735), .A2(n12879), .B1(n12880), .B2(n12752), .ZN(
        n6650) );
  AND2_X1 U8850 ( .A1(n7139), .A2(n7140), .ZN(n12743) );
  NAND2_X1 U8851 ( .A1(n7973), .A2(n7972), .ZN(n12961) );
  OR2_X1 U8852 ( .A1(n12070), .A2(n8389), .ZN(n7973) );
  NAND2_X1 U8853 ( .A1(n12754), .A2(n8495), .ZN(n12740) );
  OR2_X1 U8854 ( .A1(n12912), .A2(n12945), .ZN(n6671) );
  NAND2_X1 U8855 ( .A1(n8361), .A2(n8360), .ZN(n12968) );
  NAND2_X1 U8856 ( .A1(n6701), .A2(n6622), .ZN(n6698) );
  NAND2_X1 U8857 ( .A1(n8002), .A2(n8001), .ZN(n12974) );
  NAND2_X1 U8858 ( .A1(n8343), .A2(n8342), .ZN(n12980) );
  OR2_X1 U8859 ( .A1(n11181), .A2(n8389), .ZN(n8343) );
  NAND2_X1 U8860 ( .A1(n8328), .A2(n8327), .ZN(n12986) );
  OR2_X1 U8861 ( .A1(n11133), .A2(n8389), .ZN(n8328) );
  NAND2_X1 U8862 ( .A1(n8274), .A2(n8273), .ZN(n12993) );
  AND2_X1 U8863 ( .A1(n7152), .A2(n6488), .ZN(n12824) );
  NAND2_X1 U8864 ( .A1(n7152), .A2(n7151), .ZN(n12823) );
  NAND2_X1 U8865 ( .A1(n8251), .A2(n8250), .ZN(n13000) );
  NAND2_X1 U8866 ( .A1(n7477), .A2(n8470), .ZN(n12029) );
  OR2_X1 U8867 ( .A1(n15429), .A2(n15418), .ZN(n12949) );
  AND2_X1 U8868 ( .A1(n10558), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13013) );
  INV_X1 U8869 ( .A(n9917), .ZN(n13040) );
  MUX2_X1 U8870 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8565), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8566) );
  NAND2_X1 U8871 ( .A1(n7527), .A2(n7528), .ZN(n7988) );
  NAND2_X1 U8872 ( .A1(n7901), .A2(n6623), .ZN(n7528) );
  NAND2_X1 U8873 ( .A1(n7523), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7527) );
  INV_X1 U8874 ( .A(n6702), .ZN(n6701) );
  OAI21_X1 U8875 ( .B1(n6706), .B2(n6622), .A(n6703), .ZN(n6702) );
  NAND2_X1 U8876 ( .A1(n8358), .A2(n6704), .ZN(n6703) );
  INV_X1 U8877 ( .A(n9938), .ZN(n11134) );
  INV_X1 U8878 ( .A(SI_19_), .ZN(n12158) );
  OAI21_X1 U8879 ( .B1(n7499), .B2(n6694), .A(n6692), .ZN(n8304) );
  NAND2_X1 U8880 ( .A1(n8268), .A2(n7892), .ZN(n8302) );
  NAND2_X1 U8881 ( .A1(n8282), .A2(n8281), .ZN(n8284) );
  NAND2_X1 U8882 ( .A1(n7888), .A2(n7887), .ZN(n8282) );
  INV_X1 U8883 ( .A(SI_16_), .ZN(n10546) );
  INV_X1 U8884 ( .A(SI_15_), .ZN(n10421) );
  NAND2_X1 U8885 ( .A1(n7982), .A2(n6430), .ZN(n8247) );
  OAI21_X1 U8886 ( .B1(n7877), .B2(n7537), .A(n7535), .ZN(n8220) );
  INV_X1 U8887 ( .A(SI_13_), .ZN(n10389) );
  INV_X1 U8888 ( .A(SI_10_), .ZN(n10128) );
  NAND2_X1 U8889 ( .A1(n6711), .A2(n7511), .ZN(n8159) );
  NAND2_X1 U8890 ( .A1(n8109), .A2(n7512), .ZN(n6711) );
  OAI21_X1 U8891 ( .B1(n8109), .B2(n7516), .A(n7514), .ZN(n8138) );
  OAI21_X1 U8892 ( .B1(n8109), .B2(n7518), .A(n7871), .ZN(n8123) );
  XNOR2_X1 U8893 ( .A(n8101), .B(n8100), .ZN(n10655) );
  NAND2_X1 U8894 ( .A1(n7510), .A2(n7866), .ZN(n8099) );
  NAND2_X1 U8895 ( .A1(n8080), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U8896 ( .A1(n6685), .A2(n7862), .ZN(n8016) );
  NAND2_X1 U8897 ( .A1(n7861), .A2(n6686), .ZN(n6685) );
  INV_X1 U8898 ( .A(n6681), .ZN(n6686) );
  NAND2_X1 U8899 ( .A1(n7861), .A2(n7860), .ZN(n8061) );
  NAND2_X1 U8900 ( .A1(n7003), .A2(n7002), .ZN(n8059) );
  NAND2_X1 U8901 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8014), .ZN(n7002) );
  OAI21_X1 U8902 ( .B1(n8058), .B2(n13017), .A(P3_IR_REG_3__SCAN_IN), .ZN(
        n7003) );
  NAND2_X1 U8903 ( .A1(n8020), .A2(n7858), .ZN(n8043) );
  INV_X1 U8904 ( .A(n7857), .ZN(n8019) );
  NAND3_X1 U8905 ( .A1(n7440), .A2(n7438), .A3(n11102), .ZN(n11106) );
  NAND2_X1 U8906 ( .A1(n8831), .A2(n7439), .ZN(n7438) );
  NAND2_X1 U8907 ( .A1(n7441), .A2(n8795), .ZN(n7439) );
  NAND2_X1 U8908 ( .A1(n8967), .A2(n8966), .ZN(n13051) );
  INV_X1 U8909 ( .A(n13174), .ZN(n13183) );
  NAND2_X1 U8910 ( .A1(n11214), .A2(n8887), .ZN(n11584) );
  OAI21_X1 U8911 ( .B1(n7540), .B2(n7541), .A(n10193), .ZN(n7539) );
  AND2_X1 U8912 ( .A1(n10065), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U8913 ( .A1(n10236), .A2(n6408), .ZN(n7062) );
  NAND2_X1 U8914 ( .A1(n10678), .A2(n8795), .ZN(n10826) );
  INV_X1 U8915 ( .A(n7448), .ZN(n13127) );
  NAND2_X1 U8916 ( .A1(n6862), .A2(n11208), .ZN(n11214) );
  NAND2_X1 U8917 ( .A1(n11063), .A2(n8868), .ZN(n6862) );
  NAND2_X1 U8918 ( .A1(n13114), .A2(n9051), .ZN(n13159) );
  INV_X1 U8919 ( .A(n13187), .ZN(n13170) );
  INV_X1 U8920 ( .A(n13194), .ZN(n13173) );
  NAND2_X1 U8921 ( .A1(n10397), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13187) );
  INV_X1 U8922 ( .A(n13668), .ZN(n13594) );
  NAND2_X1 U8923 ( .A1(n8609), .A2(n8608), .ZN(n13584) );
  NAND2_X1 U8924 ( .A1(n9145), .A2(n9144), .ZN(n13631) );
  NAND2_X1 U8925 ( .A1(n9085), .A2(n9084), .ZN(n13798) );
  INV_X1 U8926 ( .A(n13608), .ZN(n13566) );
  OR2_X2 U8927 ( .A1(n10197), .A2(P2_U3088), .ZN(n13451) );
  NOR2_X1 U8928 ( .A1(n10534), .A2(n10535), .ZN(n13457) );
  NAND2_X1 U8929 ( .A1(n15285), .A2(n15286), .ZN(n15284) );
  OAI21_X1 U8930 ( .B1(n6812), .B2(n6811), .A(n10192), .ZN(n13506) );
  NAND2_X1 U8931 ( .A1(n6814), .A2(n6637), .ZN(n6811) );
  NAND2_X1 U8932 ( .A1(n10225), .A2(n10224), .ZN(n10306) );
  AOI21_X1 U8933 ( .B1(n13506), .B2(n10202), .A(n10201), .ZN(n10280) );
  OR2_X1 U8934 ( .A1(n10289), .A2(n10288), .ZN(n10665) );
  INV_X1 U8935 ( .A(n6789), .ZN(n10706) );
  OR2_X1 U8936 ( .A1(n10972), .A2(n10971), .ZN(n11506) );
  XNOR2_X1 U8937 ( .A(n11508), .B(n15312), .ZN(n15317) );
  AND2_X1 U8938 ( .A1(n6805), .A2(n7123), .ZN(n11691) );
  NAND2_X1 U8939 ( .A1(n11666), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8940 ( .A1(n6804), .A2(n6809), .ZN(n13522) );
  OAI21_X1 U8941 ( .B1(n11666), .B2(n7122), .A(n6806), .ZN(n6804) );
  NOR2_X1 U8942 ( .A1(n6796), .A2(n11690), .ZN(n6806) );
  OR2_X1 U8943 ( .A1(n10210), .A2(n13434), .ZN(n15294) );
  INV_X1 U8944 ( .A(n13386), .ZN(n13942) );
  INV_X1 U8945 ( .A(n13544), .ZN(n13945) );
  AND2_X1 U8946 ( .A1(n13344), .A2(n13343), .ZN(n13604) );
  NAND2_X1 U8947 ( .A1(n6773), .A2(n6776), .ZN(n13956) );
  AND2_X1 U8948 ( .A1(n9195), .A2(n9194), .ZN(n13692) );
  AOI21_X1 U8949 ( .B1(n13686), .B2(n13905), .A(n13685), .ZN(n13964) );
  NAND2_X1 U8950 ( .A1(n13684), .A2(n13683), .ZN(n13685) );
  OAI21_X1 U8951 ( .B1(n7711), .B2(n7328), .A(n7326), .ZN(n13698) );
  NAND2_X1 U8952 ( .A1(n7708), .A2(n13581), .ZN(n13756) );
  NAND2_X1 U8953 ( .A1(n7820), .A2(n6457), .ZN(n13763) );
  NAND2_X1 U8954 ( .A1(n7827), .A2(n7823), .ZN(n7820) );
  NAND2_X1 U8955 ( .A1(n7712), .A2(n13577), .ZN(n13778) );
  NAND2_X1 U8956 ( .A1(n7837), .A2(n7826), .ZN(n13775) );
  NAND2_X1 U8957 ( .A1(n7827), .A2(n6473), .ZN(n7826) );
  INV_X1 U8958 ( .A(n13997), .ZN(n13809) );
  NAND2_X1 U8959 ( .A1(n13834), .A2(n13625), .ZN(n13820) );
  NAND2_X1 U8960 ( .A1(n7308), .A2(n7309), .ZN(n13815) );
  AND2_X1 U8961 ( .A1(n7310), .A2(n7313), .ZN(n7308) );
  OAI21_X1 U8962 ( .B1(n13616), .B2(n6757), .A(n6756), .ZN(n13836) );
  INV_X1 U8963 ( .A(n7806), .ZN(n6757) );
  AOI21_X1 U8964 ( .B1(n7806), .B2(n7804), .A(n6761), .ZN(n6756) );
  NAND2_X1 U8965 ( .A1(n7809), .A2(n7806), .ZN(n13858) );
  NAND2_X1 U8966 ( .A1(n13616), .A2(n7803), .ZN(n7809) );
  AOI21_X1 U8967 ( .B1(n13865), .B2(n13866), .A(n7320), .ZN(n13847) );
  NAND2_X1 U8968 ( .A1(n7810), .A2(n13618), .ZN(n13863) );
  NAND2_X1 U8969 ( .A1(n13616), .A2(n7813), .ZN(n7810) );
  NAND2_X1 U8970 ( .A1(n7793), .A2(n13610), .ZN(n13934) );
  NAND2_X1 U8971 ( .A1(n13607), .A2(n13606), .ZN(n7793) );
  INV_X1 U8972 ( .A(n14036), .ZN(n13932) );
  NAND2_X1 U8973 ( .A1(n11747), .A2(n13563), .ZN(n11819) );
  NAND2_X1 U8974 ( .A1(n11786), .A2(n11746), .ZN(n11747) );
  NAND2_X1 U8975 ( .A1(n7335), .A2(n7336), .ZN(n11492) );
  NAND2_X1 U8976 ( .A1(n7339), .A2(n11081), .ZN(n11414) );
  NAND2_X1 U8977 ( .A1(n7702), .A2(n7700), .ZN(n11082) );
  NAND2_X1 U8978 ( .A1(n15359), .A2(n9304), .ZN(n13837) );
  AND2_X1 U8979 ( .A1(n6775), .A2(n6776), .ZN(n6772) );
  AND2_X1 U8980 ( .A1(n13958), .A2(n6577), .ZN(n6775) );
  INV_X1 U8981 ( .A(n15359), .ZN(n15356) );
  CLKBUF_X1 U8982 ( .A(n15338), .Z(n15354) );
  NAND2_X1 U8983 ( .A1(n14085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8600) );
  NOR2_X1 U8984 ( .A1(n7120), .A2(n7119), .ZN(n7118) );
  NOR2_X1 U8985 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7119) );
  CLKBUF_X1 U8986 ( .A(n10199), .Z(n13434) );
  XNOR2_X1 U8987 ( .A(n9234), .B(n9233), .ZN(n11785) );
  INV_X1 U8988 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9233) );
  OAI21_X1 U8989 ( .B1(n9238), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9234) );
  XNOR2_X1 U8990 ( .A(n9240), .B(n9239), .ZN(n11572) );
  INV_X1 U8991 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U8992 ( .A1(n9246), .A2(n8614), .ZN(n13373) );
  AOI21_X1 U8993 ( .B1(n8613), .B2(P2_IR_REG_22__SCAN_IN), .A(n8612), .ZN(
        n8614) );
  AND2_X1 U8994 ( .A1(n8763), .A2(n8611), .ZN(n8612) );
  NAND2_X1 U8995 ( .A1(n7343), .A2(n8610), .ZN(n8615) );
  INV_X1 U8996 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n15545) );
  INV_X1 U8997 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10241) );
  OR2_X1 U8998 ( .A1(n7457), .A2(n7454), .ZN(n8953) );
  NAND2_X1 U8999 ( .A1(n8596), .A2(n7458), .ZN(n7454) );
  INV_X1 U9000 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10237) );
  INV_X1 U9001 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10185) );
  XNOR2_X1 U9002 ( .A(n8892), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10714) );
  INV_X1 U9003 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10147) );
  INV_X1 U9004 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10112) );
  INV_X1 U9005 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10098) );
  INV_X1 U9006 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10083) );
  INV_X1 U9007 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10087) );
  INV_X1 U9008 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10085) );
  AND4_X1 U9009 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(n11826)
         );
  AOI21_X1 U9010 ( .B1(n7688), .B2(n7690), .A(n6541), .ZN(n7687) );
  NAND2_X1 U9011 ( .A1(n7694), .A2(n6433), .ZN(n12080) );
  NAND2_X1 U9012 ( .A1(n7693), .A2(n6605), .ZN(n12003) );
  NAND2_X1 U9013 ( .A1(n10111), .A2(n9845), .ZN(n7160) );
  OAI22_X1 U9014 ( .A1(n14258), .A2(n6401), .B1(n14260), .B2(n12273), .ZN(
        n10742) );
  NAND2_X1 U9015 ( .A1(n14202), .A2(n12090), .ZN(n14143) );
  NAND2_X1 U9016 ( .A1(n14202), .A2(n7697), .ZN(n14144) );
  INV_X1 U9017 ( .A(n6604), .ZN(n7008) );
  NAND2_X1 U9018 ( .A1(n7691), .A2(n6604), .ZN(n7009) );
  AOI21_X1 U9019 ( .B1(n7691), .B2(n7011), .A(n6529), .ZN(n7010) );
  NAND2_X1 U9020 ( .A1(n11350), .A2(n11349), .ZN(n11351) );
  OR2_X1 U9021 ( .A1(n12273), .A2(n15237), .ZN(n11349) );
  AND2_X1 U9022 ( .A1(n7693), .A2(n11901), .ZN(n11997) );
  NOR2_X1 U9023 ( .A1(n14198), .A2(n14933), .ZN(n14218) );
  NAND2_X1 U9024 ( .A1(n14177), .A2(n14179), .ZN(n14178) );
  INV_X1 U9025 ( .A(n7697), .ZN(n7696) );
  AOI21_X1 U9026 ( .B1(n7697), .B2(n14205), .A(n6523), .ZN(n7695) );
  NAND2_X1 U9027 ( .A1(n15109), .A2(n7116), .ZN(n9615) );
  OAI21_X1 U9028 ( .B1(n14177), .B2(n7017), .A(n7015), .ZN(n14194) );
  OR2_X1 U9029 ( .A1(n11370), .A2(P1_U3086), .ZN(n14231) );
  INV_X1 U9030 ( .A(n15254), .ZN(n11377) );
  NOR2_X1 U9031 ( .A1(n14198), .A2(n14935), .ZN(n14239) );
  NAND2_X1 U9032 ( .A1(n6892), .A2(n6891), .ZN(n7125) );
  NAND2_X1 U9033 ( .A1(n11368), .A2(n10752), .ZN(n14243) );
  NAND2_X1 U9034 ( .A1(n9686), .A2(n9685), .ZN(n14478) );
  INV_X1 U9035 ( .A(n14226), .ZN(n14479) );
  INV_X1 U9036 ( .A(n14679), .ZN(n14480) );
  INV_X1 U9037 ( .A(n14171), .ZN(n14482) );
  INV_X1 U9038 ( .A(n14784), .ZN(n14483) );
  INV_X1 U9039 ( .A(n14862), .ZN(n14896) );
  INV_X1 U9040 ( .A(n11866), .ZN(n14491) );
  INV_X1 U9041 ( .A(n11826), .ZN(n14492) );
  OR2_X1 U9042 ( .A1(n9376), .A2(n9349), .ZN(n9351) );
  OR2_X1 U9043 ( .A1(n9539), .A2(n9348), .ZN(n9352) );
  NOR2_X1 U9044 ( .A1(n10256), .A2(n10255), .ZN(n10312) );
  NAND2_X1 U9045 ( .A1(n14552), .A2(n14551), .ZN(n14550) );
  AOI21_X1 U9046 ( .B1(n14550), .B2(n10353), .A(n10352), .ZN(n10366) );
  AOI21_X1 U9047 ( .B1(n10358), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10366), .ZN(
        n10316) );
  NAND2_X1 U9048 ( .A1(n10451), .A2(n6609), .ZN(n10455) );
  NOR2_X1 U9049 ( .A1(n10771), .A2(n10770), .ZN(n14580) );
  NAND2_X1 U9050 ( .A1(n14599), .A2(n6624), .ZN(n14614) );
  INV_X1 U9051 ( .A(n14981), .ZN(n14648) );
  XNOR2_X1 U9052 ( .A(n14668), .B(n14420), .ZN(n14652) );
  AOI21_X1 U9053 ( .B1(n14710), .B2(n6976), .A(n6974), .ZN(n14713) );
  INV_X1 U9054 ( .A(n6975), .ZN(n6974) );
  AOI21_X1 U9055 ( .B1(n6976), .B2(n14750), .A(n6536), .ZN(n6975) );
  AND2_X1 U9056 ( .A1(n9628), .A2(n9627), .ZN(n15000) );
  INV_X1 U9057 ( .A(n14748), .ZN(n14692) );
  INV_X1 U9058 ( .A(n15017), .ZN(n14790) );
  AOI21_X1 U9059 ( .B1(n7778), .B2(n9770), .A(n6427), .ZN(n14781) );
  NAND2_X1 U9060 ( .A1(n9570), .A2(n7672), .ZN(n7671) );
  NAND2_X1 U9061 ( .A1(n9570), .A2(n9569), .ZN(n14810) );
  NAND2_X1 U9062 ( .A1(n14840), .A2(n9768), .ZN(n14825) );
  NAND2_X1 U9063 ( .A1(n7170), .A2(n9558), .ZN(n14823) );
  NAND2_X1 U9064 ( .A1(n14855), .A2(n7174), .ZN(n7170) );
  NAND2_X1 U9065 ( .A1(n7773), .A2(n9765), .ZN(n14842) );
  NAND2_X1 U9066 ( .A1(n14855), .A2(n9544), .ZN(n14839) );
  NAND2_X1 U9067 ( .A1(n9764), .A2(n14342), .ZN(n14852) );
  NAND2_X1 U9068 ( .A1(n14893), .A2(n9519), .ZN(n14875) );
  NAND2_X1 U9069 ( .A1(n6642), .A2(n9506), .ZN(n14891) );
  CLKBUF_X1 U9070 ( .A(n14913), .Z(n14914) );
  AND2_X1 U9071 ( .A1(n11823), .A2(n9756), .ZN(n11864) );
  NAND2_X1 U9072 ( .A1(n10093), .A2(n7401), .ZN(n7399) );
  INV_X1 U9073 ( .A(n15217), .ZN(n14974) );
  OAI21_X1 U9074 ( .B1(n14643), .B2(n15259), .A(n14979), .ZN(n9854) );
  OAI21_X1 U9075 ( .B1(n14985), .B2(n15247), .A(n6677), .ZN(n15084) );
  AND2_X1 U9076 ( .A1(n14986), .A2(n14984), .ZN(n6677) );
  AND2_X1 U9077 ( .A1(n14987), .A2(n6619), .ZN(n6662) );
  INV_X1 U9078 ( .A(n10118), .ZN(n10149) );
  XNOR2_X1 U9079 ( .A(n9843), .B(n9842), .ZN(n14087) );
  OAI21_X1 U9080 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9843) );
  NAND2_X1 U9081 ( .A1(n12219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9330) );
  XNOR2_X1 U9082 ( .A(n9271), .B(n9817), .ZN(n14094) );
  NAND2_X1 U9083 ( .A1(n7683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U9084 ( .A1(n9719), .A2(n9704), .ZN(n9709) );
  NOR2_X1 U9085 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  NAND2_X1 U9086 ( .A1(n9152), .A2(n8694), .ZN(n11335) );
  XNOR2_X1 U9087 ( .A(n9605), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15109) );
  OR2_X1 U9088 ( .A1(n9604), .A2(n6409), .ZN(n9605) );
  OAI21_X1 U9089 ( .B1(n9696), .B2(n9695), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9697) );
  INV_X1 U9090 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15495) );
  OAI21_X1 U9091 ( .B1(n7596), .B2(n7594), .A(n9106), .ZN(n11230) );
  INV_X1 U9092 ( .A(n9104), .ZN(n7596) );
  NAND2_X1 U9093 ( .A1(n7597), .A2(n9103), .ZN(n7594) );
  NAND2_X1 U9094 ( .A1(n9105), .A2(n9076), .ZN(n11130) );
  NAND2_X1 U9095 ( .A1(n7595), .A2(n9104), .ZN(n9105) );
  NAND2_X1 U9096 ( .A1(n9104), .A2(n9073), .ZN(n9075) );
  INV_X1 U9097 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11116) );
  INV_X1 U9098 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10977) );
  INV_X1 U9099 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10370) );
  INV_X1 U9100 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10494) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10394) );
  XNOR2_X1 U9102 ( .A(n9510), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11617) );
  INV_X1 U9103 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10235) );
  XNOR2_X1 U9104 ( .A(n9508), .B(P1_IR_REG_13__SCAN_IN), .ZN(n14586) );
  INV_X1 U9105 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10187) );
  INV_X1 U9106 ( .A(n10460), .ZN(n10773) );
  INV_X1 U9107 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10145) );
  INV_X1 U9108 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10114) );
  INV_X1 U9109 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8621) );
  INV_X1 U9110 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10063) );
  OR2_X1 U9111 ( .A1(n9396), .A2(n9336), .ZN(n9397) );
  INV_X1 U9112 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10060) );
  OR2_X1 U9113 ( .A1(n9360), .A2(n9336), .ZN(n9362) );
  NOR2_X1 U9114 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9360) );
  XNOR2_X1 U9115 ( .A(n10037), .B(n15498), .ZN(n10035) );
  NAND2_X1 U9116 ( .A1(n10047), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10053) );
  XNOR2_X1 U9117 ( .A(n10076), .B(n10074), .ZN(n10073) );
  XNOR2_X1 U9118 ( .A(n10716), .B(n10410), .ZN(n10411) );
  NAND2_X1 U9119 ( .A1(n7248), .A2(n7117), .ZN(n11599) );
  NOR2_X1 U9120 ( .A1(n11598), .A2(n6532), .ZN(n7117) );
  AND2_X1 U9121 ( .A1(n11248), .A2(n6475), .ZN(n7245) );
  AND2_X1 U9122 ( .A1(n11248), .A2(n6556), .ZN(n7247) );
  NAND2_X1 U9123 ( .A1(n7077), .A2(n15142), .ZN(n7076) );
  NAND2_X1 U9124 ( .A1(n6668), .A2(n6667), .ZN(n15152) );
  INV_X1 U9125 ( .A(n15150), .ZN(n6667) );
  NAND2_X1 U9126 ( .A1(n7073), .A2(n6470), .ZN(n7074) );
  INV_X1 U9127 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U9128 ( .A1(n12628), .A2(n12627), .ZN(n12652) );
  OAI21_X1 U9129 ( .B1(n6672), .B2(n12506), .A(n12340), .ZN(P3_U3154) );
  XNOR2_X1 U9130 ( .A(n12335), .B(n6673), .ZN(n6672) );
  NAND2_X1 U9131 ( .A1(n11183), .A2(n7039), .ZN(n11286) );
  INV_X1 U9132 ( .A(n7239), .ZN(n10945) );
  NAND2_X1 U9133 ( .A1(n10450), .A2(n6626), .ZN(P3_U3183) );
  AOI21_X1 U9134 ( .B1(n7216), .B2(n12707), .A(n7212), .ZN(n12662) );
  NAND2_X1 U9135 ( .A1(n7215), .A2(n7213), .ZN(n7212) );
  AOI21_X1 U9136 ( .B1(n6442), .B2(n12584), .A(n6907), .ZN(n12708) );
  OAI21_X1 U9137 ( .B1(n13039), .B2(n10095), .A(n7208), .ZN(P3_U3294) );
  NOR2_X1 U9138 ( .A1(n7210), .A2(n7209), .ZN(n7208) );
  NOR2_X1 U9139 ( .A1(P3_U3151), .A2(n7211), .ZN(n7209) );
  NOR2_X1 U9140 ( .A1(n13034), .A2(n10094), .ZN(n7210) );
  OR2_X1 U9141 ( .A1(n9285), .A2(n9287), .ZN(n9312) );
  NOR2_X1 U9142 ( .A1(n6779), .A2(n13542), .ZN(n6778) );
  NAND2_X1 U9143 ( .A1(n6786), .A2(n13428), .ZN(n6785) );
  OR2_X1 U9144 ( .A1(n15384), .A2(n7266), .ZN(n7265) );
  INV_X1 U9145 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U9146 ( .A1(n6768), .A2(n6766), .ZN(P2_U3494) );
  OR2_X1 U9147 ( .A1(n13959), .A2(n6769), .ZN(n6768) );
  AOI21_X1 U9148 ( .B1(n13666), .B2(n6607), .A(n6767), .ZN(n6766) );
  OAI21_X1 U9149 ( .B1(n15103), .B2(n14092), .A(n7329), .ZN(P2_U3297) );
  NOR2_X1 U9150 ( .A1(n7331), .A2(n7330), .ZN(n7329) );
  NOR2_X1 U9151 ( .A1(n8602), .A2(P2_U3088), .ZN(n7330) );
  NOR2_X1 U9152 ( .A1(n14097), .A2(n13368), .ZN(n7331) );
  OAI21_X1 U9153 ( .B1(n7095), .B2(n15174), .A(n7094), .ZN(P1_U3225) );
  AND2_X1 U9154 ( .A1(n14156), .A2(n14155), .ZN(n7094) );
  XNOR2_X1 U9155 ( .A(n14151), .B(n7096), .ZN(n7095) );
  AND2_X1 U9156 ( .A1(n14230), .A2(n6618), .ZN(n7097) );
  INV_X1 U9157 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10166) );
  AOI21_X1 U9158 ( .B1(n15199), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n14639), .ZN(
        n6849) );
  NAND2_X1 U9159 ( .A1(n6851), .A2(n14246), .ZN(n6850) );
  NAND2_X1 U9160 ( .A1(n6847), .A2(n14917), .ZN(n6846) );
  OAI21_X1 U9161 ( .B1(n9811), .B2(n6412), .A(n9799), .ZN(n9800) );
  MUX2_X1 U9162 ( .A(n15002), .B(n15087), .S(n15272), .Z(n15003) );
  AOI21_X1 U9163 ( .B1(n7187), .B2(n15265), .A(n6611), .ZN(n7186) );
  NAND2_X1 U9164 ( .A1(n7246), .A2(n11248), .ZN(n11589) );
  NAND2_X1 U9165 ( .A1(n11980), .A2(n7305), .ZN(n15112) );
  INV_X1 U9166 ( .A(n7303), .ZN(n15124) );
  AND2_X1 U9167 ( .A1(n7148), .A2(n6483), .ZN(n6419) );
  OR2_X1 U9168 ( .A1(n15376), .A2(n11490), .ZN(n6420) );
  XNOR2_X1 U9169 ( .A(n14476), .B(n14648), .ZN(n6421) );
  AND3_X1 U9170 ( .A1(n9779), .A2(n6446), .A3(n6421), .ZN(n6422) );
  MUX2_X1 U9171 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6639), .S(n9347), .Z(n14972)
         );
  INV_X1 U9172 ( .A(n14972), .ZN(n10837) );
  AND2_X1 U9173 ( .A1(n13301), .A2(n13303), .ZN(n6423) );
  INV_X1 U9174 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7769) );
  AND2_X1 U9175 ( .A1(n6995), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6424) );
  OR2_X1 U9176 ( .A1(n8285), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6425) );
  INV_X1 U9177 ( .A(n6833), .ZN(n11384) );
  OAI21_X1 U9178 ( .B1(n11138), .B2(n6834), .A(n11379), .ZN(n6833) );
  OR2_X1 U9179 ( .A1(n13988), .A2(n13630), .ZN(n6426) );
  NAND2_X1 U9180 ( .A1(n7982), .A2(n7910), .ZN(n8187) );
  AND2_X1 U9181 ( .A1(n7871), .A2(n7870), .ZN(n8108) );
  AND2_X1 U9182 ( .A1(n7982), .A2(n7590), .ZN(n8222) );
  NOR2_X1 U9183 ( .A1(n7847), .A2(n14801), .ZN(n6427) );
  NAND2_X1 U9184 ( .A1(n14226), .A2(n14983), .ZN(n9780) );
  AND2_X1 U9185 ( .A1(n9615), .A2(n14790), .ZN(n6428) );
  AND2_X1 U9186 ( .A1(n13878), .A2(n7553), .ZN(n6429) );
  AND2_X1 U9187 ( .A1(n7590), .A2(n8221), .ZN(n6430) );
  AND2_X1 U9188 ( .A1(n7555), .A2(n7554), .ZN(n6431) );
  AND2_X1 U9189 ( .A1(n6549), .A2(n6719), .ZN(n6432) );
  INV_X1 U9190 ( .A(n9890), .ZN(n7149) );
  INV_X1 U9191 ( .A(n6602), .ZN(n6834) );
  NAND2_X1 U9192 ( .A1(n8856), .A2(n8855), .ZN(n13246) );
  INV_X1 U9193 ( .A(n13246), .ZN(n7545) );
  INV_X1 U9194 ( .A(n12297), .ZN(n7690) );
  INV_X1 U9195 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7230) );
  NOR3_X1 U9196 ( .A1(n11902), .A2(n6530), .A3(n12002), .ZN(n6433) );
  AND2_X1 U9197 ( .A1(n12811), .A2(n12825), .ZN(n6434) );
  AND2_X1 U9198 ( .A1(n12734), .A2(n8497), .ZN(n6435) );
  NAND2_X1 U9199 ( .A1(n14178), .A2(n12255), .ZN(n14135) );
  INV_X1 U9200 ( .A(n12181), .ZN(n7569) );
  INV_X1 U9201 ( .A(n13258), .ZN(n7631) );
  AND2_X1 U9202 ( .A1(n9917), .A2(n7029), .ZN(n6436) );
  AND2_X1 U9203 ( .A1(n7321), .A2(n7315), .ZN(n6437) );
  NOR2_X1 U9204 ( .A1(n8677), .A2(n10817), .ZN(n7617) );
  AND2_X1 U9205 ( .A1(n14738), .A2(n6560), .ZN(n6438) );
  NAND2_X1 U9206 ( .A1(n10154), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6439) );
  INV_X1 U9207 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13017) );
  AND2_X1 U9208 ( .A1(n7628), .A2(n13251), .ZN(n6440) );
  NAND2_X1 U9209 ( .A1(n9315), .A2(n9314), .ZN(n9705) );
  AND2_X1 U9210 ( .A1(n7671), .A2(n9582), .ZN(n6441) );
  XOR2_X1 U9211 ( .A(n7346), .B(n7345), .Z(n6442) );
  NOR2_X1 U9212 ( .A1(n15053), .A2(n14896), .ZN(n6443) );
  AND2_X1 U9213 ( .A1(n6559), .A2(n7569), .ZN(n7567) );
  INV_X1 U9214 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9690) );
  INV_X1 U9215 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9545) );
  AOI21_X1 U9216 ( .B1(n14110), .B2(n12111), .A(n7692), .ZN(n7691) );
  AND2_X1 U9217 ( .A1(n10147), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6444) );
  INV_X1 U9218 ( .A(n9779), .ZN(n7664) );
  NAND2_X1 U9219 ( .A1(n14294), .A2(n7381), .ZN(n6445) );
  AND3_X1 U9220 ( .A1(n9679), .A2(n14656), .A3(n14456), .ZN(n6446) );
  AND2_X1 U9221 ( .A1(n7574), .A2(n12350), .ZN(n6447) );
  AND2_X1 U9222 ( .A1(n7751), .A2(n9880), .ZN(n6448) );
  NOR2_X1 U9223 ( .A1(n13575), .A2(n7314), .ZN(n6449) );
  NAND2_X1 U9224 ( .A1(n7253), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7252) );
  INV_X1 U9225 ( .A(n12046), .ZN(n6890) );
  NAND2_X1 U9226 ( .A1(n7547), .A2(n7546), .ZN(n11488) );
  NAND2_X1 U9227 ( .A1(n11857), .A2(n7733), .ZN(n11958) );
  NOR2_X1 U9228 ( .A1(n9031), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U9229 ( .A1(n7750), .A2(n6606), .ZN(n11799) );
  AND2_X1 U9230 ( .A1(n11724), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6450) );
  OR2_X1 U9231 ( .A1(n9214), .A2(SI_26_), .ZN(n6451) );
  AND2_X1 U9232 ( .A1(n10005), .A2(n13429), .ZN(n13920) );
  AND2_X1 U9233 ( .A1(n6897), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6452) );
  AND2_X1 U9234 ( .A1(n6631), .A2(n7238), .ZN(n6453) );
  OR2_X1 U9235 ( .A1(n6807), .A2(n6810), .ZN(n6454) );
  NOR2_X1 U9236 ( .A1(n7205), .A2(n6996), .ZN(n6455) );
  OR2_X1 U9237 ( .A1(n8346), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U9238 ( .A(n11501), .B(n11667), .ZN(n11666) );
  NOR2_X1 U9239 ( .A1(n8500), .A2(n7487), .ZN(n7486) );
  NAND2_X1 U9240 ( .A1(n6760), .A2(n6758), .ZN(n13834) );
  NOR2_X1 U9241 ( .A1(n12022), .A2(n12466), .ZN(n6459) );
  NAND2_X1 U9242 ( .A1(n13049), .A2(n8984), .ZN(n13105) );
  INV_X1 U9243 ( .A(n13563), .ZN(n13558) );
  NAND2_X1 U9244 ( .A1(n14107), .A2(n12111), .ZN(n12125) );
  INV_X2 U9245 ( .A(n7950), .ZN(n8395) );
  NAND2_X1 U9246 ( .A1(n7951), .A2(n7952), .ZN(n7950) );
  INV_X1 U9247 ( .A(n7950), .ZN(n8053) );
  NOR2_X1 U9248 ( .A1(n12523), .A2(n10823), .ZN(n11004) );
  NAND2_X1 U9249 ( .A1(n9770), .A2(n9769), .ZN(n14799) );
  AND2_X1 U9250 ( .A1(n7420), .A2(n12672), .ZN(n6460) );
  INV_X1 U9251 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U9252 ( .A1(n13167), .A2(n6858), .ZN(n6461) );
  NAND2_X1 U9253 ( .A1(n10145), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U9254 ( .A1(n13692), .A2(n13667), .ZN(n6463) );
  AND2_X1 U9255 ( .A1(n13600), .A2(n13599), .ZN(n6464) );
  INV_X1 U9256 ( .A(n14289), .ZN(n15260) );
  NAND2_X1 U9257 ( .A1(n9420), .A2(n9419), .ZN(n14289) );
  AND2_X1 U9258 ( .A1(n8105), .A2(n9936), .ZN(n6465) );
  NAND2_X1 U9259 ( .A1(n13912), .A2(n13614), .ZN(n6466) );
  NAND2_X1 U9260 ( .A1(n8440), .A2(n8439), .ZN(n8508) );
  AND2_X1 U9261 ( .A1(n6869), .A2(n6867), .ZN(n6467) );
  NOR2_X1 U9262 ( .A1(n11882), .A2(n12516), .ZN(n6468) );
  AND2_X1 U9263 ( .A1(n7437), .A2(n8966), .ZN(n6469) );
  AND3_X1 U9264 ( .A1(n9400), .A2(n9399), .A3(n9398), .ZN(n11357) );
  OAI21_X1 U9265 ( .B1(n10646), .B2(n7362), .A(n6478), .ZN(n7089) );
  XOR2_X1 U9266 ( .A(n15164), .B(n15159), .Z(n6470) );
  INV_X1 U9267 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7947) );
  NOR2_X1 U9268 ( .A1(n8599), .A2(n8763), .ZN(n6471) );
  XNOR2_X1 U9269 ( .A(n15005), .B(n14171), .ZN(n14750) );
  XNOR2_X1 U9270 ( .A(n13947), .B(n13391), .ZN(n13643) );
  INV_X1 U9271 ( .A(n13643), .ZN(n7603) );
  NAND4_X2 U9272 ( .A1(n8013), .A2(n8012), .A3(n8011), .A4(n8010), .ZN(n12521)
         );
  AND2_X1 U9273 ( .A1(n10313), .A2(n10244), .ZN(n6472) );
  XNOR2_X1 U9274 ( .A(n13640), .B(n6735), .ZN(n13674) );
  OAI211_X1 U9275 ( .C1(n7861), .C2(n6682), .A(n6680), .B(n7864), .ZN(n8086)
         );
  NAND2_X1 U9276 ( .A1(n9481), .A2(n9480), .ZN(n14951) );
  OR2_X1 U9277 ( .A1(n13997), .A2(n13628), .ZN(n6473) );
  NAND2_X1 U9278 ( .A1(n7711), .A2(n13585), .ZN(n13715) );
  OR2_X1 U9279 ( .A1(n15017), .A2(n12257), .ZN(n6474) );
  INV_X1 U9280 ( .A(n7123), .ZN(n7122) );
  INV_X1 U9281 ( .A(n11179), .ZN(n10983) );
  INV_X1 U9282 ( .A(n13972), .ZN(n7554) );
  NAND2_X1 U9283 ( .A1(n12856), .A2(n9888), .ZN(n12844) );
  NAND2_X1 U9284 ( .A1(n11862), .A2(n9757), .ZN(n11952) );
  NAND2_X1 U9285 ( .A1(n7311), .A2(n13572), .ZN(n13830) );
  NAND2_X1 U9286 ( .A1(n9549), .A2(n9548), .ZN(n14844) );
  INV_X1 U9287 ( .A(n14844), .ZN(n7717) );
  NAND2_X1 U9288 ( .A1(n11590), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6475) );
  INV_X1 U9289 ( .A(n8478), .ZN(n7490) );
  INV_X1 U9290 ( .A(n11776), .ZN(n7754) );
  XNOR2_X1 U9291 ( .A(n14289), .B(n14493), .ZN(n14444) );
  INV_X1 U9292 ( .A(n14444), .ZN(n9749) );
  INV_X1 U9293 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9331) );
  AND2_X1 U9294 ( .A1(n12474), .A2(n12473), .ZN(n6476) );
  AND2_X1 U9295 ( .A1(n6789), .A2(n6788), .ZN(n6477) );
  OR2_X1 U9296 ( .A1(n10636), .A2(n10655), .ZN(n6478) );
  NAND2_X1 U9297 ( .A1(n7960), .A2(n7959), .ZN(n12954) );
  OR2_X1 U9298 ( .A1(n10605), .A2(n10727), .ZN(n6479) );
  INV_X1 U9299 ( .A(n13609), .ZN(n14041) );
  INV_X1 U9300 ( .A(n12518), .ZN(n11681) );
  NAND2_X1 U9301 ( .A1(n7153), .A2(n9884), .ZN(n12030) );
  OR2_X1 U9302 ( .A1(n14697), .A2(n14983), .ZN(n6480) );
  AND2_X1 U9303 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n7049), .ZN(n6481) );
  AND3_X1 U9304 ( .A1(n10801), .A2(n9936), .A3(n8034), .ZN(n6482) );
  OR2_X1 U9305 ( .A1(n12811), .A2(n12825), .ZN(n6483) );
  AND2_X1 U9306 ( .A1(n13000), .A2(n12860), .ZN(n6484) );
  INV_X1 U9307 ( .A(n7800), .ZN(n7801) );
  NAND2_X1 U9308 ( .A1(n9524), .A2(n9523), .ZN(n15053) );
  OR2_X1 U9309 ( .A1(n8508), .A2(n12062), .ZN(n6485) );
  AND2_X1 U9310 ( .A1(n8483), .A2(n12845), .ZN(n6486) );
  INV_X1 U9311 ( .A(n13641), .ZN(n13657) );
  AND2_X1 U9312 ( .A1(n8459), .A2(n8106), .ZN(n6487) );
  NAND2_X1 U9313 ( .A1(n9036), .A2(n9035), .ZN(n14008) );
  INV_X1 U9314 ( .A(n14008), .ZN(n7552) );
  INV_X1 U9315 ( .A(n13421), .ZN(n11129) );
  NAND2_X1 U9316 ( .A1(n8047), .A2(n11004), .ZN(n10798) );
  OR2_X1 U9317 ( .A1(n12935), .A2(n12478), .ZN(n6488) );
  INV_X1 U9318 ( .A(n14750), .ZN(n14752) );
  OR2_X1 U9319 ( .A1(n12138), .A2(n12511), .ZN(n6489) );
  AND2_X1 U9320 ( .A1(n11164), .A2(n11247), .ZN(n6490) );
  NOR2_X1 U9321 ( .A1(n14815), .A2(n7847), .ZN(n6491) );
  INV_X1 U9322 ( .A(n12401), .ZN(n7028) );
  AND4_X1 U9323 ( .A1(n8597), .A2(n8596), .A3(P2_IR_REG_21__SCAN_IN), .A4(
        n8779), .ZN(n6492) );
  INV_X1 U9324 ( .A(n12208), .ZN(n7586) );
  AND2_X1 U9325 ( .A1(n13663), .A2(n13392), .ZN(n6493) );
  AND2_X1 U9326 ( .A1(n6532), .A2(n11598), .ZN(n6494) );
  AND2_X1 U9327 ( .A1(n11869), .A2(n12517), .ZN(n6495) );
  INV_X1 U9328 ( .A(n13982), .ZN(n13754) );
  NAND2_X1 U9329 ( .A1(n9136), .A2(n9135), .ZN(n13982) );
  NOR3_X1 U9330 ( .A1(n14349), .A2(n14348), .A3(n14359), .ZN(n6496) );
  AND2_X1 U9331 ( .A1(n13385), .A2(n13384), .ZN(n6497) );
  NAND2_X1 U9332 ( .A1(n9320), .A2(n9319), .ZN(n9381) );
  OR2_X1 U9333 ( .A1(n10431), .A2(n7211), .ZN(n6498) );
  NOR2_X1 U9334 ( .A1(n12243), .A2(n14215), .ZN(n6499) );
  INV_X1 U9335 ( .A(n8046), .ZN(n10949) );
  AND2_X1 U9336 ( .A1(n14650), .A2(n7663), .ZN(n6500) );
  INV_X1 U9337 ( .A(n14004), .ZN(n13824) );
  NAND2_X1 U9338 ( .A1(n9058), .A2(n9057), .ZN(n14004) );
  NOR2_X1 U9339 ( .A1(n15001), .A2(n7184), .ZN(n6501) );
  NOR2_X1 U9340 ( .A1(n12531), .A2(n12530), .ZN(n6502) );
  INV_X1 U9341 ( .A(n14248), .ZN(n10741) );
  INV_X1 U9342 ( .A(n14303), .ZN(n14302) );
  OR2_X1 U9343 ( .A1(n8484), .A2(n7490), .ZN(n6503) );
  AND2_X1 U9344 ( .A1(n13626), .A2(n13625), .ZN(n6504) );
  AND2_X1 U9345 ( .A1(n7446), .A2(n9051), .ZN(n6505) );
  AND2_X1 U9346 ( .A1(n14178), .A2(n7684), .ZN(n6506) );
  INV_X1 U9347 ( .A(n13257), .ZN(n7632) );
  AND2_X1 U9348 ( .A1(n7633), .A2(n7629), .ZN(n6507) );
  AND2_X1 U9349 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .ZN(n6508) );
  INV_X1 U9350 ( .A(n9454), .ZN(n7659) );
  AND2_X1 U9351 ( .A1(n8399), .A2(n8501), .ZN(n12725) );
  INV_X1 U9352 ( .A(n12725), .ZN(n7487) );
  AND2_X1 U9353 ( .A1(n9885), .A2(n9884), .ZN(n6509) );
  OR2_X1 U9354 ( .A1(n10821), .A2(n10501), .ZN(n6510) );
  AND2_X1 U9355 ( .A1(n7947), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6511) );
  AND2_X1 U9356 ( .A1(n14853), .A2(n14342), .ZN(n6512) );
  INV_X1 U9357 ( .A(n7151), .ZN(n7150) );
  INV_X1 U9358 ( .A(n7832), .ZN(n7822) );
  AND2_X1 U9359 ( .A1(n7664), .A2(n9678), .ZN(n6513) );
  AND2_X1 U9360 ( .A1(n14367), .A2(n14366), .ZN(n6514) );
  AND2_X1 U9361 ( .A1(n8684), .A2(n7263), .ZN(n6515) );
  OR2_X1 U9362 ( .A1(n10695), .A2(n10501), .ZN(n6516) );
  NOR2_X1 U9363 ( .A1(n13574), .A2(n7316), .ZN(n7315) );
  OR2_X1 U9364 ( .A1(n10282), .A2(n10281), .ZN(n6517) );
  INV_X1 U9365 ( .A(n11394), .ZN(n7375) );
  INV_X1 U9366 ( .A(n9753), .ZN(n7771) );
  AND2_X1 U9367 ( .A1(n6772), .A2(n6774), .ZN(n6518) );
  INV_X1 U9368 ( .A(n9880), .ZN(n7749) );
  OR2_X1 U9369 ( .A1(n9089), .A2(n8678), .ZN(n6519) );
  INV_X1 U9370 ( .A(n7670), .ZN(n7669) );
  NAND2_X1 U9371 ( .A1(n7674), .A2(n9582), .ZN(n7670) );
  NOR2_X1 U9372 ( .A1(n14303), .A2(n14936), .ZN(n6520) );
  NOR2_X1 U9373 ( .A1(n12993), .A2(n12832), .ZN(n6521) );
  NOR2_X1 U9374 ( .A1(n11577), .A2(n13256), .ZN(n6522) );
  NOR2_X1 U9375 ( .A1(n12097), .A2(n12096), .ZN(n6523) );
  INV_X1 U9376 ( .A(n8644), .ZN(n7057) );
  NAND2_X1 U9377 ( .A1(n12968), .A2(n12779), .ZN(n6524) );
  XOR2_X1 U9378 ( .A(n15167), .B(n15166), .Z(n6525) );
  AND2_X1 U9379 ( .A1(n6457), .A2(n7821), .ZN(n6526) );
  INV_X1 U9380 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U9381 ( .A1(n8499), .A2(n8396), .ZN(n9904) );
  INV_X1 U9382 ( .A(n9904), .ZN(n12734) );
  NAND2_X1 U9383 ( .A1(n9123), .A2(n13072), .ZN(n6527) );
  OR2_X1 U9384 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_30__SCAN_IN), .ZN(
        n6528) );
  OR2_X1 U9385 ( .A1(n12129), .A2(n12128), .ZN(n6529) );
  AND2_X1 U9386 ( .A1(n11996), .A2(n11995), .ZN(n6530) );
  AND4_X1 U9387 ( .A1(n7913), .A2(n7915), .A3(n7914), .A4(n7916), .ZN(n6531)
         );
  INV_X1 U9388 ( .A(n7760), .ZN(n7759) );
  AND2_X1 U9389 ( .A1(n9899), .A2(n7761), .ZN(n7760) );
  AND2_X1 U9390 ( .A1(n8997), .A2(n8707), .ZN(n9003) );
  AND2_X1 U9391 ( .A1(n11592), .A2(n11591), .ZN(n6532) );
  INV_X1 U9392 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9337) );
  AND2_X1 U9393 ( .A1(n8649), .A2(SI_9_), .ZN(n6533) );
  NAND2_X1 U9394 ( .A1(n7588), .A2(n12017), .ZN(n6534) );
  INV_X1 U9395 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7049) );
  AND2_X1 U9396 ( .A1(n13214), .A2(n13213), .ZN(n6535) );
  AND2_X1 U9397 ( .A1(n15000), .A2(n14712), .ZN(n6536) );
  OR2_X1 U9398 ( .A1(n14394), .A2(n14392), .ZN(n6537) );
  AND2_X1 U9399 ( .A1(n13932), .A2(n13611), .ZN(n6538) );
  INV_X1 U9400 ( .A(n7613), .ZN(n7612) );
  AND2_X1 U9401 ( .A1(n14380), .A2(n7849), .ZN(n6539) );
  XOR2_X1 U9402 ( .A(n14475), .B(n14643), .Z(n14457) );
  AND2_X1 U9403 ( .A1(n7286), .A2(n8100), .ZN(n6540) );
  AND3_X1 U9404 ( .A1(n8587), .A2(n8586), .A3(n8588), .ZN(n8616) );
  INV_X1 U9405 ( .A(n6735), .ZN(n13960) );
  NAND2_X1 U9406 ( .A1(n9217), .A2(n9216), .ZN(n6735) );
  AND2_X1 U9407 ( .A1(n12305), .A2(n12304), .ZN(n6541) );
  AND2_X1 U9408 ( .A1(n12261), .A2(n12260), .ZN(n6542) );
  OR2_X1 U9409 ( .A1(n8994), .A2(n8669), .ZN(n6543) );
  AND2_X1 U9410 ( .A1(n10114), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6544) );
  AND2_X1 U9411 ( .A1(n10112), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6545) );
  OR2_X1 U9412 ( .A1(n9988), .A2(n9987), .ZN(n6546) );
  AND2_X1 U9413 ( .A1(n7516), .A2(n6462), .ZN(n6547) );
  INV_X1 U9414 ( .A(n7513), .ZN(n7512) );
  NAND2_X1 U9415 ( .A1(n7514), .A2(n6462), .ZN(n7513) );
  INV_X1 U9416 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10061) );
  AND2_X1 U9417 ( .A1(n7627), .A2(n7628), .ZN(n6548) );
  INV_X1 U9418 ( .A(n7680), .ZN(n7679) );
  NAND2_X1 U9419 ( .A1(n7681), .A2(n9506), .ZN(n7680) );
  INV_X1 U9420 ( .A(n7373), .ZN(n7372) );
  OAI21_X1 U9421 ( .B1(n11394), .B2(n11395), .A(n11726), .ZN(n7373) );
  OR2_X1 U9422 ( .A1(n13303), .A2(n13301), .ZN(n6549) );
  OR2_X1 U9423 ( .A1(n7881), .A2(n7538), .ZN(n6550) );
  AND2_X1 U9424 ( .A1(n12206), .A2(n12489), .ZN(n6551) );
  OAI21_X1 U9425 ( .B1(n13736), .B2(n13633), .A(n13730), .ZN(n13632) );
  INV_X1 U9426 ( .A(n7321), .ZN(n7320) );
  NAND2_X1 U9427 ( .A1(n13878), .A2(n13886), .ZN(n7321) );
  NAND2_X1 U9428 ( .A1(n12169), .A2(n12164), .ZN(n6552) );
  NAND2_X1 U9429 ( .A1(n10061), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6553) );
  INV_X1 U9430 ( .A(n7089), .ZN(n7361) );
  INV_X1 U9431 ( .A(n7180), .ZN(n7178) );
  NAND2_X1 U9432 ( .A1(n7182), .A2(n7181), .ZN(n7180) );
  OR2_X1 U9433 ( .A1(n10607), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6554) );
  OR2_X1 U9434 ( .A1(n7633), .A2(n7629), .ZN(n6555) );
  NOR2_X1 U9435 ( .A1(n14499), .A2(n10837), .ZN(n14255) );
  AND2_X1 U9436 ( .A1(n6475), .A2(n11598), .ZN(n6556) );
  NOR3_X1 U9437 ( .A1(n13737), .A2(n13755), .A3(n13413), .ZN(n6557) );
  OR2_X1 U9438 ( .A1(n11491), .A2(n13444), .ZN(n6558) );
  OR2_X1 U9439 ( .A1(n12474), .A2(n12473), .ZN(n6559) );
  NAND2_X2 U9440 ( .A1(n9640), .A2(n9639), .ZN(n15005) );
  INV_X1 U9441 ( .A(n15005), .ZN(n7731) );
  AND2_X1 U9442 ( .A1(n7185), .A2(n14737), .ZN(n6560) );
  OR2_X1 U9443 ( .A1(n11347), .A2(n11346), .ZN(n6561) );
  AND2_X1 U9444 ( .A1(n7111), .A2(n8633), .ZN(n6562) );
  OR2_X1 U9445 ( .A1(n14331), .A2(n14330), .ZN(n6563) );
  AND2_X1 U9446 ( .A1(n6920), .A2(n6919), .ZN(n6564) );
  AND3_X1 U9447 ( .A1(n8779), .A2(n8596), .A3(n6871), .ZN(n6565) );
  OR2_X1 U9448 ( .A1(n8029), .A2(n10507), .ZN(n6566) );
  OR2_X1 U9449 ( .A1(n9054), .A2(SI_18_), .ZN(n6567) );
  OR2_X1 U9450 ( .A1(n8121), .A2(n6465), .ZN(n6568) );
  INV_X1 U9451 ( .A(n14245), .ZN(n9803) );
  XNOR2_X1 U9452 ( .A(n9697), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14245) );
  AND2_X1 U9453 ( .A1(n7718), .A2(n7717), .ZN(n6569) );
  AND2_X1 U9454 ( .A1(n7543), .A2(n13912), .ZN(n6570) );
  NOR2_X1 U9455 ( .A1(n13960), .A2(n13640), .ZN(n6571) );
  NOR2_X1 U9456 ( .A1(n11897), .A2(n11900), .ZN(n6572) );
  AND2_X1 U9457 ( .A1(n14225), .A2(n14995), .ZN(n6573) );
  OR2_X1 U9458 ( .A1(n12580), .A2(n12581), .ZN(n6574) );
  NAND2_X1 U9459 ( .A1(n7671), .A2(n7669), .ZN(n14793) );
  NOR2_X1 U9460 ( .A1(n8370), .A2(n9899), .ZN(n6575) );
  OR2_X1 U9461 ( .A1(n7728), .A2(n7634), .ZN(n6576) );
  OR2_X1 U9462 ( .A1(n13960), .A2(n14024), .ZN(n6577) );
  INV_X1 U9463 ( .A(n14350), .ZN(n6946) );
  AND2_X1 U9464 ( .A1(n7179), .A2(n9776), .ZN(n6578) );
  INV_X1 U9465 ( .A(n13708), .ZN(n13967) );
  AND2_X1 U9466 ( .A1(n9177), .A2(n9176), .ZN(n13708) );
  XNOR2_X1 U9467 ( .A(n7867), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8098) );
  AND2_X1 U9468 ( .A1(n9319), .A2(n9382), .ZN(n6579) );
  INV_X1 U9469 ( .A(n6951), .ZN(n6950) );
  OAI22_X1 U9470 ( .A1(n14424), .A2(n14425), .B1(n14423), .B2(n14422), .ZN(
        n6951) );
  AND2_X1 U9471 ( .A1(n11018), .A2(n12878), .ZN(n6580) );
  AND2_X1 U9472 ( .A1(n8496), .A2(n8376), .ZN(n6581) );
  INV_X1 U9473 ( .A(n8495), .ZN(n7472) );
  AND2_X1 U9474 ( .A1(n7660), .A2(n9454), .ZN(n6582) );
  AND2_X1 U9475 ( .A1(n7586), .A2(n7583), .ZN(n6583) );
  AND2_X1 U9476 ( .A1(n7628), .A2(n13247), .ZN(n6584) );
  AND2_X1 U9477 ( .A1(n7370), .A2(n6502), .ZN(n6585) );
  INV_X1 U9478 ( .A(n13624), .ZN(n6761) );
  AND2_X1 U9479 ( .A1(n7859), .A2(n7858), .ZN(n6586) );
  AND2_X1 U9480 ( .A1(n13578), .A2(n13577), .ZN(n6587) );
  INV_X1 U9481 ( .A(n13298), .ZN(n6720) );
  INV_X1 U9482 ( .A(n6962), .ZN(n6961) );
  OAI21_X1 U9483 ( .B1(n7772), .B2(n6963), .A(n14824), .ZN(n6962) );
  OR2_X1 U9484 ( .A1(n9877), .A2(n7137), .ZN(n6588) );
  INV_X1 U9485 ( .A(n7314), .ZN(n7313) );
  NOR2_X1 U9486 ( .A1(n7552), .A2(n13848), .ZN(n7314) );
  OR2_X1 U9487 ( .A1(n14406), .A2(n14404), .ZN(n6589) );
  NAND2_X1 U9488 ( .A1(n14650), .A2(n9687), .ZN(n9779) );
  AND2_X1 U9489 ( .A1(n8512), .A2(n8505), .ZN(n6590) );
  AND3_X1 U9490 ( .A1(n8558), .A2(n8557), .A3(n8556), .ZN(n6591) );
  OR2_X1 U9491 ( .A1(n7379), .A2(n14405), .ZN(n6592) );
  AND2_X1 U9492 ( .A1(n7809), .A2(n7805), .ZN(n6593) );
  AND2_X1 U9493 ( .A1(n7716), .A2(n7682), .ZN(n6594) );
  INV_X1 U9494 ( .A(n11379), .ZN(n11150) );
  NAND2_X1 U9495 ( .A1(n8155), .A2(n11565), .ZN(n6595) );
  INV_X1 U9496 ( .A(n8663), .ZN(n6739) );
  INV_X1 U9497 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10092) );
  INV_X1 U9498 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8246) );
  AND2_X1 U9499 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .ZN(n6596) );
  OR2_X1 U9500 ( .A1(n12909), .A2(n12767), .ZN(n6597) );
  NAND2_X1 U9501 ( .A1(n10727), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6598) );
  INV_X1 U9502 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U9503 ( .A1(n14751), .A2(n6976), .ZN(n6599) );
  AND2_X1 U9504 ( .A1(n6420), .A2(n11080), .ZN(n6600) );
  NAND2_X1 U9505 ( .A1(n14224), .A2(n14152), .ZN(n6601) );
  INV_X1 U9506 ( .A(n7391), .ZN(n7390) );
  NAND2_X1 U9507 ( .A1(n14768), .A2(n14377), .ZN(n7391) );
  INV_X1 U9508 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6871) );
  INV_X1 U9509 ( .A(n7338), .ZN(n7337) );
  NAND2_X1 U9510 ( .A1(n11081), .A2(n7340), .ZN(n7338) );
  INV_X1 U9511 ( .A(n6727), .ZN(n6726) );
  NAND2_X1 U9512 ( .A1(n7534), .A2(n6728), .ZN(n6727) );
  INV_X1 U9513 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10059) );
  INV_X1 U9514 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9515 ( .A1(n11144), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U9516 ( .A1(n14658), .A2(n15217), .ZN(n15220) );
  INV_X1 U9517 ( .A(n14804), .ZN(n7674) );
  NAND2_X1 U9518 ( .A1(n10679), .A2(n8792), .ZN(n10678) );
  NAND2_X1 U9519 ( .A1(n7720), .A2(n7722), .ZN(n11325) );
  NAND2_X1 U9520 ( .A1(n13872), .A2(n13878), .ZN(n13850) );
  NAND2_X1 U9521 ( .A1(n14900), .A2(n14888), .ZN(n14858) );
  AND2_X1 U9522 ( .A1(n13872), .A2(n7551), .ZN(n6603) );
  AND2_X1 U9523 ( .A1(n9303), .A2(n9263), .ZN(n13182) );
  INV_X1 U9524 ( .A(n13182), .ZN(n13165) );
  AND2_X1 U9525 ( .A1(n11814), .A2(n6570), .ZN(n13888) );
  AND2_X1 U9526 ( .A1(n11857), .A2(n14305), .ZN(n11858) );
  NAND2_X1 U9527 ( .A1(n11847), .A2(n7828), .ZN(n11898) );
  NAND2_X1 U9528 ( .A1(n7222), .A2(n9919), .ZN(n10796) );
  NAND2_X1 U9529 ( .A1(n6886), .A2(n9670), .ZN(n14983) );
  INV_X1 U9530 ( .A(n14983), .ZN(n7727) );
  OAI21_X1 U9531 ( .B1(n11566), .B2(n11565), .A(n9879), .ZN(n11775) );
  NAND2_X1 U9532 ( .A1(n6885), .A2(n8464), .ZN(n11774) );
  NAND2_X1 U9533 ( .A1(n13616), .A2(n13615), .ZN(n13895) );
  NAND2_X1 U9534 ( .A1(n9918), .A2(n9917), .ZN(n9920) );
  INV_X1 U9535 ( .A(n10590), .ZN(n6909) );
  XOR2_X1 U9536 ( .A(n12225), .B(n12226), .Z(n6604) );
  INV_X1 U9537 ( .A(n12536), .ZN(n7408) );
  AND2_X1 U9538 ( .A1(n8962), .A2(n8961), .ZN(n13614) );
  INV_X1 U9539 ( .A(n13614), .ZN(n13884) );
  NOR2_X1 U9540 ( .A1(n11902), .A2(n6530), .ZN(n6605) );
  OR2_X1 U9541 ( .A1(n7753), .A2(n6459), .ZN(n6606) );
  INV_X1 U9542 ( .A(n11823), .ZN(n6964) );
  AND2_X1 U9543 ( .A1(n6770), .A2(n13905), .ZN(n6607) );
  AND3_X1 U9544 ( .A1(n8978), .A2(n8977), .A3(n8976), .ZN(n13868) );
  INV_X1 U9545 ( .A(n7804), .ZN(n7803) );
  AND2_X1 U9546 ( .A1(n6750), .A2(n6451), .ZN(n6608) );
  OR2_X1 U9547 ( .A1(n10459), .A2(n10452), .ZN(n6609) );
  AND2_X1 U9548 ( .A1(n7369), .A2(n7372), .ZN(n6610) );
  INV_X1 U9549 ( .A(SI_17_), .ZN(n10817) );
  NOR2_X1 U9550 ( .A1(n15265), .A2(n15088), .ZN(n6611) );
  INV_X1 U9551 ( .A(n13621), .ZN(n7811) );
  AND2_X1 U9552 ( .A1(n9190), .A2(n12069), .ZN(n6612) );
  NOR2_X1 U9553 ( .A1(n9751), .A2(n7771), .ZN(n6613) );
  INV_X1 U9554 ( .A(n9074), .ZN(n8685) );
  NOR2_X1 U9555 ( .A1(n9154), .A2(n11529), .ZN(n6614) );
  AND2_X1 U9556 ( .A1(n7032), .A2(n12191), .ZN(n6615) );
  NAND2_X1 U9557 ( .A1(n14444), .A2(n6973), .ZN(n9750) );
  AND2_X1 U9558 ( .A1(n6903), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6616) );
  OR2_X1 U9559 ( .A1(n9158), .A2(SI_23_), .ZN(n6617) );
  OR2_X1 U9560 ( .A1(n14988), .A2(n14231), .ZN(n6618) );
  AND2_X1 U9561 ( .A1(n14989), .A2(n14988), .ZN(n6619) );
  INV_X1 U9562 ( .A(n9071), .ZN(n7445) );
  OR2_X1 U9563 ( .A1(n12579), .A2(n12568), .ZN(n6620) );
  NOR2_X1 U9564 ( .A1(n7032), .A2(n12191), .ZN(n6621) );
  INV_X1 U9565 ( .A(n6700), .ZN(n6699) );
  NAND2_X1 U9566 ( .A1(n8358), .A2(n6706), .ZN(n6700) );
  AND2_X2 U9567 ( .A1(n10384), .A2(n10383), .ZN(n15384) );
  INV_X1 U9568 ( .A(n15384), .ZN(n6771) );
  INV_X1 U9569 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6904) );
  OR2_X1 U9570 ( .A1(n8358), .A2(n6704), .ZN(n6622) );
  NOR2_X1 U9571 ( .A1(n11045), .A2(n7193), .ZN(n11044) );
  NAND2_X1 U9572 ( .A1(n7334), .A2(n7340), .ZN(n7336) );
  AND2_X1 U9573 ( .A1(n7900), .A2(n7526), .ZN(n6623) );
  OR2_X1 U9574 ( .A1(n14601), .A2(n14600), .ZN(n6624) );
  AND2_X1 U9575 ( .A1(n14612), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6625) );
  INV_X1 U9576 ( .A(n6995), .ZN(n6994) );
  NAND2_X1 U9577 ( .A1(n7205), .A2(n6996), .ZN(n6995) );
  OR2_X1 U9578 ( .A1(n12697), .A2(n7211), .ZN(n6626) );
  NOR2_X1 U9579 ( .A1(n11654), .A2(n7548), .ZN(n11418) );
  NAND2_X1 U9580 ( .A1(n10481), .A2(n10480), .ZN(n11260) );
  OR2_X1 U9581 ( .A1(n11655), .A2(n15368), .ZN(n11654) );
  INV_X1 U9582 ( .A(n11654), .ZN(n7546) );
  OR2_X1 U9583 ( .A1(n10635), .A2(n7356), .ZN(n6627) );
  OR2_X1 U9584 ( .A1(n15312), .A2(n11500), .ZN(n6628) );
  INV_X1 U9585 ( .A(n7206), .ZN(n7205) );
  NOR2_X1 U9586 ( .A1(n12653), .A2(n15575), .ZN(n7206) );
  NAND2_X1 U9587 ( .A1(n7231), .A2(n10949), .ZN(n7235) );
  INV_X1 U9588 ( .A(SI_23_), .ZN(n11529) );
  INV_X1 U9589 ( .A(n6810), .ZN(n6809) );
  NOR2_X1 U9590 ( .A1(n11688), .A2(n11689), .ZN(n6810) );
  AND2_X1 U9591 ( .A1(n6803), .A2(n6802), .ZN(n6629) );
  INV_X1 U9592 ( .A(n6992), .ZN(n6990) );
  AOI21_X1 U9593 ( .B1(n6993), .B2(n6994), .A(n6455), .ZN(n6992) );
  NAND2_X1 U9594 ( .A1(n12666), .A2(n7206), .ZN(n6630) );
  AND2_X1 U9595 ( .A1(n7236), .A2(n7235), .ZN(n6631) );
  INV_X1 U9596 ( .A(n7525), .ZN(n7524) );
  OAI21_X1 U9597 ( .B1(n7900), .B2(n7526), .A(P1_DATAO_REG_24__SCAN_IN), .ZN(
        n7525) );
  OR2_X1 U9598 ( .A1(n6990), .A2(n6987), .ZN(n6632) );
  AND2_X1 U9599 ( .A1(n11647), .A2(n13397), .ZN(n6633) );
  AND2_X1 U9600 ( .A1(n7427), .A2(n7430), .ZN(n6634) );
  INV_X1 U9601 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7526) );
  INV_X1 U9602 ( .A(n12666), .ZN(n6996) );
  XOR2_X1 U9603 ( .A(n12653), .B(P3_REG2_REG_16__SCAN_IN), .Z(n6635) );
  AND2_X1 U9604 ( .A1(n6813), .A2(n6814), .ZN(n6636) );
  INV_X1 U9605 ( .A(n13541), .ZN(n13428) );
  OR2_X1 U9606 ( .A1(n13489), .A2(n11040), .ZN(n6637) );
  INV_X1 U9607 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n7417) );
  INV_X1 U9608 ( .A(n14246), .ZN(n14917) );
  AND2_X1 U9609 ( .A1(n7433), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n6638) );
  AND2_X1 U9610 ( .A1(n9346), .A2(n9345), .ZN(n6639) );
  INV_X1 U9611 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7086) );
  INV_X1 U9612 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n6832) );
  INV_X1 U9613 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7409) );
  INV_X1 U9614 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U9615 ( .A1(n15151), .A2(n15150), .ZN(n15154) );
  NAND2_X1 U9616 ( .A1(n12041), .A2(n8474), .ZN(n12853) );
  NAND2_X1 U9617 ( .A1(n12795), .A2(n12797), .ZN(n12794) );
  NAND2_X1 U9618 ( .A1(n7467), .A2(n7466), .ZN(n11216) );
  NAND2_X1 U9619 ( .A1(n6979), .A2(n6598), .ZN(n10626) );
  NAND2_X1 U9620 ( .A1(n6908), .A2(n7109), .ZN(n6907) );
  INV_X1 U9621 ( .A(n15151), .ZN(n6668) );
  NAND2_X1 U9622 ( .A1(n13564), .A2(n6641), .ZN(n7061) );
  NAND2_X1 U9623 ( .A1(n14932), .A2(n9490), .ZN(n14920) );
  NAND2_X1 U9624 ( .A1(n15211), .A2(n9387), .ZN(n11190) );
  INV_X1 U9625 ( .A(n14436), .ZN(n11051) );
  NAND2_X1 U9626 ( .A1(n7161), .A2(n14942), .ZN(n14932) );
  NAND2_X1 U9627 ( .A1(n7164), .A2(n7165), .ZN(n14779) );
  OAI211_X1 U9628 ( .C1(n14991), .C2(n15247), .A(n14990), .B(n6662), .ZN(
        n15085) );
  NOR2_X1 U9629 ( .A1(n6660), .A2(n9892), .ZN(n6659) );
  INV_X1 U9630 ( .A(n7922), .ZN(n7463) );
  XNOR2_X1 U9631 ( .A(n7296), .B(n9951), .ZN(n7295) );
  OAI21_X1 U9632 ( .B1(n8357), .B2(n12777), .A(n6575), .ZN(n7301) );
  NAND2_X1 U9633 ( .A1(n8430), .A2(n6590), .ZN(n6658) );
  NAND2_X1 U9634 ( .A1(n8415), .A2(n6643), .ZN(n8430) );
  AOI21_X1 U9635 ( .B1(n7291), .B2(n6568), .A(n7293), .ZN(n7289) );
  NOR2_X1 U9636 ( .A1(n6487), .A2(n8121), .ZN(n7292) );
  NAND3_X1 U9637 ( .A1(n7305), .A2(n11980), .A3(n7250), .ZN(n6947) );
  NAND2_X1 U9638 ( .A1(n6648), .A2(n6645), .ZN(n8356) );
  NAND2_X1 U9639 ( .A1(n6661), .A2(n6659), .ZN(n6648) );
  AOI21_X1 U9640 ( .B1(n7289), .B2(n7290), .A(n6595), .ZN(n7288) );
  NOR2_X1 U9641 ( .A1(n7292), .A2(n7294), .ZN(n7291) );
  INV_X1 U9642 ( .A(n6853), .ZN(n6852) );
  AND3_X2 U9643 ( .A1(n8780), .A2(n8812), .A3(n8778), .ZN(n6765) );
  AND3_X2 U9644 ( .A1(n8610), .A2(n8597), .A3(n6565), .ZN(n8696) );
  NAND2_X1 U9645 ( .A1(n8492), .A2(n8371), .ZN(n9899) );
  NAND2_X4 U9646 ( .A1(n8368), .A2(n8367), .ZN(n12779) );
  NAND2_X1 U9647 ( .A1(n7141), .A2(n12776), .ZN(n7139) );
  NAND2_X1 U9648 ( .A1(n8581), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8820) );
  AOI21_X1 U9649 ( .B1(n7801), .B2(n7799), .A(n6571), .ZN(n7798) );
  NAND2_X1 U9650 ( .A1(n6464), .A2(n7268), .ZN(n6734) );
  NAND2_X1 U9651 ( .A1(n15154), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7072) );
  OAI21_X1 U9652 ( .B1(n6482), .B2(n6655), .A(n8036), .ZN(n8049) );
  NAND2_X1 U9653 ( .A1(n7295), .A2(n7504), .ZN(n8580) );
  OR2_X1 U9654 ( .A1(n8218), .A2(n8217), .ZN(n8243) );
  INV_X1 U9655 ( .A(n7297), .ZN(n7985) );
  NAND3_X1 U9656 ( .A1(n7981), .A2(n8058), .A3(n6656), .ZN(n8185) );
  AOI21_X1 U9657 ( .B1(n6676), .B2(n12734), .A(n8379), .ZN(n8401) );
  OR3_X1 U9658 ( .A1(n8073), .A2(n8072), .A3(n10987), .ZN(n8090) );
  NAND2_X1 U9659 ( .A1(n7287), .A2(n7288), .ZN(n6657) );
  NAND2_X1 U9660 ( .A1(n6658), .A2(n8507), .ZN(n8431) );
  NAND2_X1 U9661 ( .A1(n6675), .A2(n6674), .ZN(n6661) );
  OAI211_X1 U9662 ( .C1(n6960), .C2(n6962), .A(n7777), .B(n6959), .ZN(n7774)
         );
  AOI21_X2 U9663 ( .B1(n14769), .B2(n14768), .A(n9771), .ZN(n14710) );
  NAND2_X1 U9664 ( .A1(n7115), .A2(n9546), .ZN(n12219) );
  NAND2_X2 U9665 ( .A1(n9764), .A2(n6512), .ZN(n7773) );
  NAND2_X1 U9666 ( .A1(n7770), .A2(n7199), .ZN(n11708) );
  INV_X1 U9667 ( .A(n15122), .ZN(n6663) );
  OAI21_X1 U9668 ( .B1(n13539), .B2(n15294), .A(n15313), .ZN(n6783) );
  NAND2_X1 U9669 ( .A1(n6784), .A2(n6782), .ZN(n6781) );
  NAND2_X1 U9670 ( .A1(n6781), .A2(n13541), .ZN(n6780) );
  NAND2_X1 U9671 ( .A1(n13537), .A2(n13536), .ZN(n13538) );
  INV_X1 U9672 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6664) );
  INV_X1 U9673 ( .A(n13519), .ZN(n6665) );
  XNOR2_X2 U9674 ( .A(n8718), .B(n8717), .ZN(n10541) );
  NAND3_X1 U9675 ( .A1(n7305), .A2(n7254), .A3(n11980), .ZN(n6666) );
  NAND2_X1 U9676 ( .A1(n14764), .A2(n14766), .ZN(n14765) );
  NAND2_X1 U9677 ( .A1(n9546), .A2(n7083), .ZN(n7190) );
  NAND2_X1 U9678 ( .A1(n7163), .A2(n7162), .ZN(n11956) );
  OR2_X1 U9679 ( .A1(n6926), .A2(n15142), .ZN(n6925) );
  NAND2_X1 U9680 ( .A1(n7614), .A2(n6567), .ZN(n7613) );
  INV_X1 U9681 ( .A(n7187), .ZN(n7188) );
  NAND2_X1 U9682 ( .A1(n14751), .A2(n14711), .ZN(n14730) );
  AOI21_X1 U9683 ( .B1(n7608), .B2(n7610), .A(n7606), .ZN(n7605) );
  XNOR2_X1 U9684 ( .A(n9090), .B(n9089), .ZN(n11113) );
  NAND3_X1 U9685 ( .A1(n6599), .A2(n15251), .A3(n14731), .ZN(n7185) );
  NAND2_X1 U9686 ( .A1(n13758), .A2(n13582), .ZN(n13738) );
  NOR2_X1 U9687 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8588) );
  NAND2_X1 U9688 ( .A1(n7711), .A2(n7326), .ZN(n7324) );
  NAND2_X1 U9689 ( .A1(n13590), .A2(n13589), .ZN(n13665) );
  NAND2_X1 U9690 ( .A1(n13906), .A2(n7059), .ZN(n13882) );
  NAND2_X1 U9691 ( .A1(n13679), .A2(n6493), .ZN(n13662) );
  AOI21_X2 U9692 ( .B1(n13649), .B2(n13650), .A(n13651), .ZN(n13955) );
  NAND2_X1 U9693 ( .A1(n7064), .A2(n13576), .ZN(n13794) );
  NAND2_X1 U9694 ( .A1(n6924), .A2(n7076), .ZN(n6923) );
  AOI22_X1 U9695 ( .A1(n7069), .A2(n11247), .B1(n11160), .B2(n7067), .ZN(n7066) );
  NAND3_X1 U9696 ( .A1(n12911), .A2(n12910), .A3(n6671), .ZN(n12965) );
  NAND2_X1 U9697 ( .A1(n7144), .A2(n7145), .ZN(n12796) );
  OAI21_X1 U9698 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n7747) );
  NOR2_X2 U9699 ( .A1(n7073), .A2(n6470), .ZN(n6932) );
  NAND2_X1 U9700 ( .A1(n7072), .A2(n15152), .ZN(n7073) );
  NAND2_X1 U9701 ( .A1(n13803), .A2(n13809), .ZN(n13783) );
  NAND2_X1 U9702 ( .A1(n7065), .A2(n7066), .ZN(n11172) );
  INV_X1 U9703 ( .A(n7551), .ZN(n7550) );
  OAI21_X1 U9704 ( .B1(n10549), .B2(n8968), .A(n8991), .ZN(n8993) );
  INV_X1 U9705 ( .A(n11873), .ZN(n7026) );
  NAND2_X1 U9706 ( .A1(n12448), .A2(n12170), .ZN(n12173) );
  AOI21_X1 U9707 ( .B1(n10798), .B2(n10804), .A(n10895), .ZN(n10893) );
  INV_X2 U9708 ( .A(n10809), .ZN(n7223) );
  NAND2_X1 U9709 ( .A1(n10902), .A2(n10809), .ZN(n10801) );
  AND4_X2 U9710 ( .A1(n7492), .A2(n7739), .A3(n7494), .A4(n7493), .ZN(n10809)
         );
  NAND3_X1 U9711 ( .A1(n8300), .A2(n7149), .A3(n12822), .ZN(n6675) );
  NAND2_X1 U9712 ( .A1(n8432), .A2(n10430), .ZN(n7506) );
  NAND2_X1 U9713 ( .A1(n8377), .A2(n8378), .ZN(n6676) );
  INV_X1 U9714 ( .A(n6932), .ZN(n15161) );
  NAND2_X1 U9715 ( .A1(n7071), .A2(n7068), .ZN(n7065) );
  XNOR2_X1 U9716 ( .A(n6930), .B(n6525), .ZN(SUB_1596_U4) );
  NAND2_X1 U9717 ( .A1(n7129), .A2(n7941), .ZN(n7992) );
  NAND2_X1 U9718 ( .A1(n8252), .A2(n7939), .ZN(n8293) );
  NAND2_X1 U9719 ( .A1(n7107), .A2(n7940), .ZN(n8346) );
  INV_X1 U9720 ( .A(n7130), .ZN(n7962) );
  NAND2_X2 U9721 ( .A1(n7967), .A2(n7966), .ZN(n12744) );
  AND4_X2 U9722 ( .A1(n9357), .A2(n9355), .A3(n9356), .A4(n9354), .ZN(n14258)
         );
  NAND2_X1 U9723 ( .A1(n7505), .A2(n8549), .ZN(n7296) );
  NAND2_X1 U9724 ( .A1(n8431), .A2(n9936), .ZN(n7507) );
  NAND2_X1 U9725 ( .A1(n7301), .A2(n7299), .ZN(n7298) );
  NAND2_X1 U9726 ( .A1(n7298), .A2(n6581), .ZN(n8377) );
  OAI22_X1 U9727 ( .A1(n13232), .A2(n6688), .B1(n13233), .B2(n6687), .ZN(
        n13237) );
  OAI21_X1 U9728 ( .B1(n13237), .B2(n7644), .A(n7643), .ZN(n13242) );
  NAND2_X1 U9729 ( .A1(n7499), .A2(n6692), .ZN(n6689) );
  NAND2_X1 U9730 ( .A1(n7499), .A2(n7497), .ZN(n8268) );
  NAND2_X1 U9731 ( .A1(n6689), .A2(n6690), .ZN(n8324) );
  NAND2_X1 U9732 ( .A1(n8341), .A2(n6706), .ZN(n6705) );
  OAI211_X1 U9733 ( .C1(n8341), .C2(n6622), .A(n6701), .B(n6695), .ZN(n11526)
         );
  NAND2_X1 U9734 ( .A1(n8341), .A2(n6699), .ZN(n6695) );
  OAI211_X1 U9735 ( .C1(n8341), .C2(n6698), .A(n8437), .B(n6696), .ZN(n8361)
         );
  NAND2_X1 U9736 ( .A1(n8341), .A2(n6697), .ZN(n6696) );
  NAND2_X1 U9737 ( .A1(n8341), .A2(n7898), .ZN(n8000) );
  NAND4_X1 U9738 ( .A1(n7511), .A2(n7869), .A3(n7868), .A4(n6439), .ZN(n6710)
         );
  NAND3_X1 U9739 ( .A1(n6710), .A2(n6709), .A3(n6712), .ZN(n8172) );
  NAND3_X1 U9740 ( .A1(n7513), .A2(n7511), .A3(n6439), .ZN(n6709) );
  INV_X1 U9741 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U9742 ( .A1(n13299), .A2(n6432), .ZN(n6717) );
  NAND2_X1 U9743 ( .A1(n6717), .A2(n6718), .ZN(n13306) );
  OAI21_X1 U9744 ( .B1(n8184), .B2(n6727), .A(n6723), .ZN(n8245) );
  NAND3_X1 U9745 ( .A1(n12901), .A2(n7134), .A3(n7135), .ZN(n12951) );
  NAND2_X1 U9746 ( .A1(n6731), .A2(n13642), .ZN(n13644) );
  OAI21_X1 U9747 ( .B1(n13658), .B2(n13657), .A(n6731), .ZN(n13952) );
  NAND2_X1 U9748 ( .A1(n6734), .A2(n15384), .ZN(n7267) );
  NAND2_X1 U9749 ( .A1(n6733), .A2(n6732), .ZN(P2_U3528) );
  OR2_X1 U9750 ( .A1(n15390), .A2(n9292), .ZN(n6732) );
  NAND2_X1 U9751 ( .A1(n6734), .A2(n15390), .ZN(n6733) );
  NAND2_X1 U9752 ( .A1(n9002), .A2(n7848), .ZN(n8676) );
  AOI21_X1 U9753 ( .B1(n6741), .B2(n7612), .A(n7114), .ZN(n6740) );
  MUX2_X1 U9754 ( .A(n10185), .B(n10187), .S(n10065), .Z(n8658) );
  NAND2_X1 U9755 ( .A1(n9157), .A2(n7108), .ZN(n9175) );
  OAI21_X2 U9756 ( .B1(n11786), .B2(n13558), .A(n6753), .ZN(n13607) );
  NAND2_X1 U9757 ( .A1(n6755), .A2(n13616), .ZN(n6760) );
  NAND2_X1 U9758 ( .A1(n6762), .A2(n13589), .ZN(n13957) );
  AND2_X2 U9759 ( .A1(n8737), .A2(n8738), .ZN(n8779) );
  AND2_X2 U9760 ( .A1(n6765), .A2(n8593), .ZN(n8597) );
  NAND3_X1 U9761 ( .A1(n7843), .A2(n8610), .A3(n6763), .ZN(n14085) );
  NAND3_X1 U9762 ( .A1(n6773), .A2(n13959), .A3(n6772), .ZN(n14061) );
  NAND3_X1 U9763 ( .A1(n6785), .A2(n6780), .A3(n6778), .ZN(P2_U3233) );
  INV_X1 U9764 ( .A(n13520), .ZN(n6808) );
  INV_X1 U9765 ( .A(n6813), .ZN(n6812) );
  NAND3_X1 U9766 ( .A1(n15278), .A2(n6819), .A3(n15276), .ZN(n6813) );
  INV_X1 U9767 ( .A(n13493), .ZN(n6819) );
  NAND2_X1 U9768 ( .A1(n12609), .A2(n6825), .ZN(n6822) );
  NAND3_X1 U9769 ( .A1(n12595), .A2(n12608), .A3(n12549), .ZN(n6823) );
  NAND2_X1 U9770 ( .A1(n12595), .A2(n12549), .ZN(n6826) );
  OAI21_X1 U9771 ( .B1(n11932), .B2(n6839), .A(n6838), .ZN(n14622) );
  XNOR2_X1 U9772 ( .A(n14622), .B(n14628), .ZN(n14615) );
  NAND3_X1 U9773 ( .A1(n6850), .A2(n6849), .A3(n6846), .ZN(P1_U3262) );
  NAND3_X1 U9774 ( .A1(n14632), .A2(n14634), .A3(n14633), .ZN(n6851) );
  NAND2_X1 U9775 ( .A1(n13167), .A2(n9212), .ZN(n13042) );
  NAND2_X1 U9776 ( .A1(n6492), .A2(n8610), .ZN(n6869) );
  INV_X2 U9777 ( .A(n8772), .ZN(n13889) );
  NAND2_X1 U9778 ( .A1(n12521), .A2(n11024), .ZN(n6872) );
  INV_X1 U9779 ( .A(n15403), .ZN(n11024) );
  NAND2_X1 U9780 ( .A1(n8017), .A2(n15403), .ZN(n8456) );
  OAI211_X2 U9781 ( .C1(n8389), .C2(n10122), .A(n6876), .B(n6873), .ZN(n15403)
         );
  INV_X1 U9782 ( .A(n10727), .ZN(n6874) );
  NAND2_X1 U9783 ( .A1(n11441), .A2(n6878), .ZN(n6877) );
  NAND2_X1 U9784 ( .A1(n6877), .A2(n6879), .ZN(n11798) );
  NAND2_X1 U9785 ( .A1(n8473), .A2(n6888), .ZN(n12041) );
  NAND2_X1 U9786 ( .A1(n8498), .A2(n8497), .ZN(n12731) );
  NAND2_X1 U9787 ( .A1(n7485), .A2(n8499), .ZN(n6896) );
  NAND2_X1 U9788 ( .A1(n6895), .A2(n6894), .ZN(n12900) );
  NAND2_X1 U9789 ( .A1(n7485), .A2(n7486), .ZN(n6894) );
  NAND2_X1 U9790 ( .A1(n9619), .A2(n6897), .ZN(n9672) );
  NAND2_X1 U9791 ( .A1(n9619), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U9792 ( .A1(n6902), .A2(n6596), .ZN(n9423) );
  NAND2_X1 U9793 ( .A1(n9497), .A2(n6616), .ZN(n9537) );
  INV_X1 U9794 ( .A(n6916), .ZN(n6915) );
  XNOR2_X1 U9795 ( .A(n12631), .B(n12630), .ZN(n12607) );
  INV_X1 U9796 ( .A(n6920), .ZN(n12629) );
  NAND2_X1 U9797 ( .A1(n12631), .A2(n12630), .ZN(n6919) );
  NAND2_X1 U9798 ( .A1(n6923), .A2(n6922), .ZN(n6921) );
  NOR2_X1 U9799 ( .A1(n6926), .A2(n15141), .ZN(n6924) );
  OAI21_X2 U9800 ( .B1(n6932), .B2(n6931), .A(n7074), .ZN(n6930) );
  NAND2_X1 U9801 ( .A1(n9691), .A2(n6933), .ZN(n9700) );
  NAND2_X1 U9802 ( .A1(n6935), .A2(n6934), .ZN(n14382) );
  NAND3_X1 U9803 ( .A1(n6539), .A2(n7257), .A3(n7256), .ZN(n6934) );
  OAI211_X1 U9804 ( .C1(n7257), .C2(n7391), .A(n6937), .B(n14380), .ZN(n14383)
         );
  NAND2_X1 U9805 ( .A1(n7256), .A2(n7849), .ZN(n6939) );
  NAND2_X1 U9806 ( .A1(n6563), .A2(n14350), .ZN(n6944) );
  NAND2_X1 U9807 ( .A1(n14310), .A2(n6945), .ZN(n6942) );
  NAND2_X1 U9808 ( .A1(n14311), .A2(n6945), .ZN(n6943) );
  NAND4_X1 U9809 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6940), .ZN(n7258)
         );
  NOR2_X1 U9810 ( .A1(n6496), .A2(n6941), .ZN(n6940) );
  OAI211_X1 U9811 ( .C1(n6954), .C2(n6951), .A(n6948), .B(n6953), .ZN(n14459)
         );
  NAND3_X1 U9812 ( .A1(n7279), .A2(n6592), .A3(n7280), .ZN(n6954) );
  OAI211_X1 U9813 ( .C1(n6958), .C2(n14286), .A(n6957), .B(n6955), .ZN(n7393)
         );
  NAND3_X1 U9814 ( .A1(n14286), .A2(n7382), .A3(n7383), .ZN(n6956) );
  NAND2_X1 U9815 ( .A1(n7394), .A2(n14288), .ZN(n6957) );
  INV_X1 U9816 ( .A(n7773), .ZN(n6960) );
  OAI21_X1 U9817 ( .B1(n6964), .B2(n6966), .A(n6967), .ZN(n14937) );
  OAI211_X1 U9818 ( .C1(n11823), .C2(n6968), .A(n6965), .B(n9759), .ZN(n6969)
         );
  INV_X1 U9819 ( .A(n7779), .ZN(n6966) );
  NAND2_X1 U9820 ( .A1(n6969), .A2(n9760), .ZN(n14913) );
  NAND4_X1 U9821 ( .A1(n7079), .A2(n7111), .A3(n8633), .A4(n8636), .ZN(n6971)
         );
  AND2_X1 U9822 ( .A1(n6971), .A2(n6970), .ZN(n8810) );
  NAND3_X1 U9823 ( .A1(n6971), .A2(n8637), .A3(n6970), .ZN(n7159) );
  NAND2_X1 U9824 ( .A1(n6972), .A2(n8636), .ZN(n6970) );
  NAND2_X1 U9825 ( .A1(n6562), .A2(n7079), .ZN(n8777) );
  INV_X1 U9826 ( .A(n8776), .ZN(n6972) );
  NAND4_X1 U9827 ( .A1(n9428), .A2(n9426), .A3(n9429), .A4(n9427), .ZN(n14493)
         );
  NAND2_X1 U9828 ( .A1(n11378), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U9829 ( .A1(n11136), .A2(n11135), .ZN(n6978) );
  NAND2_X1 U9830 ( .A1(n6981), .A2(n10609), .ZN(n6980) );
  NAND2_X1 U9831 ( .A1(n6980), .A2(n10725), .ZN(n6979) );
  NAND2_X1 U9832 ( .A1(n6981), .A2(n10609), .ZN(n10726) );
  NAND2_X1 U9833 ( .A1(n10870), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U9834 ( .A1(n10648), .A2(n10647), .ZN(n6982) );
  NAND2_X1 U9835 ( .A1(n12628), .A2(n6984), .ZN(n6983) );
  OR2_X4 U9836 ( .A1(n14247), .A2(n14251), .ZN(n14248) );
  AND2_X2 U9837 ( .A1(n9701), .A2(n9700), .ZN(n14251) );
  XNOR2_X2 U9838 ( .A(n7004), .B(n9692), .ZN(n14247) );
  NAND3_X1 U9839 ( .A1(n7006), .A2(n7005), .A3(n11355), .ZN(n10858) );
  AND2_X1 U9840 ( .A1(n10746), .A2(n10747), .ZN(n7005) );
  INV_X1 U9841 ( .A(n7007), .ZN(n15173) );
  AOI21_X2 U9842 ( .B1(n11551), .B2(n11364), .A(n11363), .ZN(n11367) );
  AND2_X2 U9843 ( .A1(n7007), .A2(n6561), .ZN(n11551) );
  OR2_X2 U9844 ( .A1(n15175), .A2(n15176), .ZN(n7007) );
  OAI22_X1 U9845 ( .A1(n11339), .A2(n11338), .B1(n11337), .B2(n11336), .ZN(
        n15175) );
  NAND3_X1 U9846 ( .A1(n11847), .A2(n6572), .A3(n7828), .ZN(n7694) );
  NAND2_X1 U9847 ( .A1(n14177), .A2(n7015), .ZN(n7012) );
  NAND2_X1 U9848 ( .A1(n7012), .A2(n7013), .ZN(n14193) );
  NAND2_X1 U9849 ( .A1(n7023), .A2(n7021), .ZN(n7020) );
  OAI21_X1 U9850 ( .B1(n14224), .B2(n7022), .A(n7018), .ZN(n7021) );
  NAND2_X1 U9851 ( .A1(n14224), .A2(n12297), .ZN(n7018) );
  OAI211_X1 U9852 ( .C1(n14151), .C2(n7020), .A(n7019), .B(n14232), .ZN(n7098)
         );
  NAND3_X1 U9853 ( .A1(n14151), .A2(n7021), .A3(n6601), .ZN(n7019) );
  NAND3_X1 U9854 ( .A1(n7027), .A2(n10805), .A3(n7235), .ZN(n7234) );
  INV_X1 U9855 ( .A(n10893), .ZN(n7027) );
  NAND2_X1 U9856 ( .A1(n7220), .A2(n7222), .ZN(n7219) );
  NAND2_X1 U9857 ( .A1(n12437), .A2(n7574), .ZN(n12369) );
  NAND2_X1 U9858 ( .A1(n12369), .A2(n6615), .ZN(n7030) );
  NAND2_X1 U9859 ( .A1(n7031), .A2(n7030), .ZN(n12456) );
  AOI21_X1 U9860 ( .B1(n12437), .B2(n6447), .A(n6621), .ZN(n7031) );
  NAND2_X1 U9861 ( .A1(n12369), .A2(n12191), .ZN(n12351) );
  INV_X1 U9862 ( .A(n12350), .ZN(n7032) );
  INV_X1 U9863 ( .A(n7240), .ZN(n7038) );
  NAND2_X1 U9864 ( .A1(n7982), .A2(n7041), .ZN(n8555) );
  NAND2_X1 U9865 ( .A1(n7040), .A2(n7982), .ZN(n8564) );
  NAND2_X2 U9866 ( .A1(n13613), .A2(n6466), .ZN(n13616) );
  NAND2_X1 U9867 ( .A1(n7817), .A2(n7052), .ZN(n7051) );
  INV_X1 U9868 ( .A(n13636), .ZN(n7053) );
  AOI21_X1 U9869 ( .B1(n8642), .B2(n7058), .A(n7057), .ZN(n7055) );
  NAND2_X1 U9870 ( .A1(n7054), .A2(n7274), .ZN(n7271) );
  NAND2_X1 U9871 ( .A1(n7158), .A2(n8641), .ZN(n8832) );
  NAND3_X1 U9872 ( .A1(n7061), .A2(n7060), .A3(n13913), .ZN(n13906) );
  NAND3_X1 U9873 ( .A1(n7309), .A2(n6449), .A3(n7310), .ZN(n7064) );
  NAND2_X2 U9874 ( .A1(n11172), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7246) );
  INV_X1 U9875 ( .A(n11164), .ZN(n7069) );
  AND2_X1 U9876 ( .A1(n11164), .A2(n7070), .ZN(n7068) );
  NAND2_X1 U9877 ( .A1(n15161), .A2(n7074), .ZN(n15160) );
  NAND2_X1 U9878 ( .A1(n12785), .A2(n8487), .ZN(n12774) );
  NAND2_X1 U9879 ( .A1(n8462), .A2(n8461), .ZN(n11441) );
  NAND2_X1 U9880 ( .A1(n7078), .A2(n13438), .ZN(P2_U3328) );
  OAI21_X1 U9881 ( .B1(n7623), .B2(n13432), .A(n13433), .ZN(n7078) );
  NAND2_X1 U9882 ( .A1(n7453), .A2(n8596), .ZN(n7455) );
  NAND2_X1 U9883 ( .A1(n13248), .A2(n6584), .ZN(n7625) );
  OR2_X1 U9884 ( .A1(n13242), .A2(n13243), .ZN(n13244) );
  NAND2_X1 U9885 ( .A1(n13431), .A2(n13430), .ZN(n7624) );
  NAND2_X1 U9886 ( .A1(n13221), .A2(n13222), .ZN(n13220) );
  INV_X1 U9887 ( .A(n7157), .ZN(n7156) );
  NAND2_X1 U9888 ( .A1(n8623), .A2(n8622), .ZN(n7079) );
  INV_X1 U9889 ( .A(n7710), .ZN(n7709) );
  NAND2_X1 U9890 ( .A1(n7159), .A2(n8639), .ZN(n8797) );
  INV_X1 U9891 ( .A(n8693), .ZN(n7112) );
  INV_X1 U9892 ( .A(n8736), .ZN(n8625) );
  OAI21_X2 U9893 ( .B1(n12085), .B2(n7696), .A(n7695), .ZN(n14189) );
  NOR2_X1 U9894 ( .A1(n12244), .A2(n6499), .ZN(n14127) );
  NAND2_X1 U9895 ( .A1(n12080), .A2(n12079), .ZN(n14204) );
  INV_X1 U9896 ( .A(n14204), .ZN(n12085) );
  NAND2_X1 U9897 ( .A1(n14398), .A2(n14399), .ZN(n14397) );
  NAND2_X1 U9898 ( .A1(n8890), .A2(n8651), .ZN(n8908) );
  NAND4_X2 U9899 ( .A1(n7085), .A2(n9351), .A3(n9352), .A4(n9353), .ZN(n14499)
         );
  OAI21_X1 U9900 ( .B1(n8714), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7127), .ZN(
        n8736) );
  XNOR2_X1 U9901 ( .A(n14255), .B(n14414), .ZN(n14257) );
  AOI21_X1 U9902 ( .B1(n14273), .B2(n14274), .A(n14272), .ZN(n14275) );
  XNOR2_X2 U9903 ( .A(n11163), .B(n11161), .ZN(n11160) );
  NAND2_X2 U9904 ( .A1(n10718), .A2(n10717), .ZN(n11163) );
  NAND2_X1 U9905 ( .A1(n7245), .A2(n7246), .ZN(n7248) );
  AND2_X2 U9906 ( .A1(n8616), .A2(n8589), .ZN(n8610) );
  NAND2_X1 U9907 ( .A1(n15185), .A2(n15184), .ZN(n10254) );
  NAND2_X1 U9908 ( .A1(n10250), .A2(n10251), .ZN(n15185) );
  INV_X1 U9909 ( .A(n7359), .ZN(n7355) );
  NOR2_X1 U9910 ( .A1(n12582), .A2(n6574), .ZN(n12605) );
  XNOR2_X1 U9911 ( .A(n9371), .B(n9319), .ZN(n14538) );
  NAND2_X1 U9912 ( .A1(n7712), .A2(n6587), .ZN(n13776) );
  OAI211_X1 U9913 ( .C1(n8625), .C2(SI_2_), .A(n8756), .B(n8624), .ZN(n7111)
         );
  NAND2_X1 U9914 ( .A1(n8714), .A2(n10089), .ZN(n7127) );
  OR3_X1 U9915 ( .A1(n13563), .A2(n13406), .A3(n13405), .ZN(n13407) );
  NAND2_X1 U9916 ( .A1(n7271), .A2(n7272), .ZN(n8890) );
  XNOR2_X1 U9917 ( .A(n7598), .B(n13428), .ZN(n13418) );
  AOI21_X1 U9918 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n10860) );
  AOI21_X1 U9919 ( .B1(n10862), .B2(n10861), .A(n10860), .ZN(n11339) );
  NAND2_X1 U9920 ( .A1(n11541), .A2(n11540), .ZN(n11847) );
  NAND2_X1 U9921 ( .A1(n11536), .A2(n7838), .ZN(n11541) );
  NAND2_X1 U9922 ( .A1(n7098), .A2(n7097), .ZN(P1_U3240) );
  NAND2_X1 U9923 ( .A1(n7604), .A2(n7605), .ZN(n9002) );
  NOR2_X1 U9924 ( .A1(n7835), .A2(n7825), .ZN(n7824) );
  XNOR2_X1 U9925 ( .A(n9342), .B(n9341), .ZN(n14503) );
  INV_X1 U9926 ( .A(n8083), .ZN(n8084) );
  NAND2_X1 U9927 ( .A1(n7402), .A2(n7403), .ZN(n12648) );
  NAND2_X1 U9928 ( .A1(n7154), .A2(n12719), .ZN(n12724) );
  INV_X1 U9929 ( .A(n7129), .ZN(n8363) );
  INV_X1 U9930 ( .A(n7428), .ZN(n7424) );
  NOR2_X2 U9931 ( .A1(n8329), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7107) );
  AND3_X2 U9932 ( .A1(n8014), .A2(n8081), .A3(n7459), .ZN(n7738) );
  NAND2_X1 U9933 ( .A1(n7218), .A2(n7217), .ZN(n7946) );
  NAND2_X2 U9934 ( .A1(n7156), .A2(n7227), .ZN(n12055) );
  NAND2_X1 U9935 ( .A1(n8031), .A2(n8030), .ZN(n7128) );
  NAND2_X1 U9936 ( .A1(n9830), .A2(n9829), .ZN(n9833) );
  NAND2_X1 U9937 ( .A1(n9072), .A2(n8682), .ZN(n7264) );
  NAND2_X1 U9938 ( .A1(n12562), .A2(n12561), .ZN(n7204) );
  NAND2_X1 U9939 ( .A1(n12615), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12625) );
  XNOR2_X1 U9940 ( .A(n12693), .B(n12699), .ZN(n7110) );
  INV_X1 U9941 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U9942 ( .A1(n9131), .A2(n8689), .ZN(n7285) );
  NAND2_X1 U9943 ( .A1(n7324), .A2(n7322), .ZN(n13679) );
  INV_X1 U9944 ( .A(n7611), .ZN(n7114) );
  NAND2_X1 U9945 ( .A1(n11048), .A2(n14436), .ZN(n9743) );
  AND2_X1 U9946 ( .A1(n9329), .A2(n7786), .ZN(n7115) );
  NAND4_X1 U9947 ( .A1(n7196), .A2(n7840), .A3(n9359), .A4(n7195), .ZN(n7194)
         );
  NAND3_X1 U9948 ( .A1(n9328), .A2(n9545), .A3(n9396), .ZN(n9696) );
  NAND3_X1 U9949 ( .A1(n14403), .A2(n6589), .A3(n14402), .ZN(n7279) );
  NAND2_X1 U9950 ( .A1(n11668), .A2(n11667), .ZN(n7123) );
  NAND2_X1 U9951 ( .A1(n7285), .A2(n8691), .ZN(n9153) );
  NAND2_X1 U9952 ( .A1(n7267), .A2(n7265), .ZN(P2_U3496) );
  INV_X1 U9953 ( .A(n7269), .ZN(n7268) );
  NAND2_X1 U9954 ( .A1(n14382), .A2(n14381), .ZN(n7124) );
  NAND2_X1 U9955 ( .A1(n7607), .A2(n8664), .ZN(n8968) );
  NAND3_X1 U9956 ( .A1(n7126), .A2(n7125), .A3(n14467), .ZN(n14470) );
  NAND3_X1 U9957 ( .A1(n14459), .A2(n14457), .A3(n14458), .ZN(n7126) );
  NAND3_X1 U9958 ( .A1(n8033), .A2(n7128), .A3(n6566), .ZN(n10699) );
  NAND2_X1 U9959 ( .A1(n7218), .A2(n7736), .ZN(n7922) );
  NAND2_X1 U9960 ( .A1(n8032), .A2(SI_0_), .ZN(n8033) );
  NAND2_X1 U9961 ( .A1(n7919), .A2(n7918), .ZN(n7921) );
  NAND2_X1 U9962 ( .A1(n7463), .A2(n7923), .ZN(n7462) );
  XNOR2_X2 U9963 ( .A(n9362), .B(n9361), .ZN(n14522) );
  NAND2_X2 U9964 ( .A1(n9715), .A2(n9716), .ZN(n10758) );
  NAND2_X4 U9965 ( .A1(n10193), .A2(n10065), .ZN(n13369) );
  INV_X1 U9966 ( .A(n13914), .ZN(n13613) );
  NAND2_X1 U9967 ( .A1(n6526), .A2(n13793), .ZN(n7817) );
  OAI211_X1 U9968 ( .C1(n13948), .C2(n15381), .A(n7542), .B(n7270), .ZN(n7269)
         );
  NOR2_X2 U9969 ( .A1(n6456), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7129) );
  NAND2_X1 U9970 ( .A1(n12900), .A2(n15395), .ZN(n7135) );
  NAND2_X1 U9971 ( .A1(n8558), .A2(n8559), .ZN(n7735) );
  XNOR2_X2 U9972 ( .A(n10176), .B(n10174), .ZN(n10173) );
  INV_X1 U9973 ( .A(n10699), .ZN(n10823) );
  NAND2_X1 U9974 ( .A1(n11798), .A2(n11800), .ZN(n8468) );
  OR2_X1 U9975 ( .A1(n12776), .A2(n7759), .ZN(n7143) );
  NAND2_X1 U9976 ( .A1(n7143), .A2(n7757), .ZN(n12751) );
  NAND2_X1 U9977 ( .A1(n12831), .A2(n6419), .ZN(n7144) );
  NAND2_X1 U9978 ( .A1(n9883), .A2(n9882), .ZN(n7153) );
  NAND2_X1 U9979 ( .A1(n8797), .A2(n7593), .ZN(n7158) );
  NAND3_X1 U9980 ( .A1(n11704), .A2(n9439), .A3(n6582), .ZN(n7163) );
  NAND2_X1 U9981 ( .A1(n11956), .A2(n14938), .ZN(n7161) );
  NAND2_X1 U9982 ( .A1(n14854), .A2(n7167), .ZN(n7164) );
  NAND2_X1 U9983 ( .A1(n14710), .A2(n6578), .ZN(n7177) );
  NAND2_X1 U9984 ( .A1(n14710), .A2(n7179), .ZN(n7183) );
  NAND2_X1 U9985 ( .A1(n7183), .A2(n7182), .ZN(n14703) );
  AND2_X1 U9986 ( .A1(n14738), .A2(n7188), .ZN(n15087) );
  OAI21_X1 U9987 ( .B1(n14738), .B2(n15264), .A(n7186), .ZN(P1_U3520) );
  NAND2_X1 U9988 ( .A1(n14765), .A2(n9616), .ZN(n14748) );
  NAND2_X1 U9989 ( .A1(n7194), .A2(n7193), .ZN(n7852) );
  AND2_X4 U9990 ( .A1(n9332), .A2(n9333), .ZN(n9966) );
  INV_X2 U9991 ( .A(n14268), .ZN(n7193) );
  NAND3_X1 U9992 ( .A1(n7197), .A2(n7198), .A3(n8626), .ZN(n9346) );
  NAND2_X2 U9993 ( .A1(n12625), .A2(n12626), .ZN(n12628) );
  NOR2_X2 U9994 ( .A1(n7737), .A2(n7980), .ZN(n7736) );
  NOR2_X2 U9996 ( .A1(n7911), .A2(n7735), .ZN(n7734) );
  INV_X1 U9997 ( .A(n10795), .ZN(n7221) );
  NAND2_X2 U9998 ( .A1(n7219), .A2(n10797), .ZN(n10800) );
  MUX2_X1 U9999 ( .A(n10802), .B(n10801), .S(n10800), .Z(n10805) );
  NAND2_X1 U10000 ( .A1(n12495), .A2(n12493), .ZN(n7224) );
  NAND2_X1 U10001 ( .A1(n12342), .A2(n12341), .ZN(n7225) );
  INV_X1 U10002 ( .A(n7952), .ZN(n13024) );
  AND2_X2 U10003 ( .A1(n12056), .A2(n7952), .ZN(n8050) );
  NAND2_X1 U10004 ( .A1(n10944), .A2(n7235), .ZN(n7233) );
  AOI21_X1 U10005 ( .B1(n7236), .B2(n7232), .A(n6580), .ZN(n11020) );
  NAND2_X1 U10006 ( .A1(n7234), .A2(n7233), .ZN(n7232) );
  INV_X1 U10007 ( .A(n10947), .ZN(n7236) );
  INV_X1 U10008 ( .A(n10944), .ZN(n7237) );
  INV_X1 U10009 ( .A(n12018), .ZN(n12015) );
  NAND2_X1 U10010 ( .A1(n10042), .A2(n10041), .ZN(n10045) );
  NAND2_X1 U10011 ( .A1(n10067), .A2(n14531), .ZN(n10070) );
  NAND2_X1 U10012 ( .A1(n10055), .A2(n10054), .ZN(n7244) );
  AOI21_X2 U10013 ( .B1(n7246), .B2(n7247), .A(n6494), .ZN(n11938) );
  NAND3_X1 U10014 ( .A1(n7259), .A2(n7389), .A3(n7258), .ZN(n7257) );
  INV_X1 U10015 ( .A(n14374), .ZN(n7259) );
  MUX2_X1 U10016 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n10065), .Z(n8640) );
  NAND2_X2 U10017 ( .A1(n7262), .A2(n9575), .ZN(n15028) );
  OR2_X1 U10018 ( .A1(n14410), .A2(n7281), .ZN(n7278) );
  NAND2_X1 U10019 ( .A1(n14410), .A2(n7281), .ZN(n7280) );
  NAND2_X1 U10020 ( .A1(n7285), .A2(n7283), .ZN(n9157) );
  NAND2_X1 U10021 ( .A1(n8107), .A2(n7289), .ZN(n7287) );
  INV_X2 U10022 ( .A(n10430), .ZN(n9936) );
  MUX2_X1 U10023 ( .A(n8047), .B(n10801), .S(n10430), .Z(n8048) );
  AND2_X4 U10024 ( .A1(n10983), .A2(n11314), .ZN(n10430) );
  XNOR2_X2 U10025 ( .A(n7984), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11314) );
  INV_X1 U10026 ( .A(n7302), .ZN(n10079) );
  OR2_X2 U10027 ( .A1(n10080), .A2(n10081), .ZN(n7302) );
  NAND2_X1 U10028 ( .A1(n11939), .A2(n11938), .ZN(n11947) );
  NAND3_X1 U10029 ( .A1(n7702), .A2(n7700), .A3(n11080), .ZN(n7339) );
  NAND3_X1 U10030 ( .A1(n7333), .A2(n7332), .A3(n6558), .ZN(n11738) );
  NAND3_X1 U10031 ( .A1(n7338), .A2(n7336), .A3(n6420), .ZN(n7332) );
  NAND4_X1 U10032 ( .A1(n7702), .A2(n6600), .A3(n7700), .A4(n7336), .ZN(n7333)
         );
  INV_X1 U10033 ( .A(n13401), .ZN(n7334) );
  INV_X1 U10034 ( .A(n7343), .ZN(n8932) );
  AND3_X1 U10035 ( .A1(n8610), .A2(n7843), .A3(n7049), .ZN(n7342) );
  AOI21_X1 U10036 ( .B1(n10635), .B2(n10634), .A(n7367), .ZN(n10645) );
  INV_X1 U10037 ( .A(n7367), .ZN(n7362) );
  NAND2_X1 U10038 ( .A1(n10876), .A2(n10877), .ZN(n7366) );
  AND2_X1 U10039 ( .A1(n10632), .A2(n10633), .ZN(n7367) );
  NAND3_X1 U10040 ( .A1(n14257), .A2(n14437), .A3(n14256), .ZN(n7378) );
  AND2_X2 U10041 ( .A1(n9320), .A2(n6579), .ZN(n9396) );
  NAND4_X1 U10042 ( .A1(n7715), .A2(n9396), .A3(n9328), .A4(n7716), .ZN(n9710)
         );
  NOR2_X2 U10043 ( .A1(n9520), .A2(n9327), .ZN(n9328) );
  NAND4_X1 U10044 ( .A1(n9323), .A2(n9324), .A3(n9322), .A4(n9321), .ZN(n9520)
         );
  INV_X1 U10045 ( .A(n14293), .ZN(n7381) );
  NAND2_X1 U10046 ( .A1(n14282), .A2(n7384), .ZN(n7383) );
  NAND2_X1 U10047 ( .A1(n7393), .A2(n7392), .ZN(n14291) );
  OR2_X1 U10048 ( .A1(n14288), .A2(n7394), .ZN(n7392) );
  INV_X1 U10049 ( .A(n14287), .ZN(n7394) );
  NAND3_X1 U10050 ( .A1(n7399), .A2(n9347), .A3(n7398), .ZN(n7397) );
  NAND2_X1 U10051 ( .A1(n10110), .A2(n7401), .ZN(n7398) );
  NAND2_X2 U10052 ( .A1(n9347), .A2(n6410), .ZN(n9384) );
  NAND2_X1 U10053 ( .A1(n12610), .A2(n12639), .ZN(n7402) );
  NOR2_X1 U10054 ( .A1(n11723), .A2(n11732), .ZN(n7405) );
  OAI22_X1 U10055 ( .A1(n11723), .A2(n7406), .B1(n7408), .B2(n7409), .ZN(n7407) );
  NAND3_X1 U10056 ( .A1(n7416), .A2(n7415), .A3(n7414), .ZN(n11385) );
  NAND2_X1 U10057 ( .A1(n11138), .A2(n11379), .ZN(n7414) );
  AOI21_X1 U10058 ( .B1(n11379), .B2(n6834), .A(n7417), .ZN(n7415) );
  INV_X1 U10059 ( .A(n7419), .ZN(n7416) );
  NOR2_X1 U10060 ( .A1(n11138), .A2(n7418), .ZN(n7419) );
  NAND2_X1 U10061 ( .A1(n11150), .A2(n6602), .ZN(n7418) );
  INV_X1 U10062 ( .A(n12649), .ZN(n7423) );
  INV_X1 U10063 ( .A(n10650), .ZN(n7430) );
  NAND2_X1 U10064 ( .A1(n10586), .A2(n6554), .ZN(n7432) );
  NOR2_X2 U10065 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8737) );
  NAND3_X1 U10066 ( .A1(n8831), .A2(n8792), .A3(n10679), .ZN(n7440) );
  NAND2_X1 U10067 ( .A1(n7444), .A2(n7443), .ZN(n9126) );
  INV_X1 U10068 ( .A(n9102), .ZN(n13135) );
  INV_X1 U10069 ( .A(n13158), .ZN(n7446) );
  NAND2_X1 U10070 ( .A1(n8597), .A2(n8779), .ZN(n7457) );
  NOR2_X2 U10071 ( .A1(n7457), .A2(n7455), .ZN(n8706) );
  NAND2_X1 U10072 ( .A1(n7462), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7917) );
  NAND2_X1 U10073 ( .A1(n8104), .A2(n7465), .ZN(n7464) );
  NAND3_X1 U10074 ( .A1(n10980), .A2(n10982), .A3(n8104), .ZN(n7467) );
  NAND2_X1 U10075 ( .A1(n12756), .A2(n8495), .ZN(n7469) );
  NAND3_X1 U10076 ( .A1(n8530), .A2(n8529), .A3(n8573), .ZN(n7474) );
  NAND2_X1 U10077 ( .A1(n7477), .A2(n7475), .ZN(n8473) );
  INV_X1 U10078 ( .A(n8471), .ZN(n7478) );
  NAND2_X1 U10079 ( .A1(n7482), .A2(n7483), .ZN(n9943) );
  NAND2_X1 U10080 ( .A1(n12731), .A2(n7486), .ZN(n7482) );
  INV_X1 U10081 ( .A(n8485), .ZN(n7491) );
  NAND2_X1 U10082 ( .A1(n8468), .A2(n8467), .ZN(n11911) );
  NAND2_X1 U10083 ( .A1(n10798), .A2(n10801), .ZN(n12877) );
  NAND2_X1 U10084 ( .A1(n8460), .A2(n8459), .ZN(n11457) );
  NAND2_X1 U10085 ( .A1(n8453), .A2(n8452), .ZN(n10931) );
  NAND2_X1 U10086 ( .A1(n8053), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8025) );
  AOI21_X2 U10087 ( .B1(n9943), .B2(n8504), .A(n8503), .ZN(n12137) );
  NAND2_X1 U10088 ( .A1(n7496), .A2(n13007), .ZN(n12148) );
  NAND2_X1 U10089 ( .A1(n7496), .A2(n12939), .ZN(n12156) );
  AOI21_X1 U10090 ( .B1(n7496), .B2(n12855), .A(n12151), .ZN(n12152) );
  OAI21_X1 U10091 ( .B1(n7888), .B2(n7503), .A(n7500), .ZN(n8266) );
  NAND2_X1 U10092 ( .A1(n7888), .A2(n7500), .ZN(n7499) );
  NAND3_X1 U10093 ( .A1(n7507), .A2(n7506), .A3(n6485), .ZN(n7505) );
  NAND2_X1 U10094 ( .A1(n7510), .A2(n7508), .ZN(n7869) );
  NAND2_X1 U10095 ( .A1(n7901), .A2(n7521), .ZN(n7519) );
  NAND2_X1 U10096 ( .A1(n7519), .A2(n7520), .ZN(n7969) );
  NAND2_X1 U10097 ( .A1(n8020), .A2(n6586), .ZN(n7861) );
  OAI21_X1 U10098 ( .B1(n7971), .B2(n7957), .A(n7531), .ZN(n8381) );
  NAND2_X1 U10099 ( .A1(n7529), .A2(n7530), .ZN(n8383) );
  NAND2_X1 U10100 ( .A1(n7971), .A2(n7531), .ZN(n7529) );
  NAND2_X1 U10101 ( .A1(n7971), .A2(n7903), .ZN(n7958) );
  NAND2_X1 U10102 ( .A1(n12483), .A2(n12484), .ZN(n7582) );
  OAI211_X1 U10103 ( .C1(n12483), .C2(n7580), .A(n7577), .B(n7576), .ZN(n12213) );
  NAND2_X1 U10104 ( .A1(n12483), .A2(n6583), .ZN(n7576) );
  OAI22_X1 U10105 ( .A1(n7579), .A2(n7578), .B1(n7586), .B2(n7581), .ZN(n7577)
         );
  INV_X1 U10106 ( .A(n7581), .ZN(n7578) );
  NAND3_X1 U10107 ( .A1(n7592), .A2(n7925), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7926) );
  XNOR2_X1 U10108 ( .A(n7592), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U10109 ( .A1(n9073), .A2(n8685), .ZN(n7597) );
  NAND3_X1 U10110 ( .A1(n13417), .A2(n13641), .A3(n7599), .ZN(n7598) );
  NAND2_X1 U10111 ( .A1(n8908), .A2(n7608), .ZN(n7604) );
  NAND2_X1 U10112 ( .A1(n8908), .A2(n8657), .ZN(n7607) );
  NAND2_X1 U10113 ( .A1(n13217), .A2(n7618), .ZN(n7620) );
  INV_X1 U10114 ( .A(n13216), .ZN(n7618) );
  NAND2_X1 U10115 ( .A1(n7619), .A2(n7621), .ZN(n13221) );
  NAND2_X1 U10116 ( .A1(n6535), .A2(n7620), .ZN(n7619) );
  OAI21_X1 U10117 ( .B1(n13431), .B2(n13426), .A(n7624), .ZN(n7623) );
  NAND2_X1 U10118 ( .A1(n7626), .A2(n7625), .ZN(n13284) );
  AOI21_X1 U10119 ( .B1(n13252), .B2(n6440), .A(n6548), .ZN(n7626) );
  INV_X1 U10120 ( .A(n13254), .ZN(n7633) );
  NAND2_X1 U10121 ( .A1(n7637), .A2(n7635), .ZN(n13317) );
  NAND2_X1 U10122 ( .A1(n13313), .A2(n7638), .ZN(n7637) );
  NAND2_X1 U10123 ( .A1(n7642), .A2(n7640), .ZN(n13241) );
  NAND2_X1 U10124 ( .A1(n13237), .A2(n7643), .ZN(n7642) );
  NAND2_X1 U10125 ( .A1(n7645), .A2(n7646), .ZN(n13299) );
  INV_X1 U10126 ( .A(n13296), .ZN(n7649) );
  NAND2_X1 U10127 ( .A1(n13361), .A2(n7655), .ZN(n7653) );
  NAND3_X1 U10128 ( .A1(n7654), .A2(n7653), .A3(n7652), .ZN(n13420) );
  NAND3_X1 U10129 ( .A1(n13331), .A2(n7655), .A3(n7656), .ZN(n7654) );
  AND2_X1 U10130 ( .A1(n13332), .A2(n13330), .ZN(n7656) );
  NAND2_X1 U10131 ( .A1(n13306), .A2(n13307), .ZN(n13305) );
  INV_X1 U10132 ( .A(n7855), .ZN(n7660) );
  NAND2_X1 U10133 ( .A1(n9669), .A2(n9668), .ZN(n14688) );
  NAND2_X1 U10134 ( .A1(n7665), .A2(n9678), .ZN(n9688) );
  OAI21_X2 U10135 ( .B1(n14918), .B2(n7676), .A(n7675), .ZN(n14857) );
  NAND4_X1 U10136 ( .A1(n7715), .A2(n9328), .A3(n9396), .A4(n6594), .ZN(n7683)
         );
  NAND2_X1 U10137 ( .A1(n14498), .A2(n14970), .ZN(n10839) );
  INV_X1 U10138 ( .A(n14251), .ZN(n11131) );
  AND2_X4 U10139 ( .A1(n14247), .A2(n14431), .ZN(n15216) );
  NOR2_X1 U10140 ( .A1(n14251), .A2(n14245), .ZN(n14431) );
  NAND2_X1 U10141 ( .A1(n14151), .A2(n7688), .ZN(n7686) );
  NAND2_X1 U10142 ( .A1(n7686), .A2(n7687), .ZN(n14101) );
  CLKBUF_X1 U10143 ( .A(n7694), .Z(n7693) );
  NAND3_X1 U10144 ( .A1(n9328), .A2(n7699), .A3(n9396), .ZN(n9571) );
  NAND2_X1 U10145 ( .A1(n11643), .A2(n7701), .ZN(n7700) );
  NAND2_X1 U10146 ( .A1(n7705), .A2(n7703), .ZN(n7702) );
  INV_X1 U10147 ( .A(n11033), .ZN(n7704) );
  NAND2_X1 U10148 ( .A1(n11031), .A2(n11030), .ZN(n7705) );
  NAND2_X2 U10149 ( .A1(n13738), .A2(n13583), .ZN(n7711) );
  NAND2_X1 U10150 ( .A1(n13665), .A2(n13591), .ZN(n13648) );
  NAND2_X1 U10151 ( .A1(n9710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9339) );
  XNOR2_X2 U10152 ( .A(n9338), .B(n9337), .ZN(n9784) );
  INV_X1 U10153 ( .A(n14697), .ZN(n7724) );
  NAND2_X1 U10154 ( .A1(n7724), .A2(n7725), .ZN(n9976) );
  NAND2_X1 U10155 ( .A1(n8602), .A2(n14089), .ZN(n7728) );
  NAND3_X1 U10156 ( .A1(n8602), .A2(n14089), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n7729) );
  INV_X1 U10157 ( .A(n8602), .ZN(n8601) );
  NAND2_X1 U10158 ( .A1(n14785), .A2(n7730), .ZN(n14740) );
  NAND3_X2 U10159 ( .A1(n11857), .A2(n7733), .A3(n7732), .ZN(n14912) );
  NAND3_X1 U10160 ( .A1(n7733), .A2(n11857), .A3(n15071), .ZN(n14930) );
  AND3_X1 U10161 ( .A1(n7913), .A2(n7915), .A3(n7914), .ZN(n7983) );
  NAND4_X1 U10162 ( .A1(n7736), .A2(n7734), .A3(n6400), .A4(n7983), .ZN(n8562)
         );
  NAND2_X1 U10163 ( .A1(n7738), .A2(n8041), .ZN(n7737) );
  NAND2_X2 U10164 ( .A1(n10801), .A2(n8047), .ZN(n11007) );
  NAND2_X1 U10165 ( .A1(n12858), .A2(n7742), .ZN(n7741) );
  NAND2_X1 U10166 ( .A1(n7747), .A2(n7745), .ZN(n11912) );
  NAND2_X1 U10167 ( .A1(n12031), .A2(n7755), .ZN(n12050) );
  OAI21_X1 U10168 ( .B1(n12778), .B2(n9898), .A(n9897), .ZN(n12766) );
  NAND2_X1 U10169 ( .A1(n12733), .A2(n9902), .ZN(n7767) );
  INV_X1 U10170 ( .A(n9905), .ZN(n7766) );
  NAND2_X1 U10171 ( .A1(n7768), .A2(n15272), .ZN(n9992) );
  NAND2_X1 U10172 ( .A1(n7768), .A2(n15265), .ZN(n9994) );
  NAND3_X1 U10173 ( .A1(n6546), .A2(n9990), .A3(n9989), .ZN(n7768) );
  NAND2_X1 U10174 ( .A1(n9752), .A2(n7834), .ZN(n7770) );
  OAI21_X2 U10175 ( .B1(n14701), .B2(n7783), .A(n7784), .ZN(n14655) );
  INV_X1 U10176 ( .A(n14655), .ZN(n9988) );
  XNOR2_X2 U10177 ( .A(n13450), .B(n10017), .ZN(n9999) );
  NAND2_X1 U10178 ( .A1(n7802), .A2(n7801), .ZN(n13675) );
  NAND2_X1 U10179 ( .A1(n7813), .A2(n13622), .ZN(n7804) );
  NOR2_X2 U10180 ( .A1(n7808), .A2(n7807), .ZN(n7806) );
  INV_X1 U10181 ( .A(n13764), .ZN(n7821) );
  INV_X1 U10182 ( .A(n13793), .ZN(n7827) );
  NAND2_X1 U10183 ( .A1(n13764), .A2(n6426), .ZN(n7816) );
  INV_X1 U10184 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7925) );
  NAND2_X1 U10185 ( .A1(n9106), .A2(n8686), .ZN(n9131) );
  OR2_X1 U10186 ( .A1(n14704), .A2(n15050), .ZN(n14990) );
  NAND2_X1 U10187 ( .A1(n13680), .A2(n7854), .ZN(n13686) );
  INV_X1 U10188 ( .A(n13953), .ZN(n13954) );
  INV_X1 U10189 ( .A(n10758), .ZN(n10745) );
  NOR2_X1 U10190 ( .A1(n10758), .A2(n10149), .ZN(n14513) );
  AND2_X1 U10191 ( .A1(n10758), .A2(n10118), .ZN(n10752) );
  OAI21_X1 U10192 ( .B1(n13952), .B2(n15381), .A(n13951), .ZN(n13953) );
  INV_X1 U10193 ( .A(n13978), .ZN(n13736) );
  AOI21_X1 U10194 ( .B1(n9823), .B2(n9822), .A(n9821), .ZN(n9826) );
  INV_X1 U10195 ( .A(n8564), .ZN(n8560) );
  NAND2_X1 U10196 ( .A1(n13950), .A2(n6404), .ZN(n13326) );
  NAND2_X1 U10197 ( .A1(n14972), .A2(n14499), .ZN(n10843) );
  NAND2_X1 U10198 ( .A1(n13543), .A2(n13656), .ZN(n13653) );
  CLKBUF_X1 U10199 ( .A(n14854), .Z(n14855) );
  CLKBUF_X1 U10200 ( .A(n12031), .Z(n12032) );
  BUF_X4 U10201 ( .A(n8063), .Z(n8438) );
  NOR2_X1 U10202 ( .A1(n9802), .A2(n15247), .ZN(n9809) );
  CLKBUF_X1 U10203 ( .A(n11956), .Z(n14939) );
  INV_X1 U10204 ( .A(n9966), .ZN(n9535) );
  NAND2_X1 U10205 ( .A1(n9952), .A2(n11179), .ZN(n15418) );
  INV_X1 U10206 ( .A(n6417), .ZN(n9951) );
  OR2_X1 U10207 ( .A1(n11846), .A2(n11845), .ZN(n7828) );
  NAND2_X1 U10208 ( .A1(n8505), .A2(n8525), .ZN(n12140) );
  AND2_X1 U10209 ( .A1(n8577), .A2(n8576), .ZN(n7829) );
  OR2_X1 U10210 ( .A1(n7545), .A2(n13443), .ZN(n7830) );
  OR3_X1 U10211 ( .A1(n10821), .A2(P3_IR_REG_1__SCAN_IN), .A3(n10501), .ZN(
        n7831) );
  OR2_X1 U10212 ( .A1(n13993), .A2(n13798), .ZN(n7832) );
  AND2_X1 U10213 ( .A1(n12882), .A2(n10984), .ZN(n7833) );
  NOR2_X1 U10214 ( .A1(n14440), .A2(n9749), .ZN(n7834) );
  AND2_X1 U10215 ( .A1(n13993), .A2(n13798), .ZN(n7835) );
  INV_X1 U10216 ( .A(n13798), .ZN(n13629) );
  OR2_X1 U10217 ( .A1(n13809), .A2(n13781), .ZN(n7837) );
  OR2_X1 U10218 ( .A1(n11535), .A2(n11534), .ZN(n7838) );
  AND2_X1 U10219 ( .A1(n8573), .A2(n7221), .ZN(n7839) );
  INV_X1 U10220 ( .A(n12822), .ZN(n9891) );
  OR2_X1 U10221 ( .A1(n9970), .A2(n10245), .ZN(n7840) );
  AND2_X1 U10222 ( .A1(n13558), .A2(n13557), .ZN(n7841) );
  INV_X1 U10223 ( .A(n15105), .ZN(n12221) );
  AND2_X1 U10224 ( .A1(n11402), .A2(n11401), .ZN(n7842) );
  NOR2_X2 U10225 ( .A1(n14740), .A2(n14739), .ZN(n14719) );
  NAND2_X2 U10226 ( .A1(n10014), .A2(n13837), .ZN(n13880) );
  INV_X2 U10227 ( .A(n15264), .ZN(n15265) );
  OR2_X1 U10228 ( .A1(n14025), .A2(n13568), .ZN(n7844) );
  INV_X1 U10229 ( .A(n14025), .ZN(n13569) );
  XOR2_X1 U10230 ( .A(n8099), .B(n8098), .Z(n7845) );
  OR2_X1 U10231 ( .A1(n9802), .A2(n14910), .ZN(n7846) );
  INV_X1 U10232 ( .A(n13821), .ZN(n13626) );
  INV_X1 U10233 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8611) );
  OAI21_X1 U10234 ( .B1(n13635), .B2(n13978), .A(n13634), .ZN(n13636) );
  NOR2_X1 U10235 ( .A1(n15022), .A2(n14783), .ZN(n7847) );
  AND2_X1 U10236 ( .A1(n8675), .A2(n8674), .ZN(n7848) );
  AND2_X1 U10237 ( .A1(n14373), .A2(n14780), .ZN(n7849) );
  AND2_X1 U10238 ( .A1(SI_2_), .A2(SI_3_), .ZN(n7850) );
  INV_X1 U10239 ( .A(n14443), .ZN(n9754) );
  AND2_X1 U10240 ( .A1(n9286), .A2(n13182), .ZN(n7851) );
  OR2_X1 U10241 ( .A1(n10193), .A2(n10541), .ZN(n7853) );
  OR2_X1 U10242 ( .A1(n13679), .A2(n6493), .ZN(n7854) );
  OR2_X1 U10243 ( .A1(n9858), .A2(n10750), .ZN(n15270) );
  NOR2_X1 U10244 ( .A1(n9758), .A2(n11954), .ZN(n7855) );
  OR2_X1 U10245 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  INV_X1 U10246 ( .A(n9741), .ZN(n14265) );
  OR2_X1 U10247 ( .A1(n14414), .A2(n7193), .ZN(n14269) );
  AND2_X1 U10248 ( .A1(n14271), .A2(n7193), .ZN(n14273) );
  INV_X1 U10249 ( .A(n14296), .ZN(n14297) );
  AND2_X1 U10250 ( .A1(n14308), .A2(n14307), .ZN(n14309) );
  OR2_X1 U10251 ( .A1(n14339), .A2(n14338), .ZN(n14340) );
  OR2_X1 U10252 ( .A1(n14367), .A2(n14366), .ZN(n14364) );
  MUX2_X1 U10253 ( .A(n8399), .B(n8398), .S(n10430), .Z(n8400) );
  NAND2_X1 U10254 ( .A1(n13326), .A2(n13325), .ZN(n13351) );
  NAND2_X1 U10255 ( .A1(n10932), .A2(n7833), .ZN(n9868) );
  OAI21_X1 U10256 ( .B1(n15000), .B2(n14712), .A(n14711), .ZN(n9772) );
  INV_X1 U10257 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7912) );
  INV_X1 U10258 ( .A(n10843), .ZN(n10844) );
  INV_X1 U10259 ( .A(n12034), .ZN(n9885) );
  NAND2_X1 U10260 ( .A1(n9866), .A2(n10802), .ZN(n10932) );
  INV_X1 U10261 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8937) );
  INV_X1 U10262 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8708) );
  OR2_X1 U10263 ( .A1(n12279), .A2(n14170), .ZN(n12281) );
  INV_X1 U10264 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9316) );
  INV_X1 U10265 ( .A(n11443), .ZN(n9877) );
  INV_X1 U10266 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7920) );
  INV_X1 U10267 ( .A(n9210), .ZN(n9211) );
  NAND2_X1 U10268 ( .A1(n9219), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9274) );
  OR2_X1 U10269 ( .A1(n14013), .A2(n13870), .ZN(n13572) );
  INV_X1 U10270 ( .A(n14668), .ZN(n14421) );
  NAND2_X1 U10271 ( .A1(n14654), .A2(n9986), .ZN(n9987) );
  OR2_X1 U10272 ( .A1(n9818), .A2(SI_27_), .ZN(n9822) );
  INV_X1 U10273 ( .A(n9440), .ZN(n9442) );
  INV_X1 U10274 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7939) );
  INV_X1 U10275 ( .A(n8091), .ZN(n8312) );
  INV_X1 U10276 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U10277 ( .A1(n9209), .A2(n9211), .ZN(n9212) );
  AND2_X1 U10278 ( .A1(n13176), .A2(n9207), .ZN(n9208) );
  INV_X1 U10279 ( .A(n13425), .ZN(n13426) );
  INV_X1 U10280 ( .A(n13404), .ZN(n11484) );
  AND2_X1 U10281 ( .A1(n9232), .A2(n9231), .ZN(n9235) );
  INV_X1 U10282 ( .A(n14205), .ZN(n12084) );
  INV_X1 U10283 ( .A(n9750), .ZN(n9751) );
  INV_X1 U10284 ( .A(n15214), .ZN(n9794) );
  NOR3_X1 U10285 ( .A1(n14651), .A2(n15247), .A3(n14652), .ZN(n9981) );
  INV_X1 U10286 ( .A(n14439), .ZN(n14272) );
  AND2_X1 U10287 ( .A1(n14547), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10402) );
  OR2_X1 U10288 ( .A1(n11466), .A2(n11472), .ZN(n11467) );
  INV_X1 U10289 ( .A(n12016), .ZN(n12017) );
  INV_X1 U10290 ( .A(n11872), .ZN(n11871) );
  NAND2_X1 U10291 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  INV_X1 U10292 ( .A(n15391), .ZN(n12655) );
  AND2_X1 U10293 ( .A1(n10444), .A2(n10433), .ZN(n10440) );
  AND2_X1 U10294 ( .A1(n8477), .A2(n8478), .ZN(n12845) );
  OR2_X1 U10295 ( .A1(n9936), .A2(n10576), .ZN(n12144) );
  INV_X1 U10296 ( .A(n15418), .ZN(n15423) );
  AND3_X1 U10297 ( .A1(n10796), .A2(n10690), .A3(n9959), .ZN(n10808) );
  INV_X1 U10298 ( .A(n11314), .ZN(n9952) );
  OR2_X1 U10299 ( .A1(n13044), .A2(n9223), .ZN(n9229) );
  INV_X1 U10300 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11502) );
  INV_X1 U10301 ( .A(n15305), .ZN(n15313) );
  OR2_X1 U10302 ( .A1(n10195), .A2(n10205), .ZN(n13869) );
  INV_X1 U10303 ( .A(n13442), .ZN(n13556) );
  INV_X1 U10304 ( .A(n10371), .ZN(n9304) );
  OR3_X1 U10305 ( .A1(n11785), .A2(n11479), .A3(n11572), .ZN(n9995) );
  NAND2_X1 U10306 ( .A1(n9235), .A2(n9236), .ZN(n9238) );
  OAI22_X1 U10307 ( .A1(n14258), .A2(n11341), .B1(n14260), .B2(n6401), .ZN(
        n10857) );
  INV_X1 U10308 ( .A(n14712), .ZN(n14387) );
  NAND2_X1 U10309 ( .A1(n12076), .A2(n12078), .ZN(n12079) );
  INV_X1 U10310 ( .A(n14218), .ZN(n14236) );
  NAND2_X1 U10311 ( .A1(n14416), .A2(n14245), .ZN(n14432) );
  INV_X1 U10312 ( .A(n9539), .ZN(n9585) );
  INV_X1 U10313 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14531) );
  INV_X1 U10314 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14547) );
  INV_X1 U10315 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10456) );
  INV_X1 U10316 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11242) );
  INV_X1 U10317 ( .A(n14643), .ZN(n9846) );
  AOI21_X1 U10318 ( .B1(n9806), .B2(n14907), .A(n9798), .ZN(n9799) );
  INV_X1 U10319 ( .A(n14995), .ZN(n14726) );
  OR2_X1 U10320 ( .A1(n10141), .A2(n10755), .ZN(n15217) );
  NOR2_X1 U10321 ( .A1(n9982), .A2(n9981), .ZN(n9990) );
  INV_X1 U10322 ( .A(n15216), .ZN(n14929) );
  AOI21_X1 U10323 ( .B1(n11531), .B2(n9721), .A(n11840), .ZN(n9722) );
  NOR2_X1 U10324 ( .A1(n9703), .A2(n9336), .ZN(n9704) );
  NAND2_X1 U10325 ( .A1(n8625), .A2(n7850), .ZN(n8633) );
  NAND2_X1 U10326 ( .A1(n11252), .A2(n11251), .ZN(n11594) );
  AND3_X1 U10327 ( .A1(n10808), .A2(n10807), .A3(n10576), .ZN(n12497) );
  INV_X1 U10328 ( .A(n10571), .ZN(n10574) );
  INV_X1 U10329 ( .A(n12697), .ZN(n12661) );
  AND2_X1 U10330 ( .A1(n10440), .A2(n13031), .ZN(n12707) );
  INV_X1 U10331 ( .A(n12048), .ZN(n12879) );
  OR2_X1 U10332 ( .A1(n11777), .A2(n11002), .ZN(n11003) );
  NAND3_X1 U10333 ( .A1(n10574), .A2(n15423), .A3(n12889), .ZN(n12891) );
  INV_X1 U10334 ( .A(n12891), .ZN(n12873) );
  AND2_X1 U10335 ( .A1(n9934), .A2(n9933), .ZN(n10694) );
  INV_X1 U10336 ( .A(n12949), .ZN(n13007) );
  AND2_X1 U10337 ( .A1(n12889), .A2(n9952), .ZN(n15425) );
  OR2_X1 U10338 ( .A1(n11777), .A2(n15425), .ZN(n15395) );
  XNOR2_X1 U10339 ( .A(n8450), .B(n8556), .ZN(n10558) );
  INV_X1 U10340 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8139) );
  AND2_X1 U10341 ( .A1(n7866), .A2(n7865), .ZN(n8087) );
  AND2_X1 U10342 ( .A1(n9303), .A2(n13435), .ZN(n13161) );
  OR2_X1 U10343 ( .A1(n8784), .A2(n8767), .ZN(n8770) );
  AND2_X1 U10344 ( .A1(n10207), .A2(n10206), .ZN(n15305) );
  INV_X1 U10345 ( .A(n15294), .ZN(n15318) );
  AND2_X1 U10346 ( .A1(n10200), .A2(n13434), .ZN(n15315) );
  AND3_X1 U10347 ( .A1(n13653), .A2(n13889), .A3(n13652), .ZN(n13949) );
  INV_X1 U10348 ( .A(n13622), .ZN(n13866) );
  INV_X1 U10349 ( .A(n13869), .ZN(n13883) );
  INV_X1 U10350 ( .A(n13920), .ZN(n13905) );
  AND2_X1 U10351 ( .A1(n9261), .A2(n15353), .ZN(n10382) );
  NOR2_X1 U10352 ( .A1(n10373), .A2(n10372), .ZN(n10384) );
  AND2_X1 U10353 ( .A1(n9243), .A2(n9242), .ZN(n15323) );
  AND2_X1 U10354 ( .A1(n9995), .A2(n11331), .ZN(n9298) );
  INV_X1 U10355 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8738) );
  INV_X1 U10356 ( .A(n11357), .ZN(n15245) );
  INV_X1 U10357 ( .A(n15182), .ZN(n14211) );
  INV_X1 U10358 ( .A(n14198), .ZN(n15179) );
  INV_X1 U10359 ( .A(n15174), .ZN(n14232) );
  INV_X1 U10360 ( .A(n14633), .ZN(n15197) );
  INV_X1 U10361 ( .A(n14635), .ZN(n15188) );
  INV_X1 U10362 ( .A(n14637), .ZN(n15194) );
  NAND2_X1 U10363 ( .A1(n9776), .A2(n9664), .ZN(n14702) );
  INV_X1 U10364 ( .A(n14910), .ZN(n15227) );
  OAI21_X1 U10365 ( .B1(n10115), .B2(P1_D_REG_0__SCAN_IN), .A(n10148), .ZN(
        n10750) );
  INV_X1 U10366 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9863) );
  INV_X1 U10367 ( .A(n15251), .ZN(n15050) );
  AND2_X1 U10368 ( .A1(n10786), .A2(n9805), .ZN(n15255) );
  OR2_X1 U10369 ( .A1(n14243), .A2(n9814), .ZN(n9858) );
  OAI21_X1 U10370 ( .B1(P1_B_REG_SCAN_IN), .B2(n11531), .A(n9722), .ZN(n10115)
         );
  AND2_X1 U10371 ( .A1(n10444), .A2(n10443), .ZN(n15391) );
  INV_X1 U10372 ( .A(n12503), .ZN(n12451) );
  INV_X1 U10373 ( .A(n12502), .ZN(n12027) );
  NAND2_X1 U10374 ( .A1(n10570), .A2(n10574), .ZN(n12506) );
  INV_X1 U10375 ( .A(n12500), .ZN(n12859) );
  INV_X1 U10376 ( .A(n12707), .ZN(n12543) );
  INV_X1 U10377 ( .A(n12688), .ZN(n12663) );
  INV_X1 U10378 ( .A(n12896), .ZN(n12863) );
  INV_X1 U10379 ( .A(n12855), .ZN(n12867) );
  INV_X1 U10380 ( .A(n11969), .ZN(n11762) );
  NAND2_X1 U10381 ( .A1(n15589), .A2(n15395), .ZN(n12941) );
  INV_X1 U10382 ( .A(n15589), .ZN(n15440) );
  OAI21_X1 U10383 ( .B1(n12732), .B2(n12734), .A(n7485), .ZN(n12957) );
  OR2_X1 U10384 ( .A1(n15429), .A2(n12945), .ZN(n13010) );
  AND2_X2 U10385 ( .A1(n9961), .A2(n9960), .ZN(n15429) );
  AND2_X1 U10386 ( .A1(n13013), .A2(n9920), .ZN(n10132) );
  INV_X1 U10387 ( .A(n10132), .ZN(n10133) );
  INV_X1 U10388 ( .A(SI_18_), .ZN(n10819) );
  INV_X1 U10389 ( .A(SI_14_), .ZN(n10549) );
  INV_X1 U10390 ( .A(n10816), .ZN(n13036) );
  AOI21_X1 U10391 ( .B1(n6461), .B2(n9310), .A(n9309), .ZN(n9311) );
  AND2_X1 U10392 ( .A1(n9305), .A2(n13837), .ZN(n13194) );
  INV_X1 U10393 ( .A(n13868), .ZN(n13568) );
  INV_X1 U10394 ( .A(n15315), .ZN(n15300) );
  INV_X1 U10395 ( .A(n15273), .ZN(n15322) );
  AND2_X1 U10396 ( .A1(n13811), .A2(n11273), .ZN(n13935) );
  INV_X1 U10397 ( .A(n13897), .ZN(n13915) );
  INV_X1 U10398 ( .A(n15390), .ZN(n15387) );
  AND2_X2 U10399 ( .A1(n10384), .A2(n10382), .ZN(n15390) );
  NOR2_X1 U10400 ( .A1(n15323), .A2(n15356), .ZN(n15338) );
  AND2_X1 U10401 ( .A1(n9298), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15359) );
  XNOR2_X1 U10402 ( .A(n9237), .B(n9236), .ZN(n11479) );
  INV_X1 U10403 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10368) );
  INV_X1 U10404 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10154) );
  INV_X1 U10405 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10089) );
  INV_X1 U10406 ( .A(n15079), .ZN(n14305) );
  NAND2_X1 U10407 ( .A1(n10760), .A2(n10754), .ZN(n15174) );
  INV_X1 U10408 ( .A(n14225), .ZN(n14481) );
  INV_X1 U10409 ( .A(n14861), .ZN(n14486) );
  OR2_X1 U10410 ( .A1(n10261), .A2(n10257), .ZN(n14635) );
  OR2_X1 U10411 ( .A1(n10261), .A2(n14511), .ZN(n14633) );
  INV_X1 U10412 ( .A(n15223), .ZN(n14921) );
  NAND2_X1 U10413 ( .A1(n15270), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9991) );
  INV_X2 U10414 ( .A(n15270), .ZN(n15272) );
  OR2_X1 U10415 ( .A1(n9858), .A2(n9857), .ZN(n15264) );
  AND2_X1 U10416 ( .A1(n10757), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10118) );
  NAND2_X1 U10417 ( .A1(n10752), .A2(n10115), .ZN(n15230) );
  INV_X1 U10418 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10496) );
  INV_X1 U10419 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10240) );
  AND2_X2 U10420 ( .A1(n9997), .A2(n13013), .ZN(P3_U3897) );
  INV_X1 U10421 ( .A(n13451), .ZN(P2_U3947) );
  NAND2_X1 U10422 ( .A1(n8725), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8018) );
  INV_X1 U10423 ( .A(n8018), .ZN(n7856) );
  NAND2_X1 U10424 ( .A1(n10092), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10425 ( .A1(n10089), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10426 ( .A1(n10059), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10427 ( .A1(n10085), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10428 ( .A1(n10087), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10429 ( .A1(n7864), .A2(n7863), .ZN(n8015) );
  NAND2_X1 U10430 ( .A1(n10083), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10431 ( .A1(n7867), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10432 ( .A1(n10098), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7870) );
  OR2_X1 U10433 ( .A1(n8172), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10434 ( .A1(n10185), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U10435 ( .A1(n7874), .A2(n7873), .ZN(n8184) );
  NAND2_X1 U10436 ( .A1(n10240), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10437 ( .A1(n10237), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10438 ( .A1(n7876), .A2(n7875), .ZN(n8183) );
  NAND2_X1 U10439 ( .A1(n10394), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7882) );
  INV_X1 U10440 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U10441 ( .A1(n10391), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U10442 ( .A1(n7882), .A2(n7878), .ZN(n8232) );
  AND2_X1 U10443 ( .A1(n10241), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7879) );
  NOR2_X1 U10444 ( .A1(n8232), .A2(n7879), .ZN(n7880) );
  NAND2_X1 U10445 ( .A1(n10494), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U10446 ( .A1(n15545), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10447 ( .A1(n7884), .A2(n7883), .ZN(n8219) );
  NAND2_X1 U10448 ( .A1(n10370), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U10449 ( .A1(n10368), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10450 ( .A1(n7887), .A2(n7885), .ZN(n8244) );
  INV_X1 U10451 ( .A(n8244), .ZN(n7886) );
  NAND2_X1 U10452 ( .A1(n8245), .A2(n7886), .ZN(n7888) );
  NAND2_X1 U10453 ( .A1(n10496), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7890) );
  INV_X1 U10454 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U10455 ( .A1(n10497), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10456 ( .A1(n10977), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7892) );
  INV_X1 U10457 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U10458 ( .A1(n10978), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10459 ( .A1(n11116), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7894) );
  INV_X1 U10460 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11114) );
  NAND2_X1 U10461 ( .A1(n11114), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10462 ( .A1(n11132), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U10463 ( .A1(n11101), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U10464 ( .A1(n8324), .A2(n8323), .ZN(n8326) );
  NAND2_X1 U10465 ( .A1(n8326), .A2(n7896), .ZN(n8339) );
  NAND2_X1 U10466 ( .A1(n15495), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7898) );
  INV_X1 U10467 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11128) );
  NAND2_X1 U10468 ( .A1(n11128), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10469 ( .A1(n8339), .A2(n8338), .ZN(n8341) );
  XNOR2_X1 U10470 ( .A(n8687), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10471 ( .A1(n11272), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7899) );
  XNOR2_X1 U10472 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8358) );
  NAND2_X1 U10473 ( .A1(n8359), .A2(n8358), .ZN(n7901) );
  INV_X1 U10474 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10475 ( .A1(n8702), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7900) );
  INV_X1 U10476 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11478) );
  INV_X1 U10477 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U10478 ( .A1(n11576), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7903) );
  INV_X1 U10479 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U10480 ( .A1(n11573), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7902) );
  AND2_X1 U10481 ( .A1(n7903), .A2(n7902), .ZN(n7968) );
  NAND2_X1 U10482 ( .A1(n7969), .A2(n7968), .ZN(n7971) );
  INV_X1 U10483 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15483) );
  NAND2_X1 U10484 ( .A1(n15483), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7906) );
  INV_X1 U10485 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U10486 ( .A1(n11784), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10487 ( .A1(n7906), .A2(n7904), .ZN(n7957) );
  INV_X1 U10488 ( .A(n7957), .ZN(n7905) );
  INV_X1 U10489 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15108) );
  NAND2_X1 U10490 ( .A1(n15108), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8382) );
  INV_X1 U10491 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12161) );
  NAND2_X1 U10492 ( .A1(n12161), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10493 ( .A1(n8382), .A2(n7907), .ZN(n8380) );
  XNOR2_X1 U10494 ( .A(n8381), .B(n8380), .ZN(n13029) );
  NOR2_X1 U10495 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7908) );
  NAND2_X1 U10496 ( .A1(n7909), .A2(n7908), .ZN(n7980) );
  NAND4_X1 U10497 ( .A1(n7591), .A2(n7910), .A3(n8557), .A4(n7979), .ZN(n7911)
         );
  INV_X1 U10498 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10499 ( .A1(n7917), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10500 ( .A1(n7921), .A2(n7949), .ZN(n8571) );
  NAND2_X2 U10501 ( .A1(n8571), .A2(n10880), .ZN(n8029) );
  NAND2_X1 U10502 ( .A1(n13029), .A2(n8437), .ZN(n7929) );
  INV_X1 U10503 ( .A(SI_27_), .ZN(n13033) );
  OR2_X1 U10504 ( .A1(n8438), .A2(n13033), .ZN(n7928) );
  INV_X2 U10505 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8052) );
  INV_X1 U10506 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7940) );
  INV_X1 U10507 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7941) );
  INV_X1 U10508 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7942) );
  INV_X1 U10509 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10510 ( .A1(n7962), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10511 ( .A1(n8390), .A2(n7945), .ZN(n12726) );
  INV_X1 U10512 ( .A(n7946), .ZN(n7948) );
  NAND2_X1 U10513 ( .A1(n7948), .A2(n7947), .ZN(n13018) );
  INV_X1 U10514 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10515 ( .A1(n8091), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10516 ( .A1(n8442), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7953) );
  OAI211_X1 U10517 ( .C1(n7955), .C2(n8409), .A(n7954), .B(n7953), .ZN(n7956)
         );
  AOI21_X2 U10518 ( .B1(n12726), .B2(n8395), .A(n7956), .ZN(n12489) );
  OR2_X1 U10519 ( .A1(n9906), .A2(n12489), .ZN(n8399) );
  NAND2_X1 U10520 ( .A1(n9906), .A2(n12489), .ZN(n8501) );
  XNOR2_X1 U10521 ( .A(n7958), .B(n7957), .ZN(n13035) );
  NAND2_X1 U10522 ( .A1(n13035), .A2(n8437), .ZN(n7960) );
  INV_X1 U10523 ( .A(SI_26_), .ZN(n13037) );
  OR2_X1 U10524 ( .A1(n8438), .A2(n13037), .ZN(n7959) );
  NAND2_X1 U10525 ( .A1(n7975), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10526 ( .A1(n7962), .A2(n7961), .ZN(n12737) );
  NAND2_X1 U10527 ( .A1(n12737), .A2(n8395), .ZN(n7967) );
  INV_X1 U10528 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12953) );
  INV_X2 U10529 ( .A(n8312), .ZN(n8424) );
  NAND2_X1 U10530 ( .A1(n8424), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10531 ( .A1(n8347), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7963) );
  OAI211_X1 U10532 ( .C1(n12953), .C2(n8409), .A(n7964), .B(n7963), .ZN(n7965)
         );
  INV_X1 U10533 ( .A(n7965), .ZN(n7966) );
  NAND2_X1 U10534 ( .A1(n12954), .A2(n12397), .ZN(n8396) );
  OR2_X1 U10535 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U10536 ( .A1(n7971), .A2(n7970), .ZN(n12070) );
  INV_X1 U10537 ( .A(SI_25_), .ZN(n12069) );
  OR2_X1 U10538 ( .A1(n8438), .A2(n12069), .ZN(n7972) );
  NAND2_X1 U10539 ( .A1(n7992), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10540 ( .A1(n7975), .A2(n7974), .ZN(n12748) );
  INV_X1 U10541 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U10542 ( .A1(n8347), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U10543 ( .A1(n8424), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n7976) );
  OAI211_X1 U10544 ( .C1(n12959), .C2(n8409), .A(n7977), .B(n7976), .ZN(n7978)
         );
  OR2_X1 U10545 ( .A1(n12961), .A2(n12432), .ZN(n8373) );
  NAND2_X1 U10546 ( .A1(n12961), .A2(n12432), .ZN(n8497) );
  NAND2_X1 U10547 ( .A1(n8449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10548 ( .A1(n7985), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7987) );
  XNOR2_X2 U10549 ( .A(n7987), .B(n7986), .ZN(n11179) );
  MUX2_X1 U10550 ( .A(n8373), .B(n8497), .S(n10430), .Z(n8378) );
  XNOR2_X1 U10551 ( .A(n7988), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U10552 ( .A1(n12214), .A2(n8437), .ZN(n7990) );
  INV_X1 U10553 ( .A(SI_24_), .ZN(n12216) );
  OR2_X1 U10554 ( .A1(n8438), .A2(n12216), .ZN(n7989) );
  NAND2_X1 U10555 ( .A1(n8363), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U10556 ( .A1(n7992), .A2(n7991), .ZN(n12758) );
  NAND2_X1 U10557 ( .A1(n12758), .A2(n8395), .ZN(n7998) );
  INV_X1 U10558 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10559 ( .A1(n8424), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10560 ( .A1(n8442), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n7993) );
  OAI211_X1 U10561 ( .C1(n7995), .C2(n8409), .A(n7994), .B(n7993), .ZN(n7996)
         );
  INV_X1 U10562 ( .A(n7996), .ZN(n7997) );
  XNOR2_X1 U10563 ( .A(n12909), .B(n12357), .ZN(n12757) );
  XNOR2_X1 U10564 ( .A(n8000), .B(n7999), .ZN(n11313) );
  NAND2_X1 U10565 ( .A1(n11313), .A2(n8437), .ZN(n8002) );
  INV_X1 U10566 ( .A(SI_22_), .ZN(n8688) );
  OR2_X1 U10567 ( .A1(n8438), .A2(n8688), .ZN(n8001) );
  NAND2_X1 U10568 ( .A1(n8346), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10569 ( .A1(n6456), .A2(n8003), .ZN(n12782) );
  NAND2_X1 U10570 ( .A1(n12782), .A2(n8395), .ZN(n8008) );
  INV_X1 U10571 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12973) );
  NAND2_X1 U10572 ( .A1(n8442), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8005) );
  NAND2_X1 U10573 ( .A1(n8424), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8004) );
  OAI211_X1 U10574 ( .C1(n8409), .C2(n12973), .A(n8005), .B(n8004), .ZN(n8006)
         );
  INV_X1 U10575 ( .A(n8006), .ZN(n8007) );
  NAND2_X1 U10576 ( .A1(n12974), .A2(n12375), .ZN(n8489) );
  NAND2_X1 U10577 ( .A1(n8488), .A2(n8489), .ZN(n12777) );
  NAND2_X1 U10578 ( .A1(n8091), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U10579 ( .A1(n8347), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10580 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8009) );
  NAND2_X1 U10581 ( .A1(n8074), .A2(n8009), .ZN(n11016) );
  NAND2_X1 U10582 ( .A1(n8395), .A2(n11016), .ZN(n8011) );
  NAND2_X1 U10583 ( .A1(n8051), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8010) );
  INV_X1 U10584 ( .A(n12521), .ZN(n8017) );
  XNOR2_X1 U10585 ( .A(n8016), .B(n8015), .ZN(n10122) );
  INV_X1 U10586 ( .A(SI_4_), .ZN(n10123) );
  INV_X1 U10587 ( .A(SI_1_), .ZN(n10094) );
  NAND2_X1 U10588 ( .A1(n8019), .A2(n8018), .ZN(n8021) );
  AND2_X1 U10589 ( .A1(n8021), .A2(n8020), .ZN(n10095) );
  OR2_X1 U10590 ( .A1(n8062), .A2(n10095), .ZN(n8023) );
  NAND2_X1 U10591 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n10501), .ZN(n8022) );
  INV_X1 U10592 ( .A(n11005), .ZN(n10902) );
  NAND2_X1 U10593 ( .A1(n8091), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10594 ( .A1(n8050), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8027) );
  NAND4_X2 U10595 ( .A1(n8028), .A2(n8027), .A3(n8026), .A4(n8025), .ZN(n12523) );
  INV_X1 U10596 ( .A(n8062), .ZN(n8031) );
  XNOR2_X1 U10597 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .ZN(n10100) );
  INV_X1 U10598 ( .A(n10100), .ZN(n8030) );
  INV_X1 U10599 ( .A(n10501), .ZN(n10507) );
  INV_X1 U10600 ( .A(n8063), .ZN(n8032) );
  NAND2_X1 U10601 ( .A1(n12523), .A2(n10823), .ZN(n8531) );
  NAND2_X1 U10602 ( .A1(n8531), .A2(n11314), .ZN(n8035) );
  NAND2_X1 U10603 ( .A1(n8531), .A2(n10983), .ZN(n8034) );
  NAND2_X1 U10604 ( .A1(n11004), .A2(n11179), .ZN(n8036) );
  NAND2_X1 U10605 ( .A1(n8091), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8040) );
  NAND2_X1 U10606 ( .A1(n8050), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8039) );
  NAND2_X1 U10607 ( .A1(n8051), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10608 ( .A1(n8053), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8037) );
  XNOR2_X1 U10609 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8042) );
  XNOR2_X1 U10610 ( .A(n8043), .B(n8042), .ZN(n10136) );
  OR2_X1 U10611 ( .A1(n8062), .A2(n10136), .ZN(n8045) );
  OR2_X1 U10612 ( .A1(n8063), .A2(SI_2_), .ZN(n8044) );
  NAND2_X1 U10613 ( .A1(n10949), .A2(n10812), .ZN(n8452) );
  NAND2_X1 U10614 ( .A1(n8046), .A2(n12888), .ZN(n8069) );
  NAND2_X1 U10615 ( .A1(n8452), .A2(n8069), .ZN(n8533) );
  INV_X1 U10616 ( .A(n8533), .ZN(n8451) );
  NAND3_X1 U10617 ( .A1(n8049), .A2(n8451), .A3(n8048), .ZN(n8068) );
  NAND2_X1 U10618 ( .A1(n8091), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10619 ( .A1(n8050), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U10620 ( .A1(n8051), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10621 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  NAND2_X1 U10622 ( .A1(n8059), .A2(n8080), .ZN(n10607) );
  XNOR2_X1 U10623 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8060) );
  XNOR2_X1 U10624 ( .A(n8061), .B(n8060), .ZN(n10120) );
  OR2_X1 U10625 ( .A1(n8062), .A2(n10120), .ZN(n8065) );
  INV_X1 U10626 ( .A(SI_3_), .ZN(n10121) );
  OR2_X1 U10627 ( .A1(n8063), .A2(n10121), .ZN(n8064) );
  OAI211_X1 U10628 ( .C1(n10431), .C2(n10607), .A(n8065), .B(n8064), .ZN(
        n10998) );
  NAND2_X1 U10629 ( .A1(n8455), .A2(n8452), .ZN(n8066) );
  NAND2_X1 U10630 ( .A1(n8066), .A2(n9936), .ZN(n8067) );
  NAND2_X1 U10631 ( .A1(n8068), .A2(n8067), .ZN(n8071) );
  INV_X1 U10632 ( .A(n10998), .ZN(n10950) );
  NAND2_X1 U10633 ( .A1(n12878), .A2(n10950), .ZN(n8454) );
  AOI21_X1 U10634 ( .B1(n8454), .B2(n8069), .A(n9936), .ZN(n8070) );
  AOI21_X1 U10635 ( .B1(n8071), .B2(n8454), .A(n8070), .ZN(n8073) );
  NOR2_X1 U10636 ( .A1(n8455), .A2(n9936), .ZN(n8072) );
  NAND2_X1 U10637 ( .A1(n8091), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10638 ( .A1(n8347), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10639 ( .A1(n8074), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U10640 ( .A1(n8092), .A2(n8075), .ZN(n11187) );
  NAND2_X1 U10641 ( .A1(n8395), .A2(n11187), .ZN(n8077) );
  NAND2_X1 U10642 ( .A1(n8441), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10643 ( .A1(n8083), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8082) );
  MUX2_X1 U10644 ( .A(n8082), .B(P3_IR_REG_31__SCAN_IN), .S(n8081), .Z(n8085)
         );
  NAND2_X1 U10645 ( .A1(n8084), .A2(n8081), .ZN(n8110) );
  NAND2_X1 U10646 ( .A1(n8085), .A2(n8110), .ZN(n10625) );
  INV_X1 U10647 ( .A(SI_5_), .ZN(n10134) );
  OR2_X1 U10648 ( .A1(n8063), .A2(n10134), .ZN(n8089) );
  XNOR2_X1 U10649 ( .A(n8086), .B(n8087), .ZN(n10135) );
  OR2_X1 U10650 ( .A1(n8062), .A2(n10135), .ZN(n8088) );
  OAI211_X1 U10651 ( .C1(n10431), .C2(n10625), .A(n8089), .B(n8088), .ZN(
        n15408) );
  INV_X1 U10652 ( .A(n15408), .ZN(n9872) );
  NAND2_X1 U10653 ( .A1(n12520), .A2(n9872), .ZN(n8104) );
  OAI211_X1 U10654 ( .C1(n10430), .C2(n8456), .A(n8090), .B(n11094), .ZN(n8107) );
  NAND2_X1 U10655 ( .A1(n8091), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10656 ( .A1(n8442), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10657 ( .A1(n8092), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10658 ( .A1(n8114), .A2(n8093), .ZN(n11283) );
  NAND2_X1 U10659 ( .A1(n8395), .A2(n11283), .ZN(n8095) );
  NAND2_X1 U10660 ( .A1(n8441), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8094) );
  INV_X1 U10661 ( .A(SI_6_), .ZN(n10124) );
  NAND2_X1 U10662 ( .A1(n8110), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8101) );
  INV_X1 U10663 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8100) );
  OR2_X1 U10664 ( .A1(n10431), .A2(n10655), .ZN(n8102) );
  OAI211_X1 U10665 ( .C1(n8438), .C2(n10124), .A(n8103), .B(n8102), .ZN(n15413) );
  NAND2_X1 U10666 ( .A1(n12519), .A2(n11290), .ZN(n8458) );
  NAND2_X1 U10667 ( .A1(n8458), .A2(n8104), .ZN(n8105) );
  NAND2_X1 U10668 ( .A1(n11472), .A2(n15413), .ZN(n8459) );
  NAND3_X1 U10669 ( .A1(n12521), .A2(n10430), .A3(n11024), .ZN(n8106) );
  AOI21_X1 U10670 ( .B1(n8459), .B2(n8457), .A(n9936), .ZN(n8121) );
  NAND3_X1 U10671 ( .A1(n12519), .A2(n10430), .A3(n11290), .ZN(n8120) );
  XNOR2_X1 U10672 ( .A(n8109), .B(n8108), .ZN(n10125) );
  NAND2_X1 U10673 ( .A1(n10125), .A2(n8437), .ZN(n8113) );
  INV_X2 U10674 ( .A(n8438), .ZN(n8288) );
  NAND2_X1 U10675 ( .A1(n8124), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8111) );
  XNOR2_X1 U10676 ( .A(n8111), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U10677 ( .A1(n8288), .A2(SI_7_), .B1(n6875), .B2(n10877), .ZN(n8112) );
  NAND2_X1 U10678 ( .A1(n8113), .A2(n8112), .ZN(n11469) );
  NAND2_X1 U10679 ( .A1(n8424), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10680 ( .A1(n8347), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10681 ( .A1(n8114), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10682 ( .A1(n8128), .A2(n8115), .ZN(n11461) );
  NAND2_X1 U10683 ( .A1(n8395), .A2(n11461), .ZN(n8117) );
  NAND2_X1 U10684 ( .A1(n8441), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8116) );
  NAND4_X1 U10685 ( .A1(n8119), .A2(n8118), .A3(n8117), .A4(n8116), .ZN(n12518) );
  XNOR2_X1 U10686 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8122) );
  XNOR2_X1 U10687 ( .A(n8123), .B(n8122), .ZN(n10130) );
  NAND2_X1 U10688 ( .A1(n10130), .A2(n8437), .ZN(n8127) );
  INV_X1 U10689 ( .A(SI_8_), .ZN(n10131) );
  NAND2_X1 U10690 ( .A1(n8140), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8125) );
  AOI22_X1 U10691 ( .A1(n8288), .A2(n10131), .B1(n6875), .B2(n11144), .ZN(
        n8126) );
  NAND2_X1 U10692 ( .A1(n8127), .A2(n8126), .ZN(n11682) );
  NAND2_X1 U10693 ( .A1(n8091), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10694 ( .A1(n8442), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U10695 ( .A1(n8128), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U10696 ( .A1(n8148), .A2(n8129), .ZN(n11674) );
  NAND2_X1 U10697 ( .A1(n8395), .A2(n11674), .ZN(n8131) );
  NAND2_X1 U10698 ( .A1(n8441), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8130) );
  NAND4_X1 U10699 ( .A1(n8133), .A2(n8132), .A3(n8131), .A4(n8130), .ZN(n12517) );
  INV_X1 U10700 ( .A(n12517), .ZN(n11877) );
  NAND2_X1 U10701 ( .A1(n11682), .A2(n11877), .ZN(n9878) );
  OR2_X1 U10702 ( .A1(n11877), .A2(n11682), .ZN(n8134) );
  NAND2_X1 U10703 ( .A1(n9878), .A2(n8134), .ZN(n11443) );
  NAND2_X1 U10704 ( .A1(n11681), .A2(n11469), .ZN(n8461) );
  NAND2_X1 U10705 ( .A1(n15419), .A2(n12518), .ZN(n8135) );
  MUX2_X1 U10706 ( .A(n8461), .B(n8135), .S(n9936), .Z(n8136) );
  XNOR2_X1 U10707 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8137) );
  XNOR2_X1 U10708 ( .A(n8138), .B(n8137), .ZN(n10101) );
  NAND2_X1 U10709 ( .A1(n10101), .A2(n8437), .ZN(n8147) );
  INV_X1 U10710 ( .A(SI_9_), .ZN(n10102) );
  OR2_X2 U10711 ( .A1(n8140), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U10712 ( .A1(n8142), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8141) );
  MUX2_X1 U10713 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8141), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8145) );
  INV_X1 U10714 ( .A(n8142), .ZN(n8144) );
  INV_X1 U10715 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U10716 ( .A1(n8144), .A2(n8143), .ZN(n8173) );
  NAND2_X1 U10717 ( .A1(n8145), .A2(n8173), .ZN(n11379) );
  AOI22_X1 U10718 ( .A1(n8288), .A2(n10102), .B1(n11379), .B2(n6875), .ZN(
        n8146) );
  NAND2_X1 U10719 ( .A1(n8347), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10720 ( .A1(n8441), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10721 ( .A1(n8148), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U10722 ( .A1(n8164), .A2(n8149), .ZN(n11879) );
  NAND2_X1 U10723 ( .A1(n8395), .A2(n11879), .ZN(n8151) );
  NAND2_X1 U10724 ( .A1(n8091), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8150) );
  NAND4_X1 U10725 ( .A1(n8153), .A2(n8152), .A3(n8151), .A4(n8150), .ZN(n12516) );
  INV_X1 U10726 ( .A(n12516), .ZN(n12021) );
  XNOR2_X1 U10727 ( .A(n11882), .B(n12021), .ZN(n11565) );
  MUX2_X1 U10728 ( .A(n11877), .B(n11682), .S(n10430), .Z(n8154) );
  NAND2_X1 U10729 ( .A1(n8154), .A2(n9878), .ZN(n8155) );
  OR2_X1 U10730 ( .A1(n11882), .A2(n9936), .ZN(n8157) );
  NAND2_X1 U10731 ( .A1(n11882), .A2(n9936), .ZN(n8156) );
  MUX2_X1 U10732 ( .A(n8157), .B(n8156), .S(n12516), .Z(n8170) );
  XNOR2_X1 U10733 ( .A(n10154), .B(P2_DATAO_REG_10__SCAN_IN), .ZN(n8158) );
  XNOR2_X1 U10734 ( .A(n8159), .B(n8158), .ZN(n10129) );
  NAND2_X1 U10735 ( .A1(n10129), .A2(n8437), .ZN(n8163) );
  NAND2_X1 U10736 ( .A1(n8173), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8161) );
  INV_X1 U10737 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8160) );
  AOI22_X1 U10738 ( .A1(n11722), .A2(n6875), .B1(n8288), .B2(n10128), .ZN(
        n8162) );
  NAND2_X1 U10739 ( .A1(n8424), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10740 ( .A1(n8442), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10741 ( .A1(n8164), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10742 ( .A1(n8177), .A2(n8165), .ZN(n11964) );
  NAND2_X1 U10743 ( .A1(n8395), .A2(n11964), .ZN(n8167) );
  NAND2_X1 U10744 ( .A1(n8441), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8166) );
  NAND4_X1 U10745 ( .A1(n8169), .A2(n8168), .A3(n8167), .A4(n8166), .ZN(n12162) );
  OR2_X1 U10746 ( .A1(n12022), .A2(n12162), .ZN(n8466) );
  NAND2_X1 U10747 ( .A1(n12022), .A2(n12162), .ZN(n8465) );
  XNOR2_X1 U10748 ( .A(n10185), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8171) );
  XNOR2_X1 U10749 ( .A(n8172), .B(n8171), .ZN(n10156) );
  NAND2_X1 U10750 ( .A1(n10156), .A2(n8437), .ZN(n8176) );
  OAI21_X1 U10751 ( .B1(n8173), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8174) );
  XNOR2_X1 U10752 ( .A(n8174), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U10753 ( .A1(n11732), .A2(n6875), .B1(SI_11_), .B2(n8288), .ZN(
        n8175) );
  NAND2_X1 U10754 ( .A1(n8424), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10755 ( .A1(n8347), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8180) );
  XNOR2_X1 U10756 ( .A(n8177), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U10757 ( .A1(n8395), .A2(n12468), .ZN(n8179) );
  NAND2_X1 U10758 ( .A1(n8441), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8178) );
  OR2_X1 U10759 ( .A1(n12469), .A2(n12386), .ZN(n8201) );
  NAND2_X1 U10760 ( .A1(n12469), .A2(n12386), .ZN(n8467) );
  MUX2_X1 U10761 ( .A(n8466), .B(n8465), .S(n9936), .Z(n8182) );
  NAND2_X1 U10762 ( .A1(n11800), .A2(n8182), .ZN(n8199) );
  XNOR2_X1 U10763 ( .A(n8184), .B(n8183), .ZN(n10182) );
  NAND2_X1 U10764 ( .A1(n10182), .A2(n8437), .ZN(n8190) );
  INV_X1 U10765 ( .A(SI_12_), .ZN(n10183) );
  NAND2_X1 U10766 ( .A1(n8185), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8186) );
  MUX2_X1 U10767 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8186), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8188) );
  NAND2_X1 U10768 ( .A1(n8188), .A2(n8187), .ZN(n12560) );
  AOI22_X1 U10769 ( .A1(n8288), .A2(n10183), .B1(n6875), .B2(n12560), .ZN(
        n8189) );
  NAND2_X1 U10770 ( .A1(n8190), .A2(n8189), .ZN(n12387) );
  NAND2_X1 U10771 ( .A1(n8424), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10772 ( .A1(n8442), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8196) );
  INV_X1 U10773 ( .A(n8191), .ZN(n8192) );
  NAND2_X1 U10774 ( .A1(n8192), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10775 ( .A1(n8211), .A2(n8193), .ZN(n12390) );
  NAND2_X1 U10776 ( .A1(n8395), .A2(n12390), .ZN(n8195) );
  NAND2_X1 U10777 ( .A1(n8441), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8194) );
  AND2_X1 U10778 ( .A1(n8470), .A2(n8467), .ZN(n8198) );
  OAI22_X1 U10779 ( .A1(n8200), .A2(n8199), .B1(n10430), .B2(n8198), .ZN(n8203) );
  NAND2_X1 U10780 ( .A1(n12387), .A2(n12514), .ZN(n8469) );
  AOI21_X1 U10781 ( .B1(n8469), .B2(n8201), .A(n9936), .ZN(n8202) );
  AOI21_X1 U10782 ( .B1(n8203), .B2(n8469), .A(n8202), .ZN(n8218) );
  NAND2_X1 U10783 ( .A1(n8204), .A2(n10235), .ZN(n8230) );
  OR2_X1 U10784 ( .A1(n8204), .A2(n10235), .ZN(n8205) );
  NAND2_X1 U10785 ( .A1(n8230), .A2(n8205), .ZN(n8231) );
  XNOR2_X1 U10786 ( .A(n8231), .B(n10241), .ZN(n10388) );
  NAND2_X1 U10787 ( .A1(n10388), .A2(n8437), .ZN(n8210) );
  NAND2_X1 U10788 ( .A1(n8187), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8206) );
  MUX2_X1 U10789 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8206), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n8208) );
  INV_X1 U10790 ( .A(n8222), .ZN(n8207) );
  NAND2_X1 U10791 ( .A1(n8208), .A2(n8207), .ZN(n12573) );
  AOI22_X1 U10792 ( .A1(n8288), .A2(n10389), .B1(n6875), .B2(n12573), .ZN(
        n8209) );
  NAND2_X1 U10793 ( .A1(n8424), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10794 ( .A1(n8442), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U10795 ( .A1(n8211), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10796 ( .A1(n8237), .A2(n8212), .ZN(n12872) );
  NAND2_X1 U10797 ( .A1(n8395), .A2(n12872), .ZN(n8214) );
  NAND2_X1 U10798 ( .A1(n8441), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10799 ( .A1(n12868), .A2(n12513), .ZN(n8472) );
  OAI21_X1 U10800 ( .B1(n9936), .B2(n8470), .A(n12034), .ZN(n8217) );
  XNOR2_X1 U10801 ( .A(n8220), .B(n8219), .ZN(n10420) );
  NAND2_X1 U10802 ( .A1(n10420), .A2(n8437), .ZN(n8225) );
  NAND2_X1 U10803 ( .A1(n8247), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8223) );
  XNOR2_X1 U10804 ( .A(n8223), .B(n8246), .ZN(n12624) );
  INV_X1 U10805 ( .A(n12624), .ZN(n12630) );
  AOI22_X1 U10806 ( .A1(n8288), .A2(SI_15_), .B1(n12630), .B2(n6875), .ZN(
        n8224) );
  NAND2_X1 U10807 ( .A1(n8239), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10808 ( .A1(n8253), .A2(n8226), .ZN(n12854) );
  NAND2_X1 U10809 ( .A1(n12854), .A2(n8395), .ZN(n8229) );
  AOI22_X1 U10810 ( .A1(n8424), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n8347), .B2(
        P3_REG1_REG_15__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10811 ( .A1(n8441), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8227) );
  OR2_X1 U10812 ( .A1(n13006), .A2(n12405), .ZN(n8257) );
  NAND2_X1 U10813 ( .A1(n13006), .A2(n12405), .ZN(n8475) );
  NAND2_X1 U10814 ( .A1(n8257), .A2(n8475), .ZN(n12857) );
  INV_X1 U10815 ( .A(n12857), .ZN(n8540) );
  MUX2_X1 U10816 ( .A(n8471), .B(n8472), .S(n10430), .Z(n8242) );
  OAI21_X1 U10817 ( .B1(n8231), .B2(n10241), .A(n8230), .ZN(n8233) );
  XNOR2_X1 U10818 ( .A(n8233), .B(n8232), .ZN(n10548) );
  NAND2_X1 U10819 ( .A1(n10548), .A2(n8437), .ZN(n8236) );
  OR2_X1 U10820 ( .A1(n8222), .A2(n13017), .ZN(n8234) );
  XNOR2_X1 U10821 ( .A(n8234), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U10822 ( .A1(n8288), .A2(SI_14_), .B1(n6875), .B2(n12576), .ZN(
        n8235) );
  NAND2_X1 U10823 ( .A1(n8237), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10824 ( .A1(n8239), .A2(n8238), .ZN(n12346) );
  AOI22_X1 U10825 ( .A1(n12346), .A2(n8395), .B1(n8441), .B2(
        P3_REG0_REG_14__SCAN_IN), .ZN(n8241) );
  AOI22_X1 U10826 ( .A1(n8424), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n8442), .B2(
        P3_REG1_REG_14__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U10827 ( .A(n12942), .B(n12859), .ZN(n12046) );
  NAND4_X1 U10828 ( .A1(n8243), .A2(n8540), .A3(n8242), .A4(n12046), .ZN(n8261) );
  OR2_X1 U10829 ( .A1(n12942), .A2(n12500), .ZN(n8258) );
  XNOR2_X1 U10830 ( .A(n8245), .B(n8244), .ZN(n10545) );
  NAND2_X1 U10831 ( .A1(n10545), .A2(n8437), .ZN(n8251) );
  INV_X1 U10832 ( .A(n8270), .ZN(n8248) );
  NAND2_X1 U10833 ( .A1(n8248), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U10834 ( .A(n8249), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U10835 ( .A1(n8288), .A2(SI_16_), .B1(n6875), .B2(n12653), .ZN(
        n8250) );
  INV_X1 U10836 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12999) );
  INV_X1 U10837 ( .A(n8252), .ZN(n8291) );
  NAND2_X1 U10838 ( .A1(n8253), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10839 ( .A1(n8291), .A2(n8254), .ZN(n12850) );
  NAND2_X1 U10840 ( .A1(n12850), .A2(n8395), .ZN(n8256) );
  AOI22_X1 U10841 ( .A1(n8424), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n8442), .B2(
        P3_REG1_REG_16__SCAN_IN), .ZN(n8255) );
  OR2_X1 U10842 ( .A1(n13000), .A2(n12417), .ZN(n8477) );
  OAI211_X1 U10843 ( .C1(n12857), .C2(n8258), .A(n8477), .B(n8257), .ZN(n8259)
         );
  NAND2_X1 U10844 ( .A1(n8259), .A2(n9936), .ZN(n8260) );
  NAND2_X1 U10845 ( .A1(n13000), .A2(n12417), .ZN(n8478) );
  AOI21_X1 U10846 ( .B1(n8261), .B2(n8260), .A(n7490), .ZN(n8264) );
  NAND2_X1 U10847 ( .A1(n12942), .A2(n12500), .ZN(n8474) );
  OAI211_X1 U10848 ( .C1(n12857), .C2(n8474), .A(n8478), .B(n8475), .ZN(n8262)
         );
  AND2_X1 U10849 ( .A1(n8262), .A2(n10430), .ZN(n8263) );
  OAI22_X1 U10850 ( .A1(n8264), .A2(n8263), .B1(n9936), .B2(n8477), .ZN(n8300)
         );
  OR2_X1 U10851 ( .A1(n8266), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U10852 ( .A1(n8268), .A2(n8267), .ZN(n10818) );
  OR2_X1 U10853 ( .A1(n10818), .A2(n8389), .ZN(n8274) );
  NAND2_X1 U10854 ( .A1(n8270), .A2(n8269), .ZN(n8285) );
  NAND2_X1 U10855 ( .A1(n6425), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10856 ( .A(n8271), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12702) );
  NOR2_X1 U10857 ( .A1(n8438), .A2(n10819), .ZN(n8272) );
  AOI21_X1 U10858 ( .B1(n12702), .B2(n6875), .A(n8272), .ZN(n8273) );
  NAND2_X1 U10859 ( .A1(n8293), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U10860 ( .A1(n8308), .A2(n8275), .ZN(n12828) );
  NAND2_X1 U10861 ( .A1(n12828), .A2(n8395), .ZN(n8280) );
  INV_X1 U10862 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U10863 ( .A1(n8424), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10864 ( .A1(n8347), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8276) );
  OAI211_X1 U10865 ( .C1(n12992), .C2(n8409), .A(n8277), .B(n8276), .ZN(n8278)
         );
  INV_X1 U10866 ( .A(n8278), .ZN(n8279) );
  NAND2_X1 U10867 ( .A1(n12993), .A2(n12473), .ZN(n8479) );
  OR2_X1 U10868 ( .A1(n8282), .A2(n8281), .ZN(n8283) );
  NAND2_X1 U10869 ( .A1(n8284), .A2(n8283), .ZN(n10815) );
  NAND2_X1 U10870 ( .A1(n10815), .A2(n8437), .ZN(n8290) );
  NAND2_X1 U10871 ( .A1(n8285), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8286) );
  MUX2_X1 U10872 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8286), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8287) );
  NAND2_X1 U10873 ( .A1(n8287), .A2(n6425), .ZN(n12666) );
  AOI22_X1 U10874 ( .A1(n12666), .A2(n6875), .B1(n8288), .B2(n10817), .ZN(
        n8289) );
  NAND2_X1 U10875 ( .A1(n8291), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10876 ( .A1(n8293), .A2(n8292), .ZN(n12836) );
  NAND2_X1 U10877 ( .A1(n12836), .A2(n8395), .ZN(n8299) );
  INV_X1 U10878 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10879 ( .A1(n8424), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10880 ( .A1(n8442), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8294) );
  OAI211_X1 U10881 ( .C1(n8296), .C2(n8409), .A(n8295), .B(n8294), .ZN(n8297)
         );
  INV_X1 U10882 ( .A(n8297), .ZN(n8298) );
  NAND2_X1 U10883 ( .A1(n12935), .A2(n12846), .ZN(n8481) );
  NAND2_X1 U10884 ( .A1(n12812), .A2(n8481), .ZN(n9890) );
  OR2_X1 U10885 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  NAND2_X1 U10886 ( .A1(n8304), .A2(n8303), .ZN(n12159) );
  OAI22_X1 U10887 ( .A1(n9951), .A2(n10431), .B1(SI_19_), .B2(n8438), .ZN(
        n8307) );
  NAND2_X1 U10888 ( .A1(n8308), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10889 ( .A1(n8329), .A2(n8309), .ZN(n12807) );
  NAND2_X1 U10890 ( .A1(n12807), .A2(n8395), .ZN(n8315) );
  INV_X1 U10891 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U10892 ( .A1(n8441), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10893 ( .A1(n8442), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8310) );
  OAI211_X1 U10894 ( .C1(n8312), .C2(n12809), .A(n8311), .B(n8310), .ZN(n8313)
         );
  INV_X1 U10895 ( .A(n8313), .ZN(n8314) );
  NAND2_X2 U10896 ( .A1(n8315), .A2(n8314), .ZN(n12825) );
  INV_X1 U10897 ( .A(n12825), .ZN(n12441) );
  NAND2_X1 U10898 ( .A1(n12811), .A2(n12441), .ZN(n8485) );
  NAND2_X1 U10899 ( .A1(n8485), .A2(n9936), .ZN(n8320) );
  INV_X1 U10900 ( .A(n12812), .ZN(n12818) );
  NAND2_X1 U10901 ( .A1(n12822), .A2(n12818), .ZN(n8316) );
  NAND2_X1 U10902 ( .A1(n8316), .A2(n8479), .ZN(n8318) );
  OR2_X1 U10903 ( .A1(n12811), .A2(n12441), .ZN(n8480) );
  NAND3_X1 U10904 ( .A1(n8480), .A2(n10430), .A3(n12813), .ZN(n8317) );
  OAI21_X1 U10905 ( .B1(n8320), .B2(n8318), .A(n8317), .ZN(n8322) );
  INV_X1 U10906 ( .A(n8481), .ZN(n8319) );
  NAND3_X1 U10907 ( .A1(n8320), .A2(n8319), .A3(n8479), .ZN(n8321) );
  OR2_X1 U10908 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  NAND2_X1 U10909 ( .A1(n8326), .A2(n8325), .ZN(n11133) );
  INV_X1 U10910 ( .A(SI_20_), .ZN(n15447) );
  OR2_X1 U10911 ( .A1(n8438), .A2(n15447), .ZN(n8327) );
  NAND2_X1 U10912 ( .A1(n8329), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10913 ( .A1(n8344), .A2(n8330), .ZN(n12801) );
  NAND2_X1 U10914 ( .A1(n12801), .A2(n8395), .ZN(n8335) );
  INV_X1 U10915 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U10916 ( .A1(n8424), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10917 ( .A1(n8442), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8331) );
  OAI211_X1 U10918 ( .C1(n12985), .C2(n8409), .A(n8332), .B(n8331), .ZN(n8333)
         );
  INV_X1 U10919 ( .A(n8333), .ZN(n8334) );
  INV_X1 U10920 ( .A(n12805), .ZN(n8336) );
  NAND2_X1 U10921 ( .A1(n12986), .A2(n8336), .ZN(n8353) );
  NAND2_X1 U10922 ( .A1(n8486), .A2(n8353), .ZN(n9892) );
  INV_X1 U10923 ( .A(n9892), .ZN(n12797) );
  MUX2_X1 U10924 ( .A(n8480), .B(n8485), .S(n10430), .Z(n8337) );
  OR2_X1 U10925 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  NAND2_X1 U10926 ( .A1(n8341), .A2(n8340), .ZN(n11181) );
  INV_X1 U10927 ( .A(SI_21_), .ZN(n11180) );
  OR2_X1 U10928 ( .A1(n8438), .A2(n11180), .ZN(n8342) );
  NAND2_X1 U10929 ( .A1(n8344), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8345) );
  NAND2_X1 U10930 ( .A1(n8346), .A2(n8345), .ZN(n12791) );
  NAND2_X1 U10931 ( .A1(n12791), .A2(n8395), .ZN(n8352) );
  INV_X1 U10932 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U10933 ( .A1(n8424), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8349) );
  NAND2_X1 U10934 ( .A1(n8347), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8348) );
  OAI211_X1 U10935 ( .C1(n12979), .C2(n8409), .A(n8349), .B(n8348), .ZN(n8350)
         );
  INV_X1 U10936 ( .A(n8350), .ZN(n8351) );
  XNOR2_X1 U10937 ( .A(n12980), .B(n12798), .ZN(n12787) );
  MUX2_X1 U10938 ( .A(n8486), .B(n8353), .S(n9936), .Z(n8354) );
  INV_X1 U10939 ( .A(n12798), .ZN(n12189) );
  NAND2_X1 U10940 ( .A1(n12980), .A2(n12189), .ZN(n8487) );
  OR2_X1 U10941 ( .A1(n12980), .A2(n12189), .ZN(n12773) );
  MUX2_X1 U10942 ( .A(n8487), .B(n12773), .S(n9936), .Z(n8355) );
  NAND2_X1 U10943 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  OR2_X1 U10944 ( .A1(n8438), .A2(n11529), .ZN(n8360) );
  NAND2_X1 U10945 ( .A1(n6456), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10946 ( .A1(n12770), .A2(n8053), .ZN(n8368) );
  INV_X1 U10947 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U10948 ( .A1(n8424), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10949 ( .A1(n8442), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8364) );
  OAI211_X1 U10950 ( .C1(n12967), .C2(n8409), .A(n8365), .B(n8364), .ZN(n8366)
         );
  INV_X1 U10951 ( .A(n8366), .ZN(n8367) );
  NAND2_X1 U10952 ( .A1(n12968), .A2(n12459), .ZN(n8371) );
  MUX2_X1 U10953 ( .A(n8489), .B(n8488), .S(n10430), .Z(n8369) );
  INV_X1 U10954 ( .A(n8369), .ZN(n8370) );
  MUX2_X1 U10955 ( .A(n8371), .B(n8492), .S(n9936), .Z(n8372) );
  INV_X1 U10956 ( .A(n12742), .ZN(n8496) );
  NAND2_X1 U10957 ( .A1(n12909), .A2(n9936), .ZN(n8375) );
  OR2_X1 U10958 ( .A1(n12909), .A2(n9936), .ZN(n8374) );
  MUX2_X1 U10959 ( .A(n8375), .B(n8374), .S(n12767), .Z(n8376) );
  NOR2_X1 U10960 ( .A1(n8499), .A2(n10430), .ZN(n8379) );
  NAND2_X1 U10961 ( .A1(n8383), .A2(n8382), .ZN(n8386) );
  INV_X1 U10962 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U10963 ( .A1(n12218), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8402) );
  INV_X1 U10964 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U10965 ( .A1(n14098), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8384) );
  AND2_X1 U10966 ( .A1(n8402), .A2(n8384), .ZN(n8385) );
  NAND2_X1 U10967 ( .A1(n8386), .A2(n8385), .ZN(n8403) );
  OR2_X1 U10968 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  NAND2_X1 U10969 ( .A1(n8403), .A2(n8387), .ZN(n13026) );
  INV_X1 U10970 ( .A(SI_28_), .ZN(n13028) );
  OR2_X1 U10971 ( .A1(n8438), .A2(n13028), .ZN(n8388) );
  NAND2_X1 U10972 ( .A1(n8390), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10973 ( .A1(n12065), .A2(n8391), .ZN(n12714) );
  INV_X1 U10974 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n15532) );
  NAND2_X1 U10975 ( .A1(n8424), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8393) );
  NAND2_X1 U10976 ( .A1(n8442), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8392) );
  OAI211_X1 U10977 ( .C1(n15532), .C2(n8409), .A(n8393), .B(n8392), .ZN(n8394)
         );
  NAND2_X1 U10978 ( .A1(n12715), .A2(n12511), .ZN(n8502) );
  NAND2_X1 U10979 ( .A1(n8501), .A2(n8396), .ZN(n8397) );
  NAND2_X1 U10980 ( .A1(n8397), .A2(n8399), .ZN(n8398) );
  OAI211_X1 U10981 ( .C1(n7487), .C2(n8401), .A(n9907), .B(n8400), .ZN(n8415)
         );
  NAND2_X1 U10982 ( .A1(n8403), .A2(n8402), .ZN(n8418) );
  INV_X1 U10983 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12072) );
  XNOR2_X1 U10984 ( .A(n12072), .B(P1_DATAO_REG_29__SCAN_IN), .ZN(n8416) );
  XNOR2_X1 U10985 ( .A(n8418), .B(n8416), .ZN(n13022) );
  NAND2_X1 U10986 ( .A1(n13022), .A2(n8437), .ZN(n8405) );
  INV_X1 U10987 ( .A(SI_29_), .ZN(n13025) );
  OR2_X1 U10988 ( .A1(n8438), .A2(n13025), .ZN(n8404) );
  INV_X1 U10989 ( .A(n12065), .ZN(n8406) );
  NAND2_X1 U10990 ( .A1(n8406), .A2(n8395), .ZN(n8447) );
  INV_X1 U10991 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U10992 ( .A1(n8347), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10993 ( .A1(n8424), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8407) );
  OAI211_X1 U10994 ( .C1(n8409), .C2(n12147), .A(n8408), .B(n8407), .ZN(n8410)
         );
  INV_X1 U10995 ( .A(n8410), .ZN(n8411) );
  NAND2_X1 U10996 ( .A1(n8447), .A2(n8411), .ZN(n12510) );
  INV_X1 U10997 ( .A(n12510), .ZN(n8412) );
  INV_X1 U10998 ( .A(n12140), .ZN(n8414) );
  MUX2_X1 U10999 ( .A(n8502), .B(n8504), .S(n10430), .Z(n8413) );
  INV_X1 U11000 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U11001 ( .A1(n8418), .A2(n8417), .ZN(n8420) );
  NAND2_X1 U11002 ( .A1(n12072), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8419) );
  INV_X1 U11003 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15104) );
  XNOR2_X1 U11004 ( .A(n15104), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n8421) );
  XNOR2_X1 U11005 ( .A(n8434), .B(n8421), .ZN(n12057) );
  NAND2_X1 U11006 ( .A1(n12057), .A2(n8437), .ZN(n8423) );
  INV_X1 U11007 ( .A(SI_30_), .ZN(n12059) );
  OR2_X1 U11008 ( .A1(n8438), .A2(n12059), .ZN(n8422) );
  NAND2_X1 U11009 ( .A1(n8441), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U11010 ( .A1(n8424), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U11011 ( .A1(n8347), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8425) );
  AND3_X1 U11012 ( .A1(n8427), .A2(n8426), .A3(n8425), .ZN(n8428) );
  AND2_X1 U11013 ( .A1(n8447), .A2(n8428), .ZN(n12143) );
  NAND2_X1 U11014 ( .A1(n8526), .A2(n12143), .ZN(n8507) );
  AND2_X1 U11015 ( .A1(n8507), .A2(n8525), .ZN(n8429) );
  INV_X1 U11016 ( .A(n12143), .ZN(n12509) );
  AND2_X1 U11017 ( .A1(n12068), .A2(n12509), .ZN(n8550) );
  AOI21_X1 U11018 ( .B1(n8430), .B2(n8429), .A(n8550), .ZN(n8432) );
  INV_X1 U11019 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13368) );
  NOR2_X1 U11020 ( .A1(n13368), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8433) );
  OAI22_X1 U11021 ( .A1(n8434), .A2(n8433), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n15104), .ZN(n8436) );
  XNOR2_X1 U11022 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n8435) );
  XNOR2_X1 U11023 ( .A(n8436), .B(n8435), .ZN(n13015) );
  NAND2_X1 U11024 ( .A1(n13015), .A2(n8437), .ZN(n8440) );
  INV_X1 U11025 ( .A(SI_31_), .ZN(n13021) );
  OR2_X1 U11026 ( .A1(n8438), .A2(n13021), .ZN(n8439) );
  NAND2_X1 U11027 ( .A1(n8441), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U11028 ( .A1(n8424), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U11029 ( .A1(n8442), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8443) );
  AND3_X1 U11030 ( .A1(n8445), .A2(n8444), .A3(n8443), .ZN(n8446) );
  NAND2_X1 U11031 ( .A1(n8508), .A2(n12062), .ZN(n8549) );
  OR2_X1 U11032 ( .A1(n10558), .A2(P3_U3151), .ZN(n11527) );
  NAND2_X1 U11033 ( .A1(n12877), .A2(n8451), .ZN(n8453) );
  INV_X1 U11034 ( .A(n10936), .ZN(n10930) );
  NAND2_X1 U11035 ( .A1(n10929), .A2(n8455), .ZN(n10980) );
  INV_X1 U11036 ( .A(n10987), .ZN(n10982) );
  NAND2_X1 U11037 ( .A1(n8459), .A2(n8458), .ZN(n11217) );
  INV_X1 U11038 ( .A(n11217), .ZN(n11215) );
  NAND2_X1 U11039 ( .A1(n11216), .A2(n11215), .ZN(n8460) );
  NAND2_X1 U11040 ( .A1(n11457), .A2(n11456), .ZN(n8462) );
  OR2_X1 U11041 ( .A1(n11682), .A2(n12517), .ZN(n8463) );
  NAND2_X1 U11042 ( .A1(n11882), .A2(n12516), .ZN(n8464) );
  NAND2_X1 U11043 ( .A1(n12853), .A2(n8540), .ZN(n8476) );
  NAND2_X1 U11044 ( .A1(n8479), .A2(n12812), .ZN(n8484) );
  NAND2_X1 U11045 ( .A1(n8480), .A2(n8485), .ZN(n12814) );
  OAI21_X1 U11046 ( .B1(n8484), .B2(n8481), .A(n12813), .ZN(n8482) );
  NOR2_X1 U11047 ( .A1(n12814), .A2(n8482), .ZN(n8483) );
  NAND2_X1 U11048 ( .A1(n12794), .A2(n8486), .ZN(n12785) );
  AND2_X1 U11049 ( .A1(n12773), .A2(n8488), .ZN(n8491) );
  INV_X1 U11050 ( .A(n8489), .ZN(n8490) );
  NAND2_X1 U11051 ( .A1(n12764), .A2(n12765), .ZN(n8493) );
  INV_X1 U11052 ( .A(n12757), .ZN(n8494) );
  NAND2_X1 U11053 ( .A1(n12909), .A2(n12357), .ZN(n8495) );
  INV_X1 U11054 ( .A(n8499), .ZN(n8500) );
  INV_X1 U11055 ( .A(n8502), .ZN(n8503) );
  INV_X1 U11056 ( .A(n8505), .ZN(n8506) );
  NAND2_X1 U11057 ( .A1(n6485), .A2(n8507), .ZN(n8552) );
  OR2_X1 U11058 ( .A1(n8508), .A2(n6417), .ZN(n8510) );
  INV_X1 U11059 ( .A(n12062), .ZN(n12508) );
  AND2_X1 U11060 ( .A1(n12508), .A2(n9951), .ZN(n8509) );
  NAND2_X1 U11061 ( .A1(n8512), .A2(n8509), .ZN(n8515) );
  NAND2_X1 U11062 ( .A1(n8510), .A2(n8515), .ZN(n8520) );
  NAND2_X1 U11063 ( .A1(n8552), .A2(n8520), .ZN(n8519) );
  AOI21_X1 U11064 ( .B1(n12068), .B2(n8525), .A(n6417), .ZN(n8511) );
  NAND2_X1 U11065 ( .A1(n10983), .A2(n9938), .ZN(n9909) );
  AOI21_X1 U11066 ( .B1(n12950), .B2(n8511), .A(n9909), .ZN(n8518) );
  NAND2_X1 U11067 ( .A1(n8512), .A2(n12508), .ZN(n8513) );
  NAND3_X1 U11068 ( .A1(n8513), .A2(n8508), .A3(n6417), .ZN(n8514) );
  OAI21_X1 U11069 ( .B1(n8515), .B2(n8525), .A(n8514), .ZN(n8516) );
  INV_X1 U11070 ( .A(n8516), .ZN(n8517) );
  INV_X1 U11071 ( .A(n8530), .ZN(n8522) );
  OR2_X1 U11072 ( .A1(n8520), .A2(n11527), .ZN(n8521) );
  NAND2_X1 U11073 ( .A1(n8524), .A2(n8523), .ZN(n8579) );
  INV_X1 U11074 ( .A(n11527), .ZN(n8573) );
  INV_X1 U11075 ( .A(n8525), .ZN(n8528) );
  AND2_X1 U11076 ( .A1(n8526), .A2(n12062), .ZN(n8527) );
  OR4_X1 U11077 ( .A1(n8552), .A2(n9951), .A3(n8528), .A4(n8527), .ZN(n8529)
         );
  NOR2_X1 U11078 ( .A1(n11007), .A2(n9871), .ZN(n8536) );
  INV_X1 U11079 ( .A(n8531), .ZN(n8532) );
  OR2_X1 U11080 ( .A1(n8532), .A2(n11004), .ZN(n10578) );
  NOR2_X1 U11081 ( .A1(n10578), .A2(n10936), .ZN(n8535) );
  NOR2_X1 U11082 ( .A1(n12882), .A2(n10987), .ZN(n8534) );
  NAND4_X1 U11083 ( .A1(n8536), .A2(n8535), .A3(n8534), .A4(n11215), .ZN(n8537) );
  NOR3_X1 U11084 ( .A1(n8537), .A2(n11454), .A3(n9877), .ZN(n8538) );
  AND4_X1 U11085 ( .A1(n11800), .A2(n7754), .A3(n11565), .A4(n8538), .ZN(n8539) );
  NAND4_X1 U11086 ( .A1(n8540), .A2(n12034), .A3(n11913), .A4(n8539), .ZN(
        n8541) );
  NOR2_X1 U11087 ( .A1(n9890), .A2(n8541), .ZN(n8542) );
  NAND4_X1 U11088 ( .A1(n12822), .A2(n12845), .A3(n8542), .A4(n12046), .ZN(
        n8543) );
  NOR2_X1 U11089 ( .A1(n12814), .A2(n8543), .ZN(n8544) );
  NAND3_X1 U11090 ( .A1(n12787), .A2(n12797), .A3(n8544), .ZN(n8545) );
  OR3_X1 U11091 ( .A1(n9899), .A2(n12777), .A3(n8545), .ZN(n8546) );
  NOR3_X1 U11092 ( .A1(n12742), .A2(n12757), .A3(n8546), .ZN(n8547) );
  NAND4_X1 U11093 ( .A1(n9907), .A2(n12725), .A3(n12734), .A4(n8547), .ZN(
        n8548) );
  OR2_X1 U11094 ( .A1(n12140), .A2(n8548), .ZN(n8553) );
  INV_X1 U11095 ( .A(n8549), .ZN(n8551) );
  NAND2_X1 U11096 ( .A1(n11179), .A2(n9938), .ZN(n10795) );
  NAND2_X1 U11097 ( .A1(n8554), .A2(n7839), .ZN(n8577) );
  NAND2_X1 U11098 ( .A1(n6417), .A2(n11134), .ZN(n9944) );
  NAND2_X1 U11099 ( .A1(n8560), .A2(n8559), .ZN(n8567) );
  NAND2_X1 U11100 ( .A1(n8567), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8561) );
  MUX2_X1 U11101 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8561), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8563) );
  NAND2_X1 U11102 ( .A1(n8563), .A2(n8562), .ZN(n12071) );
  INV_X1 U11103 ( .A(n12071), .ZN(n8570) );
  NAND2_X1 U11104 ( .A1(n8564), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U11105 ( .A1(n8567), .A2(n8566), .ZN(n9915) );
  NAND2_X1 U11106 ( .A1(n8562), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8568) );
  NOR2_X1 U11107 ( .A1(n9915), .A2(n13040), .ZN(n8569) );
  NAND2_X1 U11108 ( .A1(n8570), .A2(n8569), .ZN(n10557) );
  INV_X1 U11109 ( .A(n13027), .ZN(n8572) );
  NAND3_X1 U11110 ( .A1(n10807), .A2(n8572), .A3(n13031), .ZN(n8575) );
  INV_X1 U11111 ( .A(P3_B_REG_SCAN_IN), .ZN(n12060) );
  AOI21_X1 U11112 ( .B1(n8573), .B2(n9952), .A(n12060), .ZN(n8574) );
  NAND2_X1 U11113 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  NAND4_X1 U11114 ( .A1(n8580), .A2(n8579), .A3(n8578), .A4(n7829), .ZN(
        P3_U3296) );
  INV_X1 U11115 ( .A(n8818), .ZN(n8581) );
  AND2_X1 U11116 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8583) );
  INV_X1 U11117 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13065) );
  NAND2_X1 U11118 ( .A1(n9139), .A2(n13065), .ZN(n8585) );
  AND2_X1 U11119 ( .A1(n9164), .A2(n8585), .ZN(n13742) );
  NOR2_X1 U11120 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8591) );
  NOR2_X1 U11121 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n8592) );
  INV_X1 U11122 ( .A(n8599), .ZN(n8701) );
  NAND2_X1 U11123 ( .A1(n13742), .A2(n9294), .ZN(n8609) );
  INV_X1 U11124 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8606) );
  INV_X4 U11125 ( .A(n9042), .ZN(n13362) );
  NAND2_X1 U11126 ( .A1(n13362), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8605) );
  INV_X1 U11127 ( .A(n8742), .ZN(n9099) );
  NAND2_X1 U11128 ( .A1(n9079), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8604) );
  OAI211_X1 U11129 ( .C1(n13365), .C2(n8606), .A(n8605), .B(n8604), .ZN(n8607)
         );
  INV_X1 U11130 ( .A(n8607), .ZN(n8608) );
  INV_X1 U11131 ( .A(n9232), .ZN(n9246) );
  NOR2_X1 U11132 ( .A1(n8696), .A2(n8763), .ZN(n8613) );
  NOR2_X2 U11133 ( .A1(n6467), .A2(n8696), .ZN(n13421) );
  INV_X1 U11134 ( .A(n8706), .ZN(n8969) );
  INV_X1 U11135 ( .A(n8616), .ZN(n8617) );
  OAI21_X1 U11136 ( .B1(n8969), .B2(n8617), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8618) );
  MUX2_X1 U11137 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8618), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8619) );
  NAND2_X1 U11138 ( .A1(n13584), .A2(n13926), .ZN(n13062) );
  INV_X1 U11139 ( .A(n13062), .ZN(n9148) );
  MUX2_X1 U11140 ( .A(n11132), .B(n11101), .S(n10093), .Z(n9074) );
  XNOR2_X1 U11141 ( .A(n8643), .B(SI_7_), .ZN(n8833) );
  INV_X1 U11142 ( .A(n8833), .ZN(n8642) );
  NAND2_X1 U11143 ( .A1(n8625), .A2(SI_2_), .ZN(n8757) );
  NAND2_X1 U11144 ( .A1(n8757), .A2(n10121), .ZN(n8623) );
  INV_X1 U11145 ( .A(n8760), .ZN(n8622) );
  NAND2_X1 U11146 ( .A1(n8760), .A2(n10121), .ZN(n8624) );
  AND2_X1 U11147 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8626) );
  AND2_X1 U11148 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8627) );
  INV_X1 U11149 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U11150 ( .A1(n8714), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U11151 ( .C1(n8714), .C2(n10109), .A(n8628), .B(n10094), .ZN(n8629) );
  NAND2_X1 U11152 ( .A1(n8713), .A2(n8629), .ZN(n8632) );
  NAND2_X1 U11153 ( .A1(n8714), .A2(n10092), .ZN(n8630) );
  OAI211_X1 U11154 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n8714), .A(n8630), .B(
        SI_1_), .ZN(n8631) );
  NAND2_X1 U11155 ( .A1(n8632), .A2(n8631), .ZN(n8756) );
  MUX2_X1 U11156 ( .A(n10060), .B(n10087), .S(n8714), .Z(n8634) );
  XNOR2_X1 U11157 ( .A(n8634), .B(SI_4_), .ZN(n8776) );
  INV_X1 U11158 ( .A(n8634), .ZN(n8635) );
  NAND2_X1 U11159 ( .A1(n8635), .A2(SI_4_), .ZN(n8636) );
  MUX2_X1 U11160 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8714), .Z(n8638) );
  XNOR2_X1 U11161 ( .A(n8638), .B(SI_5_), .ZN(n8809) );
  INV_X1 U11162 ( .A(n8809), .ZN(n8637) );
  NAND2_X1 U11163 ( .A1(n8638), .A2(SI_5_), .ZN(n8639) );
  NAND2_X1 U11164 ( .A1(n8640), .A2(SI_6_), .ZN(n8641) );
  NAND2_X1 U11165 ( .A1(n8643), .A2(SI_7_), .ZN(n8644) );
  MUX2_X1 U11166 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6410), .Z(n8646) );
  XNOR2_X1 U11167 ( .A(n8646), .B(SI_8_), .ZN(n8851) );
  INV_X1 U11168 ( .A(n8851), .ZN(n8645) );
  NAND2_X1 U11169 ( .A1(n8646), .A2(SI_8_), .ZN(n8647) );
  MUX2_X1 U11170 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6409), .Z(n8649) );
  INV_X1 U11171 ( .A(n8869), .ZN(n8648) );
  MUX2_X1 U11172 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10093), .Z(n8888) );
  INV_X1 U11173 ( .A(n8888), .ZN(n8650) );
  NAND2_X1 U11174 ( .A1(n8650), .A2(n10128), .ZN(n8651) );
  MUX2_X1 U11175 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10093), .Z(n8660) );
  NAND2_X1 U11176 ( .A1(n8660), .A2(SI_12_), .ZN(n8930) );
  INV_X1 U11177 ( .A(n8658), .ZN(n8652) );
  NAND2_X1 U11178 ( .A1(n8652), .A2(SI_11_), .ZN(n8909) );
  NAND2_X1 U11179 ( .A1(n8930), .A2(n8909), .ZN(n8949) );
  INV_X1 U11180 ( .A(n8949), .ZN(n8656) );
  MUX2_X1 U11181 ( .A(n10235), .B(n10241), .S(n7400), .Z(n8653) );
  NAND2_X1 U11182 ( .A1(n8653), .A2(n10389), .ZN(n8663) );
  INV_X1 U11183 ( .A(n8653), .ZN(n8654) );
  NAND2_X1 U11184 ( .A1(n8654), .A2(SI_13_), .ZN(n8655) );
  NAND2_X1 U11185 ( .A1(n8888), .A2(SI_10_), .ZN(n8907) );
  INV_X1 U11186 ( .A(SI_11_), .ZN(n10158) );
  NAND2_X1 U11187 ( .A1(n8659), .A2(n8930), .ZN(n8662) );
  INV_X1 U11188 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U11189 ( .A1(n8661), .A2(n10183), .ZN(n8929) );
  MUX2_X1 U11190 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6409), .Z(n8992) );
  NOR2_X1 U11191 ( .A1(n8992), .A2(SI_14_), .ZN(n8670) );
  MUX2_X1 U11192 ( .A(n10494), .B(n15545), .S(n10093), .Z(n8665) );
  NAND2_X1 U11193 ( .A1(n8665), .A2(n10421), .ZN(n8671) );
  INV_X1 U11194 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U11195 ( .A1(n8666), .A2(SI_15_), .ZN(n8667) );
  NAND2_X1 U11196 ( .A1(n8671), .A2(n8667), .ZN(n8994) );
  INV_X1 U11197 ( .A(n8992), .ZN(n8668) );
  NOR2_X1 U11198 ( .A1(n8668), .A2(n10549), .ZN(n8669) );
  MUX2_X1 U11199 ( .A(n10370), .B(n10368), .S(n6409), .Z(n8672) );
  INV_X1 U11200 ( .A(n8672), .ZN(n8673) );
  NAND2_X1 U11201 ( .A1(n8673), .A2(SI_16_), .ZN(n8674) );
  MUX2_X1 U11202 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10093), .Z(n9028) );
  INV_X1 U11203 ( .A(n9028), .ZN(n8677) );
  MUX2_X1 U11204 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6410), .Z(n9054) );
  MUX2_X1 U11205 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10093), .Z(n8679) );
  XNOR2_X1 U11206 ( .A(n8679), .B(SI_19_), .ZN(n9089) );
  INV_X1 U11207 ( .A(n9054), .ZN(n9087) );
  NOR2_X1 U11208 ( .A1(n9087), .A2(n10819), .ZN(n8678) );
  INV_X1 U11209 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U11210 ( .A1(n8680), .A2(n12158), .ZN(n8681) );
  NAND2_X1 U11211 ( .A1(n8685), .A2(SI_20_), .ZN(n8682) );
  MUX2_X1 U11212 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6409), .Z(n8683) );
  OAI21_X1 U11213 ( .B1(SI_21_), .B2(n8683), .A(n8686), .ZN(n9103) );
  INV_X1 U11214 ( .A(n9103), .ZN(n8684) );
  MUX2_X1 U11215 ( .A(n8687), .B(n11272), .S(n7400), .Z(n8690) );
  NAND2_X1 U11216 ( .A1(n8690), .A2(n8688), .ZN(n8689) );
  INV_X1 U11217 ( .A(n8690), .ZN(n9134) );
  NAND2_X1 U11218 ( .A1(n9134), .A2(SI_22_), .ZN(n8691) );
  MUX2_X1 U11219 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10093), .Z(n9158) );
  NAND2_X1 U11220 ( .A1(n9153), .A2(n9158), .ZN(n9150) );
  NAND2_X1 U11221 ( .A1(n8693), .A2(n11529), .ZN(n8694) );
  NAND2_X1 U11222 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  OR2_X1 U11223 ( .A1(n13369), .A2(n8702), .ZN(n8703) );
  NAND2_X1 U11224 ( .A1(n9003), .A2(n8708), .ZN(n9031) );
  INV_X1 U11225 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8709) );
  AOI21_X1 U11226 ( .B1(n9033), .B2(n8709), .A(n8763), .ZN(n8710) );
  AND2_X1 U11227 ( .A1(n13195), .A2(n13421), .ZN(n13203) );
  XNOR2_X1 U11228 ( .A(n6414), .B(n13203), .ZN(n8712) );
  INV_X1 U11229 ( .A(n13203), .ZN(n13424) );
  NAND2_X2 U11230 ( .A1(n10909), .A2(n13424), .ZN(n8935) );
  XNOR2_X1 U11231 ( .A(n13978), .B(n9218), .ZN(n13060) );
  INV_X1 U11232 ( .A(n13060), .ZN(n9147) );
  XNOR2_X1 U11233 ( .A(n8713), .B(n10094), .ZN(n8716) );
  MUX2_X1 U11234 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n8714), .Z(n8715) );
  XNOR2_X1 U11235 ( .A(n8716), .B(n8715), .ZN(n10110) );
  INV_X1 U11236 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11237 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8717) );
  XNOR2_X1 U11238 ( .A(n8935), .B(n10017), .ZN(n8731) );
  INV_X1 U11239 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11240 ( .A1(n8743), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U11241 ( .A1(n13450), .A2(n8772), .ZN(n8732) );
  XNOR2_X1 U11242 ( .A(n8731), .B(n8732), .ZN(n10395) );
  NAND2_X1 U11243 ( .A1(n8742), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8724) );
  INV_X1 U11244 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11245 ( .A1(n8743), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11246 ( .A1(n6409), .A2(SI_0_), .ZN(n8726) );
  NAND2_X1 U11247 ( .A1(n8726), .A2(n8725), .ZN(n8728) );
  AND2_X1 U11248 ( .A1(n8728), .A2(n8727), .ZN(n14099) );
  MUX2_X1 U11249 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14099), .S(n10193), .Z(n13200) );
  NAND2_X1 U11250 ( .A1(n13200), .A2(n13889), .ZN(n8729) );
  AND2_X1 U11251 ( .A1(n10908), .A2(n8729), .ZN(n10552) );
  INV_X1 U11252 ( .A(n13200), .ZN(n10906) );
  NAND2_X1 U11253 ( .A1(n9109), .A2(n10906), .ZN(n8730) );
  NAND2_X1 U11254 ( .A1(n10552), .A2(n8730), .ZN(n10396) );
  NAND2_X1 U11255 ( .A1(n10395), .A2(n10396), .ZN(n8735) );
  INV_X1 U11256 ( .A(n8731), .ZN(n8733) );
  NAND2_X1 U11257 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U11258 ( .A1(n8735), .A2(n8734), .ZN(n10414) );
  XNOR2_X1 U11259 ( .A(n8736), .B(SI_2_), .ZN(n8755) );
  XNOR2_X1 U11260 ( .A(n8755), .B(n8756), .ZN(n10088) );
  OR2_X1 U11261 ( .A1(n8737), .A2(n8763), .ZN(n8739) );
  OR2_X1 U11262 ( .A1(n10193), .A2(n13458), .ZN(n8740) );
  XNOR2_X1 U11263 ( .A(n15361), .B(n8935), .ZN(n8750) );
  NAND2_X1 U11264 ( .A1(n9289), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11265 ( .A1(n8742), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11266 ( .A1(n8743), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8747) );
  INV_X1 U11267 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8744) );
  OR2_X1 U11268 ( .A1(n8745), .A2(n8744), .ZN(n8746) );
  NAND2_X1 U11269 ( .A1(n13449), .A2(n8772), .ZN(n8751) );
  XNOR2_X1 U11270 ( .A(n8750), .B(n8751), .ZN(n10415) );
  NAND2_X1 U11271 ( .A1(n10414), .A2(n10415), .ZN(n8754) );
  INV_X1 U11272 ( .A(n8750), .ZN(n8752) );
  NAND2_X1 U11273 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11274 ( .A1(n8754), .A2(n8753), .ZN(n10021) );
  INV_X1 U11275 ( .A(n8755), .ZN(n8759) );
  INV_X1 U11276 ( .A(n8756), .ZN(n8758) );
  OAI21_X1 U11277 ( .B1(n8759), .B2(n8758), .A(n8757), .ZN(n8762) );
  XNOR2_X1 U11278 ( .A(n8760), .B(SI_3_), .ZN(n8761) );
  XNOR2_X1 U11279 ( .A(n8762), .B(n8761), .ZN(n10084) );
  OR2_X1 U11280 ( .A1(n13369), .A2(n10085), .ZN(n8766) );
  OR2_X1 U11281 ( .A1(n8779), .A2(n8763), .ZN(n8764) );
  XNOR2_X1 U11282 ( .A(n8778), .B(n8764), .ZN(n13468) );
  OR2_X1 U11283 ( .A1(n10193), .A2(n13468), .ZN(n8765) );
  XNOR2_X1 U11284 ( .A(n9109), .B(n13218), .ZN(n10681) );
  NAND2_X1 U11285 ( .A1(n9289), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8771) );
  INV_X1 U11286 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8767) );
  NAND2_X1 U11287 ( .A1(n13362), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8769) );
  INV_X1 U11288 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U11289 ( .A1(n8960), .A2(n10024), .ZN(n8768) );
  INV_X1 U11290 ( .A(n10681), .ZN(n8774) );
  NAND2_X1 U11291 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  NAND2_X1 U11292 ( .A1(n8791), .A2(n8775), .ZN(n10023) );
  OR2_X2 U11293 ( .A1(n10021), .A2(n10023), .ZN(n10679) );
  BUF_X1 U11294 ( .A(n8935), .Z(n9109) );
  XNOR2_X1 U11295 ( .A(n8777), .B(n8776), .ZN(n10086) );
  OR2_X1 U11296 ( .A1(n13369), .A2(n10087), .ZN(n8783) );
  NAND2_X1 U11297 ( .A1(n8779), .A2(n8778), .ZN(n8798) );
  NAND2_X1 U11298 ( .A1(n8798), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8781) );
  XNOR2_X1 U11299 ( .A(n8781), .B(n8780), .ZN(n10219) );
  OR2_X1 U11300 ( .A1(n10193), .A2(n10219), .ZN(n8782) );
  XNOR2_X1 U11301 ( .A(n9109), .B(n15368), .ZN(n10830) );
  NAND2_X1 U11302 ( .A1(n9289), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11303 ( .A1(n9079), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8789) );
  INV_X1 U11304 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11305 ( .A1(n8785), .A2(n10024), .ZN(n8786) );
  AND2_X1 U11306 ( .A1(n8786), .A2(n8818), .ZN(n11656) );
  NAND2_X1 U11307 ( .A1(n8960), .A2(n11656), .ZN(n8788) );
  NAND2_X1 U11308 ( .A1(n13362), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8787) );
  NAND4_X1 U11309 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n13447) );
  NAND2_X1 U11310 ( .A1(n13447), .A2(n13926), .ZN(n8793) );
  XNOR2_X1 U11311 ( .A(n10830), .B(n8793), .ZN(n10680) );
  AND2_X1 U11312 ( .A1(n10680), .A2(n8791), .ZN(n8792) );
  INV_X1 U11313 ( .A(n10830), .ZN(n8794) );
  NAND2_X1 U11314 ( .A1(n8794), .A2(n8793), .ZN(n8795) );
  XNOR2_X1 U11315 ( .A(n8797), .B(n8796), .ZN(n10064) );
  NAND2_X1 U11316 ( .A1(n10064), .A2(n13366), .ZN(n8802) );
  INV_X1 U11317 ( .A(n8811), .ZN(n8799) );
  NAND2_X1 U11318 ( .A1(n8799), .A2(n8812), .ZN(n8834) );
  NAND2_X1 U11319 ( .A1(n8834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8800) );
  XNOR2_X1 U11320 ( .A(n8800), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U11321 ( .A1(n9091), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9092), .B2(
        n13509), .ZN(n8801) );
  NAND2_X1 U11322 ( .A1(n8802), .A2(n8801), .ZN(n13235) );
  XNOR2_X1 U11323 ( .A(n11637), .B(n9162), .ZN(n11105) );
  NAND2_X1 U11324 ( .A1(n9079), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11325 ( .A1(n13362), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8807) );
  INV_X1 U11326 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11327 ( .A1(n8820), .A2(n8803), .ZN(n8804) );
  AND2_X1 U11328 ( .A1(n8841), .A2(n8804), .ZN(n11635) );
  NAND2_X1 U11329 ( .A1(n8960), .A2(n11635), .ZN(n8806) );
  NAND2_X1 U11330 ( .A1(n9289), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8805) );
  NAND4_X1 U11331 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n13445) );
  NAND2_X1 U11332 ( .A1(n13445), .A2(n13926), .ZN(n8827) );
  NAND2_X1 U11333 ( .A1(n11105), .A2(n8827), .ZN(n10920) );
  XNOR2_X1 U11334 ( .A(n8810), .B(n8809), .ZN(n10062) );
  NAND2_X1 U11335 ( .A1(n10062), .A2(n13366), .ZN(n8815) );
  NAND2_X1 U11336 ( .A1(n8811), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U11337 ( .A(n8813), .B(n8812), .ZN(n13489) );
  OR2_X1 U11338 ( .A1(n10193), .A2(n13489), .ZN(n8814) );
  INV_X1 U11339 ( .A(n10825), .ZN(n8825) );
  NAND2_X1 U11340 ( .A1(n9289), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11341 ( .A1(n9079), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8823) );
  INV_X1 U11342 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U11343 ( .A1(n8818), .A2(n8817), .ZN(n8819) );
  AND2_X1 U11344 ( .A1(n8820), .A2(n8819), .ZN(n11276) );
  NAND2_X1 U11345 ( .A1(n8960), .A2(n11276), .ZN(n8822) );
  NAND2_X1 U11346 ( .A1(n8743), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8821) );
  NAND4_X1 U11347 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n13446) );
  AND2_X1 U11348 ( .A1(n13446), .A2(n13926), .ZN(n8826) );
  INV_X1 U11349 ( .A(n8826), .ZN(n10824) );
  NAND2_X1 U11350 ( .A1(n8825), .A2(n10824), .ZN(n10917) );
  NAND3_X1 U11351 ( .A1(n10920), .A2(n8826), .A3(n10825), .ZN(n8830) );
  INV_X1 U11352 ( .A(n11105), .ZN(n8829) );
  INV_X1 U11353 ( .A(n8827), .ZN(n8828) );
  NAND2_X1 U11354 ( .A1(n8829), .A2(n8828), .ZN(n10919) );
  AND2_X1 U11355 ( .A1(n8830), .A2(n10919), .ZN(n8831) );
  NAND2_X1 U11356 ( .A1(n10096), .A2(n6408), .ZN(n8839) );
  INV_X1 U11357 ( .A(n8834), .ZN(n8836) );
  INV_X1 U11358 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11359 ( .A1(n8836), .A2(n8835), .ZN(n8853) );
  NAND2_X1 U11360 ( .A1(n8853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11361 ( .A(n8837), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U11362 ( .A1(n9091), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9092), .B2(
        n10283), .ZN(n8838) );
  XNOR2_X1 U11363 ( .A(n15376), .B(n9162), .ZN(n8847) );
  NAND2_X1 U11364 ( .A1(n9289), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U11365 ( .A1(n9079), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11366 ( .A1(n8841), .A2(n8840), .ZN(n8842) );
  AND2_X1 U11367 ( .A1(n8858), .A2(n8842), .ZN(n11421) );
  NAND2_X1 U11368 ( .A1(n8960), .A2(n11421), .ZN(n8844) );
  NAND2_X1 U11369 ( .A1(n13362), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8843) );
  NAND4_X1 U11370 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n13444) );
  AND2_X1 U11371 ( .A1(n13444), .A2(n13926), .ZN(n8848) );
  NAND2_X1 U11372 ( .A1(n8847), .A2(n8848), .ZN(n8864) );
  INV_X1 U11373 ( .A(n8847), .ZN(n11060) );
  INV_X1 U11374 ( .A(n8848), .ZN(n8849) );
  NAND2_X1 U11375 ( .A1(n11060), .A2(n8849), .ZN(n8850) );
  AND2_X1 U11376 ( .A1(n8864), .A2(n8850), .ZN(n11102) );
  NAND2_X1 U11377 ( .A1(n10111), .A2(n6408), .ZN(n8856) );
  NAND2_X1 U11378 ( .A1(n8871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8854) );
  XNOR2_X1 U11379 ( .A(n8854), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U11380 ( .A1(n9091), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9092), .B2(
        n10302), .ZN(n8855) );
  XNOR2_X1 U11381 ( .A(n13246), .B(n9162), .ZN(n11207) );
  NAND2_X1 U11382 ( .A1(n9289), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U11383 ( .A1(n9079), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11384 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U11385 ( .A1(n8878), .A2(n8859), .ZN(n11069) );
  INV_X1 U11386 ( .A(n11069), .ZN(n11624) );
  NAND2_X1 U11387 ( .A1(n9294), .A2(n11624), .ZN(n8861) );
  NAND2_X1 U11388 ( .A1(n13362), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8860) );
  NAND4_X1 U11389 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n13443) );
  NAND2_X1 U11390 ( .A1(n13443), .A2(n13926), .ZN(n8866) );
  XNOR2_X1 U11391 ( .A(n11207), .B(n8866), .ZN(n11073) );
  AND2_X1 U11392 ( .A1(n11073), .A2(n8864), .ZN(n8865) );
  INV_X1 U11393 ( .A(n11207), .ZN(n8867) );
  NAND2_X1 U11394 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  NAND2_X1 U11395 ( .A1(n10144), .A2(n6408), .ZN(n8876) );
  INV_X1 U11396 ( .A(n8871), .ZN(n8873) );
  INV_X1 U11397 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U11398 ( .A1(n8873), .A2(n8872), .ZN(n8891) );
  NAND2_X1 U11399 ( .A1(n8891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8874) );
  XNOR2_X1 U11400 ( .A(n8874), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U11401 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n9091), .B1(n10663), 
        .B2(n9092), .ZN(n8875) );
  XNOR2_X1 U11402 ( .A(n14051), .B(n9282), .ZN(n8884) );
  NAND2_X1 U11403 ( .A1(n9289), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U11404 ( .A1(n9079), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U11405 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  AND2_X1 U11406 ( .A1(n8896), .A2(n8879), .ZN(n11202) );
  NAND2_X1 U11407 ( .A1(n8960), .A2(n11202), .ZN(n8881) );
  NAND2_X1 U11408 ( .A1(n13362), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8880) );
  NAND4_X1 U11409 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n13442) );
  NAND2_X1 U11410 ( .A1(n13442), .A2(n13926), .ZN(n8885) );
  XNOR2_X1 U11411 ( .A(n8884), .B(n8885), .ZN(n11208) );
  INV_X1 U11412 ( .A(n8884), .ZN(n8886) );
  NAND2_X1 U11413 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  XNOR2_X1 U11414 ( .A(n8888), .B(SI_10_), .ZN(n8889) );
  XNOR2_X1 U11415 ( .A(n8890), .B(n8889), .ZN(n10151) );
  NAND2_X1 U11416 ( .A1(n10151), .A2(n6408), .ZN(n8894) );
  NAND2_X1 U11417 ( .A1(n8910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8892) );
  AOI22_X1 U11418 ( .A1(n10714), .A2(n9092), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n9091), .ZN(n8893) );
  XNOR2_X1 U11419 ( .A(n11577), .B(n9218), .ZN(n8902) );
  NAND2_X1 U11420 ( .A1(n9289), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U11421 ( .A1(n9079), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8900) );
  INV_X1 U11422 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11423 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  AND2_X1 U11424 ( .A1(n8915), .A2(n8897), .ZN(n11578) );
  NAND2_X1 U11425 ( .A1(n8960), .A2(n11578), .ZN(n8899) );
  NAND2_X1 U11426 ( .A1(n13362), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8898) );
  NOR2_X1 U11427 ( .A1(n13256), .A2(n13889), .ZN(n8903) );
  NAND2_X1 U11428 ( .A1(n8902), .A2(n8903), .ZN(n8921) );
  INV_X1 U11429 ( .A(n8902), .ZN(n11602) );
  INV_X1 U11430 ( .A(n8903), .ZN(n8904) );
  NAND2_X1 U11431 ( .A1(n11602), .A2(n8904), .ZN(n8905) );
  NAND2_X1 U11432 ( .A1(n8921), .A2(n8905), .ZN(n11585) );
  INV_X1 U11433 ( .A(n11585), .ZN(n8906) );
  NAND2_X1 U11434 ( .A1(n8908), .A2(n8907), .ZN(n8950) );
  NAND2_X1 U11435 ( .A1(n8927), .A2(n8909), .ZN(n8928) );
  XNOR2_X1 U11436 ( .A(n8950), .B(n8928), .ZN(n10184) );
  NAND2_X1 U11437 ( .A1(n10184), .A2(n6408), .ZN(n8913) );
  OAI21_X1 U11438 ( .B1(n8910), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11439 ( .A(n8911), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U11440 ( .A1(n10965), .A2(n9092), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n9091), .ZN(n8912) );
  BUF_X1 U11441 ( .A(n8935), .Z(n9162) );
  XNOR2_X1 U11442 ( .A(n13609), .B(n9162), .ZN(n8925) );
  NAND2_X1 U11443 ( .A1(n9289), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U11444 ( .A1(n9079), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U11445 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  AND2_X1 U11446 ( .A1(n8938), .A2(n8916), .ZN(n11817) );
  NAND2_X1 U11447 ( .A1(n8960), .A2(n11817), .ZN(n8918) );
  NAND2_X1 U11448 ( .A1(n13362), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8917) );
  NOR2_X1 U11449 ( .A1(n13608), .A2(n13889), .ZN(n8923) );
  XNOR2_X1 U11450 ( .A(n8925), .B(n8923), .ZN(n11612) );
  AND2_X1 U11451 ( .A1(n11612), .A2(n8921), .ZN(n8922) );
  INV_X1 U11452 ( .A(n8923), .ZN(n8924) );
  NAND2_X1 U11453 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  NAND2_X1 U11454 ( .A1(n11608), .A2(n8926), .ZN(n11520) );
  AND2_X1 U11455 ( .A1(n8930), .A2(n8929), .ZN(n8931) );
  NAND2_X1 U11456 ( .A1(n8932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8933) );
  XNOR2_X1 U11457 ( .A(n8933), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U11458 ( .A1(n9091), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9092), 
        .B2(n15304), .ZN(n8934) );
  XNOR2_X1 U11459 ( .A(n13932), .B(n9282), .ZN(n8944) );
  NAND2_X1 U11460 ( .A1(n9079), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U11461 ( .A1(n13362), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8942) );
  INV_X1 U11462 ( .A(n8936), .ZN(n8958) );
  NAND2_X1 U11463 ( .A1(n8938), .A2(n8937), .ZN(n8939) );
  AND2_X1 U11464 ( .A1(n8958), .A2(n8939), .ZN(n13929) );
  NAND2_X1 U11465 ( .A1(n9294), .A2(n13929), .ZN(n8941) );
  NAND2_X1 U11466 ( .A1(n9289), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8940) );
  OR2_X1 U11467 ( .A1(n13611), .A2(n13889), .ZN(n8945) );
  AND2_X1 U11468 ( .A1(n8944), .A2(n8945), .ZN(n11516) );
  INV_X1 U11469 ( .A(n8944), .ZN(n8947) );
  INV_X1 U11470 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11471 ( .A1(n8947), .A2(n8946), .ZN(n11517) );
  OAI21_X1 U11472 ( .B1(n11520), .B2(n11516), .A(n11517), .ZN(n11764) );
  XNOR2_X1 U11473 ( .A(n8952), .B(n8951), .ZN(n10233) );
  NAND2_X1 U11474 ( .A1(n10233), .A2(n6408), .ZN(n8956) );
  NAND2_X1 U11475 ( .A1(n8953), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8954) );
  XNOR2_X1 U11476 ( .A(n8954), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U11477 ( .A1(n9091), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9092), 
        .B2(n11504), .ZN(n8955) );
  XNOR2_X1 U11478 ( .A(n13912), .B(n9282), .ZN(n8963) );
  INV_X1 U11479 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U11480 ( .A1(n8958), .A2(n8957), .ZN(n8959) );
  AND2_X1 U11481 ( .A1(n8974), .A2(n8959), .ZN(n13910) );
  AOI22_X1 U11482 ( .A1(n13910), .A2(n8960), .B1(n13362), .B2(
        P2_REG2_REG_13__SCAN_IN), .ZN(n8962) );
  AOI22_X1 U11483 ( .A1(n9289), .A2(P2_REG0_REG_13__SCAN_IN), .B1(n9079), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n8961) );
  NOR2_X1 U11484 ( .A1(n13614), .A2(n13889), .ZN(n8964) );
  XNOR2_X1 U11485 ( .A(n8963), .B(n8964), .ZN(n11765) );
  NAND2_X1 U11486 ( .A1(n11764), .A2(n11765), .ZN(n8967) );
  INV_X1 U11487 ( .A(n8963), .ZN(n8965) );
  NAND2_X1 U11488 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U11489 ( .A1(n8968), .A2(n10549), .ZN(n8991) );
  XNOR2_X1 U11490 ( .A(n8993), .B(n8992), .ZN(n10390) );
  NAND2_X1 U11491 ( .A1(n10390), .A2(n6408), .ZN(n8972) );
  NAND2_X1 U11492 ( .A1(n8969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U11493 ( .A(n8970), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U11494 ( .A1(n9091), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9092), 
        .B2(n11507), .ZN(n8971) );
  XNOR2_X1 U11495 ( .A(n14025), .B(n9282), .ZN(n8979) );
  NAND2_X1 U11496 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  AND2_X1 U11497 ( .A1(n8986), .A2(n8975), .ZN(n13891) );
  NAND2_X1 U11498 ( .A1(n13891), .A2(n9294), .ZN(n8978) );
  AOI22_X1 U11499 ( .A1(n8742), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n13362), 
        .B2(P2_REG2_REG_14__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11500 ( .A1(n9289), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8976) );
  OR2_X1 U11501 ( .A1(n13868), .A2(n13889), .ZN(n8980) );
  NAND2_X1 U11502 ( .A1(n8979), .A2(n8980), .ZN(n8984) );
  INV_X1 U11503 ( .A(n8979), .ZN(n8982) );
  INV_X1 U11504 ( .A(n8980), .ZN(n8981) );
  NAND2_X1 U11505 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  NAND2_X1 U11506 ( .A1(n8984), .A2(n8983), .ZN(n13052) );
  INV_X1 U11507 ( .A(n8985), .ZN(n9010) );
  NAND2_X1 U11508 ( .A1(n8986), .A2(n11502), .ZN(n8987) );
  NAND2_X1 U11509 ( .A1(n9010), .A2(n8987), .ZN(n13874) );
  OR2_X1 U11510 ( .A1(n13874), .A2(n9223), .ZN(n8990) );
  AOI22_X1 U11511 ( .A1(n9289), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n9079), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11512 ( .A1(n13362), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8988) );
  NOR2_X1 U11513 ( .A1(n13620), .A2(n13889), .ZN(n9021) );
  OAI21_X1 U11514 ( .B1(n8993), .B2(n8992), .A(n8991), .ZN(n8996) );
  INV_X1 U11515 ( .A(n8994), .ZN(n8995) );
  XNOR2_X1 U11516 ( .A(n8996), .B(n8995), .ZN(n10492) );
  NAND2_X1 U11517 ( .A1(n10492), .A2(n13366), .ZN(n9001) );
  INV_X1 U11518 ( .A(n8997), .ZN(n8998) );
  NAND2_X1 U11519 ( .A1(n8998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8999) );
  XNOR2_X1 U11520 ( .A(n8999), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U11521 ( .A1(n9091), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9092), 
        .B2(n11667), .ZN(n9000) );
  XNOR2_X1 U11522 ( .A(n13878), .B(n9218), .ZN(n9019) );
  XNOR2_X1 U11523 ( .A(n9002), .B(n7848), .ZN(n10367) );
  NAND2_X1 U11524 ( .A1(n10367), .A2(n13366), .ZN(n9007) );
  INV_X1 U11525 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U11526 ( .A1(n9004), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9005) );
  XNOR2_X1 U11527 ( .A(n9005), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U11528 ( .A1(n9091), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9092), 
        .B2(n11696), .ZN(n9006) );
  XNOR2_X1 U11529 ( .A(n14013), .B(n9282), .ZN(n9022) );
  INV_X1 U11530 ( .A(n9008), .ZN(n9038) );
  INV_X1 U11531 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11532 ( .A1(n9010), .A2(n9009), .ZN(n9011) );
  NAND2_X1 U11533 ( .A1(n13854), .A2(n9294), .ZN(n9017) );
  INV_X1 U11534 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11535 ( .A1(n13362), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U11536 ( .A1(n9079), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9012) );
  OAI211_X1 U11537 ( .C1(n13365), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9015)
         );
  INV_X1 U11538 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U11539 ( .A1(n9017), .A2(n9016), .ZN(n13623) );
  AND2_X1 U11540 ( .A1(n13623), .A2(n13926), .ZN(n9023) );
  AND2_X1 U11541 ( .A1(n9022), .A2(n9023), .ZN(n9020) );
  AOI21_X1 U11542 ( .B1(n9021), .B2(n9019), .A(n9020), .ZN(n9018) );
  INV_X1 U11543 ( .A(n9019), .ZN(n13106) );
  INV_X1 U11544 ( .A(n9020), .ZN(n13104) );
  INV_X1 U11545 ( .A(n9021), .ZN(n13181) );
  NAND3_X1 U11546 ( .A1(n13106), .A2(n13104), .A3(n13181), .ZN(n9026) );
  INV_X1 U11547 ( .A(n9022), .ZN(n9025) );
  INV_X1 U11548 ( .A(n9023), .ZN(n9024) );
  NAND2_X1 U11549 ( .A1(n9025), .A2(n9024), .ZN(n13103) );
  AND2_X1 U11550 ( .A1(n9026), .A2(n13103), .ZN(n9027) );
  XNOR2_X1 U11551 ( .A(n9028), .B(n10817), .ZN(n9029) );
  XNOR2_X1 U11552 ( .A(n9030), .B(n9029), .ZN(n10495) );
  NAND2_X1 U11553 ( .A1(n10495), .A2(n6408), .ZN(n9036) );
  NAND2_X1 U11554 ( .A1(n9031), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9032) );
  MUX2_X1 U11555 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9032), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9034) );
  INV_X1 U11556 ( .A(n9033), .ZN(n9055) );
  AND2_X1 U11557 ( .A1(n9034), .A2(n9055), .ZN(n13520) );
  AOI22_X1 U11558 ( .A1(n13520), .A2(n9092), .B1(P1_DATAO_REG_17__SCAN_IN), 
        .B2(n9091), .ZN(n9035) );
  XNOR2_X1 U11559 ( .A(n14008), .B(n9218), .ZN(n9046) );
  INV_X1 U11560 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9037) );
  NAND2_X1 U11561 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NAND2_X1 U11562 ( .A1(n9059), .A2(n9039), .ZN(n13838) );
  OR2_X1 U11563 ( .A1(n13838), .A2(n9223), .ZN(n9045) );
  INV_X1 U11564 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U11565 ( .A1(n9079), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11566 ( .A1(n9289), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9040) );
  OAI211_X1 U11567 ( .C1(n13839), .C2(n9042), .A(n9041), .B(n9040), .ZN(n9043)
         );
  INV_X1 U11568 ( .A(n9043), .ZN(n9044) );
  NAND2_X1 U11569 ( .A1(n9045), .A2(n9044), .ZN(n13848) );
  NAND2_X1 U11570 ( .A1(n13848), .A2(n13926), .ZN(n9047) );
  NAND2_X1 U11571 ( .A1(n9046), .A2(n9047), .ZN(n9051) );
  INV_X1 U11572 ( .A(n9046), .ZN(n9049) );
  INV_X1 U11573 ( .A(n9047), .ZN(n9048) );
  NAND2_X1 U11574 ( .A1(n9049), .A2(n9048), .ZN(n9050) );
  AND2_X1 U11575 ( .A1(n9051), .A2(n9050), .ZN(n13116) );
  NAND2_X1 U11576 ( .A1(n9052), .A2(n10819), .ZN(n9053) );
  NAND2_X1 U11577 ( .A1(n9086), .A2(n9053), .ZN(n9088) );
  XNOR2_X1 U11578 ( .A(n9088), .B(n9054), .ZN(n10975) );
  NAND2_X1 U11579 ( .A1(n10975), .A2(n13366), .ZN(n9058) );
  NAND2_X1 U11580 ( .A1(n9055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9056) );
  XNOR2_X1 U11581 ( .A(n9056), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U11582 ( .A1(n13532), .A2(n9092), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n9091), .ZN(n9057) );
  XNOR2_X1 U11583 ( .A(n14004), .B(n9218), .ZN(n9067) );
  NAND2_X1 U11584 ( .A1(n9059), .A2(n13160), .ZN(n9060) );
  NAND2_X1 U11585 ( .A1(n9095), .A2(n9060), .ZN(n13822) );
  OR2_X1 U11586 ( .A1(n13822), .A2(n9223), .ZN(n9066) );
  INV_X1 U11587 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9063) );
  NAND2_X1 U11588 ( .A1(n9079), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U11589 ( .A1(n13362), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9061) );
  OAI211_X1 U11590 ( .C1(n13365), .C2(n9063), .A(n9062), .B(n9061), .ZN(n9064)
         );
  INV_X1 U11591 ( .A(n9064), .ZN(n9065) );
  NAND2_X1 U11592 ( .A1(n13797), .A2(n13926), .ZN(n9068) );
  XNOR2_X1 U11593 ( .A(n9067), .B(n9068), .ZN(n13158) );
  INV_X1 U11594 ( .A(n9067), .ZN(n9070) );
  INV_X1 U11595 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U11596 ( .A1(n9070), .A2(n9069), .ZN(n9071) );
  NAND2_X1 U11597 ( .A1(n9072), .A2(n15447), .ZN(n9073) );
  NAND2_X1 U11598 ( .A1(n9075), .A2(n9074), .ZN(n9076) );
  OR2_X1 U11599 ( .A1(n13369), .A2(n11101), .ZN(n9077) );
  XNOR2_X1 U11600 ( .A(n13993), .B(n9282), .ZN(n13083) );
  XNOR2_X1 U11601 ( .A(n9111), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13786) );
  NAND2_X1 U11602 ( .A1(n13786), .A2(n9294), .ZN(n9085) );
  INV_X1 U11603 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U11604 ( .A1(n13362), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U11605 ( .A1(n9079), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9080) );
  OAI211_X1 U11606 ( .C1(n13365), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9083)
         );
  INV_X1 U11607 ( .A(n9083), .ZN(n9084) );
  AND2_X1 U11608 ( .A1(n13798), .A2(n13926), .ZN(n9119) );
  NAND2_X1 U11609 ( .A1(n13083), .A2(n9119), .ZN(n9123) );
  OAI21_X1 U11610 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9090) );
  NAND2_X1 U11611 ( .A1(n11113), .A2(n6408), .ZN(n9094) );
  AOI22_X1 U11612 ( .A1(n13541), .A2(n9092), .B1(P1_DATAO_REG_19__SCAN_IN), 
        .B2(n9091), .ZN(n9093) );
  NAND2_X2 U11613 ( .A1(n9094), .A2(n9093), .ZN(n13997) );
  XNOR2_X1 U11614 ( .A(n13997), .B(n9282), .ZN(n13081) );
  NAND2_X1 U11615 ( .A1(n9095), .A2(n13075), .ZN(n9096) );
  NAND2_X1 U11616 ( .A1(n9111), .A2(n9096), .ZN(n13806) );
  INV_X1 U11617 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13534) );
  NAND2_X1 U11618 ( .A1(n9289), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11619 ( .A1(n13362), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9097) );
  OAI211_X1 U11620 ( .C1(n9099), .C2(n13534), .A(n9098), .B(n9097), .ZN(n9100)
         );
  INV_X1 U11621 ( .A(n9100), .ZN(n9101) );
  AND2_X1 U11622 ( .A1(n13628), .A2(n13926), .ZN(n9121) );
  NAND2_X1 U11623 ( .A1(n13081), .A2(n9121), .ZN(n13072) );
  OR2_X1 U11624 ( .A1(n11230), .A2(n9160), .ZN(n9108) );
  OR2_X1 U11625 ( .A1(n13369), .A2(n11128), .ZN(n9107) );
  XNOR2_X1 U11626 ( .A(n13988), .B(n9162), .ZN(n9129) );
  INV_X1 U11627 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13141) );
  INV_X1 U11628 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9110) );
  OAI21_X1 U11629 ( .B1(n9111), .B2(n13141), .A(n9110), .ZN(n9112) );
  AND2_X1 U11630 ( .A1(n9137), .A2(n9112), .ZN(n13769) );
  NAND2_X1 U11631 ( .A1(n13769), .A2(n9294), .ZN(n9118) );
  INV_X1 U11632 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U11633 ( .A1(n13362), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11634 ( .A1(n9079), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9113) );
  OAI211_X1 U11635 ( .C1(n13365), .C2(n9115), .A(n9114), .B(n9113), .ZN(n9116)
         );
  INV_X1 U11636 ( .A(n9116), .ZN(n9117) );
  NAND2_X1 U11637 ( .A1(n13630), .A2(n13926), .ZN(n9127) );
  XNOR2_X1 U11638 ( .A(n9129), .B(n9127), .ZN(n13085) );
  INV_X1 U11639 ( .A(n13083), .ZN(n9120) );
  INV_X1 U11640 ( .A(n9119), .ZN(n13082) );
  NAND2_X1 U11641 ( .A1(n9120), .A2(n13082), .ZN(n13086) );
  INV_X1 U11642 ( .A(n13081), .ZN(n9122) );
  INV_X1 U11643 ( .A(n9121), .ZN(n13084) );
  AND2_X1 U11644 ( .A1(n9122), .A2(n13084), .ZN(n13073) );
  NAND2_X1 U11645 ( .A1(n9123), .A2(n13073), .ZN(n9124) );
  AND3_X1 U11646 ( .A1(n13085), .A2(n13086), .A3(n9124), .ZN(n9125) );
  NAND2_X1 U11647 ( .A1(n9126), .A2(n9125), .ZN(n13087) );
  INV_X1 U11648 ( .A(n9127), .ZN(n9128) );
  NAND2_X1 U11649 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  OR2_X1 U11650 ( .A1(n9131), .A2(SI_22_), .ZN(n9133) );
  NAND2_X1 U11651 ( .A1(n9131), .A2(SI_22_), .ZN(n9132) );
  NAND2_X1 U11652 ( .A1(n9133), .A2(n9132), .ZN(n9604) );
  XNOR2_X1 U11653 ( .A(n9604), .B(n9134), .ZN(n11270) );
  NAND2_X1 U11654 ( .A1(n11270), .A2(n13366), .ZN(n9136) );
  OR2_X1 U11655 ( .A1(n13369), .A2(n11272), .ZN(n9135) );
  XNOR2_X1 U11656 ( .A(n13982), .B(n9282), .ZN(n9146) );
  INV_X1 U11657 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13154) );
  NAND2_X1 U11658 ( .A1(n9137), .A2(n13154), .ZN(n9138) );
  NAND2_X1 U11659 ( .A1(n9139), .A2(n9138), .ZN(n13751) );
  OR2_X1 U11660 ( .A1(n13751), .A2(n9223), .ZN(n9145) );
  INV_X1 U11661 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U11662 ( .A1(n13362), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U11663 ( .A1(n9079), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9140) );
  OAI211_X1 U11664 ( .C1(n13365), .C2(n9142), .A(n9141), .B(n9140), .ZN(n9143)
         );
  INV_X1 U11665 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U11666 ( .A1(n13631), .A2(n13926), .ZN(n13058) );
  MUX2_X1 U11667 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10093), .Z(n9149) );
  NAND2_X1 U11668 ( .A1(n9149), .A2(SI_24_), .ZN(n9174) );
  OAI21_X1 U11669 ( .B1(SI_24_), .B2(n9149), .A(n9174), .ZN(n9155) );
  AND2_X1 U11670 ( .A1(n9150), .A2(n9155), .ZN(n9151) );
  NAND2_X1 U11671 ( .A1(n9152), .A2(n9151), .ZN(n9159) );
  INV_X1 U11672 ( .A(n9158), .ZN(n9154) );
  INV_X1 U11673 ( .A(n9155), .ZN(n9156) );
  NAND2_X1 U11674 ( .A1(n9159), .A2(n9175), .ZN(n11530) );
  OR2_X1 U11675 ( .A1(n13369), .A2(n11478), .ZN(n9161) );
  XNOR2_X1 U11676 ( .A(n13972), .B(n9162), .ZN(n13094) );
  INV_X1 U11677 ( .A(n9164), .ZN(n9163) );
  INV_X1 U11678 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U11679 ( .A1(n9164), .A2(n13131), .ZN(n9165) );
  NAND2_X1 U11680 ( .A1(n9197), .A2(n9165), .ZN(n13722) );
  INV_X1 U11681 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11682 ( .A1(n13362), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11683 ( .A1(n9079), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9166) );
  OAI211_X1 U11684 ( .C1(n13365), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9169)
         );
  INV_X1 U11685 ( .A(n9169), .ZN(n9170) );
  NAND2_X2 U11686 ( .A1(n9171), .A2(n9170), .ZN(n13701) );
  AND2_X1 U11687 ( .A1(n13701), .A2(n13926), .ZN(n9172) );
  NAND2_X1 U11688 ( .A1(n13094), .A2(n9172), .ZN(n9173) );
  OAI21_X1 U11689 ( .B1(n13094), .B2(n9172), .A(n9173), .ZN(n13126) );
  INV_X1 U11690 ( .A(n9173), .ZN(n9188) );
  MUX2_X1 U11691 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6410), .Z(n9189) );
  XNOR2_X1 U11692 ( .A(n9189), .B(SI_25_), .ZN(n9191) );
  XNOR2_X1 U11693 ( .A(n9192), .B(n9191), .ZN(n11571) );
  NAND2_X1 U11694 ( .A1(n11571), .A2(n6408), .ZN(n9177) );
  OR2_X1 U11695 ( .A1(n13369), .A2(n11573), .ZN(n9176) );
  XNOR2_X1 U11696 ( .A(n13708), .B(n9218), .ZN(n9184) );
  XNOR2_X1 U11697 ( .A(n9197), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13706) );
  NAND2_X1 U11698 ( .A1(n13706), .A2(n9294), .ZN(n9183) );
  INV_X1 U11699 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11700 ( .A1(n9289), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11701 ( .A1(n9079), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9178) );
  OAI211_X1 U11702 ( .C1(n9180), .C2(n9042), .A(n9179), .B(n9178), .ZN(n9181)
         );
  INV_X1 U11703 ( .A(n9181), .ZN(n9182) );
  NOR2_X1 U11704 ( .A1(n13637), .A2(n13889), .ZN(n9185) );
  NAND2_X1 U11705 ( .A1(n9184), .A2(n9185), .ZN(n9207) );
  INV_X1 U11706 ( .A(n9184), .ZN(n13175) );
  INV_X1 U11707 ( .A(n9185), .ZN(n9186) );
  NAND2_X1 U11708 ( .A1(n13175), .A2(n9186), .ZN(n9187) );
  AND2_X1 U11709 ( .A1(n9207), .A2(n9187), .ZN(n13093) );
  INV_X1 U11710 ( .A(n9189), .ZN(n9190) );
  MUX2_X1 U11711 ( .A(n15483), .B(n11784), .S(n6409), .Z(n9213) );
  XNOR2_X1 U11712 ( .A(n9213), .B(SI_26_), .ZN(n9193) );
  NAND2_X1 U11713 ( .A1(n11783), .A2(n13366), .ZN(n9195) );
  OR2_X1 U11714 ( .A1(n13369), .A2(n11784), .ZN(n9194) );
  XNOR2_X1 U11715 ( .A(n13692), .B(n9282), .ZN(n9209) );
  INV_X1 U11716 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13098) );
  INV_X1 U11717 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9196) );
  OAI21_X1 U11718 ( .B1(n9197), .B2(n13098), .A(n9196), .ZN(n9200) );
  INV_X1 U11719 ( .A(n9197), .ZN(n9199) );
  AND2_X1 U11720 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n9198) );
  NAND2_X1 U11721 ( .A1(n13690), .A2(n9294), .ZN(n9206) );
  INV_X1 U11722 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11723 ( .A1(n9079), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11724 ( .A1(n13362), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9201) );
  OAI211_X1 U11725 ( .C1(n9203), .C2(n13365), .A(n9202), .B(n9201), .ZN(n9204)
         );
  INV_X1 U11726 ( .A(n9204), .ZN(n9205) );
  NOR2_X1 U11727 ( .A1(n13667), .A2(n13889), .ZN(n9210) );
  XNOR2_X1 U11728 ( .A(n9209), .B(n9210), .ZN(n13176) );
  INV_X1 U11729 ( .A(n9213), .ZN(n9214) );
  MUX2_X1 U11730 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6409), .Z(n9818) );
  NAND2_X1 U11731 ( .A1(n12160), .A2(n6408), .ZN(n9217) );
  OR2_X1 U11732 ( .A1(n13369), .A2(n12161), .ZN(n9216) );
  XNOR2_X1 U11733 ( .A(n13960), .B(n9218), .ZN(n9264) );
  INV_X1 U11734 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11735 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND2_X1 U11736 ( .A1(n9274), .A2(n9222), .ZN(n13044) );
  INV_X1 U11737 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U11738 ( .A1(n13362), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11739 ( .A1(n9079), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9224) );
  OAI211_X1 U11740 ( .C1(n13365), .C2(n9226), .A(n9225), .B(n9224), .ZN(n9227)
         );
  INV_X1 U11741 ( .A(n9227), .ZN(n9228) );
  NOR2_X1 U11742 ( .A1(n13640), .A2(n13889), .ZN(n9230) );
  NAND2_X1 U11743 ( .A1(n9264), .A2(n9230), .ZN(n9286) );
  OAI21_X1 U11744 ( .B1(n9264), .B2(n9230), .A(n9286), .ZN(n13041) );
  INV_X1 U11745 ( .A(n11785), .ZN(n9243) );
  NAND2_X1 U11746 ( .A1(n9248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9237) );
  XNOR2_X1 U11747 ( .A(n11479), .B(P2_B_REG_SCAN_IN), .ZN(n9241) );
  NAND2_X1 U11748 ( .A1(n9238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9240) );
  INV_X1 U11749 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11750 ( .A1(n9241), .A2(n11572), .ZN(n9242) );
  INV_X1 U11751 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15357) );
  NAND2_X1 U11752 ( .A1(n15323), .A2(n15357), .ZN(n9245) );
  NAND2_X1 U11753 ( .A1(n11785), .A2(n11572), .ZN(n9244) );
  NAND2_X1 U11754 ( .A1(n9245), .A2(n9244), .ZN(n15358) );
  INV_X1 U11755 ( .A(n15358), .ZN(n9295) );
  NAND2_X1 U11756 ( .A1(n9246), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9247) );
  MUX2_X1 U11757 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9247), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n9249) );
  NAND2_X1 U11758 ( .A1(n9249), .A2(n9248), .ZN(n11331) );
  NOR2_X1 U11759 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n9253) );
  NOR4_X1 U11760 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9252) );
  NOR4_X1 U11761 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9251) );
  NOR4_X1 U11762 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9250) );
  NAND4_X1 U11763 ( .A1(n9253), .A2(n9252), .A3(n9251), .A4(n9250), .ZN(n9259)
         );
  NOR4_X1 U11764 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9257) );
  NOR4_X1 U11765 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9256) );
  NOR4_X1 U11766 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9255) );
  NOR4_X1 U11767 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9254) );
  NAND4_X1 U11768 ( .A1(n9257), .A2(n9256), .A3(n9255), .A4(n9254), .ZN(n9258)
         );
  OAI21_X1 U11769 ( .B1(n9259), .B2(n9258), .A(n15323), .ZN(n10011) );
  AND2_X1 U11770 ( .A1(n15359), .A2(n10011), .ZN(n9262) );
  INV_X1 U11771 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11772 ( .A1(n15323), .A2(n9260), .ZN(n9261) );
  NAND2_X1 U11773 ( .A1(n11785), .A2(n11479), .ZN(n15353) );
  INV_X1 U11774 ( .A(n10195), .ZN(n9297) );
  NOR2_X1 U11775 ( .A1(n15377), .A2(n9297), .ZN(n9263) );
  INV_X1 U11776 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U11777 ( .A1(n13182), .A2(n13926), .ZN(n13174) );
  NOR3_X1 U11778 ( .A1(n9265), .A2(n13640), .A3(n13174), .ZN(n9266) );
  INV_X1 U11779 ( .A(n9267), .ZN(n9268) );
  NAND2_X1 U11780 ( .A1(n9268), .A2(SI_27_), .ZN(n9270) );
  NAND2_X1 U11781 ( .A1(n9823), .A2(n9818), .ZN(n9269) );
  NAND2_X1 U11782 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  MUX2_X1 U11783 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6410), .Z(n9824) );
  XNOR2_X1 U11784 ( .A(n9824), .B(SI_28_), .ZN(n9817) );
  NAND2_X1 U11785 ( .A1(n14094), .A2(n13366), .ZN(n9273) );
  OR2_X1 U11786 ( .A1(n13369), .A2(n14098), .ZN(n9272) );
  INV_X1 U11787 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n15559) );
  NAND2_X1 U11788 ( .A1(n9274), .A2(n15559), .ZN(n9275) );
  NAND2_X1 U11789 ( .A1(n13654), .A2(n9294), .ZN(n9281) );
  INV_X1 U11790 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11791 ( .A1(n13362), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11792 ( .A1(n9079), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U11793 ( .C1(n13365), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9279)
         );
  INV_X1 U11794 ( .A(n9279), .ZN(n9280) );
  NOR2_X1 U11795 ( .A1(n13668), .A2(n13889), .ZN(n9283) );
  XNOR2_X1 U11796 ( .A(n9283), .B(n9282), .ZN(n9284) );
  XNOR2_X1 U11797 ( .A(n13656), .B(n9284), .ZN(n9287) );
  AND2_X1 U11798 ( .A1(n9287), .A2(n7851), .ZN(n9310) );
  INV_X1 U11799 ( .A(n13423), .ZN(n13435) );
  INV_X1 U11800 ( .A(n9288), .ZN(n13602) );
  INV_X1 U11801 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11802 ( .A1(n9289), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U11803 ( .A1(n13362), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9290) );
  OAI211_X1 U11804 ( .C1(n9292), .C2(n9099), .A(n9291), .B(n9290), .ZN(n9293)
         );
  AOI21_X1 U11805 ( .B1(n13602), .B2(n9294), .A(n9293), .ZN(n13391) );
  NAND2_X1 U11806 ( .A1(n9297), .A2(n10205), .ZN(n13871) );
  OAI22_X1 U11807 ( .A1(n13391), .A2(n13871), .B1(n13640), .B2(n13869), .ZN(
        n13651) );
  INV_X1 U11808 ( .A(n13654), .ZN(n9301) );
  NAND3_X1 U11809 ( .A1(n9295), .A2(n10382), .A3(n10011), .ZN(n9296) );
  NAND2_X1 U11810 ( .A1(n13541), .A2(n13195), .ZN(n13374) );
  NAND2_X1 U11811 ( .A1(n9296), .A2(n10371), .ZN(n9300) );
  NAND2_X1 U11812 ( .A1(n13423), .A2(n9297), .ZN(n10010) );
  AND2_X1 U11813 ( .A1(n10010), .A2(n9298), .ZN(n9299) );
  NAND2_X1 U11814 ( .A1(n9300), .A2(n9299), .ZN(n10397) );
  OAI22_X1 U11815 ( .A1(n9301), .A2(n13187), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15559), .ZN(n9307) );
  NOR2_X1 U11816 ( .A1(n9302), .A2(n13195), .ZN(n10015) );
  NAND2_X1 U11817 ( .A1(n9303), .A2(n10015), .ZN(n9305) );
  NOR2_X1 U11818 ( .A1(n13656), .A2(n13194), .ZN(n9306) );
  AOI211_X1 U11819 ( .C1(n13161), .C2(n13651), .A(n9307), .B(n9306), .ZN(n9308) );
  INV_X1 U11820 ( .A(n9308), .ZN(n9309) );
  NAND2_X1 U11821 ( .A1(n9312), .A2(n9311), .ZN(P2_U3192) );
  NAND3_X1 U11822 ( .A1(n9694), .A2(n9693), .A3(n9313), .ZN(n9702) );
  INV_X1 U11823 ( .A(n9702), .ZN(n9315) );
  NAND2_X1 U11824 ( .A1(n9317), .A2(n9316), .ZN(n9318) );
  INV_X1 U11825 ( .A(n9370), .ZN(n9320) );
  NOR2_X1 U11826 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9324) );
  NOR2_X1 U11827 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n9323) );
  NOR2_X1 U11828 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9322) );
  NAND3_X1 U11829 ( .A1(n9409), .A2(n9326), .A3(n9325), .ZN(n9327) );
  XNOR2_X2 U11830 ( .A(n9330), .B(n15446), .ZN(n9333) );
  INV_X1 U11831 ( .A(n9333), .ZN(n9335) );
  INV_X1 U11832 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14964) );
  OR2_X1 U11833 ( .A1(n9539), .A2(n14964), .ZN(n9357) );
  NAND2_X1 U11834 ( .A1(n9966), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9355) );
  INV_X1 U11835 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10246) );
  INV_X1 U11836 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10263) );
  OR2_X1 U11837 ( .A1(n9376), .A2(n10263), .ZN(n9354) );
  INV_X1 U11838 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9336) );
  INV_X1 U11839 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11840 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9341) );
  OR2_X1 U11841 ( .A1(n9347), .A2(n14503), .ZN(n9343) );
  INV_X1 U11842 ( .A(SI_0_), .ZN(n10099) );
  INV_X1 U11843 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9344) );
  OAI21_X1 U11844 ( .B1(n6410), .B2(n10099), .A(n9344), .ZN(n9345) );
  NAND2_X1 U11845 ( .A1(n9966), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9353) );
  INV_X1 U11846 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9348) );
  INV_X1 U11847 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9349) );
  NAND3_X1 U11848 ( .A1(n10840), .A2(n10843), .A3(n10839), .ZN(n10842) );
  NAND2_X1 U11849 ( .A1(n10842), .A2(n10840), .ZN(n11050) );
  INV_X1 U11850 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10245) );
  INV_X1 U11851 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9358) );
  OR2_X1 U11852 ( .A1(n9539), .A2(n9358), .ZN(n9359) );
  INV_X1 U11853 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10262) );
  OR2_X1 U11854 ( .A1(n9637), .A2(n10088), .ZN(n9365) );
  OR2_X1 U11855 ( .A1(n9347), .A2(n14522), .ZN(n9363) );
  NAND2_X1 U11856 ( .A1(n11050), .A2(n11051), .ZN(n11049) );
  NAND2_X1 U11857 ( .A1(n11049), .A2(n14267), .ZN(n9374) );
  NAND2_X1 U11858 ( .A1(n9966), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9369) );
  OR2_X1 U11859 ( .A1(n9539), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9368) );
  INV_X1 U11860 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10249) );
  INV_X1 U11861 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10267) );
  OR2_X1 U11862 ( .A1(n9376), .A2(n10267), .ZN(n9366) );
  NAND2_X1 U11863 ( .A1(n9370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9371) );
  OR2_X1 U11864 ( .A1(n10084), .A2(n9637), .ZN(n9373) );
  OR2_X1 U11865 ( .A1(n9384), .A2(n10061), .ZN(n9372) );
  OAI211_X1 U11866 ( .C1(n7116), .C2(n14538), .A(n9373), .B(n9372), .ZN(n15170) );
  NAND2_X1 U11867 ( .A1(n11343), .A2(n15170), .ZN(n14277) );
  NAND2_X1 U11868 ( .A1(n14497), .A2(n11342), .ZN(n14278) );
  NAND2_X1 U11869 ( .A1(n11343), .A2(n11342), .ZN(n9375) );
  NAND2_X1 U11870 ( .A1(n11119), .A2(n9375), .ZN(n15213) );
  NAND2_X1 U11871 ( .A1(n9966), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9380) );
  OAI21_X1 U11872 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n9390), .ZN(n15218) );
  OR2_X1 U11873 ( .A1(n9539), .A2(n15218), .ZN(n9379) );
  INV_X1 U11874 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10252) );
  OR2_X1 U11875 ( .A1(n6406), .A2(n10252), .ZN(n9378) );
  INV_X1 U11876 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n15219) );
  OR2_X1 U11877 ( .A1(n9376), .A2(n15219), .ZN(n9377) );
  NAND4_X1 U11878 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n14496) );
  NAND2_X1 U11879 ( .A1(n9381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9383) );
  INV_X1 U11880 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9382) );
  XNOR2_X1 U11881 ( .A(n9383), .B(n9382), .ZN(n15195) );
  OR2_X1 U11882 ( .A1(n9347), .A2(n15195), .ZN(n9386) );
  OR2_X1 U11883 ( .A1(n9384), .A2(n10060), .ZN(n9385) );
  XNOR2_X1 U11884 ( .A(n14496), .B(n15222), .ZN(n15206) );
  INV_X1 U11885 ( .A(n15206), .ZN(n15212) );
  NAND2_X1 U11886 ( .A1(n15213), .A2(n15212), .ZN(n15211) );
  INV_X1 U11887 ( .A(n14496), .ZN(n11348) );
  NAND2_X1 U11888 ( .A1(n11348), .A2(n15237), .ZN(n9387) );
  NAND2_X1 U11889 ( .A1(n9786), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9395) );
  INV_X1 U11890 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9388) );
  OR2_X1 U11891 ( .A1(n9535), .A2(n9388), .ZN(n9394) );
  INV_X1 U11892 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11893 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  NAND2_X1 U11894 ( .A1(n9403), .A2(n9391), .ZN(n11560) );
  OR2_X1 U11895 ( .A1(n9785), .A2(n11560), .ZN(n9393) );
  INV_X1 U11896 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10244) );
  OR2_X1 U11897 ( .A1(n6405), .A2(n10244), .ZN(n9392) );
  INV_X1 U11898 ( .A(n14495), .ZN(n11358) );
  NAND2_X1 U11899 ( .A1(n9845), .A2(n10062), .ZN(n9400) );
  XNOR2_X1 U11900 ( .A(n9397), .B(n9409), .ZN(n10313) );
  OR2_X1 U11901 ( .A1(n7116), .A2(n10313), .ZN(n9399) );
  OR2_X1 U11902 ( .A1(n9384), .A2(n10063), .ZN(n9398) );
  NAND2_X1 U11903 ( .A1(n11358), .A2(n11357), .ZN(n11298) );
  NAND2_X1 U11904 ( .A1(n14495), .A2(n15245), .ZN(n9401) );
  NAND2_X1 U11905 ( .A1(n11190), .A2(n14442), .ZN(n11191) );
  NAND2_X1 U11906 ( .A1(n11191), .A2(n11298), .ZN(n9416) );
  NAND2_X1 U11907 ( .A1(n9966), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9408) );
  INV_X1 U11908 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10320) );
  OR2_X1 U11909 ( .A1(n9376), .A2(n10320), .ZN(n9407) );
  INV_X1 U11910 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U11911 ( .A1(n9403), .A2(n9402), .ZN(n9404) );
  NAND2_X1 U11912 ( .A1(n9423), .A2(n9404), .ZN(n11372) );
  OR2_X1 U11913 ( .A1(n9785), .A2(n11372), .ZN(n9406) );
  INV_X1 U11914 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10314) );
  OR2_X1 U11915 ( .A1(n6405), .A2(n10314), .ZN(n9405) );
  AND4_X2 U11916 ( .A1(n9408), .A2(n9407), .A3(n9406), .A4(n9405), .ZN(n11557)
         );
  NAND2_X1 U11917 ( .A1(n10064), .A2(n9845), .ZN(n9414) );
  NAND2_X1 U11918 ( .A1(n9411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9410) );
  MUX2_X1 U11919 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9410), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9412) );
  AND2_X1 U11920 ( .A1(n9412), .A2(n9521), .ZN(n14549) );
  AOI22_X1 U11921 ( .A1(n9844), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9574), .B2(
        n14549), .ZN(n9413) );
  NAND2_X1 U11922 ( .A1(n9414), .A2(n9413), .ZN(n15254) );
  NAND2_X1 U11923 ( .A1(n11557), .A2(n15254), .ZN(n11317) );
  INV_X1 U11924 ( .A(n11557), .ZN(n14494) );
  NAND2_X1 U11925 ( .A1(n14494), .A2(n11377), .ZN(n9415) );
  NAND2_X1 U11926 ( .A1(n11317), .A2(n9415), .ZN(n14440) );
  NAND2_X1 U11927 ( .A1(n11557), .A2(n11377), .ZN(n9417) );
  NAND2_X1 U11928 ( .A1(n11301), .A2(n9417), .ZN(n11324) );
  NAND2_X1 U11929 ( .A1(n10096), .A2(n9845), .ZN(n9420) );
  NAND2_X1 U11930 ( .A1(n9521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U11931 ( .A(n9418), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U11932 ( .A1(n9844), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9574), .B2(
        n10358), .ZN(n9419) );
  NAND2_X1 U11933 ( .A1(n9786), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9429) );
  INV_X1 U11934 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9421) );
  OR2_X1 U11935 ( .A1(n9535), .A2(n9421), .ZN(n9428) );
  NAND2_X1 U11936 ( .A1(n9423), .A2(n9422), .ZN(n9424) );
  NAND2_X1 U11937 ( .A1(n9448), .A2(n9424), .ZN(n11542) );
  OR2_X1 U11938 ( .A1(n9785), .A2(n11542), .ZN(n9427) );
  INV_X1 U11939 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9425) );
  OR2_X1 U11940 ( .A1(n6406), .A2(n9425), .ZN(n9426) );
  NAND2_X1 U11941 ( .A1(n11324), .A2(n9749), .ZN(n11323) );
  INV_X1 U11942 ( .A(n14493), .ZN(n11537) );
  NAND2_X1 U11943 ( .A1(n15260), .A2(n11537), .ZN(n9430) );
  NAND2_X1 U11944 ( .A1(n9440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9431) );
  XNOR2_X1 U11945 ( .A(n9431), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U11946 ( .A1(n9844), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9574), .B2(
        n10324), .ZN(n9432) );
  NAND2_X1 U11947 ( .A1(n9786), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9438) );
  INV_X1 U11948 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9433) );
  OR2_X1 U11949 ( .A1(n9535), .A2(n9433), .ZN(n9437) );
  INV_X1 U11950 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11849) );
  XNOR2_X1 U11951 ( .A(n9448), .B(n11849), .ZN(n14954) );
  OR2_X1 U11952 ( .A1(n9785), .A2(n14954), .ZN(n9436) );
  INV_X1 U11953 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9434) );
  OR2_X1 U11954 ( .A1(n6406), .A2(n9434), .ZN(n9435) );
  XNOR2_X1 U11955 ( .A(n14956), .B(n11826), .ZN(n14443) );
  OR2_X1 U11956 ( .A1(n14956), .A2(n14492), .ZN(n9439) );
  NAND2_X1 U11957 ( .A1(n10144), .A2(n9845), .ZN(n9445) );
  INV_X1 U11958 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U11959 ( .A1(n9442), .A2(n9441), .ZN(n9455) );
  NAND2_X1 U11960 ( .A1(n9455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9443) );
  XNOR2_X1 U11961 ( .A(n9443), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U11962 ( .A1(n9844), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9574), .B2(
        n14567), .ZN(n9444) );
  NAND2_X2 U11963 ( .A1(n9445), .A2(n9444), .ZN(n14295) );
  NAND2_X1 U11964 ( .A1(n9786), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9453) );
  INV_X1 U11965 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9446) );
  OR2_X1 U11966 ( .A1(n9535), .A2(n9446), .ZN(n9452) );
  INV_X1 U11967 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9447) );
  OAI21_X1 U11968 ( .B1(n9448), .B2(n11849), .A(n9447), .ZN(n9449) );
  NAND2_X1 U11969 ( .A1(n9449), .A2(n9463), .ZN(n11906) );
  OR2_X1 U11970 ( .A1(n9785), .A2(n11906), .ZN(n9451) );
  INV_X1 U11971 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10335) );
  OR2_X1 U11972 ( .A1(n6406), .A2(n10335), .ZN(n9450) );
  XNOR2_X1 U11973 ( .A(n14295), .B(n11866), .ZN(n14447) );
  OR2_X1 U11974 ( .A1(n14295), .A2(n14491), .ZN(n9454) );
  NAND2_X1 U11975 ( .A1(n10151), .A2(n9845), .ZN(n9460) );
  INV_X1 U11976 ( .A(n9455), .ZN(n9457) );
  INV_X1 U11977 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11978 ( .A1(n9457), .A2(n9456), .ZN(n9469) );
  NAND2_X1 U11979 ( .A1(n9469), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9458) );
  XNOR2_X1 U11980 ( .A(n9458), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U11981 ( .A1(n9574), .A2(n10343), .B1(n9844), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11982 ( .A1(n9786), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9468) );
  INV_X1 U11983 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9461) );
  OR2_X1 U11984 ( .A1(n9535), .A2(n9461), .ZN(n9467) );
  INV_X1 U11985 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U11986 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  NAND2_X1 U11987 ( .A1(n9483), .A2(n9464), .ZN(n12007) );
  OR2_X1 U11988 ( .A1(n9785), .A2(n12007), .ZN(n9466) );
  INV_X1 U11989 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10452) );
  OR2_X1 U11990 ( .A1(n6406), .A2(n10452), .ZN(n9465) );
  NAND4_X1 U11991 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n14490) );
  XNOR2_X1 U11992 ( .A(n15079), .B(n14490), .ZN(n11863) );
  INV_X1 U11993 ( .A(n11863), .ZN(n14448) );
  NAND2_X1 U11994 ( .A1(n10184), .A2(n9845), .ZN(n9472) );
  NAND2_X1 U11995 ( .A1(n9479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9470) );
  XNOR2_X1 U11996 ( .A(n9470), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U11997 ( .A1(n10460), .A2(n9574), .B1(n9844), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U11998 ( .A1(n9966), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9476) );
  INV_X1 U11999 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10453) );
  OR2_X1 U12000 ( .A1(n6405), .A2(n10453), .ZN(n9475) );
  XNOR2_X1 U12001 ( .A(n9483), .B(n10456), .ZN(n11959) );
  OR2_X1 U12002 ( .A1(n9785), .A2(n11959), .ZN(n9474) );
  INV_X1 U12003 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10772) );
  OR2_X1 U12004 ( .A1(n9376), .A2(n10772), .ZN(n9473) );
  NAND4_X1 U12005 ( .A1(n9476), .A2(n9475), .A3(n9474), .A4(n9473), .ZN(n14489) );
  NAND2_X1 U12006 ( .A1(n14303), .A2(n14489), .ZN(n9477) );
  NAND2_X1 U12007 ( .A1(n14938), .A2(n9477), .ZN(n9758) );
  INV_X1 U12008 ( .A(n9758), .ZN(n14449) );
  AND2_X1 U12009 ( .A1(n14448), .A2(n14449), .ZN(n9478) );
  OR2_X1 U12010 ( .A1(n15079), .A2(n14490), .ZN(n11954) );
  NAND2_X1 U12011 ( .A1(n10236), .A2(n9845), .ZN(n9481) );
  XNOR2_X1 U12012 ( .A(n9492), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U12013 ( .A1(n11238), .A2(n9574), .B1(n9844), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U12014 ( .A1(n9966), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9489) );
  INV_X1 U12015 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11233) );
  OR2_X1 U12016 ( .A1(n9376), .A2(n11233), .ZN(n9488) );
  OAI21_X1 U12017 ( .B1(n9483), .B2(n10456), .A(n9482), .ZN(n9484) );
  NAND2_X1 U12018 ( .A1(n9484), .A2(n9499), .ZN(n14949) );
  OR2_X1 U12019 ( .A1(n9539), .A2(n14949), .ZN(n9487) );
  INV_X1 U12020 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9485) );
  OR2_X1 U12021 ( .A1(n6406), .A2(n9485), .ZN(n9486) );
  NAND4_X1 U12022 ( .A1(n9489), .A2(n9488), .A3(n9487), .A4(n9486), .ZN(n14488) );
  XNOR2_X1 U12023 ( .A(n14951), .B(n14488), .ZN(n9759) );
  INV_X1 U12024 ( .A(n9759), .ZN(n14942) );
  OR2_X1 U12025 ( .A1(n14951), .A2(n14488), .ZN(n9490) );
  NAND2_X1 U12026 ( .A1(n10233), .A2(n9845), .ZN(n9495) );
  INV_X1 U12027 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U12028 ( .A1(n9492), .A2(n9491), .ZN(n9493) );
  NAND2_X1 U12029 ( .A1(n9493), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U12030 ( .A1(n14586), .A2(n9574), .B1(n9844), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U12031 ( .A1(n9786), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9505) );
  INV_X1 U12032 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9496) );
  OR2_X1 U12033 ( .A1(n9535), .A2(n9496), .ZN(n9504) );
  INV_X1 U12034 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U12035 ( .A1(n9499), .A2(n9498), .ZN(n9500) );
  NAND2_X1 U12036 ( .A1(n9513), .A2(n9500), .ZN(n14923) );
  OR2_X1 U12037 ( .A1(n9785), .A2(n14923), .ZN(n9503) );
  INV_X1 U12038 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9501) );
  OR2_X1 U12039 ( .A1(n6406), .A2(n9501), .ZN(n9502) );
  NAND4_X1 U12040 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n14487) );
  XNOR2_X1 U12041 ( .A(n15065), .B(n14487), .ZN(n14450) );
  OR2_X1 U12042 ( .A1(n15065), .A2(n14487), .ZN(n9506) );
  NAND2_X1 U12043 ( .A1(n10390), .A2(n9845), .ZN(n9512) );
  INV_X1 U12044 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U12045 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U12046 ( .A1(n9509), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9510) );
  AOI22_X1 U12047 ( .A1(n11617), .A2(n9574), .B1(n9844), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U12048 ( .A1(n9966), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9518) );
  INV_X1 U12049 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14904) );
  OR2_X1 U12050 ( .A1(n9376), .A2(n14904), .ZN(n9517) );
  NAND2_X1 U12051 ( .A1(n9513), .A2(n11242), .ZN(n9514) );
  NAND2_X1 U12052 ( .A1(n9526), .A2(n9514), .ZN(n14903) );
  OR2_X1 U12053 ( .A1(n9785), .A2(n14903), .ZN(n9516) );
  INV_X1 U12054 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11237) );
  OR2_X1 U12055 ( .A1(n6405), .A2(n11237), .ZN(n9515) );
  NAND4_X1 U12056 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n14879) );
  XNOR2_X1 U12057 ( .A(n14901), .B(n14879), .ZN(n14895) );
  NAND2_X1 U12058 ( .A1(n14901), .A2(n14879), .ZN(n9519) );
  NAND2_X1 U12059 ( .A1(n10492), .A2(n9845), .ZN(n9524) );
  OAI21_X1 U12060 ( .B1(n9521), .B2(n9520), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9522) );
  XNOR2_X1 U12061 ( .A(n9522), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U12062 ( .A1(n9844), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9574), 
        .B2(n11921), .ZN(n9523) );
  NAND2_X1 U12063 ( .A1(n9786), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9531) );
  INV_X1 U12064 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9525) );
  OR2_X1 U12065 ( .A1(n9535), .A2(n9525), .ZN(n9530) );
  NAND2_X1 U12066 ( .A1(n9526), .A2(n6904), .ZN(n9527) );
  NAND2_X1 U12067 ( .A1(n9537), .A2(n9527), .ZN(n14884) );
  OR2_X1 U12068 ( .A1(n9539), .A2(n14884), .ZN(n9529) );
  INV_X1 U12069 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11930) );
  OR2_X1 U12070 ( .A1(n6406), .A2(n11930), .ZN(n9528) );
  NAND2_X1 U12071 ( .A1(n10367), .A2(n9845), .ZN(n9534) );
  OR2_X1 U12072 ( .A1(n9546), .A2(n9336), .ZN(n9532) );
  XNOR2_X1 U12073 ( .A(n9532), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U12074 ( .A1(n9844), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9574), 
        .B2(n14593), .ZN(n9533) );
  NAND2_X1 U12075 ( .A1(n9786), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9543) );
  INV_X1 U12076 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15486) );
  OR2_X1 U12077 ( .A1(n9535), .A2(n15486), .ZN(n9542) );
  NAND2_X1 U12078 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  NAND2_X1 U12079 ( .A1(n9552), .A2(n9538), .ZN(n14865) );
  OR2_X1 U12080 ( .A1(n9539), .A2(n14865), .ZN(n9541) );
  INV_X1 U12081 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14600) );
  OR2_X1 U12082 ( .A1(n6406), .A2(n14600), .ZN(n9540) );
  XNOR2_X1 U12083 ( .A(n15046), .B(n14345), .ZN(n14856) );
  NAND2_X1 U12084 ( .A1(n14857), .A2(n14856), .ZN(n14854) );
  INV_X1 U12085 ( .A(n14345), .ZN(n14881) );
  OR2_X1 U12086 ( .A1(n15046), .A2(n14881), .ZN(n9544) );
  NAND2_X1 U12087 ( .A1(n10495), .A2(n9845), .ZN(n9549) );
  NAND2_X1 U12088 ( .A1(n9696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9547) );
  XNOR2_X1 U12089 ( .A(n9547), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14612) );
  AOI22_X1 U12090 ( .A1(n9844), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9574), 
        .B2(n14612), .ZN(n9548) );
  INV_X1 U12091 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U12092 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  NAND2_X1 U12093 ( .A1(n9564), .A2(n9553), .ZN(n14845) );
  OR2_X1 U12094 ( .A1(n14845), .A2(n9785), .ZN(n9557) );
  NAND2_X1 U12095 ( .A1(n9966), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12096 ( .A1(n9350), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9555) );
  INV_X1 U12097 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14609) );
  OR2_X1 U12098 ( .A1(n9376), .A2(n14609), .ZN(n9554) );
  NOR2_X1 U12099 ( .A1(n14844), .A2(n14486), .ZN(n9559) );
  NAND2_X1 U12100 ( .A1(n14844), .A2(n14486), .ZN(n9558) );
  NAND2_X1 U12101 ( .A1(n10975), .A2(n9845), .ZN(n9562) );
  NAND2_X1 U12102 ( .A1(n9571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9560) );
  XNOR2_X1 U12103 ( .A(n9560), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U12104 ( .A1(n9844), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9574), 
        .B2(n14628), .ZN(n9561) );
  INV_X1 U12105 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U12106 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  NAND2_X1 U12107 ( .A1(n9577), .A2(n9565), .ZN(n14833) );
  AOI22_X1 U12108 ( .A1(n9966), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n9786), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U12109 ( .A1(n9350), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9566) );
  OAI211_X1 U12110 ( .C1(n14833), .C2(n9785), .A(n9567), .B(n9566), .ZN(n14818) );
  OR2_X1 U12111 ( .A1(n15034), .A2(n14818), .ZN(n9568) );
  NAND2_X1 U12112 ( .A1(n15034), .A2(n14818), .ZN(n9569) );
  INV_X1 U12113 ( .A(n9691), .ZN(n9572) );
  NAND2_X1 U12114 ( .A1(n9572), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9573) );
  AOI22_X1 U12115 ( .A1(n9844), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14246), 
        .B2(n9574), .ZN(n9575) );
  INV_X1 U12116 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U12117 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  NAND2_X1 U12118 ( .A1(n9595), .A2(n9578), .ZN(n14129) );
  OR2_X1 U12119 ( .A1(n14129), .A2(n9785), .ZN(n9581) );
  AOI22_X1 U12120 ( .A1(n9966), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n9786), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9580) );
  INV_X1 U12121 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14625) );
  OR2_X1 U12122 ( .A1(n6406), .A2(n14625), .ZN(n9579) );
  OR2_X1 U12123 ( .A1(n15028), .A2(n14485), .ZN(n9582) );
  OR2_X1 U12124 ( .A1(n9384), .A2(n11132), .ZN(n9583) );
  XNOR2_X1 U12125 ( .A(n9595), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U12126 ( .A1(n14796), .A2(n9585), .ZN(n9591) );
  INV_X1 U12127 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U12128 ( .A1(n9786), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12129 ( .A1(n9966), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9586) );
  OAI211_X1 U12130 ( .C1(n9588), .C2(n6406), .A(n9587), .B(n9586), .ZN(n9589)
         );
  INV_X1 U12131 ( .A(n9589), .ZN(n9590) );
  XNOR2_X1 U12132 ( .A(n15022), .B(n14816), .ZN(n14804) );
  NAND2_X1 U12133 ( .A1(n15022), .A2(n14816), .ZN(n14371) );
  OR2_X1 U12134 ( .A1(n9384), .A2(n15495), .ZN(n9592) );
  INV_X1 U12135 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14182) );
  INV_X1 U12136 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9594) );
  OAI21_X1 U12137 ( .B1(n9595), .B2(n14182), .A(n9594), .ZN(n9596) );
  AND2_X1 U12138 ( .A1(n9596), .A2(n9607), .ZN(n14787) );
  NAND2_X1 U12139 ( .A1(n14787), .A2(n9585), .ZN(n9602) );
  INV_X1 U12140 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9599) );
  NAND2_X1 U12141 ( .A1(n9786), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9598) );
  NAND2_X1 U12142 ( .A1(n9966), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9597) );
  OAI211_X1 U12143 ( .C1(n9599), .C2(n6405), .A(n9598), .B(n9597), .ZN(n9600)
         );
  INV_X1 U12144 ( .A(n9600), .ZN(n9601) );
  OR2_X1 U12145 ( .A1(n15017), .A2(n14484), .ZN(n9603) );
  INV_X1 U12146 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15529) );
  NAND2_X1 U12147 ( .A1(n9607), .A2(n15529), .ZN(n9608) );
  NAND2_X1 U12148 ( .A1(n9642), .A2(n9608), .ZN(n14197) );
  INV_X1 U12149 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12150 ( .A1(n9966), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12151 ( .A1(n9786), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9609) );
  OAI211_X1 U12152 ( .C1(n9611), .C2(n6406), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U12153 ( .A(n9612), .ZN(n9613) );
  NAND2_X1 U12154 ( .A1(n9615), .A2(n14784), .ZN(n9616) );
  NAND2_X1 U12155 ( .A1(n11571), .A2(n9845), .ZN(n9618) );
  OR2_X1 U12156 ( .A1(n9384), .A2(n11576), .ZN(n9617) );
  INV_X1 U12157 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9641) );
  INV_X1 U12158 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9629) );
  INV_X1 U12159 ( .A(n9631), .ZN(n9619) );
  INV_X1 U12160 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U12161 ( .A1(n9631), .A2(n14153), .ZN(n9620) );
  NAND2_X1 U12162 ( .A1(n9656), .A2(n9620), .ZN(n14722) );
  INV_X1 U12163 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12164 ( .A1(n9786), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12165 ( .A1(n9966), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9621) );
  OAI211_X1 U12166 ( .C1(n9623), .C2(n6405), .A(n9622), .B(n9621), .ZN(n9624)
         );
  INV_X1 U12167 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U12168 ( .A1(n14995), .A2(n14481), .ZN(n9653) );
  OR2_X1 U12169 ( .A1(n11530), .A2(n9637), .ZN(n9628) );
  OR2_X1 U12170 ( .A1(n9384), .A2(n7526), .ZN(n9627) );
  NAND2_X1 U12171 ( .A1(n9644), .A2(n9629), .ZN(n9630) );
  NAND2_X1 U12172 ( .A1(n14743), .A2(n9585), .ZN(n9636) );
  INV_X1 U12173 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U12174 ( .A1(n9966), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U12175 ( .A1(n9786), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9632) );
  OAI211_X1 U12176 ( .C1(n6406), .C2(n15002), .A(n9633), .B(n9632), .ZN(n9634)
         );
  INV_X1 U12177 ( .A(n9634), .ZN(n9635) );
  NAND2_X1 U12178 ( .A1(n14739), .A2(n14712), .ZN(n9651) );
  INV_X1 U12179 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9638) );
  OR2_X1 U12180 ( .A1(n9384), .A2(n9638), .ZN(n9639) );
  NAND2_X1 U12181 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U12182 ( .A1(n9644), .A2(n9643), .ZN(n14757) );
  INV_X1 U12183 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9647) );
  NAND2_X1 U12184 ( .A1(n9786), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U12185 ( .A1(n9966), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9645) );
  OAI211_X1 U12186 ( .C1(n9647), .C2(n6405), .A(n9646), .B(n9645), .ZN(n9648)
         );
  INV_X1 U12187 ( .A(n9648), .ZN(n9649) );
  NAND2_X1 U12188 ( .A1(n15005), .A2(n14482), .ZN(n14733) );
  NAND2_X1 U12189 ( .A1(n14748), .A2(n9652), .ZN(n9667) );
  INV_X1 U12190 ( .A(n9652), .ZN(n14694) );
  NOR2_X1 U12191 ( .A1(n14739), .A2(n14712), .ZN(n14715) );
  AOI22_X1 U12192 ( .A1(n14715), .A2(n9653), .B1(n14225), .B2(n14726), .ZN(
        n14693) );
  NAND2_X1 U12193 ( .A1(n11783), .A2(n9845), .ZN(n9655) );
  OR2_X1 U12194 ( .A1(n9384), .A2(n15483), .ZN(n9654) );
  INV_X1 U12195 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14227) );
  NAND2_X1 U12196 ( .A1(n9656), .A2(n14227), .ZN(n9657) );
  NAND2_X1 U12197 ( .A1(n14698), .A2(n9585), .ZN(n9663) );
  INV_X1 U12198 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U12199 ( .A1(n9966), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U12200 ( .A1(n9786), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9658) );
  OAI211_X1 U12201 ( .C1(n6406), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9661)
         );
  INV_X1 U12202 ( .A(n9661), .ZN(n9662) );
  NAND2_X1 U12203 ( .A1(n14395), .A2(n14679), .ZN(n9776) );
  OR2_X1 U12204 ( .A1(n14395), .A2(n14679), .ZN(n9664) );
  OAI211_X1 U12205 ( .C1(n14750), .C2(n14694), .A(n14693), .B(n14702), .ZN(
        n9665) );
  INV_X1 U12206 ( .A(n9665), .ZN(n9666) );
  NAND2_X1 U12207 ( .A1(n9667), .A2(n9666), .ZN(n9669) );
  NAND2_X1 U12208 ( .A1(n14395), .A2(n14480), .ZN(n9668) );
  OR2_X1 U12209 ( .A1(n9384), .A2(n15108), .ZN(n9670) );
  INV_X1 U12210 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U12211 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  NAND2_X1 U12212 ( .A1(n14663), .A2(n9673), .ZN(n14684) );
  INV_X1 U12213 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U12214 ( .A1(n9786), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12215 ( .A1(n9966), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9674) );
  OAI211_X1 U12216 ( .C1(n15551), .C2(n6406), .A(n9675), .B(n9674), .ZN(n9676)
         );
  INV_X1 U12217 ( .A(n9676), .ZN(n9677) );
  INV_X1 U12218 ( .A(n14689), .ZN(n9679) );
  OR2_X1 U12219 ( .A1(n14983), .A2(n14479), .ZN(n9678) );
  NAND2_X1 U12220 ( .A1(n14094), .A2(n9845), .ZN(n9681) );
  OR2_X1 U12221 ( .A1(n9384), .A2(n12218), .ZN(n9680) );
  XNOR2_X1 U12222 ( .A(n14663), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12322) );
  NAND2_X1 U12223 ( .A1(n12322), .A2(n9585), .ZN(n9686) );
  INV_X1 U12224 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U12225 ( .A1(n9786), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U12226 ( .A1(n9966), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9682) );
  OAI211_X1 U12227 ( .C1(n15527), .C2(n6406), .A(n9683), .B(n9682), .ZN(n9684)
         );
  INV_X1 U12228 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U12229 ( .A1(n14408), .A2(n14478), .ZN(n14650) );
  NAND2_X1 U12230 ( .A1(n9688), .A2(n9779), .ZN(n9689) );
  NAND2_X1 U12231 ( .A1(n14651), .A2(n9689), .ZN(n9802) );
  NAND3_X1 U12232 ( .A1(n9694), .A2(n9693), .A3(n9692), .ZN(n9695) );
  NAND2_X1 U12233 ( .A1(n9698), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9699) );
  MUX2_X1 U12234 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9699), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9701) );
  INV_X1 U12235 ( .A(n11531), .ZN(n9716) );
  NAND2_X1 U12236 ( .A1(n9711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9712) );
  MUX2_X1 U12237 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9712), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9714) );
  NAND2_X1 U12238 ( .A1(n9717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9718) );
  MUX2_X1 U12239 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9718), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9720) );
  NAND2_X1 U12240 ( .A1(n9720), .A2(n9719), .ZN(n10757) );
  NAND2_X1 U12241 ( .A1(n11531), .A2(n11840), .ZN(n10148) );
  NAND2_X1 U12242 ( .A1(n10761), .A2(n10750), .ZN(n9735) );
  NAND2_X1 U12243 ( .A1(n11840), .A2(n11574), .ZN(n10116) );
  OAI21_X1 U12244 ( .B1(n10115), .B2(P1_D_REG_1__SCAN_IN), .A(n10116), .ZN(
        n9812) );
  INV_X1 U12245 ( .A(n9812), .ZN(n9734) );
  INV_X1 U12246 ( .A(n10115), .ZN(n9733) );
  NOR4_X1 U12247 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n9731) );
  NOR4_X1 U12248 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9730) );
  OR4_X1 U12249 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9728) );
  NOR4_X1 U12250 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9726) );
  NOR4_X1 U12251 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9725) );
  NOR4_X1 U12252 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9724) );
  NOR4_X1 U12253 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9723) );
  NAND4_X1 U12254 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n9727)
         );
  NOR4_X1 U12255 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9728), .A4(n9727), .ZN(n9729) );
  NAND3_X1 U12256 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(n9732) );
  NAND2_X1 U12257 ( .A1(n9733), .A2(n9732), .ZN(n9813) );
  NAND2_X1 U12258 ( .A1(n9734), .A2(n9813), .ZN(n10751) );
  INV_X1 U12259 ( .A(n10752), .ZN(n10141) );
  NAND2_X1 U12260 ( .A1(n15216), .A2(n14246), .ZN(n10755) );
  NAND2_X1 U12261 ( .A1(n14917), .A2(n14245), .ZN(n9736) );
  NAND2_X1 U12262 ( .A1(n14248), .A2(n9736), .ZN(n11355) );
  NAND2_X1 U12263 ( .A1(n14498), .A2(n14260), .ZN(n9738) );
  NAND2_X1 U12264 ( .A1(n9738), .A2(n14255), .ZN(n9740) );
  NAND2_X1 U12265 ( .A1(n14258), .A2(n14970), .ZN(n9739) );
  NAND2_X1 U12266 ( .A1(n9740), .A2(n9739), .ZN(n11048) );
  NAND2_X1 U12267 ( .A1(n9741), .A2(n7193), .ZN(n9742) );
  NAND2_X1 U12268 ( .A1(n9743), .A2(n9742), .ZN(n11117) );
  NAND2_X1 U12269 ( .A1(n11117), .A2(n14439), .ZN(n9744) );
  NAND2_X1 U12270 ( .A1(n9744), .A2(n14277), .ZN(n15207) );
  NAND2_X1 U12271 ( .A1(n15207), .A2(n15206), .ZN(n9746) );
  NAND2_X1 U12272 ( .A1(n11348), .A2(n15222), .ZN(n9745) );
  NAND2_X1 U12273 ( .A1(n9746), .A2(n9745), .ZN(n11199) );
  NOR2_X1 U12274 ( .A1(n14495), .A2(n11357), .ZN(n9748) );
  NAND2_X1 U12275 ( .A1(n14495), .A2(n11357), .ZN(n9747) );
  INV_X1 U12276 ( .A(n11296), .ZN(n9752) );
  NAND2_X1 U12277 ( .A1(n11537), .A2(n14289), .ZN(n9753) );
  OR2_X1 U12278 ( .A1(n14956), .A2(n11826), .ZN(n9755) );
  NAND2_X1 U12279 ( .A1(n11708), .A2(n9755), .ZN(n11824) );
  NAND2_X1 U12280 ( .A1(n14295), .A2(n11866), .ZN(n9756) );
  OR2_X1 U12281 ( .A1(n15079), .A2(n14306), .ZN(n9757) );
  INV_X1 U12282 ( .A(n14489), .ZN(n14936) );
  INV_X1 U12283 ( .A(n14488), .ZN(n14301) );
  OR2_X1 U12284 ( .A1(n14951), .A2(n14301), .ZN(n9760) );
  NAND2_X1 U12285 ( .A1(n14913), .A2(n14450), .ZN(n9762) );
  INV_X1 U12286 ( .A(n14487), .ZN(n14934) );
  OR2_X1 U12287 ( .A1(n15065), .A2(n14934), .ZN(n9761) );
  NAND2_X1 U12288 ( .A1(n9762), .A2(n9761), .ZN(n14894) );
  NAND2_X1 U12289 ( .A1(n14894), .A2(n14895), .ZN(n9763) );
  INV_X1 U12290 ( .A(n14879), .ZN(n14333) );
  OR2_X1 U12291 ( .A1(n14901), .A2(n14333), .ZN(n14341) );
  NAND2_X1 U12292 ( .A1(n15046), .A2(n14345), .ZN(n9765) );
  OR2_X1 U12293 ( .A1(n14844), .A2(n14861), .ZN(n9768) );
  NAND2_X1 U12294 ( .A1(n14844), .A2(n14861), .ZN(n9766) );
  NAND2_X1 U12295 ( .A1(n9768), .A2(n9766), .ZN(n14843) );
  INV_X1 U12296 ( .A(n14843), .ZN(n9767) );
  XNOR2_X1 U12297 ( .A(n15034), .B(n14818), .ZN(n14824) );
  INV_X1 U12298 ( .A(n14818), .ZN(n14131) );
  OR2_X1 U12299 ( .A1(n15034), .A2(n14131), .ZN(n9769) );
  INV_X1 U12300 ( .A(n14816), .ZN(n14783) );
  AND2_X1 U12301 ( .A1(n14804), .A2(n14800), .ZN(n14801) );
  INV_X1 U12302 ( .A(n14484), .ZN(n12257) );
  NOR2_X1 U12303 ( .A1(n9615), .A2(n14483), .ZN(n9771) );
  NAND2_X1 U12304 ( .A1(n15005), .A2(n14171), .ZN(n14711) );
  OAI21_X1 U12305 ( .B1(n15005), .B2(n14171), .A(n14387), .ZN(n9774) );
  NOR3_X1 U12306 ( .A1(n15005), .A2(n14171), .A3(n14387), .ZN(n9773) );
  XNOR2_X1 U12307 ( .A(n14995), .B(n14225), .ZN(n14716) );
  AOI211_X1 U12308 ( .C1(n15000), .C2(n9774), .A(n9773), .B(n14716), .ZN(n9775) );
  INV_X1 U12309 ( .A(n9776), .ZN(n9777) );
  INV_X1 U12310 ( .A(n9780), .ZN(n9778) );
  NAND2_X1 U12311 ( .A1(n7664), .A2(n9780), .ZN(n9781) );
  NAND2_X1 U12312 ( .A1(n14251), .A2(n14416), .ZN(n9783) );
  NAND2_X1 U12313 ( .A1(n14246), .A2(n14245), .ZN(n9782) );
  INV_X1 U12314 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14662) );
  INV_X1 U12315 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U12316 ( .A1(n9966), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12317 ( .A1(n9786), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9787) );
  OAI211_X1 U12318 ( .C1(n9789), .C2(n6405), .A(n9788), .B(n9787), .ZN(n9790)
         );
  INV_X1 U12319 ( .A(n9790), .ZN(n9791) );
  INV_X1 U12320 ( .A(n9784), .ZN(n14511) );
  OAI22_X1 U12321 ( .A1(n14226), .A2(n14935), .B1(n14420), .B2(n14933), .ZN(
        n9793) );
  NAND2_X1 U12322 ( .A1(n11044), .A2(n11342), .ZN(n15214) );
  NOR2_X4 U12323 ( .A1(n11829), .A2(n14295), .ZN(n11857) );
  NOR2_X4 U12324 ( .A1(n14912), .A2(n14901), .ZN(n14900) );
  INV_X1 U12325 ( .A(n15053), .ZN(n14888) );
  INV_X1 U12326 ( .A(n15034), .ZN(n14829) );
  NAND2_X1 U12327 ( .A1(n14828), .A2(n14829), .ZN(n14831) );
  NOR2_X2 U12328 ( .A1(n14831), .A2(n15028), .ZN(n9795) );
  INV_X1 U12329 ( .A(n9795), .ZN(n14811) );
  NOR2_X4 U12330 ( .A1(n14811), .A2(n15022), .ZN(n14785) );
  AND2_X2 U12331 ( .A1(n14719), .A2(n14726), .ZN(n14720) );
  AOI211_X1 U12332 ( .C1(n14408), .C2(n6480), .A(n14929), .B(n9974), .ZN(n9806) );
  NOR2_X2 U12333 ( .A1(n14658), .A2(n14246), .ZN(n14907) );
  INV_X1 U12334 ( .A(n14408), .ZN(n14254) );
  NAND2_X1 U12335 ( .A1(n14251), .A2(n14247), .ZN(n14468) );
  OR2_X1 U12336 ( .A1(n14468), .A2(n14245), .ZN(n9796) );
  NOR2_X2 U12337 ( .A1(n6412), .A2(n9796), .ZN(n15223) );
  AOI22_X1 U12338 ( .A1(n12322), .A2(n14974), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n6412), .ZN(n9797) );
  OAI21_X1 U12339 ( .B1(n14254), .B2(n14921), .A(n9797), .ZN(n9798) );
  INV_X1 U12340 ( .A(n9800), .ZN(n9801) );
  NAND2_X1 U12341 ( .A1(n7846), .A2(n9801), .ZN(P1_U3265) );
  AND2_X1 U12342 ( .A1(n9803), .A2(n14247), .ZN(n10786) );
  INV_X1 U12343 ( .A(n9804), .ZN(n9805) );
  AOI21_X1 U12344 ( .B1(n15255), .B2(n14408), .A(n9806), .ZN(n9807) );
  INV_X1 U12345 ( .A(n9807), .ZN(n9808) );
  NOR2_X1 U12346 ( .A1(n9809), .A2(n9808), .ZN(n9810) );
  NAND2_X1 U12347 ( .A1(n9811), .A2(n9810), .ZN(n9862) );
  NAND3_X1 U12348 ( .A1(n10755), .A2(n9813), .A3(n9812), .ZN(n9814) );
  NAND2_X1 U12349 ( .A1(n9862), .A2(n15272), .ZN(n9816) );
  OR2_X1 U12350 ( .A1(n15272), .A2(n15527), .ZN(n9815) );
  NAND2_X1 U12351 ( .A1(n9816), .A2(n9815), .ZN(P1_U3556) );
  INV_X1 U12352 ( .A(n9817), .ZN(n9820) );
  NAND2_X1 U12353 ( .A1(n9818), .A2(SI_27_), .ZN(n9819) );
  NAND2_X1 U12354 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  NOR2_X1 U12355 ( .A1(n9824), .A2(SI_28_), .ZN(n9825) );
  INV_X1 U12356 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14090) );
  MUX2_X1 U12357 ( .A(n12072), .B(n14090), .S(n10093), .Z(n9831) );
  XNOR2_X1 U12358 ( .A(n9831), .B(SI_29_), .ZN(n9829) );
  NAND2_X1 U12359 ( .A1(n13342), .A2(n9845), .ZN(n9828) );
  OR2_X1 U12360 ( .A1(n9384), .A2(n12072), .ZN(n9827) );
  NAND2_X1 U12361 ( .A1(n9831), .A2(n13025), .ZN(n9832) );
  MUX2_X1 U12362 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6409), .Z(n9837) );
  XNOR2_X1 U12363 ( .A(n9837), .B(SI_30_), .ZN(n9839) );
  INV_X1 U12364 ( .A(n9839), .ZN(n9834) );
  NAND2_X1 U12365 ( .A1(n13367), .A2(n9845), .ZN(n9836) );
  OR2_X1 U12366 ( .A1(n9384), .A2(n15104), .ZN(n9835) );
  NAND2_X1 U12367 ( .A1(n9837), .A2(SI_30_), .ZN(n9838) );
  MUX2_X1 U12368 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6410), .Z(n9841) );
  XNOR2_X1 U12369 ( .A(n9841), .B(SI_31_), .ZN(n9842) );
  NAND2_X1 U12370 ( .A1(n14640), .A2(n15216), .ZN(n9856) );
  INV_X1 U12371 ( .A(P1_B_REG_SCAN_IN), .ZN(n9848) );
  NOR2_X1 U12372 ( .A1(n15106), .A2(n9848), .ZN(n9849) );
  NOR2_X1 U12373 ( .A1(n14933), .A2(n9849), .ZN(n9971) );
  INV_X1 U12374 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U12375 ( .A1(n9966), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9852) );
  INV_X1 U12376 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9850) );
  OR2_X1 U12377 ( .A1(n9376), .A2(n9850), .ZN(n9851) );
  OAI211_X1 U12378 ( .C1(n6405), .C2(n9853), .A(n9852), .B(n9851), .ZN(n14475)
         );
  NAND2_X1 U12379 ( .A1(n9971), .A2(n14475), .ZN(n14979) );
  INV_X1 U12380 ( .A(n9854), .ZN(n9855) );
  NAND2_X1 U12381 ( .A1(n9856), .A2(n9855), .ZN(n14978) );
  INV_X1 U12382 ( .A(n10750), .ZN(n9857) );
  INV_X1 U12383 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U12384 ( .A1(n15265), .A2(n9859), .ZN(n9860) );
  AOI21_X1 U12385 ( .B1(n14978), .B2(n15265), .A(n9860), .ZN(n9861) );
  INV_X1 U12386 ( .A(n9861), .ZN(P1_U3527) );
  NAND2_X1 U12387 ( .A1(n9862), .A2(n15265), .ZN(n9865) );
  OR2_X1 U12388 ( .A1(n15265), .A2(n9863), .ZN(n9864) );
  NAND2_X1 U12389 ( .A1(n9865), .A2(n9864), .ZN(P1_U3524) );
  NAND2_X1 U12390 ( .A1(n12523), .A2(n10699), .ZN(n11006) );
  NAND2_X1 U12391 ( .A1(n11007), .A2(n11006), .ZN(n9866) );
  NAND2_X1 U12392 ( .A1(n12878), .A2(n10998), .ZN(n10984) );
  NAND2_X1 U12393 ( .A1(n10949), .A2(n12888), .ZN(n10933) );
  NAND2_X1 U12394 ( .A1(n10936), .A2(n10933), .ZN(n10934) );
  NAND2_X1 U12395 ( .A1(n10934), .A2(n10984), .ZN(n9867) );
  NAND3_X1 U12396 ( .A1(n9868), .A2(n10987), .A3(n9867), .ZN(n9870) );
  NAND2_X1 U12397 ( .A1(n12521), .A2(n15403), .ZN(n9869) );
  NAND2_X1 U12398 ( .A1(n9870), .A2(n9869), .ZN(n11093) );
  NAND2_X1 U12399 ( .A1(n12519), .A2(n15413), .ZN(n11452) );
  NAND2_X1 U12400 ( .A1(n9871), .A2(n11452), .ZN(n9874) );
  NAND2_X1 U12401 ( .A1(n11289), .A2(n9872), .ZN(n11218) );
  NAND2_X1 U12402 ( .A1(n11217), .A2(n11218), .ZN(n11220) );
  NAND2_X1 U12403 ( .A1(n11220), .A2(n11452), .ZN(n9873) );
  OAI211_X1 U12404 ( .C1(n11093), .C2(n9874), .A(n11454), .B(n9873), .ZN(n9876) );
  NAND2_X1 U12405 ( .A1(n12518), .A2(n11469), .ZN(n9875) );
  NAND2_X1 U12406 ( .A1(n9876), .A2(n9875), .ZN(n11442) );
  OR2_X1 U12407 ( .A1(n11882), .A2(n12021), .ZN(n9879) );
  INV_X1 U12408 ( .A(n12162), .ZN(n12466) );
  NAND2_X1 U12409 ( .A1(n12469), .A2(n12515), .ZN(n9880) );
  OR2_X1 U12410 ( .A1(n12469), .A2(n12515), .ZN(n9881) );
  INV_X1 U12411 ( .A(n11912), .ZN(n9883) );
  INV_X1 U12412 ( .A(n11913), .ZN(n9882) );
  OR2_X1 U12413 ( .A1(n12387), .A2(n12450), .ZN(n9884) );
  NAND2_X1 U12414 ( .A1(n12868), .A2(n12344), .ZN(n9886) );
  NAND2_X1 U12415 ( .A1(n12942), .A2(n12859), .ZN(n9887) );
  NAND2_X1 U12416 ( .A1(n12050), .A2(n9887), .ZN(n12858) );
  NAND2_X1 U12417 ( .A1(n13006), .A2(n12847), .ZN(n9888) );
  OR2_X1 U12418 ( .A1(n13000), .A2(n12860), .ZN(n9889) );
  INV_X1 U12419 ( .A(n12846), .ZN(n12478) );
  NAND2_X1 U12420 ( .A1(n12796), .A2(n9892), .ZN(n9894) );
  NAND2_X1 U12421 ( .A1(n12986), .A2(n12805), .ZN(n9893) );
  NAND2_X1 U12422 ( .A1(n9894), .A2(n9893), .ZN(n12786) );
  AND2_X1 U12423 ( .A1(n12980), .A2(n12798), .ZN(n9896) );
  OAI21_X2 U12424 ( .B1(n12786), .B2(n9896), .A(n9895), .ZN(n12776) );
  NOR2_X1 U12425 ( .A1(n12974), .A2(n12788), .ZN(n9898) );
  NAND2_X1 U12426 ( .A1(n12974), .A2(n12788), .ZN(n9897) );
  AND2_X1 U12427 ( .A1(n12909), .A2(n12767), .ZN(n9900) );
  NAND2_X1 U12428 ( .A1(n12961), .A2(n12752), .ZN(n9901) );
  NAND2_X1 U12429 ( .A1(n12741), .A2(n9901), .ZN(n12733) );
  OR2_X1 U12430 ( .A1(n12954), .A2(n12744), .ZN(n9902) );
  INV_X1 U12431 ( .A(n12954), .ZN(n9903) );
  INV_X1 U12432 ( .A(n12489), .ZN(n12735) );
  OR2_X1 U12433 ( .A1(n9906), .A2(n12735), .ZN(n9910) );
  NAND2_X1 U12434 ( .A1(n12719), .A2(n9910), .ZN(n9908) );
  NAND2_X1 U12435 ( .A1(n9908), .A2(n9907), .ZN(n9912) );
  NAND2_X1 U12436 ( .A1(n9951), .A2(n11314), .ZN(n9956) );
  AND2_X1 U12437 ( .A1(n12207), .A2(n9910), .ZN(n9911) );
  NAND3_X1 U12438 ( .A1(n9912), .A2(n12883), .A3(n12139), .ZN(n9914) );
  OR2_X1 U12439 ( .A1(n13027), .A2(n13031), .ZN(n10435) );
  NAND2_X1 U12440 ( .A1(n10435), .A2(n10431), .ZN(n10576) );
  INV_X1 U12441 ( .A(n10576), .ZN(n10806) );
  AOI22_X1 U12442 ( .A1(n12735), .A2(n12880), .B1(n12510), .B2(n12879), .ZN(
        n9913) );
  NAND2_X1 U12443 ( .A1(n9914), .A2(n9913), .ZN(n12712) );
  XNOR2_X1 U12444 ( .A(n9915), .B(P3_B_REG_SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12445 ( .A1(n9916), .A2(n12071), .ZN(n9918) );
  NAND2_X1 U12446 ( .A1(n9915), .A2(n13040), .ZN(n9919) );
  INV_X1 U12447 ( .A(n10796), .ZN(n13014) );
  NAND2_X1 U12448 ( .A1(n12071), .A2(n13040), .ZN(n9921) );
  XNOR2_X1 U12449 ( .A(n13014), .B(n10690), .ZN(n9934) );
  NOR2_X1 U12450 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .ZN(
        n9925) );
  NOR4_X1 U12451 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9924) );
  NOR4_X1 U12452 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9923) );
  NOR4_X1 U12453 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9922) );
  NAND4_X1 U12454 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(n9932)
         );
  NOR4_X1 U12455 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9929) );
  NOR4_X1 U12456 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9928) );
  NOR4_X1 U12457 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9927) );
  NOR4_X1 U12458 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9926) );
  NAND4_X1 U12459 ( .A1(n9929), .A2(n9928), .A3(n9927), .A4(n9926), .ZN(n9931)
         );
  INV_X1 U12460 ( .A(n9920), .ZN(n9930) );
  OAI21_X1 U12461 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9959) );
  AND2_X1 U12462 ( .A1(n10574), .A2(n9959), .ZN(n9933) );
  NAND2_X1 U12463 ( .A1(n9944), .A2(n10430), .ZN(n10559) );
  AND2_X1 U12464 ( .A1(n11314), .A2(n9938), .ZN(n9935) );
  NAND2_X1 U12465 ( .A1(n6417), .A2(n9935), .ZN(n9949) );
  NAND2_X1 U12466 ( .A1(n9949), .A2(n9936), .ZN(n10689) );
  AND2_X1 U12467 ( .A1(n10559), .A2(n10689), .ZN(n10691) );
  NAND2_X1 U12468 ( .A1(n6417), .A2(n11314), .ZN(n9937) );
  OAI21_X1 U12469 ( .B1(n9938), .B2(n15418), .A(n9937), .ZN(n9939) );
  AOI21_X1 U12470 ( .B1(n9939), .B2(n9944), .A(n10430), .ZN(n9940) );
  MUX2_X1 U12471 ( .A(n10691), .B(n9940), .S(n10690), .Z(n9941) );
  MUX2_X1 U12472 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12712), .S(n15589), .Z(
        n9942) );
  INV_X1 U12473 ( .A(n9942), .ZN(n9955) );
  XNOR2_X1 U12474 ( .A(n9943), .B(n12207), .ZN(n12718) );
  INV_X1 U12475 ( .A(n9944), .ZN(n9948) );
  NAND2_X1 U12476 ( .A1(n6417), .A2(n11179), .ZN(n9947) );
  NAND2_X1 U12477 ( .A1(n11179), .A2(n11134), .ZN(n9945) );
  XNOR2_X1 U12478 ( .A(n11314), .B(n9945), .ZN(n9946) );
  NAND2_X1 U12479 ( .A1(n9947), .A2(n9946), .ZN(n10565) );
  NAND3_X1 U12480 ( .A1(n9948), .A2(n15418), .A3(n10565), .ZN(n9950) );
  INV_X1 U12481 ( .A(n12715), .ZN(n12138) );
  OAI22_X1 U12482 ( .A1(n12718), .A2(n12941), .B1(n12138), .B2(n12905), .ZN(
        n9953) );
  INV_X1 U12483 ( .A(n9953), .ZN(n9954) );
  NAND2_X1 U12484 ( .A1(n9955), .A2(n9954), .ZN(P3_U3487) );
  INV_X1 U12485 ( .A(n10690), .ZN(n13012) );
  NAND3_X1 U12486 ( .A1(n13012), .A2(n13014), .A3(n9959), .ZN(n10569) );
  INV_X1 U12487 ( .A(n10569), .ZN(n10573) );
  OR2_X1 U12488 ( .A1(n9956), .A2(n10795), .ZN(n10566) );
  NOR2_X1 U12489 ( .A1(n10566), .A2(n10571), .ZN(n9957) );
  OR2_X1 U12490 ( .A1(n10807), .A2(n9957), .ZN(n9958) );
  NAND2_X1 U12491 ( .A1(n10573), .A2(n9958), .ZN(n9961) );
  NAND3_X1 U12492 ( .A1(n10808), .A2(n10574), .A3(n10565), .ZN(n9960) );
  MUX2_X1 U12493 ( .A(n12712), .B(P3_REG0_REG_28__SCAN_IN), .S(n15429), .Z(
        n9962) );
  INV_X1 U12494 ( .A(n9962), .ZN(n9965) );
  INV_X1 U12495 ( .A(n15395), .ZN(n12945) );
  OAI22_X1 U12496 ( .A1(n12718), .A2(n13010), .B1(n12138), .B2(n12949), .ZN(
        n9963) );
  INV_X1 U12497 ( .A(n9963), .ZN(n9964) );
  NAND2_X1 U12498 ( .A1(n9965), .A2(n9964), .ZN(P3_U3455) );
  INV_X1 U12499 ( .A(n14478), .ZN(n14680) );
  NAND2_X1 U12500 ( .A1(n14408), .A2(n14680), .ZN(n14654) );
  NOR2_X1 U12501 ( .A1(n14654), .A2(n15050), .ZN(n9979) );
  NAND4_X1 U12502 ( .A1(n14656), .A2(n15263), .A3(n14478), .A4(n14408), .ZN(
        n9973) );
  NAND2_X1 U12503 ( .A1(n14668), .A2(n15255), .ZN(n9972) );
  INV_X1 U12504 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9969) );
  INV_X1 U12505 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14645) );
  OR2_X1 U12506 ( .A1(n9376), .A2(n14645), .ZN(n9968) );
  NAND2_X1 U12507 ( .A1(n9966), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9967) );
  OAI211_X1 U12508 ( .C1(n6405), .C2(n9969), .A(n9968), .B(n9967), .ZN(n14476)
         );
  NAND2_X1 U12509 ( .A1(n9971), .A2(n14476), .ZN(n14659) );
  NAND2_X1 U12510 ( .A1(n14478), .A2(n14880), .ZN(n14666) );
  NAND4_X1 U12511 ( .A1(n9973), .A2(n9972), .A3(n14659), .A4(n14666), .ZN(
        n9978) );
  OR2_X1 U12512 ( .A1(n9974), .A2(n14421), .ZN(n9975) );
  NOR2_X1 U12513 ( .A1(n14670), .A2(n14929), .ZN(n9977) );
  AOI211_X1 U12514 ( .C1(n9979), .C2(n14656), .A(n9978), .B(n9977), .ZN(n9980)
         );
  INV_X1 U12515 ( .A(n9980), .ZN(n9982) );
  NAND2_X1 U12516 ( .A1(n14656), .A2(n15251), .ZN(n9984) );
  OAI21_X1 U12517 ( .B1(n14655), .B2(n9984), .A(n9983), .ZN(n9985) );
  INV_X1 U12518 ( .A(n9985), .ZN(n9989) );
  NAND2_X1 U12519 ( .A1(n9992), .A2(n9991), .ZN(P1_U3557) );
  NAND2_X1 U12520 ( .A1(n15264), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U12521 ( .A1(n9994), .A2(n9993), .ZN(P1_U3525) );
  INV_X1 U12522 ( .A(n9995), .ZN(n9996) );
  NAND2_X1 U12523 ( .A1(n9996), .A2(n11331), .ZN(n10197) );
  INV_X1 U12524 ( .A(n10557), .ZN(n9997) );
  INV_X1 U12525 ( .A(n9999), .ZN(n9998) );
  NAND2_X1 U12526 ( .A1(n13452), .A2(n13200), .ZN(n10000) );
  NAND2_X1 U12527 ( .A1(n9998), .A2(n10000), .ZN(n10474) );
  INV_X1 U12528 ( .A(n10000), .ZN(n10001) );
  NAND2_X1 U12529 ( .A1(n9999), .A2(n10001), .ZN(n10002) );
  AND2_X1 U12530 ( .A1(n10474), .A2(n10002), .ZN(n10379) );
  INV_X1 U12531 ( .A(n10379), .ZN(n10003) );
  INV_X1 U12532 ( .A(n10909), .ZN(n13802) );
  NAND2_X1 U12533 ( .A1(n10003), .A2(n13802), .ZN(n10009) );
  AOI22_X1 U12534 ( .A1(n13885), .A2(n13449), .B1(n13452), .B2(n13883), .ZN(
        n10008) );
  INV_X1 U12535 ( .A(n10908), .ZN(n10004) );
  OAI21_X1 U12536 ( .B1(n10004), .B2(n9999), .A(n10481), .ZN(n10006) );
  NAND2_X1 U12537 ( .A1(n13541), .A2(n6414), .ZN(n10005) );
  INV_X1 U12538 ( .A(n13195), .ZN(n13394) );
  NAND2_X1 U12539 ( .A1(n13394), .A2(n13421), .ZN(n13429) );
  NAND2_X1 U12540 ( .A1(n10006), .A2(n13905), .ZN(n10007) );
  NAND3_X1 U12541 ( .A1(n10009), .A2(n10008), .A3(n10007), .ZN(n10374) );
  NAND3_X1 U12542 ( .A1(n15359), .A2(n10011), .A3(n10010), .ZN(n10373) );
  INV_X1 U12543 ( .A(n10373), .ZN(n10013) );
  NOR2_X1 U12544 ( .A1(n10382), .A2(n15358), .ZN(n10012) );
  NAND2_X1 U12545 ( .A1(n10013), .A2(n10012), .ZN(n10014) );
  MUX2_X1 U12546 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10374), .S(n13880), .Z(
        n10020) );
  INV_X1 U12547 ( .A(n10017), .ZN(n10470) );
  OAI22_X1 U12548 ( .A1(n13931), .A2(n10470), .B1(n8719), .B2(n13837), .ZN(
        n10019) );
  NOR2_X1 U12549 ( .A1(n13374), .A2(n11129), .ZN(n10016) );
  NAND2_X1 U12550 ( .A1(n13880), .A2(n10016), .ZN(n13811) );
  NAND2_X1 U12551 ( .A1(n13880), .A2(n13428), .ZN(n13554) );
  OAI211_X1 U12552 ( .C1(n10470), .C2(n10906), .A(n13889), .B(n11265), .ZN(
        n10375) );
  OAI22_X1 U12553 ( .A1(n10379), .A2(n13811), .B1(n13554), .B2(n10375), .ZN(
        n10018) );
  OR3_X1 U12554 ( .A1(n10020), .A2(n10019), .A3(n10018), .ZN(P2_U3264) );
  INV_X1 U12555 ( .A(n10679), .ZN(n10022) );
  AOI211_X1 U12556 ( .C1(n10021), .C2(n10023), .A(n13165), .B(n10022), .ZN(
        n10027) );
  MUX2_X1 U12557 ( .A(P2_U3088), .B(n13170), .S(n10024), .Z(n10026) );
  AOI22_X1 U12558 ( .A1(n13885), .A2(n13447), .B1(n13449), .B2(n13883), .ZN(
        n10484) );
  INV_X1 U12559 ( .A(n13161), .ZN(n13120) );
  OAI22_X1 U12560 ( .A1(n10484), .A2(n13120), .B1(n13194), .B2(n11426), .ZN(
        n10025) );
  OR3_X1 U12561 ( .A1(n10027), .A2(n10026), .A3(n10025), .ZN(P2_U3190) );
  INV_X1 U12562 ( .A(n10042), .ZN(n10029) );
  INV_X1 U12563 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10502) );
  NAND2_X1 U12564 ( .A1(n10502), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10028) );
  NAND2_X1 U12565 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  INV_X1 U12566 ( .A(n10030), .ZN(n10032) );
  INV_X1 U12567 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10031) );
  AND2_X1 U12568 ( .A1(n10030), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10034) );
  AOI21_X1 U12569 ( .B1(n10032), .B2(n10031), .A(n10034), .ZN(SUB_1596_U53) );
  INV_X1 U12570 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U12571 ( .A1(n10035), .A2(n10034), .ZN(n10039) );
  OAI21_X1 U12572 ( .B1(n10035), .B2(n10034), .A(n10039), .ZN(n10036) );
  INV_X1 U12573 ( .A(n10036), .ZN(SUB_1596_U5) );
  NAND2_X1 U12574 ( .A1(n10037), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10038) );
  INV_X1 U12575 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12576 ( .A1(n10040), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n10041) );
  INV_X1 U12577 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U12578 ( .A1(n10043), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10044) );
  XNOR2_X1 U12579 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n10054) );
  INV_X1 U12580 ( .A(n10054), .ZN(n10046) );
  XNOR2_X1 U12581 ( .A(n10055), .B(n10046), .ZN(n10049) );
  OAI21_X1 U12582 ( .B1(n10047), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n10053), .ZN(
        n10048) );
  INV_X1 U12583 ( .A(n10048), .ZN(SUB_1596_U61) );
  INV_X1 U12584 ( .A(n10049), .ZN(n10050) );
  NAND2_X1 U12585 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  NAND2_X1 U12586 ( .A1(n10056), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10057) );
  XNOR2_X1 U12587 ( .A(n10067), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10074) );
  INV_X1 U12588 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10072) );
  XNOR2_X1 U12589 ( .A(n10073), .B(n10072), .ZN(SUB_1596_U60) );
  NAND2_X2 U12590 ( .A1(n7400), .A2(P1_U3086), .ZN(n15105) );
  NOR2_X1 U12591 ( .A1(n6410), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12220) );
  INV_X2 U12592 ( .A(n12220), .ZN(n10976) );
  OAI222_X1 U12593 ( .A1(n15105), .A2(n10059), .B1(n10976), .B2(n10088), .C1(
        P1_U3086), .C2(n14522), .ZN(P1_U3353) );
  OAI222_X1 U12594 ( .A1(n15105), .A2(n10060), .B1(n10976), .B2(n10086), .C1(
        P1_U3086), .C2(n15195), .ZN(P1_U3351) );
  OAI222_X1 U12595 ( .A1(n15105), .A2(n10061), .B1(n10976), .B2(n10084), .C1(
        P1_U3086), .C2(n14538), .ZN(P1_U3352) );
  INV_X1 U12596 ( .A(n10062), .ZN(n10082) );
  OAI222_X1 U12597 ( .A1(n15105), .A2(n10063), .B1(n10976), .B2(n10082), .C1(
        P1_U3086), .C2(n10313), .ZN(P1_U3350) );
  INV_X1 U12598 ( .A(n10064), .ZN(n10090) );
  AND2_X1 U12599 ( .A1(n10093), .A2(P2_U3088), .ZN(n14093) );
  INV_X2 U12600 ( .A(n14093), .ZN(n14092) );
  AND2_X1 U12601 ( .A1(n10065), .A2(P2_U3088), .ZN(n11332) );
  AOI22_X1 U12602 ( .A1(n13509), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n11332), .ZN(n10066) );
  OAI21_X1 U12603 ( .B1(n10090), .B2(n14092), .A(n10066), .ZN(P2_U3321) );
  NAND2_X1 U12604 ( .A1(n10068), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10069) );
  XNOR2_X1 U12605 ( .A(n10105), .B(n15542), .ZN(n10103) );
  XNOR2_X1 U12606 ( .A(n10103), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12607 ( .A1(n10073), .A2(n10072), .ZN(n10078) );
  INV_X1 U12608 ( .A(n10074), .ZN(n10075) );
  OR2_X1 U12609 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  NAND2_X1 U12610 ( .A1(n10078), .A2(n10077), .ZN(n10080) );
  AOI21_X1 U12611 ( .B1(n10081), .B2(n10080), .A(n10079), .ZN(SUB_1596_U59) );
  INV_X2 U12612 ( .A(n11332), .ZN(n14097) );
  OAI222_X1 U12613 ( .A1(n14097), .A2(n10083), .B1(n14092), .B2(n10082), .C1(
        P2_U3088), .C2(n13489), .ZN(P2_U3322) );
  OAI222_X1 U12614 ( .A1(n14097), .A2(n10085), .B1(n14092), .B2(n10084), .C1(
        P2_U3088), .C2(n13468), .ZN(P2_U3324) );
  OAI222_X1 U12615 ( .A1(n14097), .A2(n10087), .B1(n14092), .B2(n10086), .C1(
        P2_U3088), .C2(n10219), .ZN(P2_U3323) );
  OAI222_X1 U12616 ( .A1(n14097), .A2(n10089), .B1(n14092), .B2(n10088), .C1(
        P2_U3088), .C2(n13458), .ZN(P2_U3325) );
  INV_X1 U12617 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10091) );
  INV_X1 U12618 ( .A(n14549), .ZN(n10321) );
  OAI222_X1 U12619 ( .A1(n15105), .A2(n10091), .B1(n10976), .B2(n10090), .C1(
        P1_U3086), .C2(n10321), .ZN(P1_U3349) );
  OAI222_X1 U12620 ( .A1(n10541), .A2(P2_U3088), .B1(n14092), .B2(n10110), 
        .C1(n10092), .C2(n14097), .ZN(P2_U3326) );
  NOR2_X1 U12621 ( .A1(n6409), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13016) );
  INV_X2 U12622 ( .A(n13016), .ZN(n13039) );
  NAND2_X1 U12623 ( .A1(n10093), .A2(P3_U3151), .ZN(n13034) );
  INV_X1 U12624 ( .A(n10096), .ZN(n10140) );
  INV_X1 U12625 ( .A(n10283), .ZN(n10097) );
  OAI222_X1 U12626 ( .A1(n14097), .A2(n10098), .B1(n14092), .B2(n10140), .C1(
        P2_U3088), .C2(n10097), .ZN(P2_U3320) );
  INV_X1 U12627 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15512) );
  NOR2_X1 U12628 ( .A1(n10132), .A2(n15512), .ZN(P3_U3254) );
  INV_X1 U12629 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15471) );
  NOR2_X1 U12630 ( .A1(n10132), .A2(n15471), .ZN(P3_U3255) );
  OAI222_X1 U12631 ( .A1(n13039), .A2(n10100), .B1(n13034), .B2(n10099), .C1(
        P3_U3151), .C2(n10507), .ZN(P3_U3295) );
  OAI222_X1 U12632 ( .A1(P3_U3151), .A2(n11379), .B1(n13034), .B2(n10102), 
        .C1(n13039), .C2(n10101), .ZN(P3_U3286) );
  NAND2_X1 U12633 ( .A1(n10103), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10104) );
  NAND2_X1 U12634 ( .A1(n10105), .A2(n15542), .ZN(n10108) );
  NAND2_X1 U12635 ( .A1(n10106), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10107) );
  INV_X1 U12636 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10258) );
  XNOR2_X1 U12637 ( .A(n10167), .B(n10258), .ZN(n10174) );
  INV_X1 U12638 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n13485) );
  XNOR2_X1 U12639 ( .A(n10173), .B(n13485), .ZN(SUB_1596_U58) );
  OAI222_X1 U12640 ( .A1(n14503), .A2(P1_U3086), .B1(n10976), .B2(n10110), 
        .C1(n10109), .C2(n15105), .ZN(P1_U3354) );
  INV_X1 U12641 ( .A(n10111), .ZN(n10113) );
  INV_X1 U12642 ( .A(n10302), .ZN(n10282) );
  OAI222_X1 U12643 ( .A1(n14097), .A2(n10112), .B1(n14092), .B2(n10113), .C1(
        P2_U3088), .C2(n10282), .ZN(P2_U3319) );
  INV_X1 U12644 ( .A(n10324), .ZN(n10341) );
  OAI222_X1 U12645 ( .A1(n15105), .A2(n10114), .B1(n10976), .B2(n10113), .C1(
        P1_U3086), .C2(n10341), .ZN(P1_U3347) );
  INV_X1 U12646 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10119) );
  INV_X1 U12647 ( .A(n10116), .ZN(n10117) );
  AOI22_X1 U12648 ( .A1(n15230), .A2(n10119), .B1(n10118), .B2(n10117), .ZN(
        P1_U3446) );
  INV_X1 U12649 ( .A(n13034), .ZN(n10816) );
  OAI222_X1 U12650 ( .A1(P3_U3151), .A2(n10607), .B1(n13036), .B2(n10121), 
        .C1(n13039), .C2(n10120), .ZN(P3_U3292) );
  OAI222_X1 U12651 ( .A1(P3_U3151), .A2(n10727), .B1(n13036), .B2(n10123), 
        .C1(n13039), .C2(n10122), .ZN(P3_U3291) );
  OAI222_X1 U12652 ( .A1(P3_U3151), .A2(n10655), .B1(n13036), .B2(n10124), 
        .C1(n13039), .C2(n7845), .ZN(P3_U3289) );
  INV_X1 U12653 ( .A(n10877), .ZN(n10871) );
  INV_X1 U12654 ( .A(SI_7_), .ZN(n10127) );
  INV_X1 U12655 ( .A(n10125), .ZN(n10126) );
  OAI222_X1 U12656 ( .A1(P3_U3151), .A2(n10871), .B1(n13036), .B2(n10127), 
        .C1(n13039), .C2(n10126), .ZN(P3_U3288) );
  OAI222_X1 U12657 ( .A1(n6403), .A2(P3_U3151), .B1(n13039), .B2(n10129), .C1(
        n10128), .C2(n13034), .ZN(P3_U3285) );
  OAI222_X1 U12658 ( .A1(P3_U3151), .A2(n11144), .B1(n13036), .B2(n10131), 
        .C1(n13039), .C2(n10130), .ZN(P3_U3287) );
  AND2_X1 U12659 ( .A1(n10133), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12660 ( .A1(n10133), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12661 ( .A1(n10133), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12662 ( .A1(n10133), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12663 ( .A1(n10133), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12664 ( .A1(n10133), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12665 ( .A1(n10133), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12666 ( .A1(n10133), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12667 ( .A1(n10133), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12668 ( .A1(n10133), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12669 ( .A1(n10133), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12670 ( .A1(n10133), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12671 ( .A1(n10133), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12672 ( .A1(n10133), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12673 ( .A1(n10133), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12674 ( .A1(n10133), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12675 ( .A1(n10133), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12676 ( .A1(n10133), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12677 ( .A1(n10133), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12678 ( .A1(n10133), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12679 ( .A1(n10133), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12680 ( .A1(n10133), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12681 ( .A1(n10133), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12682 ( .A1(n10133), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12683 ( .A1(n10133), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12684 ( .A1(n10133), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12685 ( .A1(n10133), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12686 ( .A1(n10133), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  OAI222_X1 U12687 ( .A1(n10625), .A2(P3_U3151), .B1(n13039), .B2(n10135), 
        .C1(n10134), .C2(n13036), .ZN(P3_U3290) );
  INV_X1 U12688 ( .A(n10136), .ZN(n10138) );
  INV_X1 U12689 ( .A(SI_2_), .ZN(n10137) );
  OAI222_X1 U12690 ( .A1(P3_U3151), .A2(n6909), .B1(n13039), .B2(n10138), .C1(
        n10137), .C2(n13036), .ZN(P3_U3293) );
  INV_X1 U12691 ( .A(n10358), .ZN(n10139) );
  OAI222_X1 U12692 ( .A1(n15105), .A2(n8621), .B1(n10976), .B2(n10140), .C1(
        P1_U3086), .C2(n10139), .ZN(P1_U3348) );
  NOR2_X1 U12693 ( .A1(n10757), .A2(P1_U3086), .ZN(n14469) );
  INV_X1 U12694 ( .A(n14469), .ZN(n14244) );
  NAND2_X1 U12695 ( .A1(n10141), .A2(n14244), .ZN(n10161) );
  INV_X1 U12696 ( .A(n10757), .ZN(n10142) );
  OR2_X1 U12697 ( .A1(n14432), .A2(n10142), .ZN(n10143) );
  NAND2_X1 U12698 ( .A1(n10143), .A2(n7116), .ZN(n10159) );
  NOR2_X1 U12699 ( .A1(n15199), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12700 ( .A(n10144), .ZN(n10146) );
  INV_X1 U12701 ( .A(n14567), .ZN(n10336) );
  OAI222_X1 U12702 ( .A1(n15105), .A2(n10145), .B1(n10976), .B2(n10146), .C1(
        P1_U3086), .C2(n10336), .ZN(P1_U3346) );
  INV_X1 U12703 ( .A(n10663), .ZN(n10293) );
  OAI222_X1 U12704 ( .A1(n14097), .A2(n10147), .B1(n14092), .B2(n10146), .C1(
        P2_U3088), .C2(n10293), .ZN(P2_U3318) );
  INV_X1 U12705 ( .A(n15230), .ZN(n15229) );
  OAI22_X1 U12706 ( .A1(n15229), .A2(P1_D_REG_0__SCAN_IN), .B1(n10149), .B2(
        n10148), .ZN(n10150) );
  INV_X1 U12707 ( .A(n10150), .ZN(P1_U3445) );
  INV_X1 U12708 ( .A(n10151), .ZN(n10153) );
  INV_X1 U12709 ( .A(n10343), .ZN(n10459) );
  OAI222_X1 U12710 ( .A1(n15105), .A2(n6713), .B1(n10976), .B2(n10153), .C1(
        P1_U3086), .C2(n10459), .ZN(P1_U3345) );
  INV_X1 U12711 ( .A(n10714), .ZN(n10152) );
  OAI222_X1 U12712 ( .A1(n14097), .A2(n10154), .B1(n14092), .B2(n10153), .C1(
        P2_U3088), .C2(n10152), .ZN(P2_U3317) );
  INV_X1 U12713 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15530) );
  NAND2_X1 U12714 ( .A1(P3_U3897), .A2(n12162), .ZN(n10155) );
  OAI21_X1 U12715 ( .B1(P3_U3897), .B2(n15530), .A(n10155), .ZN(P3_U3501) );
  INV_X1 U12716 ( .A(n11732), .ZN(n12529) );
  INV_X1 U12717 ( .A(n10156), .ZN(n10157) );
  OAI222_X1 U12718 ( .A1(P3_U3151), .A2(n12529), .B1(n13036), .B2(n10158), 
        .C1(n13039), .C2(n10157), .ZN(P3_U3284) );
  INV_X1 U12719 ( .A(n15199), .ZN(n14583) );
  INV_X1 U12720 ( .A(n10159), .ZN(n10160) );
  NAND2_X1 U12721 ( .A1(n10161), .A2(n10160), .ZN(n10261) );
  INV_X1 U12722 ( .A(n10261), .ZN(n10164) );
  INV_X1 U12723 ( .A(n15106), .ZN(n10257) );
  AOI21_X1 U12724 ( .B1(n10257), .B2(n9349), .A(n9784), .ZN(n14515) );
  OAI21_X1 U12725 ( .B1(n10257), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14515), .ZN(
        n10162) );
  XNOR2_X1 U12726 ( .A(n10162), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U12727 ( .A1(n10164), .A2(n10163), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10165) );
  OAI21_X1 U12728 ( .B1(n10166), .B2(n14583), .A(n10165), .ZN(P1_U3243) );
  NAND2_X1 U12729 ( .A1(n10168), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10169) );
  NOR2_X1 U12730 ( .A1(n14547), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U12731 ( .A1(n10402), .A2(n10171), .ZN(n10172) );
  XNOR2_X1 U12732 ( .A(n10404), .B(n10172), .ZN(n10180) );
  NAND2_X1 U12733 ( .A1(n10173), .A2(n13485), .ZN(n10178) );
  INV_X1 U12734 ( .A(n10174), .ZN(n10175) );
  OR2_X1 U12735 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U12736 ( .A1(n10179), .A2(n10180), .ZN(n10409) );
  OAI21_X1 U12737 ( .B1(n10180), .B2(n10179), .A(n10409), .ZN(n10181) );
  INV_X1 U12738 ( .A(n10181), .ZN(SUB_1596_U57) );
  OAI222_X1 U12739 ( .A1(P3_U3151), .A2(n12560), .B1(n13036), .B2(n10183), 
        .C1(n13039), .C2(n10182), .ZN(P3_U3283) );
  INV_X1 U12740 ( .A(n10184), .ZN(n10186) );
  INV_X1 U12741 ( .A(n10965), .ZN(n10955) );
  OAI222_X1 U12742 ( .A1(n14097), .A2(n10185), .B1(n14092), .B2(n10186), .C1(
        P2_U3088), .C2(n10955), .ZN(P2_U3316) );
  OAI222_X1 U12743 ( .A1(n15105), .A2(n10187), .B1(n10976), .B2(n10186), .C1(
        P1_U3086), .C2(n10773), .ZN(P1_U3344) );
  INV_X1 U12744 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10381) );
  MUX2_X1 U12745 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10381), .S(n10541), .Z(
        n10534) );
  NAND2_X1 U12746 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10535) );
  NOR2_X1 U12747 ( .A1(n10541), .A2(n10381), .ZN(n13453) );
  INV_X1 U12748 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10188) );
  MUX2_X1 U12749 ( .A(n10188), .B(P2_REG1_REG_2__SCAN_IN), .S(n13458), .Z(
        n10189) );
  OAI21_X1 U12750 ( .B1(n13457), .B2(n13453), .A(n10189), .ZN(n13476) );
  INV_X1 U12751 ( .A(n13458), .ZN(n13463) );
  NAND2_X1 U12752 ( .A1(n13463), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13475) );
  MUX2_X1 U12753 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8767), .S(n13468), .Z(
        n13474) );
  AOI21_X1 U12754 ( .B1(n13476), .B2(n13475), .A(n13474), .ZN(n15278) );
  NOR2_X1 U12755 ( .A1(n13468), .A2(n8767), .ZN(n15277) );
  INV_X1 U12756 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U12757 ( .A(n10190), .B(P2_REG1_REG_4__SCAN_IN), .S(n10219), .Z(
        n15276) );
  INV_X1 U12758 ( .A(n10219), .ZN(n15283) );
  NAND2_X1 U12759 ( .A1(n15283), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n13494) );
  INV_X1 U12760 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11040) );
  MUX2_X1 U12761 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n11040), .S(n13489), .Z(
        n13493) );
  INV_X1 U12762 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10191) );
  MUX2_X1 U12763 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10191), .S(n13509), .Z(
        n10192) );
  NAND2_X1 U12764 ( .A1(n13509), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10202) );
  INV_X1 U12765 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15388) );
  MUX2_X1 U12766 ( .A(n15388), .B(P2_REG1_REG_7__SCAN_IN), .S(n10283), .Z(
        n10201) );
  INV_X1 U12767 ( .A(n11331), .ZN(n10194) );
  OAI21_X1 U12768 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10196) );
  AND2_X1 U12769 ( .A1(n10197), .A2(n10196), .ZN(n10204) );
  INV_X1 U12770 ( .A(n10204), .ZN(n10207) );
  OR2_X1 U12771 ( .A1(n10205), .A2(P2_U3088), .ZN(n14095) );
  INV_X1 U12772 ( .A(n14095), .ZN(n10198) );
  NAND2_X1 U12773 ( .A1(n10207), .A2(n10198), .ZN(n10210) );
  INV_X1 U12774 ( .A(n10210), .ZN(n10200) );
  NAND3_X1 U12775 ( .A1(n13506), .A2(n10202), .A3(n10201), .ZN(n10203) );
  NAND2_X1 U12776 ( .A1(n15315), .A2(n10203), .ZN(n10232) );
  AND2_X1 U12777 ( .A1(n10204), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15273) );
  NAND2_X1 U12778 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n11109) );
  INV_X1 U12779 ( .A(n11109), .ZN(n10209) );
  AND2_X1 U12780 ( .A1(n10205), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10206) );
  AND2_X1 U12781 ( .A1(n15305), .A2(n10283), .ZN(n10208) );
  AOI211_X1 U12782 ( .C1(n15273), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10209), .B(
        n10208), .ZN(n10231) );
  INV_X1 U12783 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11263) );
  MUX2_X1 U12784 ( .A(n11263), .B(P2_REG2_REG_2__SCAN_IN), .S(n13458), .Z(
        n10215) );
  INV_X1 U12785 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10211) );
  MUX2_X1 U12786 ( .A(n10211), .B(P2_REG2_REG_1__SCAN_IN), .S(n10541), .Z(
        n10213) );
  AND2_X1 U12787 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10212) );
  NAND2_X1 U12788 ( .A1(n10213), .A2(n10212), .ZN(n13460) );
  OR2_X1 U12789 ( .A1(n10541), .A2(n10211), .ZN(n13459) );
  NAND2_X1 U12790 ( .A1(n13460), .A2(n13459), .ZN(n10214) );
  NAND2_X1 U12791 ( .A1(n13463), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U12792 ( .A1(n13470), .A2(n13469), .ZN(n10217) );
  INV_X1 U12793 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11430) );
  MUX2_X1 U12794 ( .A(n11430), .B(P2_REG2_REG_3__SCAN_IN), .S(n13468), .Z(
        n10216) );
  NAND2_X1 U12795 ( .A1(n10217), .A2(n10216), .ZN(n13473) );
  INV_X1 U12796 ( .A(n13468), .ZN(n13479) );
  NAND2_X1 U12797 ( .A1(n13479), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12798 ( .A1(n13473), .A2(n10218), .ZN(n15285) );
  INV_X1 U12799 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11653) );
  MUX2_X1 U12800 ( .A(n11653), .B(P2_REG2_REG_4__SCAN_IN), .S(n10219), .Z(
        n15286) );
  OR2_X1 U12801 ( .A1(n10219), .A2(n11653), .ZN(n13491) );
  NAND2_X1 U12802 ( .A1(n15284), .A2(n13491), .ZN(n10221) );
  INV_X1 U12803 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11275) );
  MUX2_X1 U12804 ( .A(n11275), .B(P2_REG2_REG_5__SCAN_IN), .S(n13489), .Z(
        n10220) );
  NAND2_X1 U12805 ( .A1(n10221), .A2(n10220), .ZN(n13501) );
  OR2_X1 U12806 ( .A1(n13489), .A2(n11275), .ZN(n13500) );
  NAND2_X1 U12807 ( .A1(n13501), .A2(n13500), .ZN(n10223) );
  INV_X1 U12808 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11634) );
  MUX2_X1 U12809 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11634), .S(n13509), .Z(
        n10222) );
  NAND2_X1 U12810 ( .A1(n10223), .A2(n10222), .ZN(n13503) );
  NAND2_X1 U12811 ( .A1(n13509), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U12812 ( .A1(n13503), .A2(n10228), .ZN(n10225) );
  INV_X1 U12813 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U12814 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10226), .S(n10283), .Z(
        n10224) );
  MUX2_X1 U12815 ( .A(n10226), .B(P2_REG2_REG_7__SCAN_IN), .S(n10283), .Z(
        n10227) );
  NAND3_X1 U12816 ( .A1(n13503), .A2(n10228), .A3(n10227), .ZN(n10229) );
  NAND3_X1 U12817 ( .A1(n15318), .A2(n10306), .A3(n10229), .ZN(n10230) );
  OAI211_X1 U12818 ( .C1(n10280), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        P2_U3221) );
  INV_X1 U12819 ( .A(n10233), .ZN(n10242) );
  INV_X1 U12820 ( .A(n14586), .ZN(n10234) );
  OAI222_X1 U12821 ( .A1(n15105), .A2(n10235), .B1(n10976), .B2(n10242), .C1(
        n10234), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12822 ( .A(n15304), .ZN(n10238) );
  INV_X1 U12823 ( .A(n10236), .ZN(n10239) );
  OAI222_X1 U12824 ( .A1(P2_U3088), .A2(n10238), .B1(n14092), .B2(n10239), 
        .C1(n10237), .C2(n14097), .ZN(P2_U3315) );
  INV_X1 U12825 ( .A(n11238), .ZN(n11232) );
  OAI222_X1 U12826 ( .A1(n15105), .A2(n10240), .B1(n10976), .B2(n10239), .C1(
        n11232), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12827 ( .A(n11504), .ZN(n10243) );
  OAI222_X1 U12828 ( .A1(P2_U3088), .A2(n10243), .B1(n14092), .B2(n10242), 
        .C1(n10241), .C2(n14097), .ZN(P2_U3314) );
  MUX2_X1 U12829 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10244), .S(n10313), .Z(
        n10256) );
  MUX2_X1 U12830 ( .A(n10245), .B(P1_REG1_REG_2__SCAN_IN), .S(n14522), .Z(
        n10248) );
  MUX2_X1 U12831 ( .A(n10246), .B(P1_REG1_REG_1__SCAN_IN), .S(n14503), .Z(
        n14500) );
  AND2_X1 U12832 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14501) );
  OR2_X1 U12833 ( .A1(n14503), .A2(n10246), .ZN(n14516) );
  NAND2_X1 U12834 ( .A1(n14517), .A2(n14516), .ZN(n10247) );
  INV_X1 U12835 ( .A(n14522), .ZN(n10266) );
  NAND2_X1 U12836 ( .A1(n10266), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U12837 ( .A1(n14536), .A2(n14534), .ZN(n10251) );
  MUX2_X1 U12838 ( .A(n10249), .B(P1_REG1_REG_3__SCAN_IN), .S(n14538), .Z(
        n10250) );
  OR2_X1 U12839 ( .A1(n14538), .A2(n10249), .ZN(n15184) );
  MUX2_X1 U12840 ( .A(n10252), .B(P1_REG1_REG_4__SCAN_IN), .S(n15195), .Z(
        n10253) );
  NAND2_X1 U12841 ( .A1(n10254), .A2(n10253), .ZN(n15187) );
  OAI21_X1 U12842 ( .B1(n10252), .B2(n15195), .A(n15187), .ZN(n10255) );
  AOI21_X1 U12843 ( .B1(n10256), .B2(n10255), .A(n10312), .ZN(n10279) );
  INV_X1 U12844 ( .A(n10313), .ZN(n10319) );
  NAND2_X1 U12845 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11556) );
  OAI21_X1 U12846 ( .B1(n14583), .B2(n10258), .A(n11556), .ZN(n10259) );
  AOI21_X1 U12847 ( .B1(n10319), .B2(n15197), .A(n10259), .ZN(n10278) );
  OR2_X1 U12848 ( .A1(n9784), .A2(n15106), .ZN(n10260) );
  OR2_X1 U12849 ( .A1(n10261), .A2(n10260), .ZN(n14637) );
  MUX2_X1 U12850 ( .A(n10262), .B(P1_REG2_REG_2__SCAN_IN), .S(n14522), .Z(
        n10265) );
  MUX2_X1 U12851 ( .A(n10263), .B(P1_REG2_REG_1__SCAN_IN), .S(n14503), .Z(
        n14502) );
  AND2_X1 U12852 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14510) );
  NAND2_X1 U12853 ( .A1(n14502), .A2(n14510), .ZN(n14524) );
  OR2_X1 U12854 ( .A1(n14503), .A2(n10263), .ZN(n14523) );
  NAND2_X1 U12855 ( .A1(n14524), .A2(n14523), .ZN(n10264) );
  NAND2_X1 U12856 ( .A1(n10265), .A2(n10264), .ZN(n14541) );
  NAND2_X1 U12857 ( .A1(n10266), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U12858 ( .A1(n14541), .A2(n14539), .ZN(n10269) );
  MUX2_X1 U12859 ( .A(n10267), .B(P1_REG2_REG_3__SCAN_IN), .S(n14538), .Z(
        n10268) );
  NAND2_X1 U12860 ( .A1(n10269), .A2(n10268), .ZN(n15191) );
  OR2_X1 U12861 ( .A1(n14538), .A2(n10267), .ZN(n15190) );
  MUX2_X1 U12862 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n15219), .S(n15195), .Z(
        n15189) );
  AOI21_X1 U12863 ( .B1(n15191), .B2(n15190), .A(n15189), .ZN(n10271) );
  NOR2_X1 U12864 ( .A1(n15195), .A2(n15219), .ZN(n10272) );
  MUX2_X1 U12865 ( .A(n10273), .B(P1_REG2_REG_5__SCAN_IN), .S(n10313), .Z(
        n10270) );
  OAI21_X1 U12866 ( .B1(n10271), .B2(n10272), .A(n10270), .ZN(n14555) );
  INV_X1 U12867 ( .A(n10271), .ZN(n15193) );
  INV_X1 U12868 ( .A(n10272), .ZN(n10275) );
  INV_X1 U12869 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10273) );
  MUX2_X1 U12870 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10273), .S(n10313), .Z(
        n10274) );
  NAND3_X1 U12871 ( .A1(n15193), .A2(n10275), .A3(n10274), .ZN(n10276) );
  NAND3_X1 U12872 ( .A1(n15194), .A2(n14555), .A3(n10276), .ZN(n10277) );
  OAI211_X1 U12873 ( .C1(n10279), .C2(n14635), .A(n10278), .B(n10277), .ZN(
        P1_U3248) );
  XNOR2_X1 U12874 ( .A(n10663), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10660) );
  AOI21_X1 U12875 ( .B1(n10283), .B2(P2_REG1_REG_7__SCAN_IN), .A(n10280), .ZN(
        n10299) );
  XNOR2_X1 U12876 ( .A(n10302), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n10298) );
  INV_X1 U12877 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10281) );
  XOR2_X1 U12878 ( .A(n10660), .B(n10661), .Z(n10297) );
  NAND2_X1 U12879 ( .A1(n10283), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12880 ( .A1(n10306), .A2(n10305), .ZN(n10285) );
  INV_X1 U12881 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10303) );
  MUX2_X1 U12882 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10303), .S(n10302), .Z(
        n10284) );
  NAND2_X1 U12883 ( .A1(n10285), .A2(n10284), .ZN(n10308) );
  NAND2_X1 U12884 ( .A1(n10302), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U12885 ( .A1(n10308), .A2(n10286), .ZN(n10289) );
  INV_X1 U12886 ( .A(n10289), .ZN(n10291) );
  INV_X1 U12887 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10287) );
  MUX2_X1 U12888 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10287), .S(n10663), .Z(
        n10290) );
  MUX2_X1 U12889 ( .A(n10287), .B(P2_REG2_REG_9__SCAN_IN), .S(n10663), .Z(
        n10288) );
  OAI21_X1 U12890 ( .B1(n10291), .B2(n10290), .A(n10665), .ZN(n10295) );
  NAND2_X1 U12891 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U12892 ( .A1(n15273), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10292) );
  OAI211_X1 U12893 ( .C1(n15313), .C2(n10293), .A(n11205), .B(n10292), .ZN(
        n10294) );
  AOI21_X1 U12894 ( .B1(n15318), .B2(n10295), .A(n10294), .ZN(n10296) );
  OAI21_X1 U12895 ( .B1(n10297), .B2(n15300), .A(n10296), .ZN(P2_U3223) );
  XNOR2_X1 U12896 ( .A(n10299), .B(n10298), .ZN(n10311) );
  NAND2_X1 U12897 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11067) );
  INV_X1 U12898 ( .A(n11067), .ZN(n10301) );
  INV_X1 U12899 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n11159) );
  NOR2_X1 U12900 ( .A1(n15322), .A2(n11159), .ZN(n10300) );
  AOI211_X1 U12901 ( .C1(n15305), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10310) );
  MUX2_X1 U12902 ( .A(n10303), .B(P2_REG2_REG_8__SCAN_IN), .S(n10302), .Z(
        n10304) );
  NAND3_X1 U12903 ( .A1(n10306), .A2(n10305), .A3(n10304), .ZN(n10307) );
  NAND3_X1 U12904 ( .A1(n15318), .A2(n10308), .A3(n10307), .ZN(n10309) );
  OAI211_X1 U12905 ( .C1(n10311), .C2(n15300), .A(n10310), .B(n10309), .ZN(
        P2_U3222) );
  MUX2_X1 U12906 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10314), .S(n14549), .Z(
        n14551) );
  NAND2_X1 U12907 ( .A1(n14549), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10353) );
  MUX2_X1 U12908 ( .A(n9425), .B(P1_REG1_REG_7__SCAN_IN), .S(n10358), .Z(
        n10352) );
  NOR2_X1 U12909 ( .A1(n10324), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10332) );
  AOI21_X1 U12910 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10324), .A(n10332), .ZN(
        n10315) );
  NAND2_X1 U12911 ( .A1(n10316), .A2(n10315), .ZN(n10334) );
  OAI21_X1 U12912 ( .B1(n10316), .B2(n10315), .A(n10334), .ZN(n10330) );
  NAND2_X1 U12913 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10318) );
  NAND2_X1 U12914 ( .A1(n15199), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10317) );
  OAI211_X1 U12915 ( .C1(n14633), .C2(n10341), .A(n10318), .B(n10317), .ZN(
        n10329) );
  NAND2_X1 U12916 ( .A1(n10319), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14554) );
  MUX2_X1 U12917 ( .A(n10320), .B(P1_REG2_REG_6__SCAN_IN), .S(n14549), .Z(
        n14553) );
  AOI21_X1 U12918 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n10356) );
  NOR2_X1 U12919 ( .A1(n10321), .A2(n10320), .ZN(n10357) );
  INV_X1 U12920 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10322) );
  MUX2_X1 U12921 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10322), .S(n10358), .Z(
        n10323) );
  OAI21_X1 U12922 ( .B1(n10356), .B2(n10357), .A(n10323), .ZN(n10362) );
  NAND2_X1 U12923 ( .A1(n10358), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10326) );
  INV_X1 U12924 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10340) );
  MUX2_X1 U12925 ( .A(n10340), .B(P1_REG2_REG_8__SCAN_IN), .S(n10324), .Z(
        n10325) );
  AOI21_X1 U12926 ( .B1(n10362), .B2(n10326), .A(n10325), .ZN(n14573) );
  AND3_X1 U12927 ( .A1(n10362), .A2(n10326), .A3(n10325), .ZN(n10327) );
  NOR3_X1 U12928 ( .A1(n14637), .A2(n14573), .A3(n10327), .ZN(n10328) );
  AOI211_X1 U12929 ( .C1(n10330), .C2(n15188), .A(n10329), .B(n10328), .ZN(
        n10331) );
  INV_X1 U12930 ( .A(n10331), .ZN(P1_U3251) );
  INV_X1 U12931 ( .A(n10332), .ZN(n10333) );
  NAND2_X1 U12932 ( .A1(n10334), .A2(n10333), .ZN(n14562) );
  XNOR2_X1 U12933 ( .A(n14567), .B(n10335), .ZN(n14563) );
  XNOR2_X1 U12934 ( .A(n10343), .B(n10452), .ZN(n10337) );
  NAND2_X1 U12935 ( .A1(n10336), .A2(n10335), .ZN(n10338) );
  NAND2_X1 U12936 ( .A1(n10451), .A2(n15188), .ZN(n10351) );
  AOI21_X1 U12937 ( .B1(n14561), .B2(n10338), .A(n10337), .ZN(n10350) );
  INV_X1 U12938 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U12939 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12005)
         );
  OAI21_X1 U12940 ( .B1(n14583), .B2(n11253), .A(n12005), .ZN(n10339) );
  AOI21_X1 U12941 ( .B1(n10343), .B2(n15197), .A(n10339), .ZN(n10349) );
  NOR2_X1 U12942 ( .A1(n10341), .A2(n10340), .ZN(n14568) );
  INV_X1 U12943 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11833) );
  MUX2_X1 U12944 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11833), .S(n14567), .Z(
        n10342) );
  OAI21_X1 U12945 ( .B1(n14573), .B2(n14568), .A(n10342), .ZN(n14571) );
  NAND2_X1 U12946 ( .A1(n14567), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10345) );
  INV_X1 U12947 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10458) );
  MUX2_X1 U12948 ( .A(n10458), .B(P1_REG2_REG_10__SCAN_IN), .S(n10343), .Z(
        n10344) );
  AOI21_X1 U12949 ( .B1(n14571), .B2(n10345), .A(n10344), .ZN(n10466) );
  INV_X1 U12950 ( .A(n10466), .ZN(n10347) );
  NAND3_X1 U12951 ( .A1(n14571), .A2(n10345), .A3(n10344), .ZN(n10346) );
  NAND3_X1 U12952 ( .A1(n10347), .A2(n15194), .A3(n10346), .ZN(n10348) );
  OAI211_X1 U12953 ( .C1(n10351), .C2(n10350), .A(n10349), .B(n10348), .ZN(
        P1_U3253) );
  NAND3_X1 U12954 ( .A1(n14550), .A2(n10353), .A3(n10352), .ZN(n10354) );
  NAND2_X1 U12955 ( .A1(n15188), .A2(n10354), .ZN(n10365) );
  INV_X1 U12956 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U12957 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11543) );
  OAI21_X1 U12958 ( .B1(n14583), .B2(n10405), .A(n11543), .ZN(n10355) );
  AOI21_X1 U12959 ( .B1(n10358), .B2(n15197), .A(n10355), .ZN(n10364) );
  INV_X1 U12960 ( .A(n10356), .ZN(n14557) );
  INV_X1 U12961 ( .A(n10357), .ZN(n10360) );
  MUX2_X1 U12962 ( .A(n10322), .B(P1_REG2_REG_7__SCAN_IN), .S(n10358), .Z(
        n10359) );
  NAND3_X1 U12963 ( .A1(n14557), .A2(n10360), .A3(n10359), .ZN(n10361) );
  NAND3_X1 U12964 ( .A1(n15194), .A2(n10362), .A3(n10361), .ZN(n10363) );
  OAI211_X1 U12965 ( .C1(n10366), .C2(n10365), .A(n10364), .B(n10363), .ZN(
        P1_U3250) );
  INV_X1 U12966 ( .A(n11696), .ZN(n11688) );
  INV_X1 U12967 ( .A(n10367), .ZN(n10369) );
  OAI222_X1 U12968 ( .A1(P2_U3088), .A2(n11688), .B1(n14092), .B2(n10369), 
        .C1(n10368), .C2(n14097), .ZN(P2_U3311) );
  INV_X1 U12969 ( .A(n14593), .ZN(n14601) );
  OAI222_X1 U12970 ( .A1(n15105), .A2(n10370), .B1(n10976), .B2(n10369), .C1(
        n14601), .C2(P1_U3086), .ZN(P1_U3339) );
  NAND2_X1 U12971 ( .A1(n15358), .A2(n10371), .ZN(n10372) );
  OR2_X1 U12972 ( .A1(n13374), .A2(n6414), .ZN(n15371) );
  INV_X1 U12973 ( .A(n10374), .ZN(n10378) );
  INV_X1 U12974 ( .A(n10375), .ZN(n10376) );
  AOI21_X1 U12975 ( .B1(n15377), .B2(n10017), .A(n10376), .ZN(n10377) );
  OAI211_X1 U12976 ( .C1(n10379), .C2(n15371), .A(n10378), .B(n10377), .ZN(
        n10385) );
  NAND2_X1 U12977 ( .A1(n10385), .A2(n15390), .ZN(n10380) );
  OAI21_X1 U12978 ( .B1(n15390), .B2(n10381), .A(n10380), .ZN(P2_U3500) );
  INV_X1 U12979 ( .A(n10382), .ZN(n10383) );
  INV_X1 U12980 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U12981 ( .A1(n10385), .A2(n15384), .ZN(n10386) );
  OAI21_X1 U12982 ( .B1(n15384), .B2(n10387), .A(n10386), .ZN(P2_U3433) );
  OAI222_X1 U12983 ( .A1(P3_U3151), .A2(n12573), .B1(n13034), .B2(n10389), 
        .C1(n13039), .C2(n10388), .ZN(P3_U3282) );
  INV_X1 U12984 ( .A(n11507), .ZN(n15312) );
  INV_X1 U12985 ( .A(n10390), .ZN(n10393) );
  OAI222_X1 U12986 ( .A1(P2_U3088), .A2(n15312), .B1(n14092), .B2(n10393), 
        .C1(n10391), .C2(n14097), .ZN(P2_U3313) );
  INV_X1 U12987 ( .A(n11617), .ZN(n10392) );
  OAI222_X1 U12988 ( .A1(n15105), .A2(n10394), .B1(n10976), .B2(n10393), .C1(
        n10392), .C2(P1_U3086), .ZN(P1_U3341) );
  XOR2_X1 U12989 ( .A(n10396), .B(n10395), .Z(n10400) );
  NAND2_X1 U12990 ( .A1(n13161), .A2(n13883), .ZN(n13143) );
  INV_X1 U12991 ( .A(n13143), .ZN(n13191) );
  NOR2_X1 U12992 ( .A1(n10397), .A2(P2_U3088), .ZN(n10556) );
  INV_X1 U12993 ( .A(n10556), .ZN(n10416) );
  AOI22_X1 U12994 ( .A1(n13191), .A2(n13452), .B1(n10416), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10399) );
  AND2_X1 U12995 ( .A1(n13161), .A2(n13885), .ZN(n13053) );
  AOI22_X1 U12996 ( .A1(n10017), .A2(n13173), .B1(n13053), .B2(n13449), .ZN(
        n10398) );
  OAI211_X1 U12997 ( .C1(n10400), .C2(n13165), .A(n10399), .B(n10398), .ZN(
        P2_U3194) );
  INV_X1 U12998 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U12999 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10401), .ZN(n10403) );
  XNOR2_X1 U13000 ( .A(n10720), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n10719) );
  XNOR2_X1 U13001 ( .A(n10719), .B(n10405), .ZN(n10412) );
  INV_X1 U13002 ( .A(n10406), .ZN(n10407) );
  NAND2_X1 U13003 ( .A1(n10407), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10408) );
  INV_X1 U13004 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U13005 ( .A1(n10411), .A2(n10412), .ZN(n10718) );
  OAI21_X1 U13006 ( .B1(n10412), .B2(n10411), .A(n10718), .ZN(n10413) );
  INV_X1 U13007 ( .A(n10413), .ZN(SUB_1596_U56) );
  XOR2_X1 U13008 ( .A(n10414), .B(n10415), .Z(n10419) );
  AOI22_X1 U13009 ( .A1(n13191), .A2(n13450), .B1(n13173), .B2(n15361), .ZN(
        n10418) );
  AOI22_X1 U13010 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(n10416), .B1(n13053), 
        .B2(n13448), .ZN(n10417) );
  OAI211_X1 U13011 ( .C1(n10419), .C2(n13165), .A(n10418), .B(n10417), .ZN(
        P2_U3209) );
  INV_X1 U13012 ( .A(n10420), .ZN(n10422) );
  OAI222_X1 U13013 ( .A1(n12624), .A2(P3_U3151), .B1(n13039), .B2(n10422), 
        .C1(n10421), .C2(n13036), .ZN(P3_U3280) );
  AOI22_X1 U13014 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15318), .B1(n15315), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10427) );
  INV_X1 U13015 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10423) );
  NAND2_X1 U13016 ( .A1(n15315), .A2(n10423), .ZN(n10424) );
  OAI211_X1 U13017 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n15294), .A(n10424), .B(
        n15313), .ZN(n10425) );
  INV_X1 U13018 ( .A(n10425), .ZN(n10426) );
  MUX2_X1 U13019 ( .A(n10427), .B(n10426), .S(P2_IR_REG_0__SCAN_IN), .Z(n10429) );
  AOI22_X1 U13020 ( .A1(n15273), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10428) );
  NAND2_X1 U13021 ( .A1(n10429), .A2(n10428), .ZN(P2_U3214) );
  INV_X1 U13022 ( .A(P3_U3897), .ZN(n12512) );
  NAND2_X1 U13023 ( .A1(n10571), .A2(n11527), .ZN(n10444) );
  NAND2_X1 U13024 ( .A1(n10430), .A2(n10558), .ZN(n10432) );
  NAND2_X1 U13025 ( .A1(n10432), .A2(n10431), .ZN(n10443) );
  INV_X1 U13026 ( .A(n10443), .ZN(n10433) );
  INV_X1 U13027 ( .A(n10440), .ZN(n10434) );
  MUX2_X1 U13028 ( .A(n12512), .B(n10434), .S(n13027), .Z(n12697) );
  NAND2_X1 U13029 ( .A1(P3_U3897), .A2(n13027), .ZN(n12705) );
  INV_X1 U13030 ( .A(n12705), .ZN(n12584) );
  INV_X1 U13031 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10695) );
  INV_X1 U13032 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10821) );
  MUX2_X1 U13033 ( .A(n10695), .B(n10821), .S(n13031), .Z(n10500) );
  NAND2_X1 U13034 ( .A1(n10500), .A2(n10501), .ZN(n10499) );
  INV_X1 U13035 ( .A(n10499), .ZN(n10529) );
  XNOR2_X1 U13036 ( .A(n10530), .B(n10529), .ZN(n10449) );
  INV_X1 U13037 ( .A(n10435), .ZN(n10436) );
  NAND2_X1 U13038 ( .A1(n8041), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10513) );
  INV_X1 U13039 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11013) );
  OR2_X1 U13040 ( .A1(n10437), .A2(n11013), .ZN(n10514) );
  NAND2_X1 U13041 ( .A1(n10437), .A2(n11013), .ZN(n10438) );
  NAND2_X1 U13042 ( .A1(n10514), .A2(n10438), .ZN(n10439) );
  NAND2_X1 U13043 ( .A1(n12688), .A2(n10439), .ZN(n10447) );
  NAND2_X1 U13044 ( .A1(n10441), .A2(n7831), .ZN(n10519) );
  INV_X1 U13045 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10518) );
  XNOR2_X1 U13046 ( .A(n10519), .B(n10518), .ZN(n10442) );
  NAND2_X1 U13047 ( .A1(n12707), .A2(n10442), .ZN(n10446) );
  AOI22_X1 U13048 ( .A1(n15391), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10445) );
  NAND3_X1 U13049 ( .A1(n10447), .A2(n10446), .A3(n10445), .ZN(n10448) );
  AOI21_X1 U13050 ( .B1(n12584), .B2(n10449), .A(n10448), .ZN(n10450) );
  NAND2_X1 U13051 ( .A1(n10773), .A2(n10453), .ZN(n10767) );
  OAI21_X1 U13052 ( .B1(n10773), .B2(n10453), .A(n10767), .ZN(n10454) );
  AOI21_X1 U13053 ( .B1(n10455), .B2(n10454), .A(n10769), .ZN(n10469) );
  NOR2_X1 U13054 ( .A1(n10456), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14206) );
  NOR2_X1 U13055 ( .A1(n14633), .A2(n10773), .ZN(n10457) );
  AOI211_X1 U13056 ( .C1(n15199), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n14206), 
        .B(n10457), .ZN(n10468) );
  NOR2_X1 U13057 ( .A1(n10459), .A2(n10458), .ZN(n10464) );
  INV_X1 U13058 ( .A(n10464), .ZN(n10461) );
  MUX2_X1 U13059 ( .A(n10772), .B(P1_REG2_REG_11__SCAN_IN), .S(n10460), .Z(
        n10462) );
  NAND2_X1 U13060 ( .A1(n10461), .A2(n10462), .ZN(n10465) );
  INV_X1 U13061 ( .A(n10462), .ZN(n10463) );
  OAI21_X1 U13062 ( .B1(n10466), .B2(n10464), .A(n10463), .ZN(n10775) );
  OAI211_X1 U13063 ( .C1(n10466), .C2(n10465), .A(n10775), .B(n15194), .ZN(
        n10467) );
  OAI211_X1 U13064 ( .C1(n10469), .C2(n14635), .A(n10468), .B(n10467), .ZN(
        P1_U3254) );
  INV_X1 U13065 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10489) );
  INV_X1 U13066 ( .A(n13450), .ZN(n10479) );
  NAND2_X1 U13067 ( .A1(n10479), .A2(n10470), .ZN(n10472) );
  NAND2_X1 U13068 ( .A1(n10474), .A2(n10472), .ZN(n11258) );
  INV_X1 U13069 ( .A(n13396), .ZN(n11257) );
  NAND2_X1 U13070 ( .A1(n11258), .A2(n11257), .ZN(n11256) );
  XNOR2_X1 U13071 ( .A(n11426), .B(n13448), .ZN(n13399) );
  INV_X1 U13072 ( .A(n13399), .ZN(n11030) );
  NAND2_X1 U13073 ( .A1(n10482), .A2(n11266), .ZN(n10471) );
  NAND3_X1 U13074 ( .A1(n11256), .A2(n11030), .A3(n10471), .ZN(n10476) );
  AND2_X1 U13075 ( .A1(n10472), .A2(n10471), .ZN(n10473) );
  NAND2_X1 U13076 ( .A1(n10474), .A2(n10473), .ZN(n10475) );
  OAI211_X1 U13077 ( .C1(n11266), .C2(n10482), .A(n10475), .B(n13399), .ZN(
        n11403) );
  AND2_X1 U13078 ( .A1(n11403), .A2(n10476), .ZN(n11433) );
  INV_X1 U13079 ( .A(n11264), .ZN(n10478) );
  NAND2_X1 U13080 ( .A1(n11264), .A2(n11426), .ZN(n11655) );
  INV_X1 U13081 ( .A(n11655), .ZN(n10477) );
  AOI211_X1 U13082 ( .C1(n13218), .C2(n10478), .A(n13926), .B(n10477), .ZN(
        n11428) );
  AOI21_X1 U13083 ( .B1(n15377), .B2(n13218), .A(n11428), .ZN(n10487) );
  NAND2_X1 U13084 ( .A1(n10479), .A2(n10017), .ZN(n10480) );
  NAND2_X1 U13085 ( .A1(n10482), .A2(n15361), .ZN(n10483) );
  XNOR2_X1 U13086 ( .A(n11031), .B(n11030), .ZN(n10486) );
  INV_X1 U13087 ( .A(n10484), .ZN(n10485) );
  AOI21_X1 U13088 ( .B1(n10486), .B2(n13905), .A(n10485), .ZN(n11429) );
  OAI211_X1 U13089 ( .C1(n15381), .C2(n11433), .A(n10487), .B(n11429), .ZN(
        n10490) );
  NAND2_X1 U13090 ( .A1(n10490), .A2(n15384), .ZN(n10488) );
  OAI21_X1 U13091 ( .B1(n15384), .B2(n10489), .A(n10488), .ZN(P2_U3439) );
  NAND2_X1 U13092 ( .A1(n10490), .A2(n15390), .ZN(n10491) );
  OAI21_X1 U13093 ( .B1(n15390), .B2(n8767), .A(n10491), .ZN(P2_U3502) );
  INV_X1 U13094 ( .A(n11667), .ZN(n11511) );
  INV_X1 U13095 ( .A(n10492), .ZN(n10493) );
  OAI222_X1 U13096 ( .A1(P2_U3088), .A2(n11511), .B1(n14092), .B2(n10493), 
        .C1(n15545), .C2(n14097), .ZN(P2_U3312) );
  INV_X1 U13097 ( .A(n11921), .ZN(n11929) );
  OAI222_X1 U13098 ( .A1(n15105), .A2(n10494), .B1(n10976), .B2(n10493), .C1(
        n11929), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13099 ( .A(n10495), .ZN(n10498) );
  INV_X1 U13100 ( .A(n14612), .ZN(n14610) );
  OAI222_X1 U13101 ( .A1(n15105), .A2(n10496), .B1(n10976), .B2(n10498), .C1(
        n14610), .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U13102 ( .A1(P2_U3088), .A2(n6808), .B1(n14092), .B2(n10498), .C1(
        n10497), .C2(n14097), .ZN(P2_U3310) );
  NAND3_X1 U13103 ( .A1(n12663), .A2(n12543), .A3(n12705), .ZN(n10505) );
  OAI21_X1 U13104 ( .B1(n10501), .B2(n10500), .A(n10499), .ZN(n10504) );
  INV_X1 U13105 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10580) );
  OAI22_X1 U13106 ( .A1(n12655), .A2(n10502), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10580), .ZN(n10503) );
  AOI21_X1 U13107 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(n10506) );
  OAI21_X1 U13108 ( .B1(n10507), .B2(n12697), .A(n10506), .ZN(P3_U3182) );
  AND2_X1 U13109 ( .A1(n10508), .A2(n15418), .ZN(n10510) );
  NOR2_X1 U13110 ( .A1(n10809), .A2(n12048), .ZN(n10509) );
  AOI21_X1 U13111 ( .B1(n10578), .B2(n10510), .A(n10509), .ZN(n10820) );
  INV_X1 U13112 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10511) );
  MUX2_X1 U13113 ( .A(n10820), .B(n10511), .S(n15429), .Z(n10512) );
  OAI21_X1 U13114 ( .B1(n10823), .B2(n12949), .A(n10512), .ZN(P3_U3390) );
  NAND2_X1 U13115 ( .A1(n10516), .A2(n10515), .ZN(n10585) );
  OAI21_X1 U13116 ( .B1(n10516), .B2(n10515), .A(n10585), .ZN(n10526) );
  INV_X1 U13117 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10517) );
  MUX2_X1 U13118 ( .A(n10517), .B(P3_REG1_REG_2__SCAN_IN), .S(n10590), .Z(
        n10521) );
  OAI21_X1 U13119 ( .B1(n10519), .B2(n10518), .A(n7831), .ZN(n10520) );
  OAI21_X1 U13120 ( .B1(n10521), .B2(n10520), .A(n10592), .ZN(n10522) );
  AND2_X1 U13121 ( .A1(n12707), .A2(n10522), .ZN(n10525) );
  INV_X1 U13122 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10523) );
  INV_X1 U13123 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n12890) );
  OAI22_X1 U13124 ( .A1(n12655), .A2(n10523), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12890), .ZN(n10524) );
  AOI211_X1 U13125 ( .C1(n12688), .C2(n10526), .A(n10525), .B(n10524), .ZN(
        n10533) );
  AOI22_X1 U13126 ( .A1(n10530), .A2(n10529), .B1(n10528), .B2(n10527), .ZN(
        n10582) );
  XNOR2_X1 U13127 ( .A(n10582), .B(n10581), .ZN(n10531) );
  NAND2_X1 U13128 ( .A1(n12584), .A2(n10531), .ZN(n10532) );
  OAI211_X1 U13129 ( .C1(n12697), .C2(n6909), .A(n10533), .B(n10532), .ZN(
        P3_U3184) );
  AOI211_X1 U13130 ( .C1(n10535), .C2(n10534), .A(n13457), .B(n15300), .ZN(
        n10540) );
  INV_X1 U13131 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10916) );
  INV_X1 U13132 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10537) );
  MUX2_X1 U13133 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10211), .S(n10541), .Z(
        n10536) );
  OAI21_X1 U13134 ( .B1(n10916), .B2(n10537), .A(n10536), .ZN(n10538) );
  AND3_X1 U13135 ( .A1(n15318), .A2(n13460), .A3(n10538), .ZN(n10539) );
  NOR2_X1 U13136 ( .A1(n10540), .A2(n10539), .ZN(n10544) );
  INV_X1 U13137 ( .A(n10541), .ZN(n10542) );
  AOI22_X1 U13138 ( .A1(n15305), .A2(n10542), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10543) );
  OAI211_X1 U13139 ( .C1(n15498), .C2(n15322), .A(n10544), .B(n10543), .ZN(
        P2_U3215) );
  INV_X1 U13140 ( .A(n12653), .ZN(n12646) );
  INV_X1 U13141 ( .A(n10545), .ZN(n10547) );
  OAI222_X1 U13142 ( .A1(n12646), .A2(P3_U3151), .B1(n13039), .B2(n10547), 
        .C1(n10546), .C2(n13034), .ZN(P3_U3279) );
  INV_X1 U13143 ( .A(n12576), .ZN(n12590) );
  INV_X1 U13144 ( .A(n10548), .ZN(n10550) );
  OAI222_X1 U13145 ( .A1(n12590), .A2(P3_U3151), .B1(n13039), .B2(n10550), 
        .C1(n10549), .C2(n13034), .ZN(P3_U3281) );
  NAND2_X1 U13146 ( .A1(n13183), .A2(n13452), .ZN(n10551) );
  MUX2_X1 U13147 ( .A(n10551), .B(n13194), .S(n13200), .Z(n10555) );
  INV_X1 U13148 ( .A(n10552), .ZN(n10553) );
  AOI22_X1 U13149 ( .A1(n13053), .A2(n13450), .B1(n13182), .B2(n10553), .ZN(
        n10554) );
  OAI211_X1 U13150 ( .C1(n10556), .C2(n8721), .A(n10555), .B(n10554), .ZN(
        P2_U3204) );
  NAND2_X1 U13151 ( .A1(n10569), .A2(n10565), .ZN(n10561) );
  AND3_X1 U13152 ( .A1(n10559), .A2(n10558), .A3(n10557), .ZN(n10560) );
  OAI211_X1 U13153 ( .C1(n10808), .C2(n10566), .A(n10561), .B(n10560), .ZN(
        n10562) );
  NAND2_X1 U13154 ( .A1(n10562), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10564) );
  INV_X1 U13155 ( .A(n10808), .ZN(n10567) );
  NAND2_X1 U13156 ( .A1(n10807), .A2(n10567), .ZN(n10563) );
  NOR2_X1 U13157 ( .A1(n12502), .A2(P3_U3151), .ZN(n10899) );
  NAND2_X1 U13158 ( .A1(n10565), .A2(n15418), .ZN(n10568) );
  OAI22_X1 U13159 ( .A1(n10569), .A2(n10568), .B1(n10567), .B2(n10566), .ZN(
        n10570) );
  INV_X1 U13160 ( .A(n12506), .ZN(n12436) );
  NOR2_X1 U13161 ( .A1(n10571), .A2(n15418), .ZN(n10572) );
  NAND2_X1 U13162 ( .A1(n10573), .A2(n10572), .ZN(n10575) );
  OAI22_X1 U13163 ( .A1(n12451), .A2(n10823), .B1(n12488), .B2(n10809), .ZN(
        n10577) );
  AOI21_X1 U13164 ( .B1(n12436), .B2(n10578), .A(n10577), .ZN(n10579) );
  OAI21_X1 U13165 ( .B1(n10899), .B2(n10580), .A(n10579), .ZN(P3_U3172) );
  MUX2_X1 U13166 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13031), .Z(n10600) );
  XOR2_X1 U13167 ( .A(n10607), .B(n10600), .Z(n10603) );
  XOR2_X1 U13168 ( .A(n10603), .B(n10604), .Z(n10599) );
  INV_X1 U13169 ( .A(n10607), .ZN(n10602) );
  INV_X1 U13170 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10583) );
  OR2_X1 U13171 ( .A1(n10590), .A2(n10583), .ZN(n10584) );
  NAND2_X1 U13172 ( .A1(n10585), .A2(n10584), .ZN(n10586) );
  INV_X1 U13173 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U13174 ( .A1(n10587), .A2(n10997), .ZN(n10588) );
  NAND2_X1 U13175 ( .A1(n10731), .A2(n10588), .ZN(n10589) );
  NAND2_X1 U13176 ( .A1(n12688), .A2(n10589), .ZN(n10596) );
  OR2_X1 U13177 ( .A1(n10590), .A2(n10517), .ZN(n10591) );
  NAND2_X1 U13178 ( .A1(n10592), .A2(n10591), .ZN(n10608) );
  XNOR2_X1 U13179 ( .A(n10606), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10593) );
  NAND2_X1 U13180 ( .A1(n12707), .A2(n10593), .ZN(n10595) );
  NOR2_X1 U13181 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8052), .ZN(n10952) );
  AOI21_X1 U13182 ( .B1(n15391), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10952), .ZN(
        n10594) );
  NAND3_X1 U13183 ( .A1(n10596), .A2(n10595), .A3(n10594), .ZN(n10597) );
  AOI21_X1 U13184 ( .B1(n10602), .B2(n12661), .A(n10597), .ZN(n10598) );
  OAI21_X1 U13185 ( .B1(n10599), .B2(n12705), .A(n10598), .ZN(P3_U3185) );
  XOR2_X1 U13186 ( .A(n10625), .B(n10631), .Z(n10634) );
  INV_X1 U13187 ( .A(n10600), .ZN(n10601) );
  AOI22_X1 U13188 ( .A1(n10604), .A2(n10603), .B1(n10602), .B2(n10601), .ZN(
        n10723) );
  MUX2_X1 U13189 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13031), .Z(n10605) );
  XNOR2_X1 U13190 ( .A(n10605), .B(n10727), .ZN(n10724) );
  XOR2_X1 U13191 ( .A(n10634), .B(n10635), .Z(n10623) );
  NAND2_X1 U13192 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  INV_X1 U13193 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10610) );
  MUX2_X1 U13194 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10610), .S(n10727), .Z(
        n10725) );
  INV_X1 U13195 ( .A(n10625), .ZN(n10633) );
  XNOR2_X1 U13196 ( .A(n10626), .B(n10633), .ZN(n10624) );
  XNOR2_X1 U13197 ( .A(n10624), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13198 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11184) );
  INV_X1 U13199 ( .A(n11184), .ZN(n10611) );
  AOI21_X1 U13200 ( .B1(n15391), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10611), .ZN(
        n10619) );
  INV_X1 U13201 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10991) );
  XNOR2_X1 U13202 ( .A(n10727), .B(n10991), .ZN(n10728) );
  NAND2_X1 U13203 ( .A1(n10727), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13204 ( .A1(n10733), .A2(n10613), .ZN(n10614) );
  NAND2_X1 U13205 ( .A1(n10614), .A2(n10625), .ZN(n10649) );
  OAI21_X1 U13206 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n10616), .A(n10651), .ZN(
        n10617) );
  NAND2_X1 U13207 ( .A1(n12688), .A2(n10617), .ZN(n10618) );
  OAI211_X1 U13208 ( .C1(n12697), .C2(n10625), .A(n10619), .B(n10618), .ZN(
        n10620) );
  AOI21_X1 U13209 ( .B1(n12707), .B2(n10621), .A(n10620), .ZN(n10622) );
  OAI21_X1 U13210 ( .B1(n10623), .B2(n12705), .A(n10622), .ZN(P3_U3187) );
  NAND2_X1 U13211 ( .A1(n10624), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13212 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  INV_X1 U13213 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10629) );
  MUX2_X1 U13214 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10629), .S(n10655), .Z(
        n10647) );
  NAND2_X1 U13215 ( .A1(n10655), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10630) );
  XOR2_X1 U13216 ( .A(n10870), .B(P3_REG1_REG_7__SCAN_IN), .Z(n10644) );
  MUX2_X1 U13217 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13031), .Z(n10636) );
  XNOR2_X1 U13218 ( .A(n10636), .B(n10655), .ZN(n10646) );
  MUX2_X1 U13219 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13031), .Z(n10875) );
  XNOR2_X1 U13220 ( .A(n10875), .B(n10877), .ZN(n10878) );
  XNOR2_X1 U13221 ( .A(n10879), .B(n10878), .ZN(n10642) );
  XNOR2_X1 U13222 ( .A(n10655), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n10650) );
  OAI21_X1 U13223 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n10637), .A(n10884), .ZN(
        n10638) );
  NAND2_X1 U13224 ( .A1(n10638), .A2(n12688), .ZN(n10640) );
  AND2_X1 U13225 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11474) );
  AOI21_X1 U13226 ( .B1(n15391), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11474), .ZN(
        n10639) );
  OAI211_X1 U13227 ( .C1(n12697), .C2(n10871), .A(n10640), .B(n10639), .ZN(
        n10641) );
  AOI21_X1 U13228 ( .B1(n12584), .B2(n10642), .A(n10641), .ZN(n10643) );
  OAI21_X1 U13229 ( .B1(n10644), .B2(n12543), .A(n10643), .ZN(P3_U3189) );
  XOR2_X1 U13230 ( .A(n10646), .B(n10645), .Z(n10659) );
  XNOR2_X1 U13231 ( .A(n10648), .B(n10647), .ZN(n10657) );
  AND3_X1 U13232 ( .A1(n10651), .A2(n10650), .A3(n10649), .ZN(n10652) );
  OAI21_X1 U13233 ( .B1(n6634), .B2(n10652), .A(n12688), .ZN(n10654) );
  AND2_X1 U13234 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n11292) );
  AOI21_X1 U13235 ( .B1(n15391), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11292), .ZN(
        n10653) );
  OAI211_X1 U13236 ( .C1(n12697), .C2(n10655), .A(n10654), .B(n10653), .ZN(
        n10656) );
  AOI21_X1 U13237 ( .B1(n12707), .B2(n10657), .A(n10656), .ZN(n10658) );
  OAI21_X1 U13238 ( .B1(n10659), .B2(n12705), .A(n10658), .ZN(P3_U3188) );
  XNOR2_X1 U13239 ( .A(n10714), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10708) );
  XNOR2_X1 U13240 ( .A(n10965), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10957) );
  XNOR2_X1 U13241 ( .A(n6477), .B(n10957), .ZN(n10677) );
  NAND2_X1 U13242 ( .A1(n15305), .A2(n10965), .ZN(n10662) );
  NAND2_X1 U13243 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11605)
         );
  NAND2_X1 U13244 ( .A1(n10662), .A2(n11605), .ZN(n10675) );
  OR2_X1 U13245 ( .A1(n10663), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10664) );
  INV_X1 U13246 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10666) );
  MUX2_X1 U13247 ( .A(n10666), .B(P2_REG2_REG_10__SCAN_IN), .S(n10714), .Z(
        n10703) );
  NAND2_X1 U13248 ( .A1(n10714), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10667) );
  INV_X1 U13249 ( .A(n10672), .ZN(n10670) );
  INV_X1 U13250 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10668) );
  MUX2_X1 U13251 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10668), .S(n10965), .Z(
        n10671) );
  INV_X1 U13252 ( .A(n10671), .ZN(n10669) );
  NAND2_X1 U13253 ( .A1(n10670), .A2(n10669), .ZN(n10673) );
  NAND2_X1 U13254 ( .A1(n10672), .A2(n10671), .ZN(n15293) );
  AOI21_X1 U13255 ( .B1(n10673), .B2(n15293), .A(n15294), .ZN(n10674) );
  AOI211_X1 U13256 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n15273), .A(n10675), 
        .B(n10674), .ZN(n10676) );
  OAI21_X1 U13257 ( .B1(n10677), .B2(n15300), .A(n10676), .ZN(P2_U3225) );
  OAI21_X1 U13258 ( .B1(n10680), .B2(n10679), .A(n10678), .ZN(n10687) );
  INV_X1 U13259 ( .A(n10680), .ZN(n10682) );
  NAND3_X1 U13260 ( .A1(n13183), .A2(n10682), .A3(n10681), .ZN(n10683) );
  INV_X1 U13261 ( .A(n13448), .ZN(n11032) );
  AOI21_X1 U13262 ( .B1(n10683), .B2(n13143), .A(n11032), .ZN(n10686) );
  INV_X1 U13263 ( .A(n15368), .ZN(n11658) );
  AOI22_X1 U13264 ( .A1(n13053), .A2(n13446), .B1(n13170), .B2(n11656), .ZN(
        n10684) );
  NAND2_X1 U13265 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15274) );
  OAI211_X1 U13266 ( .C1(n11658), .C2(n13194), .A(n10684), .B(n15274), .ZN(
        n10685) );
  AOI211_X1 U13267 ( .C1(n13182), .C2(n10687), .A(n10686), .B(n10685), .ZN(
        n10688) );
  INV_X1 U13268 ( .A(n10688), .ZN(P2_U3202) );
  INV_X1 U13269 ( .A(n10689), .ZN(n10692) );
  MUX2_X1 U13270 ( .A(n10692), .B(n10691), .S(n10690), .Z(n10693) );
  MUX2_X1 U13271 ( .A(n10695), .B(n10820), .S(n12896), .Z(n10701) );
  INV_X1 U13272 ( .A(n10696), .ZN(n10698) );
  NOR2_X1 U13273 ( .A1(n12889), .A2(n15418), .ZN(n10697) );
  AOI22_X1 U13274 ( .A1(n12855), .A2(n10699), .B1(n12873), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10700) );
  NAND2_X1 U13275 ( .A1(n10701), .A2(n10700), .ZN(P3_U3233) );
  INV_X1 U13276 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11591) );
  NAND2_X1 U13277 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11581)
         );
  INV_X1 U13278 ( .A(n11581), .ZN(n10713) );
  AOI21_X1 U13279 ( .B1(n10703), .B2(n10702), .A(n15294), .ZN(n10705) );
  NAND2_X1 U13280 ( .A1(n10705), .A2(n10704), .ZN(n10711) );
  AOI211_X1 U13281 ( .C1(n10708), .C2(n10707), .A(n10706), .B(n15300), .ZN(
        n10709) );
  INV_X1 U13282 ( .A(n10709), .ZN(n10710) );
  NAND2_X1 U13283 ( .A1(n10711), .A2(n10710), .ZN(n10712) );
  AOI211_X1 U13284 ( .C1(n15305), .C2(n10714), .A(n10713), .B(n10712), .ZN(
        n10715) );
  OAI21_X1 U13285 ( .B1(n15322), .B2(n11591), .A(n10715), .ZN(P2_U3224) );
  NAND2_X1 U13286 ( .A1(n10716), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13287 ( .A1(n10719), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10722) );
  INV_X1 U13288 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U13289 ( .A1(n10720), .A2(n15475), .ZN(n10721) );
  NAND2_X1 U13290 ( .A1(n10722), .A2(n10721), .ZN(n11166) );
  XNOR2_X1 U13291 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n11165) );
  XNOR2_X1 U13292 ( .A(n11166), .B(n11165), .ZN(n11161) );
  XNOR2_X1 U13293 ( .A(n11160), .B(n11159), .ZN(SUB_1596_U55) );
  XOR2_X1 U13294 ( .A(n10724), .B(n10723), .Z(n10740) );
  XNOR2_X1 U13295 ( .A(n10726), .B(n10725), .ZN(n10738) );
  NOR2_X1 U13296 ( .A1(n12697), .A2(n10727), .ZN(n10737) );
  INV_X1 U13297 ( .A(n10728), .ZN(n10730) );
  NAND3_X1 U13298 ( .A1(n10731), .A2(n10730), .A3(n10729), .ZN(n10732) );
  NAND2_X1 U13299 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U13300 ( .A1(n12688), .A2(n10734), .ZN(n10735) );
  NAND2_X1 U13301 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n11022) );
  OAI211_X1 U13302 ( .C1(n10071), .C2(n12655), .A(n10735), .B(n11022), .ZN(
        n10736) );
  AOI211_X1 U13303 ( .C1(n12707), .C2(n10738), .A(n10737), .B(n10736), .ZN(
        n10739) );
  OAI21_X1 U13304 ( .B1(n10740), .B2(n12705), .A(n10739), .ZN(P3_U3186) );
  XOR2_X1 U13305 ( .A(n10742), .B(n11355), .Z(n10862) );
  XOR2_X1 U13306 ( .A(n10857), .B(n10862), .Z(n10749) );
  OAI22_X1 U13307 ( .A1(n12298), .A2(n10837), .B1(n10758), .B2(n7769), .ZN(
        n10743) );
  MUX2_X1 U13308 ( .A(n10855), .B(n12313), .S(n10783), .Z(n10748) );
  XNOR2_X1 U13309 ( .A(n10749), .B(n10748), .ZN(n10766) );
  OR2_X1 U13310 ( .A1(n10751), .A2(n10750), .ZN(n10756) );
  INV_X1 U13311 ( .A(n10756), .ZN(n10760) );
  NAND2_X1 U13312 ( .A1(n10752), .A2(n14432), .ZN(n10753) );
  NOR2_X1 U13313 ( .A1(n15255), .A2(n10753), .ZN(n10754) );
  NAND2_X1 U13314 ( .A1(n10756), .A2(n10755), .ZN(n10762) );
  AND2_X1 U13315 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  NAND2_X1 U13316 ( .A1(n10762), .A2(n10759), .ZN(n11370) );
  INV_X1 U13317 ( .A(n14499), .ZN(n10787) );
  INV_X1 U13318 ( .A(n14239), .ZN(n14216) );
  NAND2_X1 U13319 ( .A1(n10762), .A2(n10761), .ZN(n10864) );
  AOI22_X1 U13320 ( .A1(n14218), .A2(n14265), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10864), .ZN(n10763) );
  OAI21_X1 U13321 ( .B1(n10787), .B2(n14216), .A(n10763), .ZN(n10764) );
  AOI21_X1 U13322 ( .B1(n14221), .B2(n14970), .A(n10764), .ZN(n10765) );
  OAI21_X1 U13323 ( .B1(n10766), .B2(n15174), .A(n10765), .ZN(P1_U3222) );
  INV_X1 U13324 ( .A(n10767), .ZN(n10768) );
  NOR2_X1 U13325 ( .A1(n10769), .A2(n10768), .ZN(n10771) );
  XNOR2_X1 U13326 ( .A(n11238), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10770) );
  AOI21_X1 U13327 ( .B1(n10771), .B2(n10770), .A(n14580), .ZN(n10782) );
  INV_X1 U13328 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U13329 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14146)
         );
  OAI21_X1 U13330 ( .B1(n14583), .B2(n15510), .A(n14146), .ZN(n10780) );
  XNOR2_X1 U13331 ( .A(n11238), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n10777) );
  OR2_X1 U13332 ( .A1(n10773), .A2(n10772), .ZN(n10774) );
  NAND2_X1 U13333 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  NOR2_X1 U13334 ( .A1(n10776), .A2(n10777), .ZN(n11231) );
  AOI21_X1 U13335 ( .B1(n10777), .B2(n10776), .A(n11231), .ZN(n10778) );
  NOR2_X1 U13336 ( .A1(n10778), .A2(n14637), .ZN(n10779) );
  AOI211_X1 U13337 ( .C1(n15197), .C2(n11238), .A(n10780), .B(n10779), .ZN(
        n10781) );
  OAI21_X1 U13338 ( .B1(n10782), .B2(n14635), .A(n10781), .ZN(P1_U3255) );
  XNOR2_X1 U13339 ( .A(n10855), .B(n10783), .ZN(n14509) );
  AOI22_X1 U13340 ( .A1(n14218), .A2(n14498), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10864), .ZN(n10785) );
  NAND2_X1 U13341 ( .A1(n14221), .A2(n14972), .ZN(n10784) );
  OAI211_X1 U13342 ( .C1(n14509), .C2(n15174), .A(n10785), .B(n10784), .ZN(
        P1_U3232) );
  INV_X1 U13343 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10794) );
  INV_X1 U13344 ( .A(n10786), .ZN(n10792) );
  NAND2_X1 U13345 ( .A1(n10787), .A2(n10837), .ZN(n10788) );
  NAND2_X1 U13346 ( .A1(n10843), .A2(n10788), .ZN(n14438) );
  AND2_X1 U13347 ( .A1(n15247), .A2(n15050), .ZN(n10789) );
  OR2_X1 U13348 ( .A1(n14438), .A2(n10789), .ZN(n10791) );
  NAND2_X1 U13349 ( .A1(n14897), .A2(n14498), .ZN(n10790) );
  AND2_X1 U13350 ( .A1(n10791), .A2(n10790), .ZN(n14977) );
  OAI21_X1 U13351 ( .B1(n10837), .B2(n10792), .A(n14977), .ZN(n15082) );
  NAND2_X1 U13352 ( .A1(n15082), .A2(n15265), .ZN(n10793) );
  OAI21_X1 U13353 ( .B1(n15265), .B2(n10794), .A(n10793), .ZN(P1_U3459) );
  OAI21_X1 U13354 ( .B1(n12696), .B2(n10983), .A(n11134), .ZN(n10797) );
  INV_X1 U13355 ( .A(n10800), .ZN(n10799) );
  XNOR2_X1 U13356 ( .A(n10800), .B(n12888), .ZN(n10943) );
  XNOR2_X1 U13357 ( .A(n10943), .B(n12522), .ZN(n10944) );
  NAND2_X1 U13358 ( .A1(n10799), .A2(n11006), .ZN(n10804) );
  NAND2_X1 U13359 ( .A1(n7223), .A2(n10902), .ZN(n10803) );
  OAI21_X1 U13360 ( .B1(n10800), .B2(n10803), .A(n10805), .ZN(n10895) );
  XOR2_X1 U13361 ( .A(n10944), .B(n10945), .Z(n10814) );
  NAND3_X1 U13362 ( .A1(n10808), .A2(n10807), .A3(n10806), .ZN(n12499) );
  OAI22_X1 U13363 ( .A1(n12488), .A2(n11023), .B1(n10809), .B2(n12499), .ZN(
        n10811) );
  NOR2_X1 U13364 ( .A1(n10899), .A2(n12890), .ZN(n10810) );
  AOI211_X1 U13365 ( .C1(n10812), .C2(n12503), .A(n10811), .B(n10810), .ZN(
        n10813) );
  OAI21_X1 U13366 ( .B1(n10814), .B2(n12506), .A(n10813), .ZN(P3_U3177) );
  AOI222_X1 U13367 ( .A1(n12666), .A2(P3_STATE_REG_SCAN_IN), .B1(n10817), .B2(
        n10816), .C1(n10815), .C2(n13016), .ZN(P3_U3278) );
  INV_X1 U13368 ( .A(n12702), .ZN(n12690) );
  OAI222_X1 U13369 ( .A1(P3_U3151), .A2(n12690), .B1(n13034), .B2(n10819), 
        .C1(n13039), .C2(n10818), .ZN(P3_U3277) );
  MUX2_X1 U13370 ( .A(n10821), .B(n10820), .S(n15589), .Z(n10822) );
  OAI21_X1 U13371 ( .B1(n12905), .B2(n10823), .A(n10822), .ZN(P3_U3459) );
  XNOR2_X1 U13372 ( .A(n10825), .B(n10824), .ZN(n10831) );
  NAND2_X1 U13373 ( .A1(n10826), .A2(n10831), .ZN(n10918) );
  INV_X1 U13374 ( .A(n8816), .ZN(n11409) );
  NAND2_X1 U13375 ( .A1(n13445), .A2(n13885), .ZN(n10828) );
  NAND2_X1 U13376 ( .A1(n13447), .A2(n13883), .ZN(n10827) );
  NAND2_X1 U13377 ( .A1(n10828), .A2(n10827), .ZN(n11036) );
  NAND2_X1 U13378 ( .A1(n13161), .A2(n11036), .ZN(n10829) );
  NAND2_X1 U13379 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13484) );
  OAI211_X1 U13380 ( .C1(n13194), .C2(n11409), .A(n10829), .B(n13484), .ZN(
        n10835) );
  INV_X1 U13381 ( .A(n10678), .ZN(n10833) );
  AOI22_X1 U13382 ( .A1(n13183), .A2(n13447), .B1(n13182), .B2(n10830), .ZN(
        n10832) );
  NOR3_X1 U13383 ( .A1(n10833), .A2(n10832), .A3(n10831), .ZN(n10834) );
  AOI211_X1 U13384 ( .C1(n13170), .C2(n11276), .A(n10835), .B(n10834), .ZN(
        n10836) );
  OAI21_X1 U13385 ( .B1(n13165), .B2(n10918), .A(n10836), .ZN(P2_U3199) );
  INV_X1 U13386 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10852) );
  OR2_X1 U13387 ( .A1(n14260), .A2(n10837), .ZN(n10838) );
  NAND2_X1 U13388 ( .A1(n10838), .A2(n11045), .ZN(n14965) );
  XNOR2_X1 U13389 ( .A(n14258), .B(n14965), .ZN(n10841) );
  NAND2_X1 U13390 ( .A1(n10840), .A2(n10839), .ZN(n14437) );
  MUX2_X1 U13391 ( .A(n10841), .B(n14437), .S(n14499), .Z(n10849) );
  AOI22_X1 U13392 ( .A1(n14265), .A2(n14897), .B1(n14880), .B2(n14499), .ZN(
        n10848) );
  NAND2_X1 U13393 ( .A1(n14437), .A2(n10844), .ZN(n10845) );
  NAND2_X1 U13394 ( .A1(n10842), .A2(n10845), .ZN(n10846) );
  NAND2_X1 U13395 ( .A1(n10846), .A2(n15263), .ZN(n10847) );
  OAI211_X1 U13396 ( .C1(n10849), .C2(n15050), .A(n10848), .B(n10847), .ZN(
        n14967) );
  OAI22_X1 U13397 ( .A1(n15259), .A2(n14260), .B1(n14929), .B2(n14965), .ZN(
        n10850) );
  OR2_X1 U13398 ( .A1(n14967), .A2(n10850), .ZN(n10853) );
  NAND2_X1 U13399 ( .A1(n10853), .A2(n15265), .ZN(n10851) );
  OAI21_X1 U13400 ( .B1(n15265), .B2(n10852), .A(n10851), .ZN(P1_U3462) );
  NAND2_X1 U13401 ( .A1(n10853), .A2(n15272), .ZN(n10854) );
  OAI21_X1 U13402 ( .B1(n15272), .B2(n10246), .A(n10854), .ZN(P1_U3529) );
  NAND2_X1 U13403 ( .A1(n10856), .A2(n10855), .ZN(n10859) );
  NAND3_X1 U13404 ( .A1(n10858), .A2(n10859), .A3(n10857), .ZN(n10861) );
  OAI22_X1 U13405 ( .A1(n9741), .A2(n6402), .B1(n14268), .B2(n12273), .ZN(
        n10863) );
  XNOR2_X1 U13406 ( .A(n10863), .B(n11355), .ZN(n11337) );
  OAI22_X1 U13407 ( .A1(n9741), .A2(n11341), .B1(n14268), .B2(n6402), .ZN(
        n11336) );
  XNOR2_X1 U13408 ( .A(n11337), .B(n11336), .ZN(n11338) );
  XOR2_X1 U13409 ( .A(n11339), .B(n11338), .Z(n10868) );
  AOI22_X1 U13410 ( .A1(n14218), .A2(n14497), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10864), .ZN(n10865) );
  OAI21_X1 U13411 ( .B1(n14258), .B2(n14216), .A(n10865), .ZN(n10866) );
  AOI21_X1 U13412 ( .B1(n14221), .B2(n7193), .A(n10866), .ZN(n10867) );
  OAI21_X1 U13413 ( .B1(n10868), .B2(n15174), .A(n10867), .ZN(P1_U3237) );
  INV_X1 U13414 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10869) );
  MUX2_X1 U13415 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10869), .S(n11144), .Z(
        n11135) );
  NAND2_X1 U13416 ( .A1(n10872), .A2(n10871), .ZN(n10873) );
  NAND2_X1 U13417 ( .A1(n10874), .A2(n10873), .ZN(n11136) );
  XOR2_X1 U13418 ( .A(n11135), .B(n11136), .Z(n10891) );
  INV_X1 U13419 ( .A(n10875), .ZN(n10876) );
  MUX2_X1 U13420 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13031), .Z(n11145) );
  XNOR2_X1 U13421 ( .A(n11144), .B(n11145), .ZN(n11146) );
  XNOR2_X1 U13422 ( .A(n11147), .B(n11146), .ZN(n10889) );
  INV_X1 U13423 ( .A(n10881), .ZN(n10882) );
  XNOR2_X1 U13424 ( .A(n11144), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n10883) );
  AND3_X1 U13425 ( .A1(n10884), .A2(n10883), .A3(n10882), .ZN(n10885) );
  OAI21_X1 U13426 ( .B1(n11138), .B2(n10885), .A(n12688), .ZN(n10887) );
  AND2_X1 U13427 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11684) );
  AOI21_X1 U13428 ( .B1(n15391), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11684), .ZN(
        n10886) );
  OAI211_X1 U13429 ( .C1(n12697), .C2(n11144), .A(n10887), .B(n10886), .ZN(
        n10888) );
  AOI21_X1 U13430 ( .B1(n12584), .B2(n10889), .A(n10888), .ZN(n10890) );
  OAI21_X1 U13431 ( .B1(n10891), .B2(n12543), .A(n10890), .ZN(P3_U3190) );
  INV_X1 U13432 ( .A(n11006), .ZN(n10896) );
  INV_X1 U13433 ( .A(n11007), .ZN(n10892) );
  NOR3_X1 U13434 ( .A1(n10799), .A2(n10892), .A3(n11004), .ZN(n10894) );
  AOI211_X1 U13435 ( .C1(n10896), .C2(n10895), .A(n10894), .B(n10893), .ZN(
        n10904) );
  INV_X1 U13436 ( .A(n12523), .ZN(n10897) );
  OAI22_X1 U13437 ( .A1(n12488), .A2(n10949), .B1(n10897), .B2(n12499), .ZN(
        n10901) );
  INV_X1 U13438 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10898) );
  NOR2_X1 U13439 ( .A1(n10899), .A2(n10898), .ZN(n10900) );
  AOI211_X1 U13440 ( .C1(n10902), .C2(n12503), .A(n10901), .B(n10900), .ZN(
        n10903) );
  OAI21_X1 U13441 ( .B1(n10904), .B2(n12506), .A(n10903), .ZN(P3_U3162) );
  INV_X1 U13442 ( .A(n13374), .ZN(n13419) );
  NAND2_X1 U13443 ( .A1(n13200), .A2(n10905), .ZN(n14055) );
  NAND2_X1 U13444 ( .A1(n13452), .A2(n10906), .ZN(n10907) );
  AND2_X1 U13445 ( .A1(n10908), .A2(n10907), .ZN(n14057) );
  AOI21_X1 U13446 ( .B1(n13920), .B2(n10909), .A(n14057), .ZN(n10910) );
  AOI21_X1 U13447 ( .B1(n13885), .B2(n13450), .A(n10910), .ZN(n14056) );
  OAI21_X1 U13448 ( .B1(n13419), .B2(n14055), .A(n14056), .ZN(n10911) );
  INV_X1 U13449 ( .A(n13837), .ZN(n13928) );
  AOI22_X1 U13450 ( .A1(n10911), .A2(n13880), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13928), .ZN(n10915) );
  INV_X1 U13451 ( .A(n13811), .ZN(n10913) );
  INV_X1 U13452 ( .A(n14057), .ZN(n10912) );
  NAND2_X1 U13453 ( .A1(n10913), .A2(n10912), .ZN(n10914) );
  OAI211_X1 U13454 ( .C1(n10916), .C2(n13880), .A(n10915), .B(n10914), .ZN(
        P2_U3265) );
  AND2_X1 U13455 ( .A1(n10918), .A2(n10917), .ZN(n10922) );
  AND2_X1 U13456 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  NAND2_X1 U13457 ( .A1(n10922), .A2(n10921), .ZN(n11104) );
  OAI211_X1 U13458 ( .C1(n10922), .C2(n10921), .A(n11104), .B(n13182), .ZN(
        n10928) );
  NAND2_X1 U13459 ( .A1(n13444), .A2(n13885), .ZN(n10924) );
  NAND2_X1 U13460 ( .A1(n13446), .A2(n13883), .ZN(n10923) );
  NAND2_X1 U13461 ( .A1(n10924), .A2(n10923), .ZN(n11083) );
  NAND2_X1 U13462 ( .A1(n13161), .A2(n11083), .ZN(n10925) );
  NAND2_X1 U13463 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13507) );
  OAI211_X1 U13464 ( .C1(n13194), .C2(n11637), .A(n10925), .B(n13507), .ZN(
        n10926) );
  AOI21_X1 U13465 ( .B1(n11635), .B2(n13170), .A(n10926), .ZN(n10927) );
  NAND2_X1 U13466 ( .A1(n10928), .A2(n10927), .ZN(P2_U3211) );
  OAI21_X1 U13467 ( .B1(n10931), .B2(n10930), .A(n10929), .ZN(n10941) );
  NOR2_X1 U13468 ( .A1(n10950), .A2(n15418), .ZN(n10940) );
  INV_X1 U13469 ( .A(n10941), .ZN(n11001) );
  INV_X1 U13470 ( .A(n11777), .ZN(n12887) );
  AOI22_X1 U13471 ( .A1(n12879), .A2(n12521), .B1(n12880), .B2(n12522), .ZN(
        n10939) );
  NAND2_X1 U13472 ( .A1(n10932), .A2(n12882), .ZN(n12881) );
  AND2_X1 U13473 ( .A1(n12881), .A2(n10933), .ZN(n10937) );
  INV_X1 U13474 ( .A(n10934), .ZN(n10935) );
  NAND2_X1 U13475 ( .A1(n12881), .A2(n10935), .ZN(n10985) );
  OAI211_X1 U13476 ( .C1(n10937), .C2(n10936), .A(n10985), .B(n12883), .ZN(
        n10938) );
  OAI211_X1 U13477 ( .C1(n11001), .C2(n12887), .A(n10939), .B(n10938), .ZN(
        n10995) );
  AOI211_X1 U13478 ( .C1(n15425), .C2(n10941), .A(n10940), .B(n10995), .ZN(
        n15587) );
  NAND2_X1 U13479 ( .A1(n15429), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n10942) );
  OAI21_X1 U13480 ( .B1(n15587), .B2(n15429), .A(n10942), .ZN(P3_U3399) );
  XNOR2_X1 U13481 ( .A(n10800), .B(n10998), .ZN(n11017) );
  XOR2_X1 U13482 ( .A(n12878), .B(n11017), .Z(n10947) );
  AOI211_X1 U13483 ( .C1(n10947), .C2(n10946), .A(n12506), .B(n6453), .ZN(
        n10948) );
  INV_X1 U13484 ( .A(n10948), .ZN(n10954) );
  OAI22_X1 U13485 ( .A1(n12451), .A2(n10950), .B1(n10949), .B2(n12499), .ZN(
        n10951) );
  AOI211_X1 U13486 ( .C1(n12497), .C2(n12521), .A(n10952), .B(n10951), .ZN(
        n10953) );
  OAI211_X1 U13487 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12027), .A(n10954), .B(
        n10953), .ZN(P3_U3158) );
  INV_X1 U13488 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15111) );
  INV_X1 U13489 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10956) );
  OAI22_X1 U13490 ( .A1(n6477), .A2(n10957), .B1(n10956), .B2(n10955), .ZN(
        n15298) );
  XNOR2_X1 U13491 ( .A(n15304), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n15299) );
  NOR2_X1 U13492 ( .A1(n15304), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10959) );
  XNOR2_X1 U13493 ( .A(n11504), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n10958) );
  INV_X1 U13494 ( .A(n11499), .ZN(n10961) );
  OAI21_X1 U13495 ( .B1(n15297), .B2(n10959), .A(n10958), .ZN(n10960) );
  NAND3_X1 U13496 ( .A1(n10961), .A2(n15315), .A3(n10960), .ZN(n10964) );
  NAND2_X1 U13497 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n11766)
         );
  INV_X1 U13498 ( .A(n11766), .ZN(n10962) );
  AOI21_X1 U13499 ( .B1(n15305), .B2(n11504), .A(n10962), .ZN(n10963) );
  OAI211_X1 U13500 ( .C1(n15322), .C2(n15111), .A(n10964), .B(n10963), .ZN(
        n10974) );
  OR2_X1 U13501 ( .A1(n10965), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15291) );
  NAND2_X1 U13502 ( .A1(n15293), .A2(n15291), .ZN(n10967) );
  INV_X1 U13503 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10966) );
  MUX2_X1 U13504 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10966), .S(n15304), .Z(
        n15290) );
  NAND2_X1 U13505 ( .A1(n10967), .A2(n15290), .ZN(n15296) );
  OR2_X1 U13506 ( .A1(n15304), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10968) );
  NAND2_X1 U13507 ( .A1(n15296), .A2(n10968), .ZN(n10972) );
  INV_X1 U13508 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10969) );
  MUX2_X1 U13509 ( .A(n10969), .B(P2_REG2_REG_13__SCAN_IN), .S(n11504), .Z(
        n10971) );
  INV_X1 U13510 ( .A(n11506), .ZN(n10970) );
  AOI211_X1 U13511 ( .C1(n10972), .C2(n10971), .A(n15294), .B(n10970), .ZN(
        n10973) );
  OR2_X1 U13512 ( .A1(n10974), .A2(n10973), .ZN(P2_U3227) );
  INV_X1 U13513 ( .A(n10975), .ZN(n10979) );
  INV_X1 U13514 ( .A(n14628), .ZN(n14621) );
  OAI222_X1 U13515 ( .A1(n15105), .A2(n10977), .B1(n10976), .B2(n10979), .C1(
        n14621), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13516 ( .A(n13532), .ZN(n13524) );
  OAI222_X1 U13517 ( .A1(P2_U3088), .A2(n13524), .B1(n14092), .B2(n10979), 
        .C1(n10978), .C2(n14097), .ZN(P2_U3309) );
  XNOR2_X1 U13518 ( .A(n10981), .B(n10982), .ZN(n15404) );
  INV_X1 U13519 ( .A(n15404), .ZN(n10994) );
  AND2_X1 U13520 ( .A1(n12889), .A2(n10983), .ZN(n11002) );
  INV_X1 U13521 ( .A(n11002), .ZN(n12894) );
  NOR2_X1 U13522 ( .A1(n12863), .A2(n12894), .ZN(n11969) );
  NAND2_X1 U13523 ( .A1(n10985), .A2(n10984), .ZN(n10986) );
  XNOR2_X1 U13524 ( .A(n10987), .B(n10986), .ZN(n10989) );
  INV_X1 U13525 ( .A(n12883), .ZN(n12045) );
  AOI22_X1 U13526 ( .A1(n12880), .A2(n12878), .B1(n12879), .B2(n12520), .ZN(
        n10988) );
  OAI21_X1 U13527 ( .B1(n10989), .B2(n12045), .A(n10988), .ZN(n10990) );
  AOI21_X1 U13528 ( .B1(n15404), .B2(n11777), .A(n10990), .ZN(n15406) );
  MUX2_X1 U13529 ( .A(n10991), .B(n15406), .S(n12896), .Z(n10993) );
  AOI22_X1 U13530 ( .A1(n12855), .A2(n15403), .B1(n12873), .B2(n11016), .ZN(
        n10992) );
  OAI211_X1 U13531 ( .C1(n10994), .C2(n11762), .A(n10993), .B(n10992), .ZN(
        P3_U3229) );
  INV_X1 U13532 ( .A(n10995), .ZN(n10996) );
  MUX2_X1 U13533 ( .A(n10997), .B(n10996), .S(n12896), .Z(n11000) );
  AOI22_X1 U13534 ( .A1(n12855), .A2(n10998), .B1(n8052), .B2(n12873), .ZN(
        n10999) );
  OAI211_X1 U13535 ( .C1(n11001), .C2(n11762), .A(n11000), .B(n10999), .ZN(
        P3_U3230) );
  INV_X1 U13536 ( .A(n12876), .ZN(n12839) );
  XOR2_X1 U13537 ( .A(n11004), .B(n11007), .Z(n15394) );
  AOI22_X1 U13538 ( .A1(n12839), .A2(n15394), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n12873), .ZN(n11015) );
  NOR2_X1 U13539 ( .A1(n11005), .A2(n15418), .ZN(n15393) );
  INV_X1 U13540 ( .A(n12889), .ZN(n11011) );
  XNOR2_X1 U13541 ( .A(n11007), .B(n11006), .ZN(n11008) );
  NAND2_X1 U13542 ( .A1(n11008), .A2(n12883), .ZN(n11010) );
  AOI22_X1 U13543 ( .A1(n12880), .A2(n12523), .B1(n12879), .B2(n12522), .ZN(
        n11009) );
  NAND2_X1 U13544 ( .A1(n11010), .A2(n11009), .ZN(n15392) );
  AOI21_X1 U13545 ( .B1(n15393), .B2(n11011), .A(n15392), .ZN(n11012) );
  MUX2_X1 U13546 ( .A(n11013), .B(n11012), .S(n12896), .Z(n11014) );
  NAND2_X1 U13547 ( .A1(n11015), .A2(n11014), .ZN(P3_U3232) );
  INV_X1 U13548 ( .A(n11016), .ZN(n11029) );
  INV_X1 U13549 ( .A(n11017), .ZN(n11018) );
  XNOR2_X1 U13550 ( .A(n12203), .B(n15403), .ZN(n11182) );
  XNOR2_X1 U13551 ( .A(n11182), .B(n12521), .ZN(n11019) );
  OAI21_X1 U13552 ( .B1(n11020), .B2(n11019), .A(n11183), .ZN(n11021) );
  NAND2_X1 U13553 ( .A1(n11021), .A2(n12436), .ZN(n11028) );
  INV_X1 U13554 ( .A(n11022), .ZN(n11026) );
  OAI22_X1 U13555 ( .A1(n12451), .A2(n11024), .B1(n11023), .B2(n12499), .ZN(
        n11025) );
  AOI211_X1 U13556 ( .C1(n12497), .C2(n12520), .A(n11026), .B(n11025), .ZN(
        n11027) );
  OAI211_X1 U13557 ( .C1(n11029), .C2(n12027), .A(n11028), .B(n11027), .ZN(
        P3_U3170) );
  NAND2_X1 U13558 ( .A1(n11032), .A2(n11426), .ZN(n11401) );
  NAND2_X1 U13559 ( .A1(n11403), .A2(n11401), .ZN(n11644) );
  XNOR2_X1 U13560 ( .A(n13447), .B(n15368), .ZN(n13397) );
  INV_X1 U13561 ( .A(n13397), .ZN(n11643) );
  NAND2_X1 U13562 ( .A1(n11644), .A2(n11643), .ZN(n11646) );
  INV_X1 U13563 ( .A(n13447), .ZN(n11034) );
  NAND2_X1 U13564 ( .A1(n11034), .A2(n11658), .ZN(n11402) );
  NAND2_X1 U13565 ( .A1(n11646), .A2(n11402), .ZN(n11076) );
  NAND2_X1 U13566 ( .A1(n11409), .A2(n13446), .ZN(n11080) );
  INV_X1 U13567 ( .A(n13446), .ZN(n11075) );
  NAND2_X1 U13568 ( .A1(n11075), .A2(n6418), .ZN(n11081) );
  AND2_X1 U13569 ( .A1(n11080), .A2(n11081), .ZN(n13395) );
  XNOR2_X1 U13570 ( .A(n11076), .B(n13395), .ZN(n11282) );
  NAND2_X1 U13571 ( .A1(n11032), .A2(n13218), .ZN(n11033) );
  XOR2_X1 U13572 ( .A(n11082), .B(n13395), .Z(n11037) );
  AOI21_X1 U13573 ( .B1(n11037), .B2(n13905), .A(n11036), .ZN(n11274) );
  AOI211_X1 U13574 ( .C1(n6418), .C2(n11654), .A(n13926), .B(n11085), .ZN(
        n11279) );
  AOI21_X1 U13575 ( .B1(n15377), .B2(n6418), .A(n11279), .ZN(n11038) );
  OAI211_X1 U13576 ( .C1(n15381), .C2(n11282), .A(n11274), .B(n11038), .ZN(
        n11041) );
  NAND2_X1 U13577 ( .A1(n11041), .A2(n15390), .ZN(n11039) );
  OAI21_X1 U13578 ( .B1(n15390), .B2(n11040), .A(n11039), .ZN(P2_U3504) );
  INV_X1 U13579 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U13580 ( .A1(n11041), .A2(n15384), .ZN(n11042) );
  OAI21_X1 U13581 ( .B1(n15384), .B2(n11043), .A(n11042), .ZN(P2_U3445) );
  INV_X1 U13582 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11057) );
  NAND2_X1 U13583 ( .A1(n7193), .A2(n11045), .ZN(n11046) );
  NAND2_X1 U13584 ( .A1(n11046), .A2(n15216), .ZN(n11047) );
  NOR2_X1 U13585 ( .A1(n11044), .A2(n11047), .ZN(n11176) );
  XNOR2_X1 U13586 ( .A(n11051), .B(n11048), .ZN(n11055) );
  OAI21_X1 U13587 ( .B1(n11051), .B2(n11050), .A(n11049), .ZN(n11052) );
  NAND2_X1 U13588 ( .A1(n11052), .A2(n15263), .ZN(n11054) );
  AOI22_X1 U13589 ( .A1(n14497), .A2(n14897), .B1(n14880), .B2(n14498), .ZN(
        n11053) );
  OAI211_X1 U13590 ( .C1(n15050), .C2(n11055), .A(n11054), .B(n11053), .ZN(
        n11174) );
  AOI211_X1 U13591 ( .C1(n15255), .C2(n7193), .A(n11176), .B(n11174), .ZN(
        n11058) );
  OR2_X1 U13592 ( .A1(n11058), .A2(n15264), .ZN(n11056) );
  OAI21_X1 U13593 ( .B1(n15265), .B2(n11057), .A(n11056), .ZN(P1_U3465) );
  OR2_X1 U13594 ( .A1(n11058), .A2(n15270), .ZN(n11059) );
  OAI21_X1 U13595 ( .B1(n15272), .B2(n10245), .A(n11059), .ZN(P1_U3530) );
  INV_X1 U13596 ( .A(n11106), .ZN(n11062) );
  INV_X1 U13597 ( .A(n13444), .ZN(n11490) );
  NOR3_X1 U13598 ( .A1(n13174), .A2(n11490), .A3(n11060), .ZN(n11061) );
  AOI21_X1 U13599 ( .B1(n11062), .B2(n13182), .A(n11061), .ZN(n11074) );
  INV_X1 U13600 ( .A(n11063), .ZN(n11210) );
  NOR2_X1 U13601 ( .A1(n13194), .A2(n7545), .ZN(n11071) );
  NAND2_X1 U13602 ( .A1(n13442), .A2(n13885), .ZN(n11065) );
  NAND2_X1 U13603 ( .A1(n13444), .A2(n13883), .ZN(n11064) );
  AND2_X1 U13604 ( .A1(n11065), .A2(n11064), .ZN(n11493) );
  INV_X1 U13605 ( .A(n11493), .ZN(n11066) );
  NAND2_X1 U13606 ( .A1(n13161), .A2(n11066), .ZN(n11068) );
  OAI211_X1 U13607 ( .C1(n13187), .C2(n11069), .A(n11068), .B(n11067), .ZN(
        n11070) );
  AOI211_X1 U13608 ( .C1(n11210), .C2(n13182), .A(n11071), .B(n11070), .ZN(
        n11072) );
  OAI21_X1 U13609 ( .B1(n11074), .B2(n11073), .A(n11072), .ZN(P2_U3193) );
  INV_X1 U13610 ( .A(n11076), .ZN(n11078) );
  OAI21_X1 U13611 ( .B1(n11076), .B2(n11075), .A(n11409), .ZN(n11077) );
  OAI21_X1 U13612 ( .B1(n11078), .B2(n13446), .A(n11077), .ZN(n11079) );
  XNOR2_X1 U13613 ( .A(n11079), .B(n13401), .ZN(n11642) );
  XNOR2_X1 U13614 ( .A(n11414), .B(n13401), .ZN(n11084) );
  AOI21_X1 U13615 ( .B1(n11084), .B2(n13905), .A(n11083), .ZN(n11633) );
  INV_X1 U13616 ( .A(n11085), .ZN(n11086) );
  AOI211_X1 U13617 ( .C1(n13235), .C2(n11086), .A(n13926), .B(n11418), .ZN(
        n11639) );
  AOI21_X1 U13618 ( .B1(n15377), .B2(n13235), .A(n11639), .ZN(n11087) );
  OAI211_X1 U13619 ( .C1(n15381), .C2(n11642), .A(n11633), .B(n11087), .ZN(
        n11089) );
  NAND2_X1 U13620 ( .A1(n11089), .A2(n15390), .ZN(n11088) );
  OAI21_X1 U13621 ( .B1(n15390), .B2(n10191), .A(n11088), .ZN(P2_U3505) );
  INV_X1 U13622 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11091) );
  NAND2_X1 U13623 ( .A1(n11089), .A2(n15384), .ZN(n11090) );
  OAI21_X1 U13624 ( .B1(n15384), .B2(n11091), .A(n11090), .ZN(P2_U3448) );
  XNOR2_X1 U13625 ( .A(n11092), .B(n11094), .ZN(n15409) );
  INV_X1 U13626 ( .A(n15409), .ZN(n11100) );
  NOR2_X1 U13627 ( .A1(n11093), .A2(n11094), .ZN(n11221) );
  AOI21_X1 U13628 ( .B1(n11094), .B2(n11093), .A(n11221), .ZN(n11096) );
  AOI22_X1 U13629 ( .A1(n12880), .A2(n12521), .B1(n12879), .B2(n12519), .ZN(
        n11095) );
  OAI21_X1 U13630 ( .B1(n11096), .B2(n12045), .A(n11095), .ZN(n11097) );
  AOI21_X1 U13631 ( .B1(n15409), .B2(n11777), .A(n11097), .ZN(n15411) );
  MUX2_X1 U13632 ( .A(n6832), .B(n15411), .S(n12896), .Z(n11099) );
  AOI22_X1 U13633 ( .A1(n12855), .A2(n15408), .B1(n12873), .B2(n11187), .ZN(
        n11098) );
  OAI211_X1 U13634 ( .C1(n11100), .C2(n11762), .A(n11099), .B(n11098), .ZN(
        P3_U3228) );
  OAI222_X1 U13635 ( .A1(P2_U3088), .A2(n13195), .B1(n14092), .B2(n11130), 
        .C1(n11101), .C2(n14097), .ZN(P2_U3307) );
  INV_X1 U13636 ( .A(n15376), .ZN(n11491) );
  INV_X1 U13637 ( .A(n11102), .ZN(n11103) );
  AOI21_X1 U13638 ( .B1(n11104), .B2(n11103), .A(n13165), .ZN(n11108) );
  INV_X1 U13639 ( .A(n13445), .ZN(n11413) );
  NOR3_X1 U13640 ( .A1(n13174), .A2(n11413), .A3(n11105), .ZN(n11107) );
  OAI21_X1 U13641 ( .B1(n11108), .B2(n11107), .A(n11106), .ZN(n11112) );
  AOI22_X1 U13642 ( .A1(n13885), .A2(n13443), .B1(n13445), .B2(n13883), .ZN(
        n11415) );
  OAI21_X1 U13643 ( .B1(n13120), .B2(n11415), .A(n11109), .ZN(n11110) );
  AOI21_X1 U13644 ( .B1(n11421), .B2(n13170), .A(n11110), .ZN(n11111) );
  OAI211_X1 U13645 ( .C1(n11491), .C2(n13194), .A(n11112), .B(n11111), .ZN(
        P2_U3185) );
  INV_X1 U13646 ( .A(n11113), .ZN(n11115) );
  OAI222_X1 U13647 ( .A1(n14097), .A2(n11114), .B1(n14092), .B2(n11115), .C1(
        P2_U3088), .C2(n13428), .ZN(P2_U3308) );
  OAI222_X1 U13648 ( .A1(n15105), .A2(n11116), .B1(n10976), .B2(n11115), .C1(
        n14917), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U13649 ( .A(n14907), .ZN(n15225) );
  OAI211_X1 U13650 ( .C1(n11044), .C2(n11342), .A(n15214), .B(n15216), .ZN(
        n15231) );
  XNOR2_X1 U13651 ( .A(n11117), .B(n14272), .ZN(n11124) );
  NAND3_X1 U13652 ( .A1(n11049), .A2(n14439), .A3(n14267), .ZN(n11118) );
  NAND2_X1 U13653 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  NAND2_X1 U13654 ( .A1(n11120), .A2(n15263), .ZN(n11123) );
  OR2_X1 U13655 ( .A1(n9741), .A2(n14935), .ZN(n11122) );
  NAND2_X1 U13656 ( .A1(n14897), .A2(n14496), .ZN(n11121) );
  AND2_X1 U13657 ( .A1(n11122), .A2(n11121), .ZN(n15172) );
  OAI211_X1 U13658 ( .C1(n15050), .C2(n11124), .A(n11123), .B(n15172), .ZN(
        n15234) );
  MUX2_X1 U13659 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n15234), .S(n15220), .Z(
        n11125) );
  INV_X1 U13660 ( .A(n11125), .ZN(n11127) );
  INV_X1 U13661 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U13662 ( .A1(n15223), .A2(n15170), .B1(n14530), .B2(n14974), .ZN(
        n11126) );
  OAI211_X1 U13663 ( .C1(n15225), .C2(n15231), .A(n11127), .B(n11126), .ZN(
        P1_U3290) );
  OAI222_X1 U13664 ( .A1(P2_U3088), .A2(n11129), .B1(n14092), .B2(n11230), 
        .C1(n11128), .C2(n14097), .ZN(P2_U3306) );
  OAI222_X1 U13665 ( .A1(n15105), .A2(n11132), .B1(P1_U3086), .B2(n11131), 
        .C1(n10976), .C2(n11130), .ZN(P1_U3335) );
  OAI222_X1 U13666 ( .A1(n11134), .A2(P3_U3151), .B1(n13034), .B2(n15447), 
        .C1(n13039), .C2(n11133), .ZN(P3_U3275) );
  NAND2_X1 U13667 ( .A1(n11144), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11137) );
  INV_X1 U13668 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11772) );
  XNOR2_X1 U13669 ( .A(n11378), .B(n11772), .ZN(n11158) );
  OAI21_X1 U13670 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11139), .A(n11385), .ZN(
        n11143) );
  NAND2_X1 U13671 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11875) );
  INV_X1 U13672 ( .A(n11875), .ZN(n11140) );
  AOI21_X1 U13673 ( .B1(n15391), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11140), .ZN(
        n11141) );
  OAI21_X1 U13674 ( .B1(n12697), .B2(n11379), .A(n11141), .ZN(n11142) );
  AOI21_X1 U13675 ( .B1(n11143), .B2(n12688), .A(n11142), .ZN(n11157) );
  MUX2_X1 U13676 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13031), .Z(n11148) );
  NAND2_X1 U13677 ( .A1(n11379), .A2(n11148), .ZN(n11153) );
  INV_X1 U13678 ( .A(n11148), .ZN(n11149) );
  NAND2_X1 U13679 ( .A1(n11150), .A2(n11149), .ZN(n11395) );
  INV_X1 U13680 ( .A(n11395), .ZN(n11151) );
  NOR2_X1 U13681 ( .A1(n11396), .A2(n11151), .ZN(n11155) );
  AOI21_X1 U13682 ( .B1(n11395), .B2(n11153), .A(n11152), .ZN(n11154) );
  OAI21_X1 U13683 ( .B1(n11155), .B2(n11154), .A(n12584), .ZN(n11156) );
  OAI211_X1 U13684 ( .C1(n11158), .C2(n12543), .A(n11157), .B(n11156), .ZN(
        P3_U3191) );
  INV_X1 U13685 ( .A(n11161), .ZN(n11162) );
  NAND2_X1 U13686 ( .A1(n11166), .A2(n11165), .ZN(n11169) );
  INV_X1 U13687 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U13688 ( .A1(n11167), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11168) );
  INV_X1 U13689 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15548) );
  NAND2_X1 U13690 ( .A1(n15548), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11251) );
  INV_X1 U13691 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U13692 ( .A1(n11170), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U13693 ( .A1(n11251), .A2(n11171), .ZN(n11249) );
  XNOR2_X1 U13694 ( .A(n11250), .B(n11249), .ZN(n11247) );
  OAI21_X1 U13695 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n11172), .A(n7246), .ZN(
        n11173) );
  INV_X1 U13696 ( .A(n11173), .ZN(SUB_1596_U54) );
  MUX2_X1 U13697 ( .A(n11174), .B(P1_REG2_REG_2__SCAN_IN), .S(n6412), .Z(
        n11175) );
  INV_X1 U13698 ( .A(n11175), .ZN(n11178) );
  AOI22_X1 U13699 ( .A1(n14907), .A2(n11176), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14974), .ZN(n11177) );
  OAI211_X1 U13700 ( .C1(n14268), .C2(n14921), .A(n11178), .B(n11177), .ZN(
        P1_U3291) );
  OAI222_X1 U13701 ( .A1(n13039), .A2(n11181), .B1(n13036), .B2(n11180), .C1(
        P3_U3151), .C2(n11179), .ZN(P3_U3274) );
  XNOR2_X1 U13702 ( .A(n12203), .B(n15408), .ZN(n11284) );
  XNOR2_X1 U13703 ( .A(n11284), .B(n12520), .ZN(n11285) );
  XOR2_X1 U13704 ( .A(n11285), .B(n11286), .Z(n11189) );
  INV_X1 U13705 ( .A(n12499), .ZN(n12485) );
  AOI22_X1 U13706 ( .A1(n12485), .A2(n12521), .B1(n12503), .B2(n15408), .ZN(
        n11185) );
  OAI211_X1 U13707 ( .C1(n11472), .C2(n12488), .A(n11185), .B(n11184), .ZN(
        n11186) );
  AOI21_X1 U13708 ( .B1(n11187), .B2(n12502), .A(n11186), .ZN(n11188) );
  OAI21_X1 U13709 ( .B1(n11189), .B2(n12506), .A(n11188), .ZN(P3_U3167) );
  INV_X1 U13710 ( .A(n11190), .ZN(n11193) );
  INV_X1 U13711 ( .A(n14442), .ZN(n11192) );
  INV_X1 U13712 ( .A(n11191), .ZN(n11300) );
  AOI21_X1 U13713 ( .B1(n11193), .B2(n11192), .A(n11300), .ZN(n15248) );
  AOI211_X1 U13714 ( .C1(n15245), .C2(n15215), .A(n14929), .B(n11307), .ZN(
        n15243) );
  OR2_X1 U13715 ( .A1(n11557), .A2(n14933), .ZN(n11195) );
  NAND2_X1 U13716 ( .A1(n14880), .A2(n14496), .ZN(n11194) );
  NAND2_X1 U13717 ( .A1(n11195), .A2(n11194), .ZN(n15244) );
  MUX2_X1 U13718 ( .A(n15244), .B(P1_REG2_REG_5__SCAN_IN), .S(n6412), .Z(
        n11198) );
  NAND2_X1 U13719 ( .A1(n15223), .A2(n15245), .ZN(n11196) );
  OAI21_X1 U13720 ( .B1(n15217), .B2(n11560), .A(n11196), .ZN(n11197) );
  AOI211_X1 U13721 ( .C1(n15243), .C2(n14907), .A(n11198), .B(n11197), .ZN(
        n11201) );
  XOR2_X1 U13722 ( .A(n11199), .B(n14442), .Z(n15250) );
  NOR2_X1 U13723 ( .A1(n6412), .A2(n15050), .ZN(n14850) );
  NAND2_X1 U13724 ( .A1(n15250), .A2(n14850), .ZN(n11200) );
  OAI211_X1 U13725 ( .C1(n15248), .C2(n14910), .A(n11201), .B(n11200), .ZN(
        P1_U3288) );
  INV_X1 U13726 ( .A(n11202), .ZN(n11794) );
  OR2_X1 U13727 ( .A1(n13256), .A2(n13871), .ZN(n11204) );
  NAND2_X1 U13728 ( .A1(n13443), .A2(n13883), .ZN(n11203) );
  NAND2_X1 U13729 ( .A1(n11204), .A2(n11203), .ZN(n11789) );
  NAND2_X1 U13730 ( .A1(n13161), .A2(n11789), .ZN(n11206) );
  OAI211_X1 U13731 ( .C1(n13187), .C2(n11794), .A(n11206), .B(n11205), .ZN(
        n11212) );
  AOI22_X1 U13732 ( .A1(n13183), .A2(n13443), .B1(n13182), .B2(n11207), .ZN(
        n11209) );
  NOR3_X1 U13733 ( .A1(n11210), .A2(n11209), .A3(n11208), .ZN(n11211) );
  AOI211_X1 U13734 ( .C1(n14051), .C2(n13173), .A(n11212), .B(n11211), .ZN(
        n11213) );
  OAI21_X1 U13735 ( .B1(n13165), .B2(n11214), .A(n11213), .ZN(P2_U3203) );
  XNOR2_X1 U13736 ( .A(n11216), .B(n11215), .ZN(n15414) );
  INV_X1 U13737 ( .A(n15414), .ZN(n11229) );
  INV_X1 U13738 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11226) );
  OAI22_X1 U13739 ( .A1(n11681), .A2(n12048), .B1(n11289), .B2(n12144), .ZN(
        n11225) );
  INV_X1 U13740 ( .A(n11221), .ZN(n11219) );
  AOI21_X1 U13741 ( .B1(n11219), .B2(n11218), .A(n11217), .ZN(n11223) );
  OR2_X1 U13742 ( .A1(n11221), .A2(n11220), .ZN(n11453) );
  INV_X1 U13743 ( .A(n11453), .ZN(n11222) );
  NOR3_X1 U13744 ( .A1(n11223), .A2(n11222), .A3(n12045), .ZN(n11224) );
  AOI211_X1 U13745 ( .C1(n15414), .C2(n11777), .A(n11225), .B(n11224), .ZN(
        n15416) );
  MUX2_X1 U13746 ( .A(n11226), .B(n15416), .S(n12896), .Z(n11228) );
  AOI22_X1 U13747 ( .A1(n12855), .A2(n15413), .B1(n12873), .B2(n11283), .ZN(
        n11227) );
  OAI211_X1 U13748 ( .C1(n11229), .C2(n11762), .A(n11228), .B(n11227), .ZN(
        P3_U3227) );
  OAI222_X1 U13749 ( .A1(n15105), .A2(n15495), .B1(P1_U3086), .B2(n14247), 
        .C1(n10976), .C2(n11230), .ZN(P1_U3334) );
  AOI21_X1 U13750 ( .B1(n11233), .B2(n11232), .A(n11231), .ZN(n14589) );
  INV_X1 U13751 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n14924) );
  MUX2_X1 U13752 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n14924), .S(n14586), .Z(
        n14588) );
  NAND2_X1 U13753 ( .A1(n14589), .A2(n14588), .ZN(n14587) );
  NAND2_X1 U13754 ( .A1(n14586), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11235) );
  MUX2_X1 U13755 ( .A(n14904), .B(P1_REG2_REG_14__SCAN_IN), .S(n11617), .Z(
        n11234) );
  AOI21_X1 U13756 ( .B1(n14587), .B2(n11235), .A(n11234), .ZN(n11614) );
  NAND3_X1 U13757 ( .A1(n14587), .A2(n11235), .A3(n11234), .ZN(n11236) );
  NAND2_X1 U13758 ( .A1(n11236), .A2(n15194), .ZN(n11246) );
  XNOR2_X1 U13759 ( .A(n11617), .B(n11237), .ZN(n11240) );
  NOR2_X1 U13760 ( .A1(n11238), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n14579) );
  XNOR2_X1 U13761 ( .A(n14586), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n14578) );
  OAI21_X1 U13762 ( .B1(n11240), .B2(n11239), .A(n11616), .ZN(n11241) );
  NAND2_X1 U13763 ( .A1(n11241), .A2(n15188), .ZN(n11245) );
  NOR2_X1 U13764 ( .A1(n11242), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14112) );
  INV_X1 U13765 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15125) );
  NOR2_X1 U13766 ( .A1(n14583), .A2(n15125), .ZN(n11243) );
  AOI211_X1 U13767 ( .C1(n15197), .C2(n11617), .A(n14112), .B(n11243), .ZN(
        n11244) );
  OAI211_X1 U13768 ( .C1(n11614), .C2(n11246), .A(n11245), .B(n11244), .ZN(
        P1_U3257) );
  XNOR2_X1 U13769 ( .A(n11253), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n11593) );
  INV_X1 U13770 ( .A(n11593), .ZN(n11254) );
  XNOR2_X1 U13771 ( .A(n11594), .B(n11254), .ZN(n11590) );
  XNOR2_X1 U13772 ( .A(n11590), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n11255) );
  XNOR2_X1 U13773 ( .A(n11589), .B(n11255), .ZN(SUB_1596_U70) );
  NAND2_X1 U13774 ( .A1(n13880), .A2(n13802), .ZN(n11273) );
  NAND2_X1 U13775 ( .A1(n11273), .A2(n13811), .ZN(n13897) );
  OAI21_X1 U13776 ( .B1(n11258), .B2(n11257), .A(n11256), .ZN(n11259) );
  INV_X1 U13777 ( .A(n11259), .ZN(n15364) );
  OAI21_X1 U13778 ( .B1(n11260), .B2(n13396), .A(n11261), .ZN(n11262) );
  AOI222_X1 U13779 ( .A1(n13905), .A2(n11262), .B1(n13448), .B2(n13885), .C1(
        n13450), .C2(n13883), .ZN(n15363) );
  MUX2_X1 U13780 ( .A(n11263), .B(n15363), .S(n13880), .Z(n11269) );
  AOI211_X1 U13781 ( .C1(n15361), .C2(n11265), .A(n13926), .B(n11264), .ZN(
        n15360) );
  OAI22_X1 U13782 ( .A1(n13931), .A2(n11266), .B1(n13837), .B2(n8744), .ZN(
        n11267) );
  AOI21_X1 U13783 ( .B1(n13938), .B2(n15360), .A(n11267), .ZN(n11268) );
  OAI211_X1 U13784 ( .C1(n13915), .C2(n15364), .A(n11269), .B(n11268), .ZN(
        P2_U3263) );
  INV_X1 U13785 ( .A(n11270), .ZN(n11271) );
  OAI222_X1 U13786 ( .A1(n14097), .A2(n11272), .B1(P2_U3088), .B2(n13373), 
        .C1(n14092), .C2(n11271), .ZN(P2_U3305) );
  MUX2_X1 U13787 ( .A(n11275), .B(n11274), .S(n13880), .Z(n11281) );
  INV_X1 U13788 ( .A(n11276), .ZN(n11277) );
  OAI22_X1 U13789 ( .A1(n13931), .A2(n11409), .B1(n11277), .B2(n13837), .ZN(
        n11278) );
  AOI21_X1 U13790 ( .B1(n11279), .B2(n13938), .A(n11278), .ZN(n11280) );
  OAI211_X1 U13791 ( .C1(n13935), .C2(n11282), .A(n11281), .B(n11280), .ZN(
        P2_U3260) );
  INV_X1 U13792 ( .A(n11283), .ZN(n11295) );
  XNOR2_X1 U13793 ( .A(n12203), .B(n15413), .ZN(n11466) );
  XNOR2_X1 U13794 ( .A(n11466), .B(n12519), .ZN(n11287) );
  OAI211_X1 U13795 ( .C1(n11288), .C2(n11287), .A(n11468), .B(n12436), .ZN(
        n11294) );
  OAI22_X1 U13796 ( .A1(n12451), .A2(n11290), .B1(n11289), .B2(n12499), .ZN(
        n11291) );
  AOI211_X1 U13797 ( .C1(n12497), .C2(n12518), .A(n11292), .B(n11291), .ZN(
        n11293) );
  OAI211_X1 U13798 ( .C1(n11295), .C2(n12027), .A(n11294), .B(n11293), .ZN(
        P3_U3179) );
  OR2_X1 U13799 ( .A1(n11296), .A2(n14440), .ZN(n11318) );
  INV_X1 U13800 ( .A(n11318), .ZN(n11297) );
  AOI21_X1 U13801 ( .B1(n14440), .B2(n11296), .A(n11297), .ZN(n11306) );
  INV_X1 U13802 ( .A(n11298), .ZN(n11299) );
  NOR3_X1 U13803 ( .A1(n11300), .A2(n11299), .A3(n14440), .ZN(n11303) );
  INV_X1 U13804 ( .A(n11301), .ZN(n11302) );
  OAI21_X1 U13805 ( .B1(n11303), .B2(n11302), .A(n15263), .ZN(n11305) );
  AOI22_X1 U13806 ( .A1(n14897), .A2(n14493), .B1(n14880), .B2(n14495), .ZN(
        n11304) );
  OAI211_X1 U13807 ( .C1(n15050), .C2(n11306), .A(n11305), .B(n11304), .ZN(
        n15252) );
  INV_X1 U13808 ( .A(n15252), .ZN(n11312) );
  INV_X1 U13809 ( .A(n11307), .ZN(n11308) );
  AOI211_X1 U13810 ( .C1(n15254), .C2(n11308), .A(n14929), .B(n11326), .ZN(
        n15253) );
  NOR2_X1 U13811 ( .A1(n14921), .A2(n11377), .ZN(n11310) );
  OAI22_X1 U13812 ( .A1(n15220), .A2(n10320), .B1(n11372), .B2(n15217), .ZN(
        n11309) );
  AOI211_X1 U13813 ( .C1(n15253), .C2(n14907), .A(n11310), .B(n11309), .ZN(
        n11311) );
  OAI21_X1 U13814 ( .B1(n11312), .B2(n6412), .A(n11311), .ZN(P1_U3287) );
  INV_X1 U13815 ( .A(n11313), .ZN(n11316) );
  OAI22_X1 U13816 ( .A1(n11314), .A2(P3_U3151), .B1(SI_22_), .B2(n13036), .ZN(
        n11315) );
  AOI21_X1 U13817 ( .B1(n11316), .B2(n13016), .A(n11315), .ZN(P3_U3273) );
  NAND3_X1 U13818 ( .A1(n11318), .A2(n9749), .A3(n11317), .ZN(n11319) );
  NAND2_X1 U13819 ( .A1(n11320), .A2(n11319), .ZN(n11322) );
  OAI22_X1 U13820 ( .A1(n11557), .A2(n14935), .B1(n11826), .B2(n14933), .ZN(
        n11321) );
  AOI21_X1 U13821 ( .B1(n11322), .B2(n15251), .A(n11321), .ZN(n15258) );
  OAI21_X1 U13822 ( .B1(n11324), .B2(n9749), .A(n11323), .ZN(n15262) );
  OAI211_X1 U13823 ( .C1(n11326), .C2(n15260), .A(n15216), .B(n11325), .ZN(
        n15257) );
  OAI22_X1 U13824 ( .A1(n15220), .A2(n10322), .B1(n11542), .B2(n15217), .ZN(
        n11327) );
  AOI21_X1 U13825 ( .B1(n15223), .B2(n14289), .A(n11327), .ZN(n11328) );
  OAI21_X1 U13826 ( .B1(n15225), .B2(n15257), .A(n11328), .ZN(n11329) );
  AOI21_X1 U13827 ( .B1(n15262), .B2(n15227), .A(n11329), .ZN(n11330) );
  OAI21_X1 U13828 ( .B1(n6412), .B2(n15258), .A(n11330), .ZN(P1_U3286) );
  NOR2_X1 U13829 ( .A1(n11331), .A2(P2_U3088), .ZN(n13433) );
  AOI21_X1 U13830 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n11332), .A(n13433), 
        .ZN(n11333) );
  OAI21_X1 U13831 ( .B1(n11335), .B2(n14092), .A(n11333), .ZN(P2_U3304) );
  AOI21_X1 U13832 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n12221), .A(n14469), 
        .ZN(n11334) );
  OAI21_X1 U13833 ( .B1(n11335), .B2(n10976), .A(n11334), .ZN(P1_U3332) );
  INV_X1 U13834 ( .A(n14221), .ZN(n14242) );
  OAI22_X1 U13835 ( .A1(n11343), .A2(n6402), .B1(n11342), .B2(n12273), .ZN(
        n11340) );
  XNOR2_X1 U13836 ( .A(n11340), .B(n11355), .ZN(n11344) );
  OAI22_X1 U13837 ( .A1(n11343), .A2(n6416), .B1(n11342), .B2(n6401), .ZN(
        n11345) );
  XNOR2_X1 U13838 ( .A(n11344), .B(n11345), .ZN(n15176) );
  INV_X1 U13839 ( .A(n11344), .ZN(n11347) );
  INV_X1 U13840 ( .A(n11345), .ZN(n11346) );
  OAI22_X1 U13841 ( .A1(n11348), .A2(n6416), .B1(n15237), .B2(n6402), .ZN(
        n11548) );
  NAND2_X1 U13842 ( .A1(n12315), .A2(n14496), .ZN(n11350) );
  XNOR2_X1 U13843 ( .A(n11351), .B(n12313), .ZN(n11434) );
  NAND2_X1 U13844 ( .A1(n12315), .A2(n14495), .ZN(n11354) );
  OR2_X1 U13845 ( .A1(n12273), .A2(n11357), .ZN(n11353) );
  NAND2_X1 U13846 ( .A1(n11354), .A2(n11353), .ZN(n11356) );
  XNOR2_X1 U13847 ( .A(n11356), .B(n11538), .ZN(n11553) );
  INV_X1 U13848 ( .A(n11553), .ZN(n11359) );
  OAI22_X1 U13849 ( .A1(n11358), .A2(n6416), .B1(n11357), .B2(n6401), .ZN(
        n11552) );
  AOI22_X1 U13850 ( .A1(n11548), .A2(n11434), .B1(n11359), .B2(n11552), .ZN(
        n11364) );
  OAI21_X1 U13851 ( .B1(n11434), .B2(n11548), .A(n11552), .ZN(n11361) );
  NOR3_X1 U13852 ( .A1(n11434), .A2(n11548), .A3(n11552), .ZN(n11360) );
  AOI21_X1 U13853 ( .B1(n11553), .B2(n11361), .A(n11360), .ZN(n11362) );
  INV_X1 U13854 ( .A(n11362), .ZN(n11363) );
  OAI22_X1 U13855 ( .A1(n11557), .A2(n6416), .B1(n11377), .B2(n6401), .ZN(
        n11533) );
  OAI22_X1 U13856 ( .A1(n11557), .A2(n6402), .B1(n11377), .B2(n12273), .ZN(
        n11365) );
  XNOR2_X1 U13857 ( .A(n11365), .B(n12313), .ZN(n11532) );
  XOR2_X1 U13858 ( .A(n11533), .B(n11532), .Z(n11366) );
  NAND2_X1 U13859 ( .A1(n11367), .A2(n11366), .ZN(n11536) );
  OAI211_X1 U13860 ( .C1(n11367), .C2(n11366), .A(n11536), .B(n14232), .ZN(
        n11376) );
  INV_X1 U13861 ( .A(n11368), .ZN(n11369) );
  OR2_X1 U13862 ( .A1(n11370), .A2(n11369), .ZN(n11371) );
  NOR2_X1 U13863 ( .A1(n15182), .A2(n11372), .ZN(n11374) );
  NAND2_X1 U13864 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14546) );
  OAI21_X1 U13865 ( .B1(n14236), .B2(n11537), .A(n14546), .ZN(n11373) );
  AOI211_X1 U13866 ( .C1(n14239), .C2(n14495), .A(n11374), .B(n11373), .ZN(
        n11375) );
  OAI211_X1 U13867 ( .C1(n11377), .C2(n14242), .A(n11376), .B(n11375), .ZN(
        P1_U3239) );
  INV_X1 U13868 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11950) );
  XNOR2_X1 U13869 ( .A(n6403), .B(n11950), .ZN(n11717) );
  NAND2_X1 U13870 ( .A1(n11380), .A2(n11379), .ZN(n11381) );
  XOR2_X1 U13871 ( .A(n11717), .B(n11718), .Z(n11400) );
  INV_X1 U13872 ( .A(n6403), .ZN(n11391) );
  NAND2_X1 U13873 ( .A1(n15391), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U13874 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12020)
         );
  NAND2_X1 U13875 ( .A1(n11383), .A2(n12020), .ZN(n11390) );
  XNOR2_X1 U13876 ( .A(n6403), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11386) );
  INV_X1 U13877 ( .A(n11721), .ZN(n11388) );
  NAND3_X1 U13878 ( .A1(n11385), .A2(n11386), .A3(n6833), .ZN(n11387) );
  AOI21_X1 U13879 ( .B1(n11388), .B2(n11387), .A(n12663), .ZN(n11389) );
  AOI211_X1 U13880 ( .C1(n12661), .C2(n11391), .A(n11390), .B(n11389), .ZN(
        n11399) );
  MUX2_X1 U13881 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13031), .Z(n11392) );
  OR2_X1 U13882 ( .A1(n6403), .A2(n11392), .ZN(n11726) );
  NAND2_X1 U13883 ( .A1(n6403), .A2(n11392), .ZN(n11393) );
  NAND2_X1 U13884 ( .A1(n11726), .A2(n11393), .ZN(n11394) );
  AND3_X1 U13885 ( .A1(n11396), .A2(n11395), .A3(n11394), .ZN(n11397) );
  OAI21_X1 U13886 ( .B1(n11727), .B2(n11397), .A(n12584), .ZN(n11398) );
  OAI211_X1 U13887 ( .C1(n11400), .C2(n12543), .A(n11399), .B(n11398), .ZN(
        P3_U3192) );
  NAND2_X1 U13888 ( .A1(n11403), .A2(n7842), .ZN(n11407) );
  AOI22_X1 U13889 ( .A1(n6418), .A2(n13446), .B1(n13447), .B2(n15368), .ZN(
        n11405) );
  NAND2_X1 U13890 ( .A1(n13235), .A2(n13445), .ZN(n11404) );
  AND2_X1 U13891 ( .A1(n11405), .A2(n11404), .ZN(n11406) );
  NAND2_X1 U13892 ( .A1(n11407), .A2(n11406), .ZN(n11412) );
  OAI21_X1 U13893 ( .B1(n6418), .B2(n13446), .A(n13445), .ZN(n11410) );
  NOR2_X1 U13894 ( .A1(n13445), .A2(n13446), .ZN(n11408) );
  AOI22_X1 U13895 ( .A1(n11637), .A2(n11410), .B1(n11409), .B2(n11408), .ZN(
        n11411) );
  NAND2_X1 U13896 ( .A1(n11412), .A2(n11411), .ZN(n11481) );
  XNOR2_X1 U13897 ( .A(n15376), .B(n13444), .ZN(n13402) );
  XNOR2_X1 U13898 ( .A(n11481), .B(n13402), .ZN(n15380) );
  INV_X1 U13899 ( .A(n13402), .ZN(n11480) );
  XNOR2_X1 U13900 ( .A(n11480), .B(n11492), .ZN(n11417) );
  INV_X1 U13901 ( .A(n11415), .ZN(n11416) );
  AOI21_X1 U13902 ( .B1(n11417), .B2(n13905), .A(n11416), .ZN(n15379) );
  MUX2_X1 U13903 ( .A(n10226), .B(n15379), .S(n13880), .Z(n11425) );
  INV_X1 U13904 ( .A(n11418), .ZN(n11420) );
  INV_X1 U13905 ( .A(n11488), .ZN(n11419) );
  AOI211_X1 U13906 ( .C1(n15376), .C2(n11420), .A(n13926), .B(n11419), .ZN(
        n15375) );
  INV_X1 U13907 ( .A(n11421), .ZN(n11422) );
  OAI22_X1 U13908 ( .A1(n13931), .A2(n11491), .B1(n11422), .B2(n13837), .ZN(
        n11423) );
  AOI21_X1 U13909 ( .B1(n15375), .B2(n13938), .A(n11423), .ZN(n11424) );
  OAI211_X1 U13910 ( .C1(n13915), .C2(n15380), .A(n11425), .B(n11424), .ZN(
        P2_U3258) );
  OAI22_X1 U13911 ( .A1(n13931), .A2(n11426), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13837), .ZN(n11427) );
  AOI21_X1 U13912 ( .B1(n13938), .B2(n11428), .A(n11427), .ZN(n11432) );
  MUX2_X1 U13913 ( .A(n11430), .B(n11429), .S(n13880), .Z(n11431) );
  OAI211_X1 U13914 ( .C1(n13915), .C2(n11433), .A(n11432), .B(n11431), .ZN(
        P2_U3262) );
  XNOR2_X1 U13915 ( .A(n11551), .B(n11548), .ZN(n11435) );
  NAND2_X1 U13916 ( .A1(n11435), .A2(n11434), .ZN(n11549) );
  OAI211_X1 U13917 ( .C1(n11435), .C2(n11434), .A(n11549), .B(n14232), .ZN(
        n11440) );
  INV_X1 U13918 ( .A(n15218), .ZN(n11438) );
  AOI22_X1 U13919 ( .A1(n14497), .A2(n14880), .B1(n14897), .B2(n14495), .ZN(
        n15208) );
  INV_X1 U13920 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n11436) );
  OAI22_X1 U13921 ( .A1(n14198), .A2(n15208), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11436), .ZN(n11437) );
  AOI21_X1 U13922 ( .B1(n14211), .B2(n11438), .A(n11437), .ZN(n11439) );
  OAI211_X1 U13923 ( .C1(n15237), .C2(n14242), .A(n11440), .B(n11439), .ZN(
        P1_U3230) );
  XNOR2_X1 U13924 ( .A(n11441), .B(n11443), .ZN(n15426) );
  INV_X1 U13925 ( .A(n15426), .ZN(n11451) );
  INV_X1 U13926 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U13927 ( .A1(n11442), .A2(n11443), .ZN(n11444) );
  AOI21_X1 U13928 ( .B1(n11445), .B2(n11444), .A(n12045), .ZN(n11447) );
  OAI22_X1 U13929 ( .A1(n12021), .A2(n12048), .B1(n11681), .B2(n12144), .ZN(
        n11446) );
  AOI211_X1 U13930 ( .C1(n15426), .C2(n11777), .A(n11447), .B(n11446), .ZN(
        n15428) );
  MUX2_X1 U13931 ( .A(n11448), .B(n15428), .S(n12896), .Z(n11450) );
  INV_X1 U13932 ( .A(n11682), .ZN(n15424) );
  AOI22_X1 U13933 ( .A1(n12855), .A2(n15424), .B1(n12873), .B2(n11674), .ZN(
        n11449) );
  OAI211_X1 U13934 ( .C1(n11451), .C2(n11762), .A(n11450), .B(n11449), .ZN(
        P3_U3225) );
  INV_X1 U13935 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15474) );
  NAND2_X1 U13936 ( .A1(n11453), .A2(n11452), .ZN(n11455) );
  XNOR2_X1 U13937 ( .A(n11454), .B(n11455), .ZN(n11460) );
  XNOR2_X1 U13938 ( .A(n11457), .B(n11456), .ZN(n15422) );
  NAND2_X1 U13939 ( .A1(n15422), .A2(n11777), .ZN(n11459) );
  AOI22_X1 U13940 ( .A1(n12879), .A2(n12517), .B1(n12880), .B2(n12519), .ZN(
        n11458) );
  OAI211_X1 U13941 ( .C1(n12045), .C2(n11460), .A(n11459), .B(n11458), .ZN(
        n15420) );
  INV_X1 U13942 ( .A(n15422), .ZN(n11462) );
  INV_X1 U13943 ( .A(n11461), .ZN(n11477) );
  OAI22_X1 U13944 ( .A1(n11462), .A2(n12894), .B1(n11477), .B2(n12891), .ZN(
        n11463) );
  NOR2_X1 U13945 ( .A1(n15420), .A2(n11463), .ZN(n11464) );
  MUX2_X1 U13946 ( .A(n15474), .B(n11464), .S(n12896), .Z(n11465) );
  OAI21_X1 U13947 ( .B1(n15419), .B2(n12867), .A(n11465), .ZN(P3_U3226) );
  XNOR2_X1 U13948 ( .A(n12203), .B(n11469), .ZN(n11675) );
  XNOR2_X1 U13949 ( .A(n11675), .B(n12518), .ZN(n11470) );
  OAI211_X1 U13950 ( .C1(n11471), .C2(n11470), .A(n11678), .B(n12436), .ZN(
        n11476) );
  OAI22_X1 U13951 ( .A1(n12451), .A2(n15419), .B1(n11472), .B2(n12499), .ZN(
        n11473) );
  AOI211_X1 U13952 ( .C1(n12497), .C2(n12517), .A(n11474), .B(n11473), .ZN(
        n11475) );
  OAI211_X1 U13953 ( .C1(n11477), .C2(n12027), .A(n11476), .B(n11475), .ZN(
        P3_U3153) );
  OAI222_X1 U13954 ( .A1(P2_U3088), .A2(n11479), .B1(n14092), .B2(n11530), 
        .C1(n11478), .C2(n14097), .ZN(P2_U3303) );
  NAND2_X1 U13955 ( .A1(n11481), .A2(n11480), .ZN(n11483) );
  OR2_X1 U13956 ( .A1(n15376), .A2(n13444), .ZN(n11482) );
  NAND2_X1 U13957 ( .A1(n11483), .A2(n11482), .ZN(n11486) );
  INV_X1 U13958 ( .A(n11486), .ZN(n11485) );
  XNOR2_X1 U13959 ( .A(n13246), .B(n13443), .ZN(n13404) );
  NAND2_X1 U13960 ( .A1(n11485), .A2(n11484), .ZN(n11745) );
  NAND2_X1 U13961 ( .A1(n11486), .A2(n13404), .ZN(n11487) );
  AND2_X1 U13962 ( .A1(n11745), .A2(n11487), .ZN(n11631) );
  INV_X1 U13963 ( .A(n15381), .ZN(n14028) );
  AOI21_X1 U13964 ( .B1(n11488), .B2(n13246), .A(n13926), .ZN(n11489) );
  NAND2_X1 U13965 ( .A1(n11489), .A2(n11793), .ZN(n11626) );
  OAI21_X1 U13966 ( .B1(n7545), .B2(n14024), .A(n11626), .ZN(n11495) );
  XOR2_X1 U13967 ( .A(n11738), .B(n13404), .Z(n11494) );
  OAI21_X1 U13968 ( .B1(n11494), .B2(n13920), .A(n11493), .ZN(n11627) );
  AOI211_X1 U13969 ( .C1(n11631), .C2(n14028), .A(n11495), .B(n11627), .ZN(
        n11498) );
  NAND2_X1 U13970 ( .A1(n6771), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n11496) );
  OAI21_X1 U13971 ( .B1(n11498), .B2(n6771), .A(n11496), .ZN(P2_U3454) );
  NAND2_X1 U13972 ( .A1(n15387), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11497) );
  OAI21_X1 U13973 ( .B1(n11498), .B2(n15387), .A(n11497), .ZN(P2_U3507) );
  XNOR2_X1 U13974 ( .A(n11507), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15310) );
  INV_X1 U13975 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11500) );
  INV_X1 U13976 ( .A(n11668), .ZN(n11501) );
  XNOR2_X1 U13977 ( .A(n11666), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n11515) );
  NOR2_X1 U13978 ( .A1(n11502), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13190) );
  NOR2_X1 U13979 ( .A1(n15313), .A2(n11511), .ZN(n11503) );
  AOI211_X1 U13980 ( .C1(n15273), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n13190), 
        .B(n11503), .ZN(n11514) );
  NAND2_X1 U13981 ( .A1(n11504), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U13982 ( .A1(n11506), .A2(n11505), .ZN(n11508) );
  NAND2_X1 U13983 ( .A1(n15317), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U13984 ( .A1(n11508), .A2(n11507), .ZN(n11509) );
  NAND2_X1 U13985 ( .A1(n11510), .A2(n11509), .ZN(n11663) );
  XNOR2_X1 U13986 ( .A(n11663), .B(n11511), .ZN(n11662) );
  XOR2_X1 U13987 ( .A(P2_REG2_REG_15__SCAN_IN), .B(n11662), .Z(n11512) );
  NAND2_X1 U13988 ( .A1(n11512), .A2(n15318), .ZN(n11513) );
  OAI211_X1 U13989 ( .C1(n11515), .C2(n15300), .A(n11514), .B(n11513), .ZN(
        P2_U3229) );
  INV_X1 U13990 ( .A(n11516), .ZN(n11518) );
  NAND2_X1 U13991 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  XNOR2_X1 U13992 ( .A(n11520), .B(n11519), .ZN(n11525) );
  INV_X1 U13993 ( .A(n13929), .ZN(n11522) );
  OAI22_X1 U13994 ( .A1(n13614), .A2(n13871), .B1(n13608), .B2(n13869), .ZN(
        n13922) );
  AOI22_X1 U13995 ( .A1(n13161), .A2(n13922), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11521) );
  OAI21_X1 U13996 ( .B1(n11522), .B2(n13187), .A(n11521), .ZN(n11523) );
  AOI21_X1 U13997 ( .B1(n14036), .B2(n13173), .A(n11523), .ZN(n11524) );
  OAI21_X1 U13998 ( .B1(n11525), .B2(n13165), .A(n11524), .ZN(P2_U3196) );
  NAND2_X1 U13999 ( .A1(n11526), .A2(n13016), .ZN(n11528) );
  OAI211_X1 U14000 ( .C1(n11529), .C2(n13036), .A(n11528), .B(n11527), .ZN(
        P3_U3272) );
  OAI222_X1 U14001 ( .A1(n15105), .A2(n7526), .B1(P1_U3086), .B2(n11531), .C1(
        n10976), .C2(n11530), .ZN(P1_U3331) );
  INV_X1 U14002 ( .A(n11532), .ZN(n11535) );
  INV_X1 U14003 ( .A(n11533), .ZN(n11534) );
  OAI22_X1 U14004 ( .A1(n15260), .A2(n12273), .B1(n11537), .B2(n6402), .ZN(
        n11539) );
  XNOR2_X1 U14005 ( .A(n11539), .B(n12313), .ZN(n11844) );
  AOI22_X1 U14006 ( .A1(n10744), .A2(n14493), .B1(n12315), .B2(n14289), .ZN(
        n11845) );
  XNOR2_X1 U14007 ( .A(n11844), .B(n11845), .ZN(n11540) );
  OAI211_X1 U14008 ( .C1(n11541), .C2(n11540), .A(n11847), .B(n14232), .ZN(
        n11547) );
  NOR2_X1 U14009 ( .A1(n15182), .A2(n11542), .ZN(n11545) );
  OAI21_X1 U14010 ( .B1(n14236), .B2(n11826), .A(n11543), .ZN(n11544) );
  AOI211_X1 U14011 ( .C1(n14239), .C2(n14494), .A(n11545), .B(n11544), .ZN(
        n11546) );
  OAI211_X1 U14012 ( .C1(n15260), .C2(n14242), .A(n11547), .B(n11546), .ZN(
        P1_U3213) );
  INV_X1 U14013 ( .A(n11548), .ZN(n11550) );
  OAI21_X1 U14014 ( .B1(n11551), .B2(n11550), .A(n11549), .ZN(n11555) );
  XNOR2_X1 U14015 ( .A(n11553), .B(n11552), .ZN(n11554) );
  XNOR2_X1 U14016 ( .A(n11555), .B(n11554), .ZN(n11563) );
  OAI21_X1 U14017 ( .B1(n14236), .B2(n11557), .A(n11556), .ZN(n11558) );
  AOI21_X1 U14018 ( .B1(n14239), .B2(n14496), .A(n11558), .ZN(n11559) );
  OAI21_X1 U14019 ( .B1(n11560), .B2(n15182), .A(n11559), .ZN(n11561) );
  AOI21_X1 U14020 ( .B1(n14221), .B2(n15245), .A(n11561), .ZN(n11562) );
  OAI21_X1 U14021 ( .B1(n11563), .B2(n15174), .A(n11562), .ZN(P1_U3227) );
  XNOR2_X1 U14022 ( .A(n11564), .B(n11565), .ZN(n11756) );
  XNOR2_X1 U14023 ( .A(n11566), .B(n11565), .ZN(n11569) );
  NAND2_X1 U14024 ( .A1(n11756), .A2(n11777), .ZN(n11568) );
  AOI22_X1 U14025 ( .A1(n12880), .A2(n12517), .B1(n12879), .B2(n12162), .ZN(
        n11567) );
  OAI211_X1 U14026 ( .C1(n12045), .C2(n11569), .A(n11568), .B(n11567), .ZN(
        n11757) );
  AOI21_X1 U14027 ( .B1(n15425), .B2(n11756), .A(n11757), .ZN(n11771) );
  INV_X1 U14028 ( .A(n11882), .ZN(n11759) );
  AOI22_X1 U14029 ( .A1(n13007), .A2(n11759), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15429), .ZN(n11570) );
  OAI21_X1 U14030 ( .B1(n11771), .B2(n15429), .A(n11570), .ZN(P3_U3417) );
  INV_X1 U14031 ( .A(n11571), .ZN(n11575) );
  OAI222_X1 U14032 ( .A1(n14097), .A2(n11573), .B1(n14092), .B2(n11575), .C1(
        P2_U3088), .C2(n11572), .ZN(P2_U3302) );
  OAI222_X1 U14033 ( .A1(n15105), .A2(n11576), .B1(n10976), .B2(n11575), .C1(
        n11574), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U14034 ( .A(n11578), .ZN(n11748) );
  OR2_X1 U14035 ( .A1(n13608), .A2(n13871), .ZN(n11580) );
  NAND2_X1 U14036 ( .A1(n13442), .A2(n13883), .ZN(n11579) );
  NAND2_X1 U14037 ( .A1(n11580), .A2(n11579), .ZN(n11742) );
  NAND2_X1 U14038 ( .A1(n13161), .A2(n11742), .ZN(n11582) );
  OAI211_X1 U14039 ( .C1(n13187), .C2(n11748), .A(n11582), .B(n11581), .ZN(
        n11587) );
  INV_X1 U14040 ( .A(n11583), .ZN(n11604) );
  AOI211_X1 U14041 ( .C1(n11585), .C2(n11584), .A(n13165), .B(n11604), .ZN(
        n11586) );
  AOI211_X1 U14042 ( .C1(n14046), .C2(n13173), .A(n11587), .B(n11586), .ZN(
        n11588) );
  INV_X1 U14043 ( .A(n11588), .ZN(P2_U3189) );
  INV_X1 U14044 ( .A(n11590), .ZN(n11592) );
  INV_X1 U14045 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U14046 ( .A1(n11595), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n11596) );
  XNOR2_X1 U14047 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n11940) );
  XNOR2_X1 U14048 ( .A(n11941), .B(n11940), .ZN(n11598) );
  AND2_X1 U14049 ( .A1(n11938), .A2(n11599), .ZN(n11601) );
  INV_X1 U14050 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15549) );
  INV_X1 U14051 ( .A(n11938), .ZN(n11600) );
  OAI22_X1 U14052 ( .A1(n11601), .A2(n15549), .B1(n11939), .B2(n11600), .ZN(
        SUB_1596_U69) );
  NOR3_X1 U14053 ( .A1(n11602), .A2(n13256), .A3(n13174), .ZN(n11603) );
  AOI21_X1 U14054 ( .B1(n11604), .B2(n13182), .A(n11603), .ZN(n11613) );
  INV_X1 U14055 ( .A(n11817), .ZN(n11607) );
  OAI22_X1 U14056 ( .A1(n13256), .A2(n13869), .B1(n13611), .B2(n13871), .ZN(
        n11812) );
  NAND2_X1 U14057 ( .A1(n13161), .A2(n11812), .ZN(n11606) );
  OAI211_X1 U14058 ( .C1(n13187), .C2(n11607), .A(n11606), .B(n11605), .ZN(
        n11610) );
  NOR2_X1 U14059 ( .A1(n11608), .A2(n13165), .ZN(n11609) );
  AOI211_X1 U14060 ( .C1(n14041), .C2(n13173), .A(n11610), .B(n11609), .ZN(
        n11611) );
  OAI21_X1 U14061 ( .B1(n11613), .B2(n11612), .A(n11611), .ZN(P2_U3208) );
  AOI21_X1 U14062 ( .B1(n11617), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11614), 
        .ZN(n11920) );
  XNOR2_X1 U14063 ( .A(n11920), .B(n11929), .ZN(n11615) );
  NOR2_X1 U14064 ( .A1(n11615), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11925) );
  AOI21_X1 U14065 ( .B1(n11615), .B2(P1_REG2_REG_15__SCAN_IN), .A(n11925), 
        .ZN(n11623) );
  XNOR2_X1 U14066 ( .A(n11928), .B(n11921), .ZN(n11931) );
  XNOR2_X1 U14067 ( .A(n11931), .B(n11930), .ZN(n11618) );
  NAND2_X1 U14068 ( .A1(n11618), .A2(n15188), .ZN(n11622) );
  NOR2_X1 U14069 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6904), .ZN(n11620) );
  NOR2_X1 U14070 ( .A1(n14633), .A2(n11929), .ZN(n11619) );
  AOI211_X1 U14071 ( .C1(n15199), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11620), 
        .B(n11619), .ZN(n11621) );
  OAI211_X1 U14072 ( .C1(n11623), .C2(n14637), .A(n11622), .B(n11621), .ZN(
        P1_U3258) );
  INV_X1 U14073 ( .A(n13935), .ZN(n11630) );
  INV_X1 U14074 ( .A(n13931), .ZN(n13853) );
  AOI22_X1 U14075 ( .A1(n13853), .A2(n13246), .B1(n13928), .B2(n11624), .ZN(
        n11625) );
  OAI21_X1 U14076 ( .B1(n11626), .B2(n13554), .A(n11625), .ZN(n11629) );
  MUX2_X1 U14077 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11627), .S(n13880), .Z(
        n11628) );
  AOI211_X1 U14078 ( .C1(n11631), .C2(n11630), .A(n11629), .B(n11628), .ZN(
        n11632) );
  INV_X1 U14079 ( .A(n11632), .ZN(P2_U3257) );
  MUX2_X1 U14080 ( .A(n11634), .B(n11633), .S(n13880), .Z(n11641) );
  INV_X1 U14081 ( .A(n11635), .ZN(n11636) );
  OAI22_X1 U14082 ( .A1(n13931), .A2(n11637), .B1(n13837), .B2(n11636), .ZN(
        n11638) );
  AOI21_X1 U14083 ( .B1(n11639), .B2(n13938), .A(n11638), .ZN(n11640) );
  OAI211_X1 U14084 ( .C1(n13935), .C2(n11642), .A(n11641), .B(n11640), .ZN(
        P2_U3259) );
  OR2_X1 U14085 ( .A1(n11644), .A2(n11643), .ZN(n11645) );
  NAND2_X1 U14086 ( .A1(n11646), .A2(n11645), .ZN(n11649) );
  INV_X1 U14087 ( .A(n11649), .ZN(n15372) );
  NOR2_X1 U14088 ( .A1(n11647), .A2(n13397), .ZN(n11648) );
  OAI21_X1 U14089 ( .B1(n6633), .B2(n11648), .A(n13905), .ZN(n11652) );
  AOI22_X1 U14090 ( .A1(n13885), .A2(n13446), .B1(n13448), .B2(n13883), .ZN(
        n11651) );
  NAND2_X1 U14091 ( .A1(n11649), .A2(n13802), .ZN(n11650) );
  AND3_X1 U14092 ( .A1(n11652), .A2(n11651), .A3(n11650), .ZN(n15370) );
  MUX2_X1 U14093 ( .A(n11653), .B(n15370), .S(n13880), .Z(n11661) );
  AOI211_X1 U14094 ( .C1(n15368), .C2(n11655), .A(n13926), .B(n7546), .ZN(
        n15367) );
  INV_X1 U14095 ( .A(n11656), .ZN(n11657) );
  OAI22_X1 U14096 ( .A1(n13931), .A2(n11658), .B1(n13837), .B2(n11657), .ZN(
        n11659) );
  AOI21_X1 U14097 ( .B1(n15367), .B2(n13938), .A(n11659), .ZN(n11660) );
  OAI211_X1 U14098 ( .C1(n15372), .C2(n13811), .A(n11661), .B(n11660), .ZN(
        P2_U3261) );
  NAND2_X1 U14099 ( .A1(n11662), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U14100 ( .A1(n11663), .A2(n11667), .ZN(n11664) );
  NAND2_X1 U14101 ( .A1(n11665), .A2(n11664), .ZN(n11695) );
  INV_X1 U14102 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13857) );
  XNOR2_X1 U14103 ( .A(n11696), .B(n13857), .ZN(n11694) );
  XNOR2_X1 U14104 ( .A(n11695), .B(n11694), .ZN(n11673) );
  XNOR2_X1 U14105 ( .A(n11696), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11690) );
  XOR2_X1 U14106 ( .A(n11690), .B(n11691), .Z(n11671) );
  NAND2_X1 U14107 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13109)
         );
  NAND2_X1 U14108 ( .A1(n15273), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n11669) );
  OAI211_X1 U14109 ( .C1(n15313), .C2(n11688), .A(n13109), .B(n11669), .ZN(
        n11670) );
  AOI21_X1 U14110 ( .B1(n11671), .B2(n15315), .A(n11670), .ZN(n11672) );
  OAI21_X1 U14111 ( .B1(n11673), .B2(n15294), .A(n11672), .ZN(P2_U3230) );
  INV_X1 U14112 ( .A(n11674), .ZN(n11687) );
  INV_X1 U14113 ( .A(n11675), .ZN(n11676) );
  NAND2_X1 U14114 ( .A1(n11676), .A2(n12518), .ZN(n11677) );
  XNOR2_X1 U14115 ( .A(n12203), .B(n11682), .ZN(n11869) );
  XOR2_X1 U14116 ( .A(n12517), .B(n11869), .Z(n11679) );
  OAI211_X1 U14117 ( .C1(n11680), .C2(n11679), .A(n11870), .B(n12436), .ZN(
        n11686) );
  OAI22_X1 U14118 ( .A1(n12451), .A2(n11682), .B1(n11681), .B2(n12499), .ZN(
        n11683) );
  AOI211_X1 U14119 ( .C1(n12497), .C2(n12516), .A(n11684), .B(n11683), .ZN(
        n11685) );
  OAI211_X1 U14120 ( .C1(n11687), .C2(n12027), .A(n11686), .B(n11685), .ZN(
        P3_U3161) );
  INV_X1 U14121 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11689) );
  INV_X1 U14122 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11692) );
  XNOR2_X1 U14123 ( .A(n13520), .B(n11692), .ZN(n13521) );
  XNOR2_X1 U14124 ( .A(n13522), .B(n13521), .ZN(n11703) );
  NAND2_X1 U14125 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13119)
         );
  OAI21_X1 U14126 ( .B1(n15313), .B2(n6808), .A(n13119), .ZN(n11693) );
  AOI21_X1 U14127 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15273), .A(n11693), 
        .ZN(n11702) );
  NAND2_X1 U14128 ( .A1(n11695), .A2(n11694), .ZN(n11698) );
  NAND2_X1 U14129 ( .A1(n11696), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11697) );
  NAND2_X1 U14130 ( .A1(n11698), .A2(n11697), .ZN(n11700) );
  MUX2_X1 U14131 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n13839), .S(n13520), .Z(
        n11699) );
  NAND2_X1 U14132 ( .A1(n11700), .A2(n11699), .ZN(n13515) );
  OAI211_X1 U14133 ( .C1(n11700), .C2(n11699), .A(n13515), .B(n15318), .ZN(
        n11701) );
  OAI211_X1 U14134 ( .C1(n11703), .C2(n15300), .A(n11702), .B(n11701), .ZN(
        P2_U3231) );
  OAI21_X1 U14135 ( .B1(n11705), .B2(n14443), .A(n11704), .ZN(n14962) );
  INV_X1 U14136 ( .A(n11325), .ZN(n11706) );
  INV_X1 U14137 ( .A(n14956), .ZN(n11707) );
  OAI21_X1 U14138 ( .B1(n11706), .B2(n11707), .A(n11829), .ZN(n14958) );
  OAI22_X1 U14139 ( .A1(n14958), .A2(n14929), .B1(n11707), .B2(n15259), .ZN(
        n11713) );
  NAND2_X1 U14140 ( .A1(n11709), .A2(n14443), .ZN(n11710) );
  NAND3_X1 U14141 ( .A1(n11708), .A2(n15251), .A3(n11710), .ZN(n11712) );
  AOI22_X1 U14142 ( .A1(n14491), .A2(n14897), .B1(n14880), .B2(n14493), .ZN(
        n11711) );
  NAND2_X1 U14143 ( .A1(n11712), .A2(n11711), .ZN(n14959) );
  AOI211_X1 U14144 ( .C1(n15263), .C2(n14962), .A(n11713), .B(n14959), .ZN(
        n11716) );
  NAND2_X1 U14145 ( .A1(n15264), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11714) );
  OAI21_X1 U14146 ( .B1(n11716), .B2(n15264), .A(n11714), .ZN(P1_U3483) );
  NAND2_X1 U14147 ( .A1(n15270), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11715) );
  OAI21_X1 U14148 ( .B1(n11716), .B2(n15270), .A(n11715), .ZN(P1_U3536) );
  NAND2_X1 U14149 ( .A1(n11718), .A2(n11717), .ZN(n11720) );
  NAND2_X1 U14150 ( .A1(n6403), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11719) );
  XOR2_X1 U14151 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n12524), .Z(n11735) );
  NOR2_X1 U14152 ( .A1(n11724), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n11725) );
  OAI21_X1 U14153 ( .B1(n11725), .B2(n6450), .A(n12688), .ZN(n11734) );
  INV_X1 U14154 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11942) );
  NAND2_X1 U14155 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12464)
         );
  OAI21_X1 U14156 ( .B1(n12655), .B2(n11942), .A(n12464), .ZN(n11731) );
  MUX2_X1 U14157 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13031), .Z(n12528) );
  XOR2_X1 U14158 ( .A(n12528), .B(n11732), .Z(n11728) );
  AOI21_X1 U14159 ( .B1(n6610), .B2(n11728), .A(n12532), .ZN(n11729) );
  NOR2_X1 U14160 ( .A1(n11729), .A2(n12705), .ZN(n11730) );
  AOI211_X1 U14161 ( .C1(n12661), .C2(n11732), .A(n11731), .B(n11730), .ZN(
        n11733) );
  OAI211_X1 U14162 ( .C1(n11735), .C2(n12543), .A(n11734), .B(n11733), .ZN(
        P3_U3193) );
  XNOR2_X2 U14163 ( .A(n14046), .B(n13256), .ZN(n13563) );
  INV_X1 U14164 ( .A(n13443), .ZN(n11736) );
  OR2_X1 U14165 ( .A1(n13246), .A2(n11736), .ZN(n11737) );
  NAND2_X1 U14166 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  NAND2_X1 U14167 ( .A1(n11739), .A2(n7830), .ZN(n13555) );
  XNOR2_X1 U14168 ( .A(n14051), .B(n13556), .ZN(n13406) );
  NOR2_X1 U14169 ( .A1(n13555), .A2(n13406), .ZN(n11788) );
  OR2_X1 U14170 ( .A1(n14051), .A2(n13556), .ZN(n13562) );
  INV_X1 U14171 ( .A(n13562), .ZN(n11740) );
  NOR2_X1 U14172 ( .A1(n11788), .A2(n11740), .ZN(n11741) );
  NOR2_X1 U14173 ( .A1(n11741), .A2(n13563), .ZN(n11810) );
  AOI211_X1 U14174 ( .C1(n13563), .C2(n11741), .A(n13920), .B(n11810), .ZN(
        n11743) );
  NOR2_X1 U14175 ( .A1(n11743), .A2(n11742), .ZN(n14048) );
  NAND2_X1 U14176 ( .A1(n13246), .A2(n13443), .ZN(n11744) );
  NAND2_X1 U14177 ( .A1(n11745), .A2(n11744), .ZN(n11787) );
  NAND2_X1 U14178 ( .A1(n11787), .A2(n13406), .ZN(n11786) );
  NAND2_X1 U14179 ( .A1(n14051), .A2(n13442), .ZN(n11746) );
  OAI21_X1 U14180 ( .B1(n11747), .B2(n13563), .A(n11819), .ZN(n14049) );
  OAI22_X1 U14181 ( .A1(n13880), .A2(n10666), .B1(n11748), .B2(n13837), .ZN(
        n11749) );
  AOI21_X1 U14182 ( .B1(n14046), .B2(n13853), .A(n11749), .ZN(n11753) );
  OR2_X2 U14183 ( .A1(n11793), .A2(n14051), .ZN(n11791) );
  NOR2_X4 U14184 ( .A1(n11791), .A2(n14046), .ZN(n11814) );
  NAND2_X1 U14185 ( .A1(n11791), .A2(n14046), .ZN(n11750) );
  NAND2_X1 U14186 ( .A1(n11750), .A2(n13889), .ZN(n11751) );
  NOR2_X1 U14187 ( .A1(n11814), .A2(n11751), .ZN(n14045) );
  NAND2_X1 U14188 ( .A1(n14045), .A2(n13938), .ZN(n11752) );
  OAI211_X1 U14189 ( .C1(n14049), .C2(n13935), .A(n11753), .B(n11752), .ZN(
        n11754) );
  INV_X1 U14190 ( .A(n11754), .ZN(n11755) );
  OAI21_X1 U14191 ( .B1(n14048), .B2(n13940), .A(n11755), .ZN(P2_U3255) );
  INV_X1 U14192 ( .A(n11756), .ZN(n11763) );
  INV_X1 U14193 ( .A(n11757), .ZN(n11758) );
  MUX2_X1 U14194 ( .A(n7417), .B(n11758), .S(n12896), .Z(n11761) );
  AOI22_X1 U14195 ( .A1(n12855), .A2(n11759), .B1(n12873), .B2(n11879), .ZN(
        n11760) );
  OAI211_X1 U14196 ( .C1(n11763), .C2(n11762), .A(n11761), .B(n11760), .ZN(
        P3_U3224) );
  XNOR2_X1 U14197 ( .A(n11764), .B(n11765), .ZN(n11770) );
  INV_X1 U14198 ( .A(n13611), .ZN(n13440) );
  AOI22_X1 U14199 ( .A1(n13568), .A2(n13885), .B1(n13883), .B2(n13440), .ZN(
        n13908) );
  NAND2_X1 U14200 ( .A1(n13170), .A2(n13910), .ZN(n11767) );
  OAI211_X1 U14201 ( .C1(n13120), .C2(n13908), .A(n11767), .B(n11766), .ZN(
        n11768) );
  AOI21_X1 U14202 ( .B1(n14031), .B2(n13173), .A(n11768), .ZN(n11769) );
  OAI21_X1 U14203 ( .B1(n11770), .B2(n13165), .A(n11769), .ZN(P2_U3206) );
  MUX2_X1 U14204 ( .A(n11772), .B(n11771), .S(n15589), .Z(n11773) );
  OAI21_X1 U14205 ( .B1(n12905), .B2(n11882), .A(n11773), .ZN(P3_U3468) );
  XNOR2_X1 U14206 ( .A(n11774), .B(n11776), .ZN(n11968) );
  XNOR2_X1 U14207 ( .A(n11775), .B(n11776), .ZN(n11780) );
  NAND2_X1 U14208 ( .A1(n11968), .A2(n11777), .ZN(n11779) );
  AOI22_X1 U14209 ( .A1(n12515), .A2(n12879), .B1(n12880), .B2(n12516), .ZN(
        n11778) );
  OAI211_X1 U14210 ( .C1(n12045), .C2(n11780), .A(n11779), .B(n11778), .ZN(
        n11965) );
  AOI21_X1 U14211 ( .B1(n15425), .B2(n11968), .A(n11965), .ZN(n11949) );
  INV_X1 U14212 ( .A(n12022), .ZN(n11781) );
  AOI22_X1 U14213 ( .A1(n13007), .A2(n11781), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15429), .ZN(n11782) );
  OAI21_X1 U14214 ( .B1(n11949), .B2(n15429), .A(n11782), .ZN(P3_U3420) );
  INV_X1 U14215 ( .A(n11783), .ZN(n11839) );
  OAI222_X1 U14216 ( .A1(P2_U3088), .A2(n11785), .B1(n14092), .B2(n11839), 
        .C1(n11784), .C2(n14097), .ZN(P2_U3301) );
  OAI21_X1 U14217 ( .B1(n13406), .B2(n11787), .A(n11786), .ZN(n14054) );
  AOI211_X1 U14218 ( .C1(n13406), .C2(n13555), .A(n13920), .B(n11788), .ZN(
        n11790) );
  NOR2_X1 U14219 ( .A1(n11790), .A2(n11789), .ZN(n14053) );
  MUX2_X1 U14220 ( .A(n10287), .B(n14053), .S(n13880), .Z(n11797) );
  INV_X1 U14221 ( .A(n11791), .ZN(n11792) );
  AOI211_X1 U14222 ( .C1(n14051), .C2(n11793), .A(n11792), .B(n13926), .ZN(
        n14050) );
  INV_X1 U14223 ( .A(n14051), .ZN(n13253) );
  OAI22_X1 U14224 ( .A1(n13931), .A2(n13253), .B1(n11794), .B2(n13837), .ZN(
        n11795) );
  AOI21_X1 U14225 ( .B1(n14050), .B2(n13938), .A(n11795), .ZN(n11796) );
  OAI211_X1 U14226 ( .C1(n13935), .C2(n14054), .A(n11797), .B(n11796), .ZN(
        P2_U3256) );
  XOR2_X1 U14227 ( .A(n11798), .B(n11800), .Z(n11885) );
  AOI22_X1 U14228 ( .A1(n12855), .A2(n12469), .B1(n12873), .B2(n12468), .ZN(
        n11806) );
  INV_X1 U14229 ( .A(n11800), .ZN(n11801) );
  XNOR2_X1 U14230 ( .A(n11799), .B(n11801), .ZN(n11804) );
  NAND2_X1 U14231 ( .A1(n12880), .A2(n12162), .ZN(n11802) );
  OAI21_X1 U14232 ( .B1(n12450), .B2(n12048), .A(n11802), .ZN(n11803) );
  AOI21_X1 U14233 ( .B1(n11804), .B2(n12883), .A(n11803), .ZN(n11889) );
  MUX2_X1 U14234 ( .A(n7409), .B(n11889), .S(n12896), .Z(n11805) );
  OAI211_X1 U14235 ( .C1(n11885), .C2(n12876), .A(n11806), .B(n11805), .ZN(
        P3_U3222) );
  INV_X1 U14236 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11807) );
  MUX2_X1 U14237 ( .A(n11807), .B(n11889), .S(n15589), .Z(n11809) );
  NAND2_X1 U14238 ( .A1(n12939), .A2(n12469), .ZN(n11808) );
  OAI211_X1 U14239 ( .C1(n11885), .C2(n12941), .A(n11809), .B(n11808), .ZN(
        P3_U3470) );
  INV_X1 U14240 ( .A(n13256), .ZN(n13441) );
  AND2_X1 U14241 ( .A1(n11577), .A2(n13441), .ZN(n13560) );
  NOR2_X1 U14242 ( .A1(n11810), .A2(n13560), .ZN(n11811) );
  XNOR2_X1 U14243 ( .A(n14041), .B(n13566), .ZN(n13408) );
  NAND2_X1 U14244 ( .A1(n11811), .A2(n13408), .ZN(n13902) );
  OAI21_X1 U14245 ( .B1(n11811), .B2(n13408), .A(n13902), .ZN(n11813) );
  AOI21_X1 U14246 ( .B1(n11813), .B2(n13905), .A(n11812), .ZN(n14043) );
  INV_X1 U14247 ( .A(n11814), .ZN(n11816) );
  INV_X1 U14248 ( .A(n13927), .ZN(n11815) );
  AOI211_X1 U14249 ( .C1(n14041), .C2(n11816), .A(n13926), .B(n11815), .ZN(
        n14040) );
  AOI22_X1 U14250 ( .A1(n13940), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11817), 
        .B2(n13928), .ZN(n11818) );
  OAI21_X1 U14251 ( .B1(n13609), .B2(n13931), .A(n11818), .ZN(n11821) );
  XOR2_X1 U14252 ( .A(n13607), .B(n13408), .Z(n14044) );
  NOR2_X1 U14253 ( .A1(n14044), .A2(n13915), .ZN(n11820) );
  AOI211_X1 U14254 ( .C1(n14040), .C2(n13938), .A(n11821), .B(n11820), .ZN(
        n11822) );
  OAI21_X1 U14255 ( .B1(n14043), .B2(n13940), .A(n11822), .ZN(P2_U3254) );
  AOI21_X1 U14256 ( .B1(n14447), .B2(n11824), .A(n6964), .ZN(n11825) );
  OAI222_X1 U14257 ( .A1(n14933), .A2(n14306), .B1(n14935), .B2(n11826), .C1(
        n15050), .C2(n11825), .ZN(n11973) );
  INV_X1 U14258 ( .A(n11973), .ZN(n11838) );
  OAI21_X1 U14259 ( .B1(n11828), .B2(n14447), .A(n11827), .ZN(n11975) );
  INV_X1 U14260 ( .A(n14295), .ZN(n11832) );
  INV_X1 U14261 ( .A(n11829), .ZN(n11831) );
  INV_X1 U14262 ( .A(n11857), .ZN(n11830) );
  OAI211_X1 U14263 ( .C1(n11832), .C2(n11831), .A(n11830), .B(n15216), .ZN(
        n11972) );
  OAI22_X1 U14264 ( .A1(n15220), .A2(n11833), .B1(n11906), .B2(n15217), .ZN(
        n11834) );
  AOI21_X1 U14265 ( .B1(n15223), .B2(n14295), .A(n11834), .ZN(n11835) );
  OAI21_X1 U14266 ( .B1(n11972), .B2(n15225), .A(n11835), .ZN(n11836) );
  AOI21_X1 U14267 ( .B1(n11975), .B2(n15227), .A(n11836), .ZN(n11837) );
  OAI21_X1 U14268 ( .B1(n11838), .B2(n6412), .A(n11837), .ZN(P1_U3284) );
  OAI222_X1 U14269 ( .A1(n15105), .A2(n15483), .B1(P1_U3086), .B2(n11840), 
        .C1(n10976), .C2(n11839), .ZN(P1_U3329) );
  AOI22_X1 U14270 ( .A1(n14956), .A2(n12315), .B1(n14492), .B2(n10744), .ZN(
        n11894) );
  NAND2_X1 U14271 ( .A1(n14956), .A2(n12316), .ZN(n11842) );
  NAND2_X1 U14272 ( .A1(n14492), .A2(n12315), .ZN(n11841) );
  NAND2_X1 U14273 ( .A1(n11842), .A2(n11841), .ZN(n11843) );
  XNOR2_X1 U14274 ( .A(n11843), .B(n12313), .ZN(n11893) );
  XOR2_X1 U14275 ( .A(n11894), .B(n11893), .Z(n11897) );
  INV_X1 U14276 ( .A(n11844), .ZN(n11846) );
  OR2_X1 U14277 ( .A1(n11898), .A2(n11897), .ZN(n11896) );
  INV_X1 U14278 ( .A(n11896), .ZN(n11848) );
  AOI21_X1 U14279 ( .B1(n11897), .B2(n11898), .A(n11848), .ZN(n11854) );
  OAI22_X1 U14280 ( .A1(n14236), .A2(n11866), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11849), .ZN(n11850) );
  AOI21_X1 U14281 ( .B1(n14239), .B2(n14493), .A(n11850), .ZN(n11851) );
  OAI21_X1 U14282 ( .B1(n14954), .B2(n15182), .A(n11851), .ZN(n11852) );
  AOI21_X1 U14283 ( .B1(n14221), .B2(n14956), .A(n11852), .ZN(n11853) );
  OAI21_X1 U14284 ( .B1(n11854), .B2(n15174), .A(n11853), .ZN(P1_U3221) );
  NAND2_X1 U14285 ( .A1(n11855), .A2(n14448), .ZN(n11955) );
  OAI21_X1 U14286 ( .B1(n11855), .B2(n14448), .A(n11955), .ZN(n11856) );
  INV_X1 U14287 ( .A(n11856), .ZN(n15081) );
  OAI21_X1 U14288 ( .B1(n11857), .B2(n14305), .A(n15216), .ZN(n11859) );
  NAND2_X1 U14289 ( .A1(n14897), .A2(n14489), .ZN(n12006) );
  OAI21_X1 U14290 ( .B1(n11859), .B2(n11858), .A(n12006), .ZN(n15078) );
  NOR2_X1 U14291 ( .A1(n14921), .A2(n14305), .ZN(n11861) );
  OAI22_X1 U14292 ( .A1(n15220), .A2(n10458), .B1(n12007), .B2(n15217), .ZN(
        n11860) );
  AOI211_X1 U14293 ( .C1(n15078), .C2(n14907), .A(n11861), .B(n11860), .ZN(
        n11868) );
  OAI211_X1 U14294 ( .C1(n11864), .C2(n11863), .A(n11862), .B(n15251), .ZN(
        n11865) );
  OAI21_X1 U14295 ( .B1(n11866), .B2(n14935), .A(n11865), .ZN(n15077) );
  NAND2_X1 U14296 ( .A1(n15077), .A2(n15220), .ZN(n11867) );
  OAI211_X1 U14297 ( .C1(n15081), .C2(n14910), .A(n11868), .B(n11867), .ZN(
        P1_U3283) );
  XNOR2_X1 U14298 ( .A(n12203), .B(n11882), .ZN(n12012) );
  XNOR2_X1 U14299 ( .A(n12012), .B(n12516), .ZN(n11872) );
  NAND2_X1 U14300 ( .A1(n11873), .A2(n11872), .ZN(n11874) );
  AOI21_X1 U14301 ( .B1(n12014), .B2(n11874), .A(n12506), .ZN(n11884) );
  NAND2_X1 U14302 ( .A1(n12497), .A2(n12162), .ZN(n11876) );
  OAI211_X1 U14303 ( .C1(n11877), .C2(n12499), .A(n11876), .B(n11875), .ZN(
        n11878) );
  INV_X1 U14304 ( .A(n11878), .ZN(n11881) );
  NAND2_X1 U14305 ( .A1(n12502), .A2(n11879), .ZN(n11880) );
  OAI211_X1 U14306 ( .C1(n12451), .C2(n11882), .A(n11881), .B(n11880), .ZN(
        n11883) );
  OR2_X1 U14307 ( .A1(n11884), .A2(n11883), .ZN(P3_U3171) );
  INV_X1 U14308 ( .A(n11885), .ZN(n11886) );
  INV_X1 U14309 ( .A(n13010), .ZN(n11988) );
  NAND2_X1 U14310 ( .A1(n11886), .A2(n11988), .ZN(n11888) );
  AOI22_X1 U14311 ( .A1(n13007), .A2(n12469), .B1(n15429), .B2(
        P3_REG0_REG_11__SCAN_IN), .ZN(n11887) );
  OAI211_X1 U14312 ( .C1(n15429), .C2(n11889), .A(n11888), .B(n11887), .ZN(
        P3_U3423) );
  NAND2_X1 U14313 ( .A1(n14295), .A2(n15255), .ZN(n11971) );
  NAND2_X1 U14314 ( .A1(n14295), .A2(n12316), .ZN(n11891) );
  NAND2_X1 U14315 ( .A1(n14491), .A2(n12315), .ZN(n11890) );
  NAND2_X1 U14316 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  XNOR2_X1 U14317 ( .A(n11892), .B(n12313), .ZN(n11994) );
  AOI22_X1 U14318 ( .A1(n14295), .A2(n12315), .B1(n10744), .B2(n14491), .ZN(
        n11995) );
  XNOR2_X1 U14319 ( .A(n11994), .B(n11995), .ZN(n11904) );
  INV_X1 U14320 ( .A(n11893), .ZN(n11895) );
  NAND2_X1 U14321 ( .A1(n11895), .A2(n11894), .ZN(n11899) );
  NAND2_X1 U14322 ( .A1(n11896), .A2(n11899), .ZN(n11903) );
  INV_X1 U14323 ( .A(n11904), .ZN(n11900) );
  OR2_X1 U14324 ( .A1(n11900), .A2(n11899), .ZN(n11901) );
  INV_X1 U14325 ( .A(n11901), .ZN(n11902) );
  OAI21_X1 U14326 ( .B1(n11904), .B2(n11903), .A(n11997), .ZN(n11905) );
  NAND2_X1 U14327 ( .A1(n11905), .A2(n14232), .ZN(n11910) );
  NOR2_X1 U14328 ( .A1(n15182), .A2(n11906), .ZN(n11908) );
  NAND2_X1 U14329 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14565) );
  OAI21_X1 U14330 ( .B1(n14236), .B2(n14306), .A(n14565), .ZN(n11907) );
  AOI211_X1 U14331 ( .C1(n14239), .C2(n14492), .A(n11908), .B(n11907), .ZN(
        n11909) );
  OAI211_X1 U14332 ( .C1(n14231), .C2(n11971), .A(n11910), .B(n11909), .ZN(
        P1_U3231) );
  XOR2_X1 U14333 ( .A(n11911), .B(n11913), .Z(n11987) );
  INV_X1 U14334 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15452) );
  XNOR2_X1 U14335 ( .A(n11912), .B(n9882), .ZN(n11915) );
  OAI22_X1 U14336 ( .A1(n12386), .A2(n12144), .B1(n12344), .B2(n12048), .ZN(
        n11914) );
  AOI21_X1 U14337 ( .B1(n11915), .B2(n12883), .A(n11914), .ZN(n11993) );
  MUX2_X1 U14338 ( .A(n15452), .B(n11993), .S(n15589), .Z(n11917) );
  INV_X1 U14339 ( .A(n12387), .ZN(n11990) );
  NAND2_X1 U14340 ( .A1(n11990), .A2(n12939), .ZN(n11916) );
  OAI211_X1 U14341 ( .C1(n11987), .C2(n12941), .A(n11917), .B(n11916), .ZN(
        P3_U3471) );
  AOI22_X1 U14342 ( .A1(n11990), .A2(n12855), .B1(n12873), .B2(n12390), .ZN(
        n11919) );
  INV_X1 U14343 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12546) );
  MUX2_X1 U14344 ( .A(n12546), .B(n11993), .S(n12896), .Z(n11918) );
  OAI211_X1 U14345 ( .C1(n11987), .C2(n12876), .A(n11919), .B(n11918), .ZN(
        P3_U3221) );
  INV_X1 U14346 ( .A(n11920), .ZN(n11922) );
  NOR2_X1 U14347 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  XNOR2_X1 U14348 ( .A(n14593), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n11923) );
  NOR3_X1 U14349 ( .A1(n11925), .A2(n11924), .A3(n11923), .ZN(n14596) );
  INV_X1 U14350 ( .A(n14596), .ZN(n11927) );
  OAI21_X1 U14351 ( .B1(n11925), .B2(n11924), .A(n11923), .ZN(n11926) );
  NAND3_X1 U14352 ( .A1(n11927), .A2(n15194), .A3(n11926), .ZN(n11937) );
  NAND2_X1 U14353 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14160)
         );
  XOR2_X1 U14354 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14593), .Z(n11933) );
  AOI22_X1 U14355 ( .A1(n11931), .A2(n11930), .B1(n11929), .B2(n11928), .ZN(
        n11932) );
  OAI211_X1 U14356 ( .C1(n11933), .C2(n11932), .A(n15188), .B(n14599), .ZN(
        n11934) );
  NAND2_X1 U14357 ( .A1(n14160), .A2(n11934), .ZN(n11935) );
  AOI21_X1 U14358 ( .B1(n15199), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11935), 
        .ZN(n11936) );
  OAI211_X1 U14359 ( .C1(n14633), .C2(n14601), .A(n11937), .B(n11936), .ZN(
        P1_U3259) );
  NAND2_X1 U14360 ( .A1(n11941), .A2(n11940), .ZN(n11944) );
  NAND2_X1 U14361 ( .A1(n11942), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U14362 ( .A1(n11944), .A2(n11943), .ZN(n11982) );
  XNOR2_X1 U14363 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n11945) );
  XNOR2_X1 U14364 ( .A(n11982), .B(n11945), .ZN(n11946) );
  NAND2_X1 U14365 ( .A1(n11979), .A2(n11980), .ZN(n11948) );
  XNOR2_X1 U14366 ( .A(n11948), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  MUX2_X1 U14367 ( .A(n11950), .B(n11949), .S(n15589), .Z(n11951) );
  OAI21_X1 U14368 ( .B1(n12905), .B2(n12022), .A(n11951), .ZN(P3_U3469) );
  XNOR2_X1 U14369 ( .A(n11952), .B(n14449), .ZN(n11953) );
  AOI222_X1 U14370 ( .A1(n15251), .A2(n11953), .B1(n14488), .B2(n14897), .C1(
        n14490), .C2(n14880), .ZN(n15076) );
  NAND2_X1 U14371 ( .A1(n11955), .A2(n11954), .ZN(n11957) );
  OAI21_X1 U14372 ( .B1(n11957), .B2(n14449), .A(n14939), .ZN(n15072) );
  OAI211_X1 U14373 ( .C1(n11858), .C2(n14302), .A(n15216), .B(n11958), .ZN(
        n15073) );
  INV_X1 U14374 ( .A(n11959), .ZN(n14210) );
  AOI22_X1 U14375 ( .A1(n6412), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n14210), 
        .B2(n14974), .ZN(n11961) );
  NAND2_X1 U14376 ( .A1(n14303), .A2(n15223), .ZN(n11960) );
  OAI211_X1 U14377 ( .C1(n15073), .C2(n15225), .A(n11961), .B(n11960), .ZN(
        n11962) );
  AOI21_X1 U14378 ( .B1(n15072), .B2(n15227), .A(n11962), .ZN(n11963) );
  OAI21_X1 U14379 ( .B1(n15076), .B2(n6412), .A(n11963), .ZN(P1_U3282) );
  INV_X1 U14380 ( .A(n11964), .ZN(n12028) );
  OAI22_X1 U14381 ( .A1(n12867), .A2(n12022), .B1(n12028), .B2(n12891), .ZN(
        n11967) );
  MUX2_X1 U14382 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n11965), .S(n12896), .Z(
        n11966) );
  AOI211_X1 U14383 ( .C1(n11969), .C2(n11968), .A(n11967), .B(n11966), .ZN(
        n11970) );
  INV_X1 U14384 ( .A(n11970), .ZN(P3_U3223) );
  NAND2_X1 U14385 ( .A1(n11972), .A2(n11971), .ZN(n11974) );
  AOI211_X1 U14386 ( .C1(n15263), .C2(n11975), .A(n11974), .B(n11973), .ZN(
        n11978) );
  NAND2_X1 U14387 ( .A1(n15270), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11976) );
  OAI21_X1 U14388 ( .B1(n11978), .B2(n15270), .A(n11976), .ZN(P1_U3537) );
  NAND2_X1 U14389 ( .A1(n15264), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11977) );
  OAI21_X1 U14390 ( .B1(n11978), .B2(n15264), .A(n11977), .ZN(P1_U3486) );
  INV_X1 U14391 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15308) );
  NOR2_X1 U14392 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n15510), .ZN(n11981) );
  NAND2_X1 U14393 ( .A1(n15510), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11983) );
  INV_X1 U14394 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15113) );
  XNOR2_X1 U14395 ( .A(n15113), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n11985) );
  XNOR2_X1 U14396 ( .A(n15115), .B(n11985), .ZN(n15110) );
  XNOR2_X1 U14397 ( .A(n15110), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(n11986) );
  XNOR2_X1 U14398 ( .A(n15112), .B(n11986), .ZN(SUB_1596_U67) );
  INV_X1 U14399 ( .A(n11987), .ZN(n11989) );
  NAND2_X1 U14400 ( .A1(n11989), .A2(n11988), .ZN(n11992) );
  AOI22_X1 U14401 ( .A1(n11990), .A2(n13007), .B1(P3_REG0_REG_12__SCAN_IN), 
        .B2(n15429), .ZN(n11991) );
  OAI211_X1 U14402 ( .C1(n15429), .C2(n11993), .A(n11992), .B(n11991), .ZN(
        P3_U3426) );
  INV_X1 U14403 ( .A(n11994), .ZN(n11996) );
  NOR2_X1 U14404 ( .A1(n14306), .A2(n6416), .ZN(n11998) );
  AOI21_X1 U14405 ( .B1(n15079), .B2(n12315), .A(n11998), .ZN(n12077) );
  NAND2_X1 U14406 ( .A1(n15079), .A2(n12316), .ZN(n12000) );
  NAND2_X1 U14407 ( .A1(n12315), .A2(n14490), .ZN(n11999) );
  NAND2_X1 U14408 ( .A1(n12000), .A2(n11999), .ZN(n12001) );
  XNOR2_X1 U14409 ( .A(n12001), .B(n12313), .ZN(n12076) );
  XOR2_X1 U14410 ( .A(n12077), .B(n12076), .Z(n12002) );
  AOI21_X1 U14411 ( .B1(n12003), .B2(n12002), .A(n15174), .ZN(n12004) );
  NAND2_X1 U14412 ( .A1(n12004), .A2(n12080), .ZN(n12011) );
  OAI21_X1 U14413 ( .B1(n14198), .B2(n12006), .A(n12005), .ZN(n12009) );
  NOR2_X1 U14414 ( .A1(n15182), .A2(n12007), .ZN(n12008) );
  AOI211_X1 U14415 ( .C1(n14239), .C2(n14491), .A(n12009), .B(n12008), .ZN(
        n12010) );
  OAI211_X1 U14416 ( .C1(n14305), .C2(n14242), .A(n12011), .B(n12010), .ZN(
        P1_U3217) );
  XNOR2_X1 U14417 ( .A(n12022), .B(n12203), .ZN(n12163) );
  XNOR2_X1 U14418 ( .A(n12163), .B(n12162), .ZN(n12016) );
  AOI21_X1 U14419 ( .B1(n12015), .B2(n12016), .A(n12506), .ZN(n12019) );
  NAND2_X1 U14420 ( .A1(n12019), .A2(n12165), .ZN(n12026) );
  OAI21_X1 U14421 ( .B1(n12499), .B2(n12021), .A(n12020), .ZN(n12024) );
  NOR2_X1 U14422 ( .A1(n12451), .A2(n12022), .ZN(n12023) );
  AOI211_X1 U14423 ( .C1(n12497), .C2(n12515), .A(n12024), .B(n12023), .ZN(
        n12025) );
  OAI211_X1 U14424 ( .C1(n12028), .C2(n12027), .A(n12026), .B(n12025), .ZN(
        P3_U3157) );
  XOR2_X1 U14425 ( .A(n12029), .B(n12034), .Z(n12875) );
  INV_X1 U14426 ( .A(n12868), .ZN(n12039) );
  INV_X1 U14427 ( .A(n12032), .ZN(n12033) );
  AOI21_X1 U14428 ( .B1(n12034), .B2(n12030), .A(n12033), .ZN(n12035) );
  OAI222_X1 U14429 ( .A1(n12048), .A2(n12500), .B1(n12144), .B2(n12450), .C1(
        n12045), .C2(n12035), .ZN(n12869) );
  MUX2_X1 U14430 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12869), .S(n15589), .Z(
        n12036) );
  AOI21_X1 U14431 ( .B1(n12939), .B2(n12039), .A(n12036), .ZN(n12037) );
  OAI21_X1 U14432 ( .B1(n12941), .B2(n12875), .A(n12037), .ZN(P3_U3472) );
  MUX2_X1 U14433 ( .A(P3_REG0_REG_13__SCAN_IN), .B(n12869), .S(n15431), .Z(
        n12038) );
  AOI21_X1 U14434 ( .B1(n13007), .B2(n12039), .A(n12038), .ZN(n12040) );
  OAI21_X1 U14435 ( .B1(n13010), .B2(n12875), .A(n12040), .ZN(P3_U3429) );
  INV_X1 U14436 ( .A(n12041), .ZN(n12042) );
  AOI21_X1 U14437 ( .B1(n6890), .B2(n12043), .A(n12042), .ZN(n12946) );
  INV_X1 U14438 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12575) );
  INV_X1 U14439 ( .A(n12346), .ZN(n12044) );
  OAI22_X1 U14440 ( .A1(n12896), .A2(n12575), .B1(n12044), .B2(n12891), .ZN(
        n12053) );
  AOI21_X1 U14441 ( .B1(n12047), .B2(n12046), .A(n12045), .ZN(n12051) );
  OAI22_X1 U14442 ( .A1(n12405), .A2(n12048), .B1(n12344), .B2(n12144), .ZN(
        n12049) );
  AOI21_X1 U14443 ( .B1(n12051), .B2(n12050), .A(n12049), .ZN(n12944) );
  NOR2_X1 U14444 ( .A1(n12944), .A2(n12863), .ZN(n12052) );
  AOI211_X1 U14445 ( .C1(n12855), .C2(n12942), .A(n12053), .B(n12052), .ZN(
        n12054) );
  OAI21_X1 U14446 ( .B1(n12946), .B2(n12876), .A(n12054), .ZN(P3_U3219) );
  INV_X1 U14448 ( .A(n12057), .ZN(n12058) );
  OAI222_X1 U14449 ( .A1(n13034), .A2(n12059), .B1(P3_U3151), .B2(n12056), 
        .C1(n13039), .C2(n12058), .ZN(P3_U3265) );
  NAND2_X1 U14450 ( .A1(n15429), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12063) );
  OR2_X1 U14451 ( .A1(n13027), .A2(n12060), .ZN(n12061) );
  NAND2_X1 U14452 ( .A1(n12879), .A2(n12061), .ZN(n12142) );
  NAND2_X1 U14453 ( .A1(n12066), .A2(n15431), .ZN(n12948) );
  OAI211_X1 U14454 ( .C1(n12068), .C2(n12949), .A(n12063), .B(n12948), .ZN(
        P3_U3457) );
  NAND2_X1 U14455 ( .A1(n15440), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U14456 ( .A1(n12066), .A2(n15589), .ZN(n12899) );
  OAI211_X1 U14457 ( .C1(n12068), .C2(n12905), .A(n12064), .B(n12899), .ZN(
        P3_U3489) );
  NOR2_X1 U14458 ( .A1(n12065), .A2(n12891), .ZN(n12151) );
  AOI21_X1 U14459 ( .B1(n12066), .B2(n12896), .A(n12151), .ZN(n12711) );
  NAND2_X1 U14460 ( .A1(n12863), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12067) );
  OAI211_X1 U14461 ( .C1(n12068), .C2(n12867), .A(n12711), .B(n12067), .ZN(
        P3_U3203) );
  OAI222_X1 U14462 ( .A1(n12071), .A2(P3_U3151), .B1(n13039), .B2(n12070), 
        .C1(n12069), .C2(n13034), .ZN(P3_U3270) );
  INV_X1 U14463 ( .A(n13342), .ZN(n14091) );
  OAI222_X1 U14464 ( .A1(n10976), .A2(n14091), .B1(P1_U3086), .B2(n9332), .C1(
        n12072), .C2(n15105), .ZN(P1_U3326) );
  NAND2_X1 U14465 ( .A1(n15053), .A2(n12316), .ZN(n12074) );
  NAND2_X1 U14466 ( .A1(n14896), .A2(n12315), .ZN(n12073) );
  NAND2_X1 U14467 ( .A1(n12074), .A2(n12073), .ZN(n12075) );
  XNOR2_X1 U14468 ( .A(n12075), .B(n12313), .ZN(n12126) );
  INV_X1 U14469 ( .A(n12126), .ZN(n12114) );
  INV_X1 U14470 ( .A(n12077), .ZN(n12078) );
  NAND2_X1 U14471 ( .A1(n14303), .A2(n12316), .ZN(n12082) );
  NAND2_X1 U14472 ( .A1(n12315), .A2(n14489), .ZN(n12081) );
  NAND2_X1 U14473 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  XNOR2_X1 U14474 ( .A(n12083), .B(n12313), .ZN(n12086) );
  OAI22_X1 U14475 ( .A1(n14302), .A2(n6401), .B1(n14936), .B2(n6416), .ZN(
        n12087) );
  XNOR2_X1 U14476 ( .A(n12086), .B(n12087), .ZN(n14205) );
  INV_X1 U14477 ( .A(n12086), .ZN(n12089) );
  INV_X1 U14478 ( .A(n12087), .ZN(n12088) );
  NAND2_X1 U14479 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  NOR2_X1 U14480 ( .A1(n14301), .A2(n6416), .ZN(n12091) );
  AOI21_X1 U14481 ( .B1(n14951), .B2(n12315), .A(n12091), .ZN(n12096) );
  NAND2_X1 U14482 ( .A1(n14951), .A2(n12316), .ZN(n12093) );
  NAND2_X1 U14483 ( .A1(n12315), .A2(n14488), .ZN(n12092) );
  NAND2_X1 U14484 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  XNOR2_X1 U14485 ( .A(n12094), .B(n12313), .ZN(n12095) );
  XOR2_X1 U14486 ( .A(n12096), .B(n12095), .Z(n14142) );
  INV_X1 U14487 ( .A(n12095), .ZN(n12097) );
  NOR2_X1 U14488 ( .A1(n14934), .A2(n6416), .ZN(n12098) );
  AOI21_X1 U14489 ( .B1(n15065), .B2(n12315), .A(n12098), .ZN(n12101) );
  AOI22_X1 U14490 ( .A1(n15065), .A2(n12316), .B1(n12315), .B2(n14487), .ZN(
        n12099) );
  XNOR2_X1 U14491 ( .A(n12099), .B(n12313), .ZN(n12100) );
  XOR2_X1 U14492 ( .A(n12101), .B(n12100), .Z(n14188) );
  NAND2_X1 U14493 ( .A1(n14189), .A2(n14188), .ZN(n14187) );
  INV_X1 U14494 ( .A(n12100), .ZN(n12103) );
  INV_X1 U14495 ( .A(n12101), .ZN(n12102) );
  NAND2_X1 U14496 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  AOI22_X1 U14497 ( .A1(n14901), .A2(n12315), .B1(n10744), .B2(n14879), .ZN(
        n12109) );
  NAND2_X1 U14498 ( .A1(n14901), .A2(n12316), .ZN(n12106) );
  NAND2_X1 U14499 ( .A1(n12315), .A2(n14879), .ZN(n12105) );
  NAND2_X1 U14500 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  XNOR2_X1 U14501 ( .A(n12107), .B(n12313), .ZN(n12108) );
  XOR2_X1 U14502 ( .A(n12109), .B(n12108), .Z(n14110) );
  INV_X1 U14503 ( .A(n12108), .ZN(n12110) );
  NAND2_X1 U14504 ( .A1(n12110), .A2(n12109), .ZN(n12111) );
  XNOR2_X1 U14505 ( .A(n12125), .B(n12126), .ZN(n14235) );
  NAND2_X1 U14506 ( .A1(n15053), .A2(n12315), .ZN(n12113) );
  NAND2_X1 U14507 ( .A1(n14896), .A2(n10744), .ZN(n12112) );
  NAND2_X1 U14508 ( .A1(n12113), .A2(n12112), .ZN(n14234) );
  NAND2_X1 U14509 ( .A1(n14235), .A2(n14234), .ZN(n14233) );
  OAI21_X1 U14510 ( .B1(n12114), .B2(n12125), .A(n14233), .ZN(n14158) );
  NAND2_X1 U14511 ( .A1(n15046), .A2(n12316), .ZN(n12116) );
  NAND2_X1 U14512 ( .A1(n14881), .A2(n12315), .ZN(n12115) );
  NAND2_X1 U14513 ( .A1(n12116), .A2(n12115), .ZN(n12117) );
  XNOR2_X1 U14514 ( .A(n12117), .B(n11538), .ZN(n12123) );
  NOR2_X1 U14515 ( .A1(n14345), .A2(n6416), .ZN(n12118) );
  AOI21_X1 U14516 ( .B1(n15046), .B2(n12315), .A(n12118), .ZN(n12122) );
  XNOR2_X1 U14517 ( .A(n12123), .B(n12122), .ZN(n14159) );
  NOR2_X1 U14518 ( .A1(n14158), .A2(n14159), .ZN(n14157) );
  INV_X1 U14519 ( .A(n12123), .ZN(n12120) );
  INV_X1 U14520 ( .A(n12122), .ZN(n12119) );
  NOR2_X1 U14521 ( .A1(n12120), .A2(n12119), .ZN(n12128) );
  AOI22_X1 U14522 ( .A1(n14844), .A2(n12316), .B1(n12315), .B2(n14486), .ZN(
        n12121) );
  XNOR2_X1 U14523 ( .A(n12121), .B(n12313), .ZN(n12225) );
  AOI22_X1 U14524 ( .A1(n14844), .A2(n12315), .B1(n10744), .B2(n14486), .ZN(
        n12226) );
  NOR3_X1 U14525 ( .A1(n14157), .A2(n12128), .A3(n6604), .ZN(n12130) );
  NOR2_X1 U14526 ( .A1(n12123), .A2(n12122), .ZN(n12127) );
  AOI21_X1 U14527 ( .B1(n14234), .B2(n12126), .A(n12127), .ZN(n12124) );
  NOR3_X1 U14528 ( .A1(n12127), .A2(n12126), .A3(n14234), .ZN(n12129) );
  OAI21_X1 U14529 ( .B1(n12130), .B2(n12240), .A(n14232), .ZN(n12136) );
  INV_X1 U14530 ( .A(n14845), .ZN(n12134) );
  OR2_X1 U14531 ( .A1(n14345), .A2(n14935), .ZN(n12132) );
  NAND2_X1 U14532 ( .A1(n14818), .A2(n14897), .ZN(n12131) );
  AND2_X1 U14533 ( .A1(n12132), .A2(n12131), .ZN(n15037) );
  NAND2_X1 U14534 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14604)
         );
  OAI21_X1 U14535 ( .B1(n14198), .B2(n15037), .A(n14604), .ZN(n12133) );
  AOI21_X1 U14536 ( .B1(n14211), .B2(n12134), .A(n12133), .ZN(n12135) );
  OAI211_X1 U14537 ( .C1(n7717), .C2(n14242), .A(n12136), .B(n12135), .ZN(
        P1_U3228) );
  NAND2_X1 U14538 ( .A1(n12139), .A2(n6489), .ZN(n12141) );
  XNOR2_X1 U14539 ( .A(n12141), .B(n8414), .ZN(n12146) );
  OAI22_X1 U14540 ( .A1(n12511), .A2(n12144), .B1(n12143), .B2(n12142), .ZN(
        n12145) );
  AOI21_X1 U14541 ( .B1(n12146), .B2(n12883), .A(n12145), .ZN(n12155) );
  MUX2_X1 U14542 ( .A(n12155), .B(n12147), .S(n15429), .Z(n12149) );
  OAI211_X1 U14543 ( .C1(n6458), .C2(n13010), .A(n12149), .B(n12148), .ZN(
        P3_U3456) );
  INV_X1 U14544 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12150) );
  MUX2_X1 U14545 ( .A(n12150), .B(n12155), .S(n12896), .Z(n12153) );
  OAI211_X1 U14546 ( .C1(n6458), .C2(n12876), .A(n12153), .B(n12152), .ZN(
        P3_U3204) );
  INV_X1 U14547 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12154) );
  MUX2_X1 U14548 ( .A(n12155), .B(n12154), .S(n15440), .Z(n12157) );
  OAI211_X1 U14549 ( .C1(n6458), .C2(n12941), .A(n12157), .B(n12156), .ZN(
        P3_U3488) );
  OAI222_X1 U14550 ( .A1(n13039), .A2(n12159), .B1(n13036), .B2(n12158), .C1(
        P3_U3151), .C2(n6417), .ZN(P3_U3276) );
  INV_X1 U14551 ( .A(n13367), .ZN(n15103) );
  INV_X1 U14552 ( .A(n12160), .ZN(n15107) );
  OAI222_X1 U14553 ( .A1(n14097), .A2(n12161), .B1(n14092), .B2(n15107), .C1(
        P2_U3088), .C2(n13434), .ZN(P2_U3300) );
  NAND2_X1 U14554 ( .A1(n12163), .A2(n12162), .ZN(n12164) );
  XNOR2_X1 U14555 ( .A(n12387), .B(n12203), .ZN(n12382) );
  XNOR2_X1 U14556 ( .A(n12469), .B(n12203), .ZN(n12380) );
  INV_X1 U14557 ( .A(n12380), .ZN(n12379) );
  AOI22_X1 U14558 ( .A1(n12382), .A2(n12514), .B1(n12379), .B2(n12515), .ZN(
        n12169) );
  AOI21_X1 U14559 ( .B1(n12380), .B2(n12386), .A(n12450), .ZN(n12167) );
  NAND3_X1 U14560 ( .A1(n12380), .A2(n12386), .A3(n12450), .ZN(n12166) );
  OAI21_X1 U14561 ( .B1(n12167), .B2(n12382), .A(n12166), .ZN(n12168) );
  XNOR2_X1 U14562 ( .A(n12868), .B(n10799), .ZN(n12446) );
  NAND2_X1 U14563 ( .A1(n12446), .A2(n12344), .ZN(n12170) );
  INV_X1 U14564 ( .A(n12446), .ZN(n12171) );
  NAND2_X1 U14565 ( .A1(n12171), .A2(n12513), .ZN(n12172) );
  NAND2_X1 U14566 ( .A1(n12173), .A2(n12172), .ZN(n12342) );
  XNOR2_X1 U14567 ( .A(n12942), .B(n12203), .ZN(n12174) );
  XOR2_X1 U14568 ( .A(n12500), .B(n12174), .Z(n12341) );
  INV_X1 U14569 ( .A(n12174), .ZN(n12175) );
  NAND2_X1 U14570 ( .A1(n12175), .A2(n12859), .ZN(n12176) );
  XNOR2_X1 U14571 ( .A(n13006), .B(n12203), .ZN(n12177) );
  NAND2_X1 U14572 ( .A1(n12177), .A2(n12405), .ZN(n12493) );
  INV_X1 U14573 ( .A(n12177), .ZN(n12178) );
  NAND2_X1 U14574 ( .A1(n12178), .A2(n12847), .ZN(n12494) );
  XNOR2_X1 U14575 ( .A(n12935), .B(n10799), .ZN(n12413) );
  XNOR2_X1 U14576 ( .A(n13000), .B(n10799), .ZN(n12410) );
  INV_X1 U14577 ( .A(n12410), .ZN(n12412) );
  AOI22_X1 U14578 ( .A1(n12413), .A2(n12478), .B1(n12417), .B2(n12412), .ZN(
        n12182) );
  AOI21_X1 U14579 ( .B1(n12410), .B2(n12860), .A(n12846), .ZN(n12180) );
  NAND2_X1 U14580 ( .A1(n12846), .A2(n12860), .ZN(n12179) );
  OAI22_X1 U14581 ( .A1(n12180), .A2(n12413), .B1(n12412), .B2(n12179), .ZN(
        n12181) );
  XNOR2_X1 U14582 ( .A(n12993), .B(n12203), .ZN(n12474) );
  XNOR2_X1 U14583 ( .A(n12811), .B(n12203), .ZN(n12183) );
  XOR2_X1 U14584 ( .A(n12825), .B(n12183), .Z(n12361) );
  INV_X1 U14585 ( .A(n12183), .ZN(n12184) );
  NAND2_X1 U14586 ( .A1(n12184), .A2(n12825), .ZN(n12185) );
  XNOR2_X1 U14587 ( .A(n12986), .B(n12203), .ZN(n12186) );
  XNOR2_X1 U14588 ( .A(n12186), .B(n12805), .ZN(n12438) );
  INV_X1 U14589 ( .A(n12186), .ZN(n12187) );
  NAND2_X1 U14590 ( .A1(n12187), .A2(n12805), .ZN(n12188) );
  XNOR2_X1 U14591 ( .A(n12980), .B(n12203), .ZN(n12190) );
  XOR2_X1 U14592 ( .A(n12798), .B(n12190), .Z(n12372) );
  NAND2_X1 U14593 ( .A1(n12190), .A2(n12189), .ZN(n12191) );
  XNOR2_X1 U14594 ( .A(n12974), .B(n10799), .ZN(n12350) );
  XNOR2_X1 U14595 ( .A(n12909), .B(n12203), .ZN(n12427) );
  XNOR2_X1 U14596 ( .A(n12968), .B(n10799), .ZN(n12352) );
  NAND2_X1 U14597 ( .A1(n12352), .A2(n12779), .ZN(n12425) );
  OAI21_X1 U14598 ( .B1(n12427), .B2(n12357), .A(n12425), .ZN(n12194) );
  AOI21_X1 U14599 ( .B1(n12350), .B2(n12788), .A(n12194), .ZN(n12192) );
  INV_X1 U14600 ( .A(n12352), .ZN(n12193) );
  NAND2_X1 U14601 ( .A1(n12193), .A2(n12459), .ZN(n12423) );
  NAND2_X1 U14602 ( .A1(n12423), .A2(n12767), .ZN(n12197) );
  NOR3_X1 U14603 ( .A1(n12352), .A2(n12779), .A3(n12767), .ZN(n12196) );
  NOR3_X1 U14604 ( .A1(n12194), .A2(n12350), .A3(n12788), .ZN(n12195) );
  AOI211_X1 U14605 ( .C1(n12427), .C2(n12197), .A(n12196), .B(n12195), .ZN(
        n12198) );
  NAND2_X1 U14606 ( .A1(n12199), .A2(n12198), .ZN(n12393) );
  XNOR2_X1 U14607 ( .A(n12961), .B(n12203), .ZN(n12200) );
  XOR2_X1 U14608 ( .A(n12432), .B(n12200), .Z(n12394) );
  NAND2_X1 U14609 ( .A1(n12393), .A2(n12394), .ZN(n12202) );
  NAND2_X1 U14610 ( .A1(n12200), .A2(n12432), .ZN(n12201) );
  NAND2_X1 U14611 ( .A1(n12202), .A2(n12201), .ZN(n12483) );
  XNOR2_X1 U14612 ( .A(n12954), .B(n12203), .ZN(n12204) );
  XNOR2_X1 U14613 ( .A(n12204), .B(n12744), .ZN(n12484) );
  NAND2_X1 U14614 ( .A1(n12204), .A2(n12397), .ZN(n12205) );
  XNOR2_X1 U14615 ( .A(n9906), .B(n12203), .ZN(n12206) );
  XOR2_X1 U14616 ( .A(n12489), .B(n12206), .Z(n12336) );
  XOR2_X1 U14617 ( .A(n12207), .B(n12203), .Z(n12208) );
  NAND2_X1 U14618 ( .A1(n12510), .A2(n12497), .ZN(n12210) );
  AOI22_X1 U14619 ( .A1(n12714), .A2(n12502), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12209) );
  OAI211_X1 U14620 ( .C1(n12489), .C2(n12499), .A(n12210), .B(n12209), .ZN(
        n12211) );
  AOI21_X1 U14621 ( .B1(n12715), .B2(n12503), .A(n12211), .ZN(n12212) );
  OAI21_X1 U14622 ( .B1(n12213), .B2(n12506), .A(n12212), .ZN(P3_U3160) );
  INV_X1 U14623 ( .A(n12214), .ZN(n12215) );
  OAI222_X1 U14624 ( .A1(n9915), .A2(P3_U3151), .B1(n13034), .B2(n12216), .C1(
        n13039), .C2(n12215), .ZN(P3_U3271) );
  INV_X1 U14625 ( .A(n14094), .ZN(n12217) );
  OAI222_X1 U14626 ( .A1(n15105), .A2(n12218), .B1(n10976), .B2(n12217), .C1(
        n9784), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND3_X1 U14627 ( .A1(n15446), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n12224) );
  NAND2_X1 U14628 ( .A1(n14087), .A2(n12220), .ZN(n12223) );
  NAND2_X1 U14629 ( .A1(n12221), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n12222) );
  OAI211_X1 U14630 ( .C1(n12219), .C2(n12224), .A(n12223), .B(n12222), .ZN(
        P1_U3324) );
  INV_X1 U14631 ( .A(n12225), .ZN(n12228) );
  INV_X1 U14632 ( .A(n12226), .ZN(n12227) );
  NOR2_X1 U14633 ( .A1(n12228), .A2(n12227), .ZN(n14122) );
  NAND2_X1 U14634 ( .A1(n15034), .A2(n12316), .ZN(n12230) );
  NAND2_X1 U14635 ( .A1(n14818), .A2(n12315), .ZN(n12229) );
  NAND2_X1 U14636 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  XNOR2_X1 U14637 ( .A(n12231), .B(n12313), .ZN(n12241) );
  INV_X1 U14638 ( .A(n12241), .ZN(n12233) );
  OAI22_X1 U14639 ( .A1(n14829), .A2(n6402), .B1(n14131), .B2(n6416), .ZN(
        n12242) );
  INV_X1 U14640 ( .A(n12242), .ZN(n12232) );
  NAND2_X1 U14641 ( .A1(n12233), .A2(n12232), .ZN(n14123) );
  NOR2_X1 U14642 ( .A1(n14827), .A2(n6416), .ZN(n12234) );
  AOI21_X1 U14643 ( .B1(n15028), .B2(n12315), .A(n12234), .ZN(n12246) );
  NAND2_X1 U14644 ( .A1(n15028), .A2(n12316), .ZN(n12236) );
  NAND2_X1 U14645 ( .A1(n14485), .A2(n12315), .ZN(n12235) );
  NAND2_X1 U14646 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  XNOR2_X1 U14647 ( .A(n12237), .B(n12313), .ZN(n12245) );
  XOR2_X1 U14648 ( .A(n12246), .B(n12245), .Z(n14125) );
  INV_X1 U14649 ( .A(n14125), .ZN(n12238) );
  NAND2_X1 U14650 ( .A1(n14123), .A2(n12238), .ZN(n12243) );
  OR2_X1 U14651 ( .A1(n14122), .A2(n12243), .ZN(n12239) );
  XOR2_X1 U14652 ( .A(n12242), .B(n12241), .Z(n14215) );
  INV_X1 U14653 ( .A(n12245), .ZN(n12247) );
  OR2_X1 U14654 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  NAND2_X1 U14655 ( .A1(n14127), .A2(n12248), .ZN(n14177) );
  AND2_X1 U14656 ( .A1(n14816), .A2(n10744), .ZN(n12249) );
  AOI21_X1 U14657 ( .B1(n15022), .B2(n12315), .A(n12249), .ZN(n12252) );
  AOI22_X1 U14658 ( .A1(n15022), .A2(n12316), .B1(n12315), .B2(n14816), .ZN(
        n12250) );
  XNOR2_X1 U14659 ( .A(n12250), .B(n12313), .ZN(n12251) );
  XOR2_X1 U14660 ( .A(n12252), .B(n12251), .Z(n14179) );
  INV_X1 U14661 ( .A(n12251), .ZN(n12254) );
  INV_X1 U14662 ( .A(n12252), .ZN(n12253) );
  NAND2_X1 U14663 ( .A1(n12254), .A2(n12253), .ZN(n12255) );
  OAI22_X1 U14664 ( .A1(n14790), .A2(n12273), .B1(n12257), .B2(n6401), .ZN(
        n12256) );
  XNOR2_X1 U14665 ( .A(n12256), .B(n12313), .ZN(n12258) );
  OAI22_X1 U14666 ( .A1(n14790), .A2(n6401), .B1(n12257), .B2(n6416), .ZN(
        n12259) );
  XNOR2_X1 U14667 ( .A(n12258), .B(n12259), .ZN(n14136) );
  INV_X1 U14668 ( .A(n12258), .ZN(n12261) );
  INV_X1 U14669 ( .A(n12259), .ZN(n12260) );
  OR2_X1 U14670 ( .A1(n9615), .A2(n6402), .ZN(n12263) );
  NAND2_X1 U14671 ( .A1(n14483), .A2(n10744), .ZN(n12262) );
  NAND2_X1 U14672 ( .A1(n12263), .A2(n12262), .ZN(n12266) );
  OAI22_X1 U14673 ( .A1(n9615), .A2(n12273), .B1(n14784), .B2(n6402), .ZN(
        n12264) );
  XNOR2_X1 U14674 ( .A(n12264), .B(n12313), .ZN(n12265) );
  XOR2_X1 U14675 ( .A(n12266), .B(n12265), .Z(n14195) );
  INV_X1 U14676 ( .A(n12265), .ZN(n12268) );
  INV_X1 U14677 ( .A(n12266), .ZN(n12267) );
  NAND2_X1 U14678 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  NAND2_X1 U14679 ( .A1(n14193), .A2(n12269), .ZN(n14117) );
  NAND2_X1 U14680 ( .A1(n15005), .A2(n12316), .ZN(n12271) );
  NAND2_X1 U14681 ( .A1(n14482), .A2(n12315), .ZN(n12270) );
  NAND2_X1 U14682 ( .A1(n12271), .A2(n12270), .ZN(n12272) );
  XNOR2_X1 U14683 ( .A(n12272), .B(n12313), .ZN(n12282) );
  AOI22_X1 U14684 ( .A1(n15005), .A2(n12315), .B1(n10744), .B2(n14482), .ZN(
        n12283) );
  XNOR2_X1 U14685 ( .A(n12282), .B(n12283), .ZN(n14166) );
  OAI22_X1 U14686 ( .A1(n15000), .A2(n12273), .B1(n14387), .B2(n6402), .ZN(
        n12274) );
  XNOR2_X1 U14687 ( .A(n12274), .B(n12313), .ZN(n12277) );
  INV_X1 U14688 ( .A(n12277), .ZN(n12276) );
  OAI22_X1 U14689 ( .A1(n15000), .A2(n6401), .B1(n14387), .B2(n6416), .ZN(
        n12278) );
  INV_X1 U14690 ( .A(n12278), .ZN(n12275) );
  NAND2_X1 U14691 ( .A1(n12276), .A2(n12275), .ZN(n12285) );
  INV_X1 U14692 ( .A(n12285), .ZN(n12279) );
  XOR2_X1 U14693 ( .A(n12278), .B(n12277), .Z(n14170) );
  AND2_X1 U14694 ( .A1(n14166), .A2(n12281), .ZN(n12280) );
  NAND2_X1 U14695 ( .A1(n14117), .A2(n12280), .ZN(n12289) );
  INV_X1 U14696 ( .A(n12281), .ZN(n12287) );
  INV_X1 U14697 ( .A(n12282), .ZN(n12284) );
  NAND2_X1 U14698 ( .A1(n12284), .A2(n12283), .ZN(n14167) );
  AND2_X1 U14699 ( .A1(n14167), .A2(n12285), .ZN(n12286) );
  OAI22_X1 U14700 ( .A1(n14726), .A2(n6401), .B1(n14225), .B2(n6416), .ZN(
        n12294) );
  NAND2_X1 U14701 ( .A1(n14995), .A2(n12316), .ZN(n12291) );
  NAND2_X1 U14702 ( .A1(n14481), .A2(n12315), .ZN(n12290) );
  NAND2_X1 U14703 ( .A1(n12291), .A2(n12290), .ZN(n12292) );
  XNOR2_X1 U14704 ( .A(n12292), .B(n12313), .ZN(n12293) );
  XOR2_X1 U14705 ( .A(n12294), .B(n12293), .Z(n14152) );
  INV_X1 U14706 ( .A(n12293), .ZN(n12296) );
  INV_X1 U14707 ( .A(n12294), .ZN(n12295) );
  NAND2_X1 U14708 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  OAI22_X1 U14709 ( .A1(n14700), .A2(n6402), .B1(n14679), .B2(n6416), .ZN(
        n12303) );
  NAND2_X1 U14710 ( .A1(n14395), .A2(n12316), .ZN(n12300) );
  NAND2_X1 U14711 ( .A1(n14480), .A2(n12315), .ZN(n12299) );
  NAND2_X1 U14712 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  XNOR2_X1 U14713 ( .A(n12301), .B(n12313), .ZN(n12302) );
  XOR2_X1 U14714 ( .A(n12303), .B(n12302), .Z(n14224) );
  INV_X1 U14715 ( .A(n12302), .ZN(n12305) );
  INV_X1 U14716 ( .A(n12303), .ZN(n12304) );
  NAND2_X1 U14717 ( .A1(n14983), .A2(n12316), .ZN(n12307) );
  NAND2_X1 U14718 ( .A1(n14479), .A2(n12315), .ZN(n12306) );
  NAND2_X1 U14719 ( .A1(n12307), .A2(n12306), .ZN(n12308) );
  XNOR2_X1 U14720 ( .A(n12308), .B(n11538), .ZN(n12320) );
  NOR2_X1 U14721 ( .A1(n14226), .A2(n6416), .ZN(n12309) );
  AOI21_X1 U14722 ( .B1(n14983), .B2(n12315), .A(n12309), .ZN(n12319) );
  XNOR2_X1 U14723 ( .A(n12320), .B(n12319), .ZN(n14100) );
  INV_X1 U14724 ( .A(n14100), .ZN(n12310) );
  NAND2_X1 U14725 ( .A1(n14101), .A2(n12310), .ZN(n12334) );
  NAND2_X1 U14726 ( .A1(n14408), .A2(n12315), .ZN(n12312) );
  NAND2_X1 U14727 ( .A1(n14478), .A2(n10744), .ZN(n12311) );
  NAND2_X1 U14728 ( .A1(n12312), .A2(n12311), .ZN(n12314) );
  XNOR2_X1 U14729 ( .A(n12314), .B(n12313), .ZN(n12318) );
  AOI22_X1 U14730 ( .A1(n14408), .A2(n12316), .B1(n12315), .B2(n14478), .ZN(
        n12317) );
  XNOR2_X1 U14731 ( .A(n12318), .B(n12317), .ZN(n12325) );
  NAND2_X1 U14732 ( .A1(n12325), .A2(n14232), .ZN(n12333) );
  AND2_X1 U14733 ( .A1(n12320), .A2(n12319), .ZN(n12326) );
  NOR3_X1 U14734 ( .A1(n12325), .A2(n12326), .A3(n15174), .ZN(n12321) );
  NAND2_X1 U14735 ( .A1(n12334), .A2(n12321), .ZN(n12332) );
  INV_X1 U14736 ( .A(n14420), .ZN(n14477) );
  AOI22_X1 U14737 ( .A1(n14477), .A2(n14218), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12324) );
  NAND2_X1 U14738 ( .A1(n12322), .A2(n14211), .ZN(n12323) );
  OAI211_X1 U14739 ( .C1(n14226), .C2(n14216), .A(n12324), .B(n12323), .ZN(
        n12330) );
  INV_X1 U14740 ( .A(n12325), .ZN(n12328) );
  INV_X1 U14741 ( .A(n12326), .ZN(n12327) );
  NOR3_X1 U14742 ( .A1(n12328), .A2(n15174), .A3(n12327), .ZN(n12329) );
  AOI211_X1 U14743 ( .C1(n14221), .C2(n14408), .A(n12330), .B(n12329), .ZN(
        n12331) );
  OAI211_X1 U14744 ( .C1(n12334), .C2(n12333), .A(n12332), .B(n12331), .ZN(
        P1_U3220) );
  NOR2_X1 U14745 ( .A1(n12511), .A2(n12488), .ZN(n12339) );
  AOI22_X1 U14746 ( .A1(n12726), .A2(n12502), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12337) );
  OAI21_X1 U14747 ( .B1(n12397), .B2(n12499), .A(n12337), .ZN(n12338) );
  AOI211_X1 U14748 ( .C1(n9906), .C2(n12503), .A(n12339), .B(n12338), .ZN(
        n12340) );
  XNOR2_X1 U14749 ( .A(n12342), .B(n12341), .ZN(n12349) );
  NAND2_X1 U14750 ( .A1(n12497), .A2(n12847), .ZN(n12343) );
  NAND2_X1 U14751 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12586)
         );
  OAI211_X1 U14752 ( .C1(n12344), .C2(n12499), .A(n12343), .B(n12586), .ZN(
        n12345) );
  AOI21_X1 U14753 ( .B1(n12346), .B2(n12502), .A(n12345), .ZN(n12348) );
  NAND2_X1 U14754 ( .A1(n12942), .A2(n12503), .ZN(n12347) );
  OAI211_X1 U14755 ( .C1(n12349), .C2(n12506), .A(n12348), .B(n12347), .ZN(
        P3_U3155) );
  NAND2_X1 U14756 ( .A1(n12351), .A2(n7032), .ZN(n12422) );
  NAND2_X1 U14757 ( .A1(n12424), .A2(n12422), .ZN(n12354) );
  XNOR2_X1 U14758 ( .A(n12352), .B(n12779), .ZN(n12353) );
  XNOR2_X1 U14759 ( .A(n12354), .B(n12353), .ZN(n12360) );
  AOI22_X1 U14760 ( .A1(n12788), .A2(n12485), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12356) );
  NAND2_X1 U14761 ( .A1(n12770), .A2(n12502), .ZN(n12355) );
  OAI211_X1 U14762 ( .C1(n12357), .C2(n12488), .A(n12356), .B(n12355), .ZN(
        n12358) );
  AOI21_X1 U14763 ( .B1(n12968), .B2(n12503), .A(n12358), .ZN(n12359) );
  OAI21_X1 U14764 ( .B1(n12360), .B2(n12506), .A(n12359), .ZN(P3_U3156) );
  INV_X1 U14765 ( .A(n12811), .ZN(n12928) );
  AOI21_X1 U14766 ( .B1(n12362), .B2(n12361), .A(n12506), .ZN(n12364) );
  NAND2_X1 U14767 ( .A1(n12364), .A2(n12363), .ZN(n12368) );
  NAND2_X1 U14768 ( .A1(n12805), .A2(n12497), .ZN(n12365) );
  NAND2_X1 U14769 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12695)
         );
  OAI211_X1 U14770 ( .C1(n12473), .C2(n12499), .A(n12365), .B(n12695), .ZN(
        n12366) );
  AOI21_X1 U14771 ( .B1(n12807), .B2(n12502), .A(n12366), .ZN(n12367) );
  OAI211_X1 U14772 ( .C1(n12451), .C2(n12928), .A(n12368), .B(n12367), .ZN(
        P3_U3159) );
  INV_X1 U14773 ( .A(n12369), .ZN(n12370) );
  AOI21_X1 U14774 ( .B1(n12372), .B2(n12371), .A(n12370), .ZN(n12378) );
  AOI22_X1 U14775 ( .A1(n12805), .A2(n12485), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12374) );
  NAND2_X1 U14776 ( .A1(n12791), .A2(n12502), .ZN(n12373) );
  OAI211_X1 U14777 ( .C1(n12375), .C2(n12488), .A(n12374), .B(n12373), .ZN(
        n12376) );
  AOI21_X1 U14778 ( .B1(n12980), .B2(n12503), .A(n12376), .ZN(n12377) );
  OAI21_X1 U14779 ( .B1(n12378), .B2(n12506), .A(n12377), .ZN(P3_U3163) );
  XNOR2_X1 U14780 ( .A(n12381), .B(n12379), .ZN(n12463) );
  AOI22_X1 U14781 ( .A1(n12463), .A2(n12386), .B1(n12381), .B2(n12380), .ZN(
        n12384) );
  XNOR2_X1 U14782 ( .A(n12382), .B(n12450), .ZN(n12383) );
  XNOR2_X1 U14783 ( .A(n12384), .B(n12383), .ZN(n12392) );
  NAND2_X1 U14784 ( .A1(n12497), .A2(n12513), .ZN(n12385) );
  NAND2_X1 U14785 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12533)
         );
  OAI211_X1 U14786 ( .C1(n12386), .C2(n12499), .A(n12385), .B(n12533), .ZN(
        n12389) );
  NOR2_X1 U14787 ( .A1(n12387), .A2(n12451), .ZN(n12388) );
  AOI211_X1 U14788 ( .C1(n12390), .C2(n12502), .A(n12389), .B(n12388), .ZN(
        n12391) );
  OAI21_X1 U14789 ( .B1(n12392), .B2(n12506), .A(n12391), .ZN(P3_U3164) );
  XOR2_X1 U14790 ( .A(n12394), .B(n12393), .Z(n12400) );
  AOI22_X1 U14791 ( .A1(n12767), .A2(n12485), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12396) );
  NAND2_X1 U14792 ( .A1(n12748), .A2(n12502), .ZN(n12395) );
  OAI211_X1 U14793 ( .C1(n12397), .C2(n12488), .A(n12396), .B(n12395), .ZN(
        n12398) );
  AOI21_X1 U14794 ( .B1(n12961), .B2(n12503), .A(n12398), .ZN(n12399) );
  OAI21_X1 U14795 ( .B1(n12400), .B2(n12506), .A(n12399), .ZN(P3_U3165) );
  XNOR2_X1 U14796 ( .A(n12410), .B(n12417), .ZN(n12403) );
  XNOR2_X1 U14797 ( .A(n12402), .B(n12403), .ZN(n12409) );
  NAND2_X1 U14798 ( .A1(n12497), .A2(n12846), .ZN(n12404) );
  NAND2_X1 U14799 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12635)
         );
  OAI211_X1 U14800 ( .C1(n12405), .C2(n12499), .A(n12404), .B(n12635), .ZN(
        n12406) );
  AOI21_X1 U14801 ( .B1(n12850), .B2(n12502), .A(n12406), .ZN(n12408) );
  NAND2_X1 U14802 ( .A1(n13000), .A2(n12503), .ZN(n12407) );
  OAI211_X1 U14803 ( .C1(n12409), .C2(n12506), .A(n12408), .B(n12407), .ZN(
        P3_U3166) );
  OAI21_X1 U14804 ( .B1(n12402), .B2(n12410), .A(n12860), .ZN(n12411) );
  OAI21_X1 U14805 ( .B1(n7028), .B2(n12412), .A(n12411), .ZN(n12415) );
  XNOR2_X1 U14806 ( .A(n12413), .B(n12846), .ZN(n12414) );
  XNOR2_X1 U14807 ( .A(n12415), .B(n12414), .ZN(n12421) );
  NAND2_X1 U14808 ( .A1(n12832), .A2(n12497), .ZN(n12416) );
  NAND2_X1 U14809 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12654)
         );
  OAI211_X1 U14810 ( .C1(n12417), .C2(n12499), .A(n12416), .B(n12654), .ZN(
        n12419) );
  NOR2_X1 U14811 ( .A1(n12935), .A2(n12451), .ZN(n12418) );
  AOI211_X1 U14812 ( .C1(n12836), .C2(n12502), .A(n12419), .B(n12418), .ZN(
        n12420) );
  OAI21_X1 U14813 ( .B1(n12421), .B2(n12506), .A(n12420), .ZN(P3_U3168) );
  NAND3_X1 U14814 ( .A1(n12424), .A2(n12423), .A3(n12422), .ZN(n12426) );
  NAND2_X1 U14815 ( .A1(n12426), .A2(n12425), .ZN(n12429) );
  XNOR2_X1 U14816 ( .A(n12427), .B(n12767), .ZN(n12428) );
  XNOR2_X1 U14817 ( .A(n12429), .B(n12428), .ZN(n12435) );
  AOI22_X1 U14818 ( .A1(n12779), .A2(n12485), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12431) );
  NAND2_X1 U14819 ( .A1(n12758), .A2(n12502), .ZN(n12430) );
  OAI211_X1 U14820 ( .C1(n12432), .C2(n12488), .A(n12431), .B(n12430), .ZN(
        n12433) );
  AOI21_X1 U14821 ( .B1(n12909), .B2(n12503), .A(n12433), .ZN(n12434) );
  OAI21_X1 U14822 ( .B1(n12435), .B2(n12506), .A(n12434), .ZN(P3_U3169) );
  INV_X1 U14823 ( .A(n12986), .ZN(n12445) );
  OAI211_X1 U14824 ( .C1(n12439), .C2(n12438), .A(n12437), .B(n12436), .ZN(
        n12444) );
  AOI22_X1 U14825 ( .A1(n12798), .A2(n12497), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12440) );
  OAI21_X1 U14826 ( .B1(n12441), .B2(n12499), .A(n12440), .ZN(n12442) );
  AOI21_X1 U14827 ( .B1(n12801), .B2(n12502), .A(n12442), .ZN(n12443) );
  OAI211_X1 U14828 ( .C1(n12445), .C2(n12451), .A(n12444), .B(n12443), .ZN(
        P3_U3173) );
  XNOR2_X1 U14829 ( .A(n12446), .B(n12513), .ZN(n12447) );
  XNOR2_X1 U14830 ( .A(n12448), .B(n12447), .ZN(n12455) );
  NAND2_X1 U14831 ( .A1(n12497), .A2(n12859), .ZN(n12449) );
  NAND2_X1 U14832 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12551)
         );
  OAI211_X1 U14833 ( .C1(n12450), .C2(n12499), .A(n12449), .B(n12551), .ZN(
        n12453) );
  NOR2_X1 U14834 ( .A1(n12868), .A2(n12451), .ZN(n12452) );
  AOI211_X1 U14835 ( .C1(n12872), .C2(n12502), .A(n12453), .B(n12452), .ZN(
        n12454) );
  OAI21_X1 U14836 ( .B1(n12455), .B2(n12506), .A(n12454), .ZN(P3_U3174) );
  XNOR2_X1 U14837 ( .A(n12456), .B(n12788), .ZN(n12462) );
  AOI22_X1 U14838 ( .A1(n12798), .A2(n12485), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12458) );
  NAND2_X1 U14839 ( .A1(n12782), .A2(n12502), .ZN(n12457) );
  OAI211_X1 U14840 ( .C1(n12459), .C2(n12488), .A(n12458), .B(n12457), .ZN(
        n12460) );
  AOI21_X1 U14841 ( .B1(n12974), .B2(n12503), .A(n12460), .ZN(n12461) );
  OAI21_X1 U14842 ( .B1(n12462), .B2(n12506), .A(n12461), .ZN(P3_U3175) );
  XNOR2_X1 U14843 ( .A(n12463), .B(n12515), .ZN(n12472) );
  NAND2_X1 U14844 ( .A1(n12497), .A2(n12514), .ZN(n12465) );
  OAI211_X1 U14845 ( .C1(n12466), .C2(n12499), .A(n12465), .B(n12464), .ZN(
        n12467) );
  AOI21_X1 U14846 ( .B1(n12468), .B2(n12502), .A(n12467), .ZN(n12471) );
  NAND2_X1 U14847 ( .A1(n12469), .A2(n12503), .ZN(n12470) );
  OAI211_X1 U14848 ( .C1(n12472), .C2(n12506), .A(n12471), .B(n12470), .ZN(
        P3_U3176) );
  XNOR2_X1 U14849 ( .A(n12474), .B(n12473), .ZN(n12475) );
  XNOR2_X1 U14850 ( .A(n12476), .B(n12475), .ZN(n12482) );
  NAND2_X1 U14851 ( .A1(n12825), .A2(n12497), .ZN(n12477) );
  NAND2_X1 U14852 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12680)
         );
  OAI211_X1 U14853 ( .C1(n12478), .C2(n12499), .A(n12477), .B(n12680), .ZN(
        n12479) );
  AOI21_X1 U14854 ( .B1(n12828), .B2(n12502), .A(n12479), .ZN(n12481) );
  NAND2_X1 U14855 ( .A1(n12993), .A2(n12503), .ZN(n12480) );
  OAI211_X1 U14856 ( .C1(n12482), .C2(n12506), .A(n12481), .B(n12480), .ZN(
        P3_U3178) );
  XOR2_X1 U14857 ( .A(n12484), .B(n12483), .Z(n12492) );
  AOI22_X1 U14858 ( .A1(n12752), .A2(n12485), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12487) );
  NAND2_X1 U14859 ( .A1(n12737), .A2(n12502), .ZN(n12486) );
  OAI211_X1 U14860 ( .C1(n12489), .C2(n12488), .A(n12487), .B(n12486), .ZN(
        n12490) );
  AOI21_X1 U14861 ( .B1(n12954), .B2(n12503), .A(n12490), .ZN(n12491) );
  OAI21_X1 U14862 ( .B1(n12492), .B2(n12506), .A(n12491), .ZN(P3_U3180) );
  NAND2_X1 U14863 ( .A1(n12494), .A2(n12493), .ZN(n12496) );
  XOR2_X1 U14864 ( .A(n12496), .B(n12495), .Z(n12507) );
  NAND2_X1 U14865 ( .A1(n12497), .A2(n12860), .ZN(n12498) );
  NAND2_X1 U14866 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12617)
         );
  OAI211_X1 U14867 ( .C1(n12500), .C2(n12499), .A(n12498), .B(n12617), .ZN(
        n12501) );
  AOI21_X1 U14868 ( .B1(n12854), .B2(n12502), .A(n12501), .ZN(n12505) );
  NAND2_X1 U14869 ( .A1(n13006), .A2(n12503), .ZN(n12504) );
  OAI211_X1 U14870 ( .C1(n12507), .C2(n12506), .A(n12505), .B(n12504), .ZN(
        P3_U3181) );
  MUX2_X1 U14871 ( .A(n12508), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12512), .Z(
        P3_U3522) );
  MUX2_X1 U14872 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12509), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14873 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12510), .S(P3_U3897), .Z(
        P3_U3520) );
  INV_X1 U14874 ( .A(n12511), .ZN(n12720) );
  MUX2_X1 U14875 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12720), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14876 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12735), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14877 ( .A(n12744), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12512), .Z(
        P3_U3517) );
  MUX2_X1 U14878 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12752), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14879 ( .A(n12767), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12512), .Z(
        P3_U3515) );
  MUX2_X1 U14880 ( .A(n12779), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12512), .Z(
        P3_U3514) );
  MUX2_X1 U14881 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12788), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14882 ( .A(n12798), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12512), .Z(
        P3_U3512) );
  MUX2_X1 U14883 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12805), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14884 ( .A(n12825), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12512), .Z(
        P3_U3510) );
  MUX2_X1 U14885 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12832), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14886 ( .A(n12846), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12512), .Z(
        P3_U3508) );
  MUX2_X1 U14887 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12860), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14888 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12847), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14889 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12859), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12513), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14891 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12514), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12515), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14893 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12516), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12517), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14895 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12518), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12519), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12520), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12521), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12878), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14900 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12522), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n7223), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12523), .S(P3_U3897), .Z(
        P3_U3491) );
  XNOR2_X1 U14903 ( .A(n12560), .B(n15452), .ZN(n12561) );
  NAND2_X1 U14904 ( .A1(n12524), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U14905 ( .A1(n12525), .A2(n12529), .ZN(n12526) );
  XOR2_X1 U14906 ( .A(n12561), .B(n12562), .Z(n12544) );
  NOR2_X1 U14907 ( .A1(n12529), .A2(n12528), .ZN(n12531) );
  MUX2_X1 U14908 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13031), .Z(n12552) );
  XNOR2_X1 U14909 ( .A(n12552), .B(n12560), .ZN(n12530) );
  NOR2_X1 U14910 ( .A1(n12555), .A2(n12705), .ZN(n12541) );
  OAI21_X1 U14911 ( .B1(n12532), .B2(n12531), .A(n12530), .ZN(n12540) );
  INV_X1 U14912 ( .A(n12533), .ZN(n12534) );
  AOI21_X1 U14913 ( .B1(n15391), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12534), 
        .ZN(n12535) );
  OAI21_X1 U14914 ( .B1(n12697), .B2(n12560), .A(n12535), .ZN(n12539) );
  XNOR2_X1 U14915 ( .A(n12560), .B(n12546), .ZN(n12536) );
  OR3_X1 U14916 ( .A1(n6450), .A2(n7405), .A3(n12536), .ZN(n12537) );
  AOI21_X1 U14917 ( .B1(n12545), .B2(n12537), .A(n12663), .ZN(n12538) );
  AOI211_X1 U14918 ( .C1(n12541), .C2(n12540), .A(n12539), .B(n12538), .ZN(
        n12542) );
  OAI21_X1 U14919 ( .B1(n12544), .B2(n12543), .A(n12542), .ZN(P3_U3194) );
  INV_X1 U14920 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12550) );
  INV_X1 U14921 ( .A(n12560), .ZN(n12547) );
  OAI21_X1 U14922 ( .B1(n12547), .B2(n12546), .A(n12545), .ZN(n12548) );
  NAND2_X1 U14923 ( .A1(n12548), .A2(n12573), .ZN(n12595) );
  OAI21_X1 U14924 ( .B1(n12548), .B2(n12573), .A(n12595), .ZN(n12549) );
  AOI21_X1 U14925 ( .B1(n12550), .B2(n12549), .A(n12593), .ZN(n12566) );
  INV_X1 U14926 ( .A(n12573), .ZN(n12567) );
  OAI21_X1 U14927 ( .B1(n12655), .B2(n15113), .A(n12551), .ZN(n12559) );
  AND2_X1 U14928 ( .A1(n12552), .A2(n12560), .ZN(n12554) );
  MUX2_X1 U14929 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13031), .Z(n12574) );
  XNOR2_X1 U14930 ( .A(n12574), .B(n12573), .ZN(n12553) );
  INV_X1 U14931 ( .A(n12582), .ZN(n12557) );
  OAI21_X1 U14932 ( .B1(n12555), .B2(n12554), .A(n12553), .ZN(n12556) );
  AOI21_X1 U14933 ( .B1(n12557), .B2(n12556), .A(n12705), .ZN(n12558) );
  AOI211_X1 U14934 ( .C1(n12661), .C2(n12567), .A(n12559), .B(n12558), .ZN(
        n12565) );
  XOR2_X1 U14935 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12569), .Z(n12563) );
  NAND2_X1 U14936 ( .A1(n12563), .A2(n12707), .ZN(n12564) );
  OAI211_X1 U14937 ( .C1(n12566), .C2(n12663), .A(n12565), .B(n12564), .ZN(
        P3_U3195) );
  INV_X1 U14938 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U14939 ( .A1(n12590), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12614) );
  INV_X1 U14940 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U14941 ( .A1(n12576), .A2(n12570), .ZN(n12571) );
  AND2_X1 U14942 ( .A1(n12614), .A2(n12571), .ZN(n12578) );
  OAI21_X1 U14943 ( .B1(n12572), .B2(n12578), .A(n12613), .ZN(n12600) );
  NOR2_X1 U14944 ( .A1(n12574), .A2(n12573), .ZN(n12581) );
  NAND2_X1 U14945 ( .A1(n12590), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U14946 ( .A1(n12576), .A2(n12575), .ZN(n12577) );
  AND2_X1 U14947 ( .A1(n12608), .A2(n12577), .ZN(n12591) );
  INV_X1 U14948 ( .A(n12591), .ZN(n12594) );
  INV_X1 U14949 ( .A(n12578), .ZN(n12579) );
  MUX2_X1 U14950 ( .A(n12594), .B(n12579), .S(n13031), .Z(n12580) );
  INV_X1 U14951 ( .A(n12605), .ZN(n12585) );
  OAI21_X1 U14952 ( .B1(n12582), .B2(n12581), .A(n12580), .ZN(n12583) );
  NAND3_X1 U14953 ( .A1(n12585), .A2(n12584), .A3(n12583), .ZN(n12589) );
  INV_X1 U14954 ( .A(n12586), .ZN(n12587) );
  AOI21_X1 U14955 ( .B1(n15391), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12587), 
        .ZN(n12588) );
  OAI211_X1 U14956 ( .C1(n12697), .C2(n12590), .A(n12589), .B(n12588), .ZN(
        n12599) );
  INV_X1 U14957 ( .A(n12595), .ZN(n12592) );
  INV_X1 U14958 ( .A(n12593), .ZN(n12596) );
  NAND3_X1 U14959 ( .A1(n12596), .A2(n12595), .A3(n12594), .ZN(n12597) );
  AOI21_X1 U14960 ( .B1(n12609), .B2(n12597), .A(n12663), .ZN(n12598) );
  AOI211_X1 U14961 ( .C1(n12707), .C2(n12600), .A(n12599), .B(n12598), .ZN(
        n12601) );
  INV_X1 U14962 ( .A(n12601), .ZN(P3_U3196) );
  INV_X1 U14963 ( .A(n12608), .ZN(n12603) );
  INV_X1 U14964 ( .A(n12614), .ZN(n12602) );
  MUX2_X1 U14965 ( .A(n12603), .B(n12602), .S(n13031), .Z(n12604) );
  MUX2_X1 U14966 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13031), .Z(n12606) );
  AOI21_X1 U14967 ( .B1(n12607), .B2(n12606), .A(n12629), .ZN(n12622) );
  OAI21_X1 U14968 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n12611), .A(n12640), 
        .ZN(n12612) );
  NAND2_X1 U14969 ( .A1(n12612), .A2(n12688), .ZN(n12621) );
  INV_X1 U14970 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15130) );
  OAI21_X1 U14971 ( .B1(n12615), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12625), 
        .ZN(n12616) );
  NAND2_X1 U14972 ( .A1(n12707), .A2(n12616), .ZN(n12618) );
  OAI211_X1 U14973 ( .C1(n12655), .C2(n15130), .A(n12618), .B(n12617), .ZN(
        n12619) );
  AOI21_X1 U14974 ( .B1(n12630), .B2(n12661), .A(n12619), .ZN(n12620) );
  OAI211_X1 U14975 ( .C1(n12622), .C2(n12705), .A(n12621), .B(n12620), .ZN(
        P3_U3197) );
  NAND2_X1 U14976 ( .A1(n12624), .A2(n12623), .ZN(n12626) );
  XNOR2_X1 U14977 ( .A(n12653), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U14978 ( .B1(n12628), .B2(n12627), .A(n12652), .ZN(n12644) );
  INV_X1 U14979 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12849) );
  INV_X1 U14980 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n15575) );
  MUX2_X1 U14981 ( .A(n12849), .B(n15575), .S(n13031), .Z(n12632) );
  NOR2_X1 U14982 ( .A1(n12653), .A2(n12632), .ZN(n12657) );
  NAND2_X1 U14983 ( .A1(n12653), .A2(n12632), .ZN(n12656) );
  INV_X1 U14984 ( .A(n12656), .ZN(n12633) );
  NOR2_X1 U14985 ( .A1(n12657), .A2(n12633), .ZN(n12634) );
  XNOR2_X1 U14986 ( .A(n6564), .B(n12634), .ZN(n12638) );
  INV_X1 U14987 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U14988 ( .B1(n12655), .B2(n15147), .A(n12635), .ZN(n12636) );
  AOI21_X1 U14989 ( .B1(n12653), .B2(n12661), .A(n12636), .ZN(n12637) );
  OAI21_X1 U14990 ( .B1(n12638), .B2(n12705), .A(n12637), .ZN(n12643) );
  NAND3_X1 U14991 ( .A1(n12640), .A2(n6635), .A3(n12639), .ZN(n12641) );
  AOI21_X1 U14992 ( .B1(n12648), .B2(n12641), .A(n12663), .ZN(n12642) );
  AOI211_X1 U14993 ( .C1(n12707), .C2(n12644), .A(n12643), .B(n12642), .ZN(
        n12645) );
  INV_X1 U14994 ( .A(n12645), .ZN(P3_U3198) );
  INV_X1 U14995 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U14996 ( .A1(n12646), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U14997 ( .A1(n12648), .A2(n12647), .ZN(n12649) );
  AOI21_X1 U14998 ( .B1(n12651), .B2(n12650), .A(n6460), .ZN(n12664) );
  INV_X1 U14999 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15497) );
  MUX2_X1 U15000 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13031), .Z(n12667) );
  XNOR2_X1 U15001 ( .A(n12666), .B(n12667), .ZN(n12659) );
  NOR2_X1 U15002 ( .A1(n12658), .A2(n12659), .ZN(n12665) );
  AOI211_X1 U15003 ( .C1(n12659), .C2(n12658), .A(n12705), .B(n12665), .ZN(
        n12660) );
  OAI21_X1 U15004 ( .B1(n12664), .B2(n12663), .A(n12662), .ZN(P3_U3199) );
  MUX2_X1 U15005 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13031), .Z(n12669) );
  AOI21_X1 U15006 ( .B1(n12667), .B2(n12666), .A(n12665), .ZN(n12703) );
  AOI21_X1 U15007 ( .B1(n12669), .B2(n12668), .A(n12701), .ZN(n12685) );
  INV_X1 U15008 ( .A(n12672), .ZN(n12671) );
  NAND2_X1 U15009 ( .A1(n12690), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12686) );
  INV_X1 U15010 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U15011 ( .A1(n12702), .A2(n12827), .ZN(n12670) );
  AND2_X1 U15012 ( .A1(n12686), .A2(n12670), .ZN(n12673) );
  NOR3_X1 U15013 ( .A1(n6460), .A2(n12671), .A3(n12673), .ZN(n12676) );
  INV_X1 U15014 ( .A(n12674), .ZN(n12675) );
  OAI21_X1 U15015 ( .B1(n12676), .B2(n12675), .A(n12688), .ZN(n12684) );
  INV_X1 U15016 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12677) );
  XNOR2_X1 U15017 ( .A(n12702), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12691) );
  XNOR2_X1 U15018 ( .A(n12692), .B(n12691), .ZN(n12682) );
  NAND2_X1 U15019 ( .A1(n15391), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12679) );
  OAI211_X1 U15020 ( .C1(n12697), .C2(n12690), .A(n12680), .B(n12679), .ZN(
        n12681) );
  AOI21_X1 U15021 ( .B1(n12707), .B2(n12682), .A(n12681), .ZN(n12683) );
  OAI211_X1 U15022 ( .C1(n12685), .C2(n12705), .A(n12684), .B(n12683), .ZN(
        P3_U3200) );
  NAND2_X1 U15023 ( .A1(n12674), .A2(n12686), .ZN(n12687) );
  XNOR2_X1 U15024 ( .A(n6417), .B(n12809), .ZN(n12698) );
  XNOR2_X1 U15025 ( .A(n12687), .B(n12698), .ZN(n12689) );
  NAND2_X1 U15026 ( .A1(n12689), .A2(n12688), .ZN(n12709) );
  AOI22_X1 U15027 ( .A1(n12692), .A2(n12691), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12690), .ZN(n12693) );
  XNOR2_X1 U15028 ( .A(n6417), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12699) );
  NAND2_X1 U15029 ( .A1(n15391), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12694) );
  OAI211_X1 U15030 ( .C1(n12697), .C2(n6417), .A(n12695), .B(n12694), .ZN(
        n12706) );
  INV_X1 U15031 ( .A(n12698), .ZN(n12700) );
  MUX2_X1 U15032 ( .A(n12700), .B(n12699), .S(n13031), .Z(n12704) );
  NAND2_X1 U15033 ( .A1(n12709), .A2(n12708), .ZN(P3_U3201) );
  NAND2_X1 U15034 ( .A1(n12863), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12710) );
  OAI211_X1 U15035 ( .C1(n12950), .C2(n12867), .A(n12711), .B(n12710), .ZN(
        P3_U3202) );
  MUX2_X1 U15036 ( .A(P3_REG2_REG_28__SCAN_IN), .B(n12712), .S(n12896), .Z(
        n12713) );
  INV_X1 U15037 ( .A(n12713), .ZN(n12717) );
  AOI22_X1 U15038 ( .A1(n12715), .A2(n12855), .B1(n12873), .B2(n12714), .ZN(
        n12716) );
  OAI211_X1 U15039 ( .C1(n12718), .C2(n12876), .A(n12717), .B(n12716), .ZN(
        P3_U3205) );
  NAND2_X1 U15040 ( .A1(n12720), .A2(n12879), .ZN(n12722) );
  INV_X1 U15041 ( .A(n9906), .ZN(n12728) );
  AOI22_X1 U15042 ( .A1(n12726), .A2(n12873), .B1(n12863), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12727) );
  OAI21_X1 U15043 ( .B1(n12728), .B2(n12867), .A(n12727), .ZN(n12729) );
  AOI21_X1 U15044 ( .B1(n12900), .B2(n12839), .A(n12729), .ZN(n12730) );
  OAI21_X1 U15045 ( .B1(n12901), .B2(n12863), .A(n12730), .ZN(P3_U3206) );
  INV_X1 U15046 ( .A(n12731), .ZN(n12732) );
  INV_X1 U15047 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12736) );
  MUX2_X1 U15048 ( .A(n12736), .B(n12952), .S(n12896), .Z(n12739) );
  AOI22_X1 U15049 ( .A1(n12954), .A2(n12855), .B1(n12873), .B2(n12737), .ZN(
        n12738) );
  OAI211_X1 U15050 ( .C1(n12957), .C2(n12876), .A(n12739), .B(n12738), .ZN(
        P3_U3207) );
  XNOR2_X1 U15051 ( .A(n12740), .B(n12742), .ZN(n12964) );
  OAI211_X1 U15052 ( .C1(n12743), .C2(n12742), .A(n12741), .B(n12883), .ZN(
        n12746) );
  AOI22_X1 U15053 ( .A1(n12744), .A2(n12879), .B1(n12767), .B2(n12880), .ZN(
        n12745) );
  NAND2_X1 U15054 ( .A1(n12746), .A2(n12745), .ZN(n12958) );
  MUX2_X1 U15055 ( .A(n12958), .B(P3_REG2_REG_25__SCAN_IN), .S(n12863), .Z(
        n12747) );
  INV_X1 U15056 ( .A(n12747), .ZN(n12750) );
  AOI22_X1 U15057 ( .A1(n12961), .A2(n12855), .B1(n12873), .B2(n12748), .ZN(
        n12749) );
  OAI211_X1 U15058 ( .C1(n12964), .C2(n12876), .A(n12750), .B(n12749), .ZN(
        P3_U3208) );
  XOR2_X1 U15059 ( .A(n12757), .B(n12751), .Z(n12753) );
  AOI222_X1 U15060 ( .A1(n12883), .A2(n12753), .B1(n12779), .B2(n12880), .C1(
        n12752), .C2(n12879), .ZN(n12911) );
  INV_X1 U15061 ( .A(n12754), .ZN(n12755) );
  AOI21_X1 U15062 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(n12912) );
  INV_X1 U15063 ( .A(n12912), .ZN(n12762) );
  INV_X1 U15064 ( .A(n12909), .ZN(n12760) );
  AOI22_X1 U15065 ( .A1(n12758), .A2(n12873), .B1(n12863), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12759) );
  OAI21_X1 U15066 ( .B1(n12760), .B2(n12867), .A(n12759), .ZN(n12761) );
  AOI21_X1 U15067 ( .B1(n12762), .B2(n12839), .A(n12761), .ZN(n12763) );
  OAI21_X1 U15068 ( .B1(n12911), .B2(n12863), .A(n12763), .ZN(P3_U3209) );
  XNOR2_X1 U15069 ( .A(n12764), .B(n12765), .ZN(n12971) );
  INV_X1 U15070 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12769) );
  XNOR2_X1 U15071 ( .A(n12766), .B(n12765), .ZN(n12768) );
  AOI222_X1 U15072 ( .A1(n12883), .A2(n12768), .B1(n12767), .B2(n12879), .C1(
        n12788), .C2(n12880), .ZN(n12966) );
  MUX2_X1 U15073 ( .A(n12769), .B(n12966), .S(n12896), .Z(n12772) );
  AOI22_X1 U15074 ( .A1(n12968), .A2(n12855), .B1(n12873), .B2(n12770), .ZN(
        n12771) );
  OAI211_X1 U15075 ( .C1(n12971), .C2(n12876), .A(n12772), .B(n12771), .ZN(
        P3_U3210) );
  NAND2_X1 U15076 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  XOR2_X1 U15077 ( .A(n12777), .B(n12775), .Z(n12977) );
  INV_X1 U15078 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12781) );
  XNOR2_X1 U15079 ( .A(n12778), .B(n12777), .ZN(n12780) );
  AOI222_X1 U15080 ( .A1(n12883), .A2(n12780), .B1(n12779), .B2(n12879), .C1(
        n12798), .C2(n12880), .ZN(n12972) );
  MUX2_X1 U15081 ( .A(n12781), .B(n12972), .S(n12896), .Z(n12784) );
  AOI22_X1 U15082 ( .A1(n12974), .A2(n12855), .B1(n12873), .B2(n12782), .ZN(
        n12783) );
  OAI211_X1 U15083 ( .C1(n12977), .C2(n12876), .A(n12784), .B(n12783), .ZN(
        P3_U3211) );
  XNOR2_X1 U15084 ( .A(n12785), .B(n12787), .ZN(n12983) );
  INV_X1 U15085 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12790) );
  XNOR2_X1 U15086 ( .A(n12786), .B(n12787), .ZN(n12789) );
  AOI222_X1 U15087 ( .A1(n12883), .A2(n12789), .B1(n12788), .B2(n12879), .C1(
        n12805), .C2(n12880), .ZN(n12978) );
  MUX2_X1 U15088 ( .A(n12790), .B(n12978), .S(n12896), .Z(n12793) );
  AOI22_X1 U15089 ( .A1(n12980), .A2(n12855), .B1(n12873), .B2(n12791), .ZN(
        n12792) );
  OAI211_X1 U15090 ( .C1(n12983), .C2(n12876), .A(n12793), .B(n12792), .ZN(
        P3_U3212) );
  OAI21_X1 U15091 ( .B1(n12795), .B2(n12797), .A(n12794), .ZN(n12989) );
  INV_X1 U15092 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12800) );
  XNOR2_X1 U15093 ( .A(n12796), .B(n12797), .ZN(n12799) );
  AOI222_X1 U15094 ( .A1(n12883), .A2(n12799), .B1(n12798), .B2(n12879), .C1(
        n12825), .C2(n12880), .ZN(n12984) );
  MUX2_X1 U15095 ( .A(n12800), .B(n12984), .S(n12896), .Z(n12803) );
  AOI22_X1 U15096 ( .A1(n12986), .A2(n12855), .B1(n12873), .B2(n12801), .ZN(
        n12802) );
  OAI211_X1 U15097 ( .C1(n12989), .C2(n12876), .A(n12803), .B(n12802), .ZN(
        P3_U3213) );
  XNOR2_X1 U15098 ( .A(n12804), .B(n12814), .ZN(n12806) );
  AOI222_X1 U15099 ( .A1(n12883), .A2(n12806), .B1(n12805), .B2(n12879), .C1(
        n12832), .C2(n12880), .ZN(n12927) );
  INV_X1 U15100 ( .A(n12807), .ZN(n12808) );
  OAI22_X1 U15101 ( .A1(n12896), .A2(n12809), .B1(n12808), .B2(n12891), .ZN(
        n12810) );
  AOI21_X1 U15102 ( .B1(n12811), .B2(n12855), .A(n12810), .ZN(n12817) );
  NAND2_X1 U15103 ( .A1(n12835), .A2(n7149), .ZN(n12834) );
  NAND3_X1 U15104 ( .A1(n12834), .A2(n12822), .A3(n12812), .ZN(n12820) );
  NAND2_X1 U15105 ( .A1(n12820), .A2(n12813), .ZN(n12815) );
  XNOR2_X1 U15106 ( .A(n12815), .B(n12814), .ZN(n12925) );
  NAND2_X1 U15107 ( .A1(n12925), .A2(n12839), .ZN(n12816) );
  OAI211_X1 U15108 ( .C1(n12927), .C2(n12863), .A(n12817), .B(n12816), .ZN(
        P3_U3214) );
  INV_X1 U15109 ( .A(n12834), .ZN(n12819) );
  NOR2_X1 U15110 ( .A1(n12819), .A2(n12818), .ZN(n12821) );
  OAI21_X1 U15111 ( .B1(n12821), .B2(n12822), .A(n12820), .ZN(n12996) );
  OAI21_X1 U15112 ( .B1(n12824), .B2(n9891), .A(n12823), .ZN(n12826) );
  AOI222_X1 U15113 ( .A1(n12883), .A2(n12826), .B1(n12846), .B2(n12880), .C1(
        n12825), .C2(n12879), .ZN(n12991) );
  MUX2_X1 U15114 ( .A(n12827), .B(n12991), .S(n12896), .Z(n12830) );
  AOI22_X1 U15115 ( .A1(n12993), .A2(n12855), .B1(n12873), .B2(n12828), .ZN(
        n12829) );
  OAI211_X1 U15116 ( .C1(n12996), .C2(n12876), .A(n12830), .B(n12829), .ZN(
        P3_U3215) );
  XNOR2_X1 U15117 ( .A(n12831), .B(n7149), .ZN(n12833) );
  AOI222_X1 U15118 ( .A1(n12883), .A2(n12833), .B1(n12860), .B2(n12880), .C1(
        n12832), .C2(n12879), .ZN(n12934) );
  OAI21_X1 U15119 ( .B1(n12835), .B2(n7149), .A(n12834), .ZN(n12932) );
  AOI22_X1 U15120 ( .A1(n12863), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n12873), 
        .B2(n12836), .ZN(n12837) );
  OAI21_X1 U15121 ( .B1(n12935), .B2(n12867), .A(n12837), .ZN(n12838) );
  AOI21_X1 U15122 ( .B1(n12932), .B2(n12839), .A(n12838), .ZN(n12840) );
  OAI21_X1 U15123 ( .B1(n12934), .B2(n12863), .A(n12840), .ZN(P3_U3216) );
  OAI21_X1 U15124 ( .B1(n12842), .B2(n12845), .A(n12841), .ZN(n12843) );
  INV_X1 U15125 ( .A(n12843), .ZN(n13003) );
  XNOR2_X1 U15126 ( .A(n12844), .B(n12845), .ZN(n12848) );
  AOI222_X1 U15127 ( .A1(n12883), .A2(n12848), .B1(n12847), .B2(n12880), .C1(
        n12846), .C2(n12879), .ZN(n12998) );
  MUX2_X1 U15128 ( .A(n12849), .B(n12998), .S(n12896), .Z(n12852) );
  AOI22_X1 U15129 ( .A1(n13000), .A2(n12855), .B1(n12873), .B2(n12850), .ZN(
        n12851) );
  OAI211_X1 U15130 ( .C1(n13003), .C2(n12876), .A(n12852), .B(n12851), .ZN(
        P3_U3217) );
  XNOR2_X1 U15131 ( .A(n12853), .B(n12857), .ZN(n13009) );
  AOI22_X1 U15132 ( .A1(n13006), .A2(n12855), .B1(n12873), .B2(n12854), .ZN(
        n12866) );
  OAI211_X1 U15133 ( .C1(n12858), .C2(n12857), .A(n12856), .B(n12883), .ZN(
        n12862) );
  AOI22_X1 U15134 ( .A1(n12860), .A2(n12879), .B1(n12859), .B2(n12880), .ZN(
        n12861) );
  NAND2_X1 U15135 ( .A1(n12862), .A2(n12861), .ZN(n13004) );
  INV_X1 U15136 ( .A(n13004), .ZN(n12864) );
  MUX2_X1 U15137 ( .A(n12864), .B(n7404), .S(n12863), .Z(n12865) );
  OAI211_X1 U15138 ( .C1(n13009), .C2(n12876), .A(n12866), .B(n12865), .ZN(
        P3_U3218) );
  NOR2_X1 U15139 ( .A1(n12868), .A2(n12867), .ZN(n12871) );
  MUX2_X1 U15140 ( .A(P3_REG2_REG_13__SCAN_IN), .B(n12869), .S(n12896), .Z(
        n12870) );
  AOI211_X1 U15141 ( .C1(n12873), .C2(n12872), .A(n12871), .B(n12870), .ZN(
        n12874) );
  OAI21_X1 U15142 ( .B1(n12876), .B2(n12875), .A(n12874), .ZN(P3_U3220) );
  XNOR2_X1 U15143 ( .A(n12877), .B(n12882), .ZN(n15399) );
  AOI22_X1 U15144 ( .A1(n7223), .A2(n12880), .B1(n12879), .B2(n12878), .ZN(
        n12886) );
  OAI21_X1 U15145 ( .B1(n10932), .B2(n12882), .A(n12881), .ZN(n12884) );
  NAND2_X1 U15146 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  OAI211_X1 U15147 ( .C1(n15399), .C2(n12887), .A(n12886), .B(n12885), .ZN(
        n15401) );
  OR2_X1 U15148 ( .A1(n12888), .A2(n15418), .ZN(n15397) );
  OAI22_X1 U15149 ( .A1(n12891), .A2(n12890), .B1(n12889), .B2(n15397), .ZN(
        n12892) );
  INV_X1 U15150 ( .A(n12892), .ZN(n12893) );
  OAI21_X1 U15151 ( .B1(n15399), .B2(n12894), .A(n12893), .ZN(n12895) );
  OR2_X1 U15152 ( .A1(n15401), .A2(n12895), .ZN(n12897) );
  MUX2_X1 U15153 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n12897), .S(n12896), .Z(
        P3_U3231) );
  NAND2_X1 U15154 ( .A1(n15440), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12898) );
  OAI211_X1 U15155 ( .C1(n12950), .C2(n12905), .A(n12899), .B(n12898), .ZN(
        P3_U3490) );
  MUX2_X1 U15156 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12951), .S(n15589), .Z(
        P3_U3486) );
  INV_X1 U15157 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12902) );
  MUX2_X1 U15158 ( .A(n12902), .B(n12952), .S(n15589), .Z(n12904) );
  NAND2_X1 U15159 ( .A1(n12954), .A2(n12939), .ZN(n12903) );
  OAI211_X1 U15160 ( .C1(n12941), .C2(n12957), .A(n12904), .B(n12903), .ZN(
        P3_U3485) );
  MUX2_X1 U15161 ( .A(n12958), .B(P3_REG1_REG_25__SCAN_IN), .S(n15440), .Z(
        n12908) );
  INV_X1 U15162 ( .A(n12961), .ZN(n12906) );
  OAI22_X1 U15163 ( .A1(n12964), .A2(n12941), .B1(n12906), .B2(n12905), .ZN(
        n12907) );
  OR2_X1 U15164 ( .A1(n12908), .A2(n12907), .ZN(P3_U3484) );
  NAND2_X1 U15165 ( .A1(n12909), .A2(n15423), .ZN(n12910) );
  MUX2_X1 U15166 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12965), .S(n15589), .Z(
        P3_U3483) );
  INV_X1 U15167 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12913) );
  MUX2_X1 U15168 ( .A(n12913), .B(n12966), .S(n15589), .Z(n12915) );
  NAND2_X1 U15169 ( .A1(n12968), .A2(n12939), .ZN(n12914) );
  OAI211_X1 U15170 ( .C1(n12971), .C2(n12941), .A(n12915), .B(n12914), .ZN(
        P3_U3482) );
  INV_X1 U15171 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12916) );
  MUX2_X1 U15172 ( .A(n12916), .B(n12972), .S(n15589), .Z(n12918) );
  NAND2_X1 U15173 ( .A1(n12974), .A2(n12939), .ZN(n12917) );
  OAI211_X1 U15174 ( .C1(n12977), .C2(n12941), .A(n12918), .B(n12917), .ZN(
        P3_U3481) );
  INV_X1 U15175 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12919) );
  MUX2_X1 U15176 ( .A(n12919), .B(n12978), .S(n15589), .Z(n12921) );
  NAND2_X1 U15177 ( .A1(n12980), .A2(n12939), .ZN(n12920) );
  OAI211_X1 U15178 ( .C1(n12941), .C2(n12983), .A(n12921), .B(n12920), .ZN(
        P3_U3480) );
  INV_X1 U15179 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12922) );
  MUX2_X1 U15180 ( .A(n12922), .B(n12984), .S(n15589), .Z(n12924) );
  NAND2_X1 U15181 ( .A1(n12986), .A2(n12939), .ZN(n12923) );
  OAI211_X1 U15182 ( .C1(n12941), .C2(n12989), .A(n12924), .B(n12923), .ZN(
        P3_U3479) );
  NAND2_X1 U15183 ( .A1(n12925), .A2(n15395), .ZN(n12926) );
  OAI211_X1 U15184 ( .C1(n15418), .C2(n12928), .A(n12927), .B(n12926), .ZN(
        n12990) );
  MUX2_X1 U15185 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12990), .S(n15589), .Z(
        P3_U3478) );
  INV_X1 U15186 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12929) );
  MUX2_X1 U15187 ( .A(n12929), .B(n12991), .S(n15589), .Z(n12931) );
  NAND2_X1 U15188 ( .A1(n12993), .A2(n12939), .ZN(n12930) );
  OAI211_X1 U15189 ( .C1(n12941), .C2(n12996), .A(n12931), .B(n12930), .ZN(
        P3_U3477) );
  NAND2_X1 U15190 ( .A1(n12932), .A2(n15395), .ZN(n12933) );
  OAI211_X1 U15191 ( .C1(n15418), .C2(n12935), .A(n12934), .B(n12933), .ZN(
        n12997) );
  MUX2_X1 U15192 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12997), .S(n15589), .Z(
        P3_U3476) );
  MUX2_X1 U15193 ( .A(n15575), .B(n12998), .S(n15589), .Z(n12937) );
  NAND2_X1 U15194 ( .A1(n13000), .A2(n12939), .ZN(n12936) );
  OAI211_X1 U15195 ( .C1(n13003), .C2(n12941), .A(n12937), .B(n12936), .ZN(
        P3_U3475) );
  MUX2_X1 U15196 ( .A(n13004), .B(P3_REG1_REG_15__SCAN_IN), .S(n15440), .Z(
        n12938) );
  AOI21_X1 U15197 ( .B1(n12939), .B2(n13006), .A(n12938), .ZN(n12940) );
  OAI21_X1 U15198 ( .B1(n12941), .B2(n13009), .A(n12940), .ZN(P3_U3474) );
  NAND2_X1 U15199 ( .A1(n12942), .A2(n15423), .ZN(n12943) );
  OAI211_X1 U15200 ( .C1(n12946), .C2(n12945), .A(n12944), .B(n12943), .ZN(
        n13011) );
  MUX2_X1 U15201 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13011), .S(n15589), .Z(
        P3_U3473) );
  NAND2_X1 U15202 ( .A1(n15429), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12947) );
  OAI211_X1 U15203 ( .C1(n12950), .C2(n12949), .A(n12948), .B(n12947), .ZN(
        P3_U3458) );
  MUX2_X1 U15204 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12951), .S(n15431), .Z(
        P3_U3454) );
  MUX2_X1 U15205 ( .A(n12953), .B(n12952), .S(n15431), .Z(n12956) );
  NAND2_X1 U15206 ( .A1(n12954), .A2(n13007), .ZN(n12955) );
  OAI211_X1 U15207 ( .C1(n12957), .C2(n13010), .A(n12956), .B(n12955), .ZN(
        P3_U3453) );
  INV_X1 U15208 ( .A(n12958), .ZN(n12960) );
  MUX2_X1 U15209 ( .A(n12960), .B(n12959), .S(n15429), .Z(n12963) );
  NAND2_X1 U15210 ( .A1(n12961), .A2(n13007), .ZN(n12962) );
  OAI211_X1 U15211 ( .C1(n12964), .C2(n13010), .A(n12963), .B(n12962), .ZN(
        P3_U3452) );
  MUX2_X1 U15212 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12965), .S(n15431), .Z(
        P3_U3451) );
  MUX2_X1 U15213 ( .A(n12967), .B(n12966), .S(n15431), .Z(n12970) );
  NAND2_X1 U15214 ( .A1(n12968), .A2(n13007), .ZN(n12969) );
  OAI211_X1 U15215 ( .C1(n12971), .C2(n13010), .A(n12970), .B(n12969), .ZN(
        P3_U3450) );
  MUX2_X1 U15216 ( .A(n12973), .B(n12972), .S(n15431), .Z(n12976) );
  NAND2_X1 U15217 ( .A1(n12974), .A2(n13007), .ZN(n12975) );
  OAI211_X1 U15218 ( .C1(n12977), .C2(n13010), .A(n12976), .B(n12975), .ZN(
        P3_U3449) );
  MUX2_X1 U15219 ( .A(n12979), .B(n12978), .S(n15431), .Z(n12982) );
  NAND2_X1 U15220 ( .A1(n12980), .A2(n13007), .ZN(n12981) );
  OAI211_X1 U15221 ( .C1(n12983), .C2(n13010), .A(n12982), .B(n12981), .ZN(
        P3_U3448) );
  MUX2_X1 U15222 ( .A(n12985), .B(n12984), .S(n15431), .Z(n12988) );
  NAND2_X1 U15223 ( .A1(n12986), .A2(n13007), .ZN(n12987) );
  OAI211_X1 U15224 ( .C1(n12989), .C2(n13010), .A(n12988), .B(n12987), .ZN(
        P3_U3447) );
  MUX2_X1 U15225 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12990), .S(n15431), .Z(
        P3_U3446) );
  MUX2_X1 U15226 ( .A(n12992), .B(n12991), .S(n15431), .Z(n12995) );
  NAND2_X1 U15227 ( .A1(n12993), .A2(n13007), .ZN(n12994) );
  OAI211_X1 U15228 ( .C1(n12996), .C2(n13010), .A(n12995), .B(n12994), .ZN(
        P3_U3444) );
  MUX2_X1 U15229 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12997), .S(n15431), .Z(
        P3_U3441) );
  MUX2_X1 U15230 ( .A(n12999), .B(n12998), .S(n15431), .Z(n13002) );
  NAND2_X1 U15231 ( .A1(n13000), .A2(n13007), .ZN(n13001) );
  OAI211_X1 U15232 ( .C1(n13003), .C2(n13010), .A(n13002), .B(n13001), .ZN(
        P3_U3438) );
  MUX2_X1 U15233 ( .A(n13004), .B(P3_REG0_REG_15__SCAN_IN), .S(n15429), .Z(
        n13005) );
  AOI21_X1 U15234 ( .B1(n13007), .B2(n13006), .A(n13005), .ZN(n13008) );
  OAI21_X1 U15235 ( .B1(n13010), .B2(n13009), .A(n13008), .ZN(P3_U3435) );
  MUX2_X1 U15236 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13011), .S(n15431), .Z(
        P3_U3432) );
  MUX2_X1 U15237 ( .A(P3_D_REG_1__SCAN_IN), .B(n13012), .S(n13013), .Z(
        P3_U3377) );
  MUX2_X1 U15238 ( .A(P3_D_REG_0__SCAN_IN), .B(n13014), .S(n13013), .Z(
        P3_U3376) );
  NAND2_X1 U15239 ( .A1(n13015), .A2(n13016), .ZN(n13020) );
  OR4_X1 U15240 ( .A1(n13018), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13017), .A4(
        P3_U3151), .ZN(n13019) );
  OAI211_X1 U15241 ( .C1(n13021), .C2(n13036), .A(n13020), .B(n13019), .ZN(
        P3_U3264) );
  INV_X1 U15242 ( .A(n13022), .ZN(n13023) );
  OAI222_X1 U15243 ( .A1(n13034), .A2(n13025), .B1(P3_U3151), .B2(n13024), 
        .C1(n13039), .C2(n13023), .ZN(P3_U3266) );
  OAI222_X1 U15244 ( .A1(n13034), .A2(n13028), .B1(P3_U3151), .B2(n13027), 
        .C1(n13039), .C2(n13026), .ZN(P3_U3267) );
  INV_X1 U15245 ( .A(n13029), .ZN(n13032) );
  OAI222_X1 U15246 ( .A1(n13034), .A2(n13033), .B1(n13039), .B2(n13032), .C1(
        n13031), .C2(P3_U3151), .ZN(P3_U3268) );
  INV_X1 U15247 ( .A(n13035), .ZN(n13038) );
  OAI222_X1 U15248 ( .A1(P3_U3151), .A2(n13040), .B1(n13039), .B2(n13038), 
        .C1(n13037), .C2(n13036), .ZN(P3_U3269) );
  NAND2_X1 U15249 ( .A1(n13042), .A2(n13041), .ZN(n13043) );
  NAND3_X1 U15250 ( .A1(n6461), .A2(n13182), .A3(n13043), .ZN(n13048) );
  INV_X1 U15251 ( .A(n13044), .ZN(n13670) );
  AOI22_X1 U15252 ( .A1(n13670), .A2(n13170), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13045) );
  OAI21_X1 U15253 ( .B1(n13667), .B2(n13143), .A(n13045), .ZN(n13046) );
  AOI21_X1 U15254 ( .B1(n13594), .B2(n13053), .A(n13046), .ZN(n13047) );
  OAI211_X1 U15255 ( .C1(n13960), .C2(n13194), .A(n13048), .B(n13047), .ZN(
        P2_U3186) );
  INV_X1 U15256 ( .A(n13049), .ZN(n13050) );
  AOI21_X1 U15257 ( .B1(n13052), .B2(n13051), .A(n13050), .ZN(n13057) );
  INV_X1 U15258 ( .A(n13053), .ZN(n13188) );
  AOI22_X1 U15259 ( .A1(n13191), .A2(n13884), .B1(n13891), .B2(n13170), .ZN(
        n13054) );
  NAND2_X1 U15260 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15311)
         );
  OAI211_X1 U15261 ( .C1(n13620), .C2(n13188), .A(n13054), .B(n15311), .ZN(
        n13055) );
  AOI21_X1 U15262 ( .B1(n13569), .B2(n13173), .A(n13055), .ZN(n13056) );
  OAI21_X1 U15263 ( .B1(n13057), .B2(n13165), .A(n13056), .ZN(P2_U3187) );
  OR2_X1 U15264 ( .A1(n13149), .A2(n13058), .ZN(n13150) );
  NAND2_X1 U15265 ( .A1(n13150), .A2(n13059), .ZN(n13061) );
  XNOR2_X1 U15266 ( .A(n13061), .B(n13060), .ZN(n13063) );
  NAND3_X1 U15267 ( .A1(n13063), .A2(n13182), .A3(n13062), .ZN(n13071) );
  INV_X1 U15268 ( .A(n13063), .ZN(n13064) );
  NAND3_X1 U15269 ( .A1(n13064), .A2(n13183), .A3(n13584), .ZN(n13070) );
  OAI22_X1 U15270 ( .A1(n13740), .A2(n13143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13065), .ZN(n13068) );
  INV_X1 U15271 ( .A(n13742), .ZN(n13066) );
  OAI22_X1 U15272 ( .A1(n13741), .A2(n13188), .B1(n13187), .B2(n13066), .ZN(
        n13067) );
  AOI211_X1 U15273 ( .C1(n13978), .C2(n13173), .A(n13068), .B(n13067), .ZN(
        n13069) );
  NAND3_X1 U15274 ( .A1(n13071), .A2(n13070), .A3(n13069), .ZN(P2_U3188) );
  INV_X1 U15275 ( .A(n13072), .ZN(n13080) );
  NOR2_X1 U15276 ( .A1(n13080), .A2(n13073), .ZN(n13074) );
  XNOR2_X1 U15277 ( .A(n13135), .B(n13074), .ZN(n13079) );
  NOR2_X1 U15278 ( .A1(n13075), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13542) );
  OAI22_X1 U15279 ( .A1(n13188), .A2(n13629), .B1(n13187), .B2(n13806), .ZN(
        n13076) );
  AOI211_X1 U15280 ( .C1(n13191), .C2(n13797), .A(n13542), .B(n13076), .ZN(
        n13078) );
  NAND2_X1 U15281 ( .A1(n13997), .A2(n13173), .ZN(n13077) );
  OAI211_X1 U15282 ( .C1(n13079), .C2(n13165), .A(n13078), .B(n13077), .ZN(
        P2_U3191) );
  AOI21_X1 U15283 ( .B1(n13135), .B2(n13081), .A(n13080), .ZN(n13137) );
  XNOR2_X1 U15284 ( .A(n13083), .B(n13082), .ZN(n13138) );
  OAI211_X1 U15285 ( .C1(n9102), .C2(n13084), .A(n13137), .B(n13138), .ZN(
        n13148) );
  AOI21_X1 U15286 ( .B1(n13148), .B2(n13086), .A(n13085), .ZN(n13092) );
  NAND2_X1 U15287 ( .A1(n13087), .A2(n13182), .ZN(n13091) );
  AOI22_X1 U15288 ( .A1(n13631), .A2(n13885), .B1(n13883), .B2(n13798), .ZN(
        n13766) );
  AOI22_X1 U15289 ( .A1(n13170), .A2(n13769), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13088) );
  OAI21_X1 U15290 ( .B1(n13766), .B2(n13120), .A(n13088), .ZN(n13089) );
  AOI21_X1 U15291 ( .B1(n13988), .B2(n13173), .A(n13089), .ZN(n13090) );
  OAI21_X1 U15292 ( .B1(n13092), .B2(n13091), .A(n13090), .ZN(P2_U3195) );
  OAI21_X1 U15293 ( .B1(n13125), .B2(n13093), .A(n13182), .ZN(n13096) );
  NAND3_X1 U15294 ( .A1(n13094), .A2(n13183), .A3(n13701), .ZN(n13095) );
  NAND2_X1 U15295 ( .A1(n13096), .A2(n13095), .ZN(n13097) );
  NAND2_X1 U15296 ( .A1(n13168), .A2(n13097), .ZN(n13102) );
  OAI22_X1 U15297 ( .A1(n13741), .A2(n13143), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13098), .ZN(n13100) );
  NOR2_X1 U15298 ( .A1(n13667), .A2(n13188), .ZN(n13099) );
  AOI211_X1 U15299 ( .C1(n13170), .C2(n13706), .A(n13100), .B(n13099), .ZN(
        n13101) );
  OAI211_X1 U15300 ( .C1(n13708), .C2(n13194), .A(n13102), .B(n13101), .ZN(
        P2_U3197) );
  NAND2_X1 U15301 ( .A1(n13104), .A2(n13103), .ZN(n13108) );
  XNOR2_X1 U15302 ( .A(n13105), .B(n13106), .ZN(n13184) );
  OAI22_X1 U15303 ( .A1(n13184), .A2(n13181), .B1(n13106), .B2(n13105), .ZN(
        n13107) );
  XOR2_X1 U15304 ( .A(n13108), .B(n13107), .Z(n13113) );
  INV_X1 U15305 ( .A(n13848), .ZN(n13573) );
  AOI22_X1 U15306 ( .A1(n13191), .A2(n13886), .B1(n13854), .B2(n13170), .ZN(
        n13110) );
  OAI211_X1 U15307 ( .C1(n13573), .C2(n13188), .A(n13110), .B(n13109), .ZN(
        n13111) );
  AOI21_X1 U15308 ( .B1(n14013), .B2(n13173), .A(n13111), .ZN(n13112) );
  OAI21_X1 U15309 ( .B1(n13113), .B2(n13165), .A(n13112), .ZN(P2_U3198) );
  OAI21_X1 U15310 ( .B1(n13116), .B2(n13115), .A(n13114), .ZN(n13117) );
  NAND2_X1 U15311 ( .A1(n13117), .A2(n13182), .ZN(n13124) );
  INV_X1 U15312 ( .A(n13838), .ZN(n13122) );
  AND2_X1 U15313 ( .A1(n13623), .A2(n13883), .ZN(n13118) );
  AOI21_X1 U15314 ( .B1(n13797), .B2(n13885), .A(n13118), .ZN(n13831) );
  OAI21_X1 U15315 ( .B1(n13120), .B2(n13831), .A(n13119), .ZN(n13121) );
  AOI21_X1 U15316 ( .B1(n13122), .B2(n13170), .A(n13121), .ZN(n13123) );
  OAI211_X1 U15317 ( .C1(n7552), .C2(n13194), .A(n13124), .B(n13123), .ZN(
        P2_U3200) );
  AOI211_X1 U15318 ( .C1(n13127), .C2(n13126), .A(n13165), .B(n13125), .ZN(
        n13128) );
  INV_X1 U15319 ( .A(n13128), .ZN(n13134) );
  OR2_X1 U15320 ( .A1(n13637), .A2(n13871), .ZN(n13130) );
  NAND2_X1 U15321 ( .A1(n13584), .A2(n13883), .ZN(n13129) );
  NAND2_X1 U15322 ( .A1(n13130), .A2(n13129), .ZN(n13716) );
  OAI22_X1 U15323 ( .A1(n13722), .A2(n13187), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13131), .ZN(n13132) );
  AOI21_X1 U15324 ( .B1(n13716), .B2(n13161), .A(n13132), .ZN(n13133) );
  OAI211_X1 U15325 ( .C1(n7554), .C2(n13194), .A(n13134), .B(n13133), .ZN(
        P2_U3201) );
  NAND3_X1 U15326 ( .A1(n13135), .A2(n13183), .A3(n13628), .ZN(n13136) );
  OAI21_X1 U15327 ( .B1(n13137), .B2(n13165), .A(n13136), .ZN(n13140) );
  INV_X1 U15328 ( .A(n13138), .ZN(n13139) );
  NAND2_X1 U15329 ( .A1(n13140), .A2(n13139), .ZN(n13147) );
  INV_X1 U15330 ( .A(n13630), .ZN(n13782) );
  OAI22_X1 U15331 ( .A1(n13188), .A2(n13782), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13141), .ZN(n13145) );
  INV_X1 U15332 ( .A(n13628), .ZN(n13781) );
  INV_X1 U15333 ( .A(n13786), .ZN(n13142) );
  OAI22_X1 U15334 ( .A1(n13143), .A2(n13781), .B1(n13142), .B2(n13187), .ZN(
        n13144) );
  AOI211_X1 U15335 ( .C1(n13993), .C2(n13173), .A(n13145), .B(n13144), .ZN(
        n13146) );
  OAI211_X1 U15336 ( .C1(n13148), .C2(n13165), .A(n13147), .B(n13146), .ZN(
        P2_U3205) );
  OAI22_X1 U15337 ( .A1(n13149), .A2(n13165), .B1(n13740), .B2(n13174), .ZN(
        n13151) );
  NAND2_X1 U15338 ( .A1(n13151), .A2(n13150), .ZN(n13157) );
  NAND2_X1 U15339 ( .A1(n13584), .A2(n13885), .ZN(n13153) );
  NAND2_X1 U15340 ( .A1(n13630), .A2(n13883), .ZN(n13152) );
  NAND2_X1 U15341 ( .A1(n13153), .A2(n13152), .ZN(n13757) );
  OAI22_X1 U15342 ( .A1(n13751), .A2(n13187), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13154), .ZN(n13155) );
  AOI21_X1 U15343 ( .B1(n13757), .B2(n13161), .A(n13155), .ZN(n13156) );
  OAI211_X1 U15344 ( .C1(n13754), .C2(n13194), .A(n13157), .B(n13156), .ZN(
        P2_U3207) );
  XNOR2_X1 U15345 ( .A(n13159), .B(n13158), .ZN(n13166) );
  OAI22_X1 U15346 ( .A1(n13781), .A2(n13871), .B1(n13573), .B2(n13869), .ZN(
        n13816) );
  NOR2_X1 U15347 ( .A1(n13160), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13526) );
  AOI21_X1 U15348 ( .B1(n13816), .B2(n13161), .A(n13526), .ZN(n13162) );
  OAI21_X1 U15349 ( .B1(n13822), .B2(n13187), .A(n13162), .ZN(n13163) );
  AOI21_X1 U15350 ( .B1(n14004), .B2(n13173), .A(n13163), .ZN(n13164) );
  OAI21_X1 U15351 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(P2_U3210) );
  OAI21_X1 U15352 ( .B1(n13176), .B2(n13168), .A(n13167), .ZN(n13169) );
  NAND2_X1 U15353 ( .A1(n13169), .A2(n13182), .ZN(n13180) );
  AOI22_X1 U15354 ( .A1(n13690), .A2(n13170), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13171) );
  OAI21_X1 U15355 ( .B1(n13640), .B2(n13188), .A(n13171), .ZN(n13172) );
  AOI21_X1 U15356 ( .B1(n13962), .B2(n13173), .A(n13172), .ZN(n13179) );
  NOR3_X1 U15357 ( .A1(n13176), .A2(n13175), .A3(n13174), .ZN(n13177) );
  OAI21_X1 U15358 ( .B1(n13177), .B2(n13191), .A(n13682), .ZN(n13178) );
  NAND3_X1 U15359 ( .A1(n13180), .A2(n13179), .A3(n13178), .ZN(P2_U3212) );
  NAND2_X1 U15360 ( .A1(n13182), .A2(n13181), .ZN(n13186) );
  NAND2_X1 U15361 ( .A1(n13183), .A2(n13886), .ZN(n13185) );
  MUX2_X1 U15362 ( .A(n13186), .B(n13185), .S(n13184), .Z(n13193) );
  OAI22_X1 U15363 ( .A1(n13188), .A2(n13870), .B1(n13187), .B2(n13874), .ZN(
        n13189) );
  AOI211_X1 U15364 ( .C1(n13191), .C2(n13568), .A(n13190), .B(n13189), .ZN(
        n13192) );
  OAI211_X1 U15365 ( .C1(n13878), .C2(n13194), .A(n13193), .B(n13192), .ZN(
        P2_U3213) );
  AND3_X1 U15366 ( .A1(n13373), .A2(n13421), .A3(n13195), .ZN(n13196) );
  NAND2_X1 U15367 ( .A1(n13215), .A2(n13198), .ZN(n13199) );
  NAND2_X1 U15368 ( .A1(n13199), .A2(n13200), .ZN(n13202) );
  AOI21_X1 U15369 ( .B1(n13377), .B2(n13452), .A(n13200), .ZN(n13206) );
  INV_X1 U15370 ( .A(n13206), .ZN(n13201) );
  NAND2_X1 U15371 ( .A1(n13202), .A2(n13201), .ZN(n13205) );
  OAI21_X1 U15372 ( .B1(n13428), .B2(n6414), .A(n13203), .ZN(n13204) );
  NAND2_X1 U15373 ( .A1(n13205), .A2(n13204), .ZN(n13208) );
  NAND2_X1 U15374 ( .A1(n13206), .A2(n13452), .ZN(n13207) );
  NAND2_X1 U15375 ( .A1(n13208), .A2(n13207), .ZN(n13212) );
  MUX2_X1 U15376 ( .A(n10017), .B(n13450), .S(n13215), .Z(n13211) );
  NAND2_X1 U15377 ( .A1(n13212), .A2(n13211), .ZN(n13210) );
  MUX2_X1 U15378 ( .A(n13450), .B(n10017), .S(n13372), .Z(n13209) );
  NAND2_X1 U15379 ( .A1(n13210), .A2(n13209), .ZN(n13214) );
  MUX2_X1 U15380 ( .A(n13449), .B(n15361), .S(n13372), .Z(n13217) );
  MUX2_X1 U15381 ( .A(n15361), .B(n13449), .S(n6407), .Z(n13216) );
  MUX2_X1 U15382 ( .A(n13218), .B(n13448), .S(n13372), .Z(n13222) );
  MUX2_X1 U15383 ( .A(n13448), .B(n13218), .S(n13372), .Z(n13219) );
  NAND2_X1 U15384 ( .A1(n13220), .A2(n13219), .ZN(n13226) );
  INV_X1 U15385 ( .A(n13221), .ZN(n13224) );
  INV_X1 U15386 ( .A(n13222), .ZN(n13223) );
  NAND2_X1 U15387 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  NAND2_X1 U15388 ( .A1(n13226), .A2(n13225), .ZN(n13228) );
  MUX2_X1 U15389 ( .A(n13447), .B(n15368), .S(n13372), .Z(n13229) );
  MUX2_X1 U15390 ( .A(n15368), .B(n13447), .S(n13372), .Z(n13227) );
  INV_X1 U15391 ( .A(n13229), .ZN(n13230) );
  MUX2_X1 U15392 ( .A(n6418), .B(n13446), .S(n13372), .Z(n13233) );
  MUX2_X1 U15393 ( .A(n13446), .B(n6418), .S(n13372), .Z(n13231) );
  INV_X1 U15394 ( .A(n13233), .ZN(n13234) );
  MUX2_X1 U15395 ( .A(n13445), .B(n13235), .S(n6407), .Z(n13238) );
  MUX2_X1 U15396 ( .A(n13235), .B(n13445), .S(n13372), .Z(n13236) );
  INV_X1 U15397 ( .A(n13238), .ZN(n13239) );
  MUX2_X1 U15398 ( .A(n13444), .B(n15376), .S(n6404), .Z(n13243) );
  MUX2_X1 U15399 ( .A(n13444), .B(n15376), .S(n13372), .Z(n13240) );
  NAND2_X1 U15400 ( .A1(n13241), .A2(n13240), .ZN(n13245) );
  NAND2_X1 U15401 ( .A1(n13245), .A2(n13244), .ZN(n13249) );
  MUX2_X1 U15402 ( .A(n13443), .B(n13246), .S(n13372), .Z(n13250) );
  NAND2_X1 U15403 ( .A1(n13249), .A2(n13250), .ZN(n13248) );
  MUX2_X1 U15404 ( .A(n13443), .B(n13246), .S(n6404), .Z(n13247) );
  INV_X1 U15405 ( .A(n13249), .ZN(n13252) );
  INV_X1 U15406 ( .A(n13250), .ZN(n13251) );
  MUX2_X1 U15407 ( .A(n13442), .B(n14051), .S(n6404), .Z(n13255) );
  MUX2_X1 U15408 ( .A(n13556), .B(n13253), .S(n13372), .Z(n13254) );
  MUX2_X1 U15409 ( .A(n13256), .B(n11577), .S(n6404), .Z(n13258) );
  MUX2_X1 U15410 ( .A(n13441), .B(n14046), .S(n13372), .Z(n13257) );
  MUX2_X1 U15411 ( .A(n13611), .B(n13932), .S(n6407), .Z(n13264) );
  MUX2_X1 U15412 ( .A(n13440), .B(n14036), .S(n6404), .Z(n13263) );
  MUX2_X1 U15413 ( .A(n13868), .B(n14025), .S(n6404), .Z(n13270) );
  MUX2_X1 U15414 ( .A(n13568), .B(n13569), .S(n13372), .Z(n13269) );
  NAND2_X1 U15415 ( .A1(n13270), .A2(n13269), .ZN(n13273) );
  MUX2_X1 U15416 ( .A(n13614), .B(n13912), .S(n6404), .Z(n13268) );
  MUX2_X1 U15417 ( .A(n13884), .B(n14031), .S(n13372), .Z(n13267) );
  NAND2_X1 U15418 ( .A1(n13268), .A2(n13267), .ZN(n13265) );
  OAI211_X1 U15419 ( .C1(n13264), .C2(n13263), .A(n13273), .B(n13265), .ZN(
        n13278) );
  MUX2_X1 U15420 ( .A(n13608), .B(n13609), .S(n6407), .Z(n13276) );
  MUX2_X1 U15421 ( .A(n13566), .B(n14041), .S(n6404), .Z(n13275) );
  OAI22_X1 U15422 ( .A1(n13276), .A2(n13275), .B1(n7632), .B2(n7631), .ZN(
        n13259) );
  NOR2_X1 U15423 ( .A1(n13278), .A2(n13259), .ZN(n13283) );
  MUX2_X1 U15424 ( .A(n13848), .B(n14008), .S(n6404), .Z(n13290) );
  NAND2_X1 U15425 ( .A1(n14008), .A2(n13848), .ZN(n13625) );
  AND2_X1 U15426 ( .A1(n13623), .A2(n13372), .ZN(n13261) );
  NOR2_X1 U15427 ( .A1(n13623), .A2(n6407), .ZN(n13260) );
  MUX2_X1 U15428 ( .A(n13261), .B(n13260), .S(n14013), .Z(n13262) );
  AOI21_X1 U15429 ( .B1(n13290), .B2(n13625), .A(n13262), .ZN(n13285) );
  NAND3_X1 U15430 ( .A1(n13265), .A2(n13264), .A3(n13263), .ZN(n13266) );
  OAI21_X1 U15431 ( .B1(n13268), .B2(n13267), .A(n13266), .ZN(n13274) );
  INV_X1 U15432 ( .A(n13269), .ZN(n13272) );
  INV_X1 U15433 ( .A(n13270), .ZN(n13271) );
  AOI22_X1 U15434 ( .A1(n13274), .A2(n13273), .B1(n13272), .B2(n13271), .ZN(
        n13281) );
  NAND2_X1 U15435 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  OR2_X1 U15436 ( .A1(n13278), .A2(n13277), .ZN(n13280) );
  MUX2_X1 U15437 ( .A(n13620), .B(n13878), .S(n13372), .Z(n13287) );
  INV_X2 U15438 ( .A(n13878), .ZN(n14019) );
  MUX2_X1 U15439 ( .A(n13886), .B(n14019), .S(n6404), .Z(n13286) );
  NAND2_X1 U15440 ( .A1(n13287), .A2(n13286), .ZN(n13279) );
  NAND4_X1 U15441 ( .A1(n13285), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13282) );
  AOI21_X1 U15442 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(n13295) );
  INV_X1 U15443 ( .A(n13285), .ZN(n13293) );
  INV_X1 U15444 ( .A(n13286), .ZN(n13289) );
  INV_X1 U15445 ( .A(n13287), .ZN(n13288) );
  XNOR2_X1 U15446 ( .A(n14013), .B(n13870), .ZN(n13859) );
  AOI21_X1 U15447 ( .B1(n13289), .B2(n13288), .A(n13859), .ZN(n13292) );
  NOR2_X1 U15448 ( .A1(n14008), .A2(n13848), .ZN(n13291) );
  OAI22_X1 U15449 ( .A1(n13293), .A2(n13292), .B1(n13291), .B2(n13290), .ZN(
        n13294) );
  MUX2_X1 U15450 ( .A(n13797), .B(n14004), .S(n13372), .Z(n13296) );
  MUX2_X1 U15451 ( .A(n13797), .B(n14004), .S(n6404), .Z(n13297) );
  MUX2_X1 U15452 ( .A(n13628), .B(n13997), .S(n6404), .Z(n13298) );
  MUX2_X1 U15453 ( .A(n13628), .B(n13997), .S(n13372), .Z(n13300) );
  MUX2_X1 U15454 ( .A(n13798), .B(n13993), .S(n6407), .Z(n13302) );
  MUX2_X1 U15455 ( .A(n13798), .B(n13993), .S(n6404), .Z(n13301) );
  INV_X1 U15456 ( .A(n13302), .ZN(n13303) );
  MUX2_X1 U15457 ( .A(n13630), .B(n13988), .S(n6404), .Z(n13307) );
  MUX2_X1 U15458 ( .A(n13630), .B(n13988), .S(n6407), .Z(n13304) );
  NAND2_X1 U15459 ( .A1(n13305), .A2(n13304), .ZN(n13311) );
  INV_X1 U15460 ( .A(n13306), .ZN(n13309) );
  INV_X1 U15461 ( .A(n13307), .ZN(n13308) );
  NAND2_X1 U15462 ( .A1(n13309), .A2(n13308), .ZN(n13310) );
  NAND2_X1 U15463 ( .A1(n13311), .A2(n13310), .ZN(n13313) );
  MUX2_X1 U15464 ( .A(n13631), .B(n13982), .S(n6407), .Z(n13314) );
  MUX2_X1 U15465 ( .A(n13631), .B(n13982), .S(n6404), .Z(n13312) );
  INV_X1 U15466 ( .A(n13314), .ZN(n13315) );
  MUX2_X1 U15467 ( .A(n13584), .B(n13978), .S(n6404), .Z(n13318) );
  MUX2_X1 U15468 ( .A(n13584), .B(n13978), .S(n6407), .Z(n13316) );
  NAND2_X1 U15469 ( .A1(n13317), .A2(n13316), .ZN(n13319) );
  MUX2_X1 U15470 ( .A(n13701), .B(n13972), .S(n13372), .Z(n13321) );
  MUX2_X1 U15471 ( .A(n13741), .B(n7554), .S(n6404), .Z(n13320) );
  NOR2_X1 U15472 ( .A1(n13322), .A2(n13321), .ZN(n13323) );
  MUX2_X1 U15473 ( .A(n13637), .B(n13708), .S(n13372), .Z(n13329) );
  MUX2_X1 U15474 ( .A(n13682), .B(n13967), .S(n6404), .Z(n13328) );
  OAI22_X1 U15475 ( .A1(n13324), .A2(n13323), .B1(n13329), .B2(n13328), .ZN(
        n13331) );
  MUX2_X1 U15476 ( .A(n13668), .B(n13656), .S(n13372), .Z(n13352) );
  NAND2_X1 U15477 ( .A1(n13594), .A2(n13372), .ZN(n13325) );
  NAND2_X1 U15478 ( .A1(n13352), .A2(n13351), .ZN(n13341) );
  MUX2_X1 U15479 ( .A(n13640), .B(n13960), .S(n6407), .Z(n13338) );
  INV_X1 U15480 ( .A(n13640), .ZN(n13681) );
  MUX2_X1 U15481 ( .A(n6735), .B(n13681), .S(n13372), .Z(n13337) );
  NAND2_X1 U15482 ( .A1(n13338), .A2(n13337), .ZN(n13327) );
  MUX2_X1 U15483 ( .A(n13667), .B(n13692), .S(n6407), .Z(n13334) );
  MUX2_X1 U15484 ( .A(n13702), .B(n13962), .S(n6404), .Z(n13333) );
  AOI22_X1 U15485 ( .A1(n13334), .A2(n13333), .B1(n13329), .B2(n13328), .ZN(
        n13330) );
  INV_X1 U15486 ( .A(n13332), .ZN(n13360) );
  INV_X1 U15487 ( .A(n13333), .ZN(n13336) );
  INV_X1 U15488 ( .A(n13334), .ZN(n13335) );
  NAND2_X1 U15489 ( .A1(n13336), .A2(n13335), .ZN(n13359) );
  INV_X1 U15490 ( .A(n13337), .ZN(n13340) );
  INV_X1 U15491 ( .A(n13338), .ZN(n13339) );
  NAND3_X1 U15492 ( .A1(n13341), .A2(n13340), .A3(n13339), .ZN(n13358) );
  NAND2_X1 U15493 ( .A1(n13342), .A2(n6408), .ZN(n13344) );
  OR2_X1 U15494 ( .A1(n13369), .A2(n14090), .ZN(n13343) );
  MUX2_X1 U15495 ( .A(n13391), .B(n13604), .S(n6407), .Z(n13379) );
  INV_X1 U15496 ( .A(n13391), .ZN(n13439) );
  MUX2_X1 U15497 ( .A(n13439), .B(n13947), .S(n6404), .Z(n13378) );
  NAND2_X1 U15498 ( .A1(n14087), .A2(n6408), .ZN(n13346) );
  INV_X1 U15499 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14083) );
  OR2_X1 U15500 ( .A1(n13369), .A2(n14083), .ZN(n13345) );
  INV_X1 U15501 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13349) );
  NAND2_X1 U15502 ( .A1(n13362), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13348) );
  NAND2_X1 U15503 ( .A1(n9079), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n13347) );
  OAI211_X1 U15504 ( .C1(n13365), .C2(n13349), .A(n13348), .B(n13347), .ZN(
        n13547) );
  OR2_X1 U15505 ( .A1(n13386), .A2(n13547), .ZN(n13387) );
  NAND2_X1 U15506 ( .A1(n13386), .A2(n13547), .ZN(n13350) );
  NAND2_X1 U15507 ( .A1(n13387), .A2(n13350), .ZN(n13417) );
  INV_X1 U15508 ( .A(n13351), .ZN(n13354) );
  INV_X1 U15509 ( .A(n13352), .ZN(n13353) );
  NAND2_X1 U15510 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  OAI211_X1 U15511 ( .C1(n13379), .C2(n13378), .A(n13417), .B(n13355), .ZN(
        n13356) );
  INV_X1 U15512 ( .A(n13356), .ZN(n13357) );
  INV_X1 U15513 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U15514 ( .A1(n13362), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U15515 ( .A1(n9079), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n13363) );
  OAI211_X1 U15516 ( .C1(n13365), .C2(n15569), .A(n13364), .B(n13363), .ZN(
        n13592) );
  NAND2_X1 U15517 ( .A1(n13367), .A2(n13366), .ZN(n13371) );
  OR2_X1 U15518 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  MUX2_X1 U15519 ( .A(n13592), .B(n13544), .S(n6407), .Z(n13385) );
  OR2_X1 U15520 ( .A1(n13374), .A2(n13373), .ZN(n13427) );
  NAND2_X1 U15521 ( .A1(n13372), .A2(n13547), .ZN(n13388) );
  NAND4_X1 U15522 ( .A1(n13427), .A2(n13388), .A3(n13421), .A4(n13423), .ZN(
        n13375) );
  AND2_X1 U15523 ( .A1(n13375), .A2(n13592), .ZN(n13376) );
  AOI21_X1 U15524 ( .B1(n13544), .B2(n6404), .A(n13376), .ZN(n13384) );
  INV_X1 U15525 ( .A(n13378), .ZN(n13381) );
  INV_X1 U15526 ( .A(n13379), .ZN(n13380) );
  OAI22_X1 U15527 ( .A1(n13385), .A2(n13384), .B1(n13381), .B2(n13380), .ZN(
        n13382) );
  NAND2_X1 U15528 ( .A1(n13382), .A2(n13417), .ZN(n13383) );
  OAI211_X1 U15529 ( .C1(n13942), .C2(n6407), .A(n13388), .B(n13387), .ZN(
        n13389) );
  INV_X1 U15530 ( .A(n13592), .ZN(n13390) );
  XNOR2_X1 U15531 ( .A(n13544), .B(n13390), .ZN(n13415) );
  NAND2_X1 U15532 ( .A1(n13962), .A2(n13667), .ZN(n13663) );
  XNOR2_X1 U15533 ( .A(n13978), .B(n13633), .ZN(n13737) );
  XNOR2_X1 U15534 ( .A(n13982), .B(n13740), .ZN(n13755) );
  NAND2_X1 U15535 ( .A1(n13993), .A2(n13629), .ZN(n13579) );
  OR2_X1 U15536 ( .A1(n13993), .A2(n13629), .ZN(n13393) );
  NAND2_X1 U15537 ( .A1(n13579), .A2(n13393), .ZN(n13779) );
  NAND2_X1 U15538 ( .A1(n14036), .A2(n13611), .ZN(n13565) );
  NAND2_X1 U15539 ( .A1(n13903), .A2(n13565), .ZN(n13933) );
  NAND4_X1 U15540 ( .A1(n14057), .A2(n13395), .A3(n13394), .A4(n9999), .ZN(
        n13400) );
  NAND2_X1 U15541 ( .A1(n13397), .A2(n13396), .ZN(n13398) );
  NAND4_X1 U15542 ( .A1(n13404), .A2(n13403), .A3(n13402), .A4(n13401), .ZN(
        n13405) );
  NOR2_X1 U15543 ( .A1(n13933), .A2(n13407), .ZN(n13409) );
  NAND2_X1 U15544 ( .A1(n13569), .A2(n13568), .ZN(n13617) );
  NAND2_X1 U15545 ( .A1(n13618), .A2(n13617), .ZN(n13896) );
  NAND4_X1 U15546 ( .A1(n13409), .A2(n13913), .A3(n13896), .A4(n13408), .ZN(
        n13410) );
  XNOR2_X1 U15547 ( .A(n14008), .B(n13573), .ZN(n13835) );
  NOR2_X1 U15548 ( .A1(n13779), .A2(n13411), .ZN(n13412) );
  XNOR2_X1 U15549 ( .A(n13988), .B(n13630), .ZN(n13764) );
  XNOR2_X1 U15550 ( .A(n14004), .B(n13797), .ZN(n13821) );
  NAND4_X1 U15551 ( .A1(n13412), .A2(n13764), .A3(n13821), .A4(n13796), .ZN(
        n13413) );
  NAND2_X1 U15552 ( .A1(n13967), .A2(n13637), .ZN(n13588) );
  OR2_X1 U15553 ( .A1(n13967), .A2(n13637), .ZN(n13414) );
  NAND2_X1 U15554 ( .A1(n13588), .A2(n13414), .ZN(n13711) );
  NAND2_X1 U15555 ( .A1(n13950), .A2(n13594), .ZN(n13642) );
  OR2_X1 U15556 ( .A1(n13950), .A2(n13594), .ZN(n13416) );
  NAND2_X1 U15557 ( .A1(n13642), .A2(n13416), .ZN(n13641) );
  AOI211_X1 U15558 ( .C1(n13420), .C2(n13419), .A(n13421), .B(n13418), .ZN(
        n13432) );
  INV_X1 U15559 ( .A(n13420), .ZN(n13431) );
  NAND2_X1 U15560 ( .A1(n13428), .A2(n13421), .ZN(n13422) );
  OAI211_X1 U15561 ( .C1(n6414), .C2(n13424), .A(n13423), .B(n13422), .ZN(
        n13425) );
  OAI21_X1 U15562 ( .B1(n13429), .B2(n13428), .A(n13427), .ZN(n13430) );
  INV_X1 U15563 ( .A(n13433), .ZN(n13437) );
  INV_X1 U15564 ( .A(n13434), .ZN(n13546) );
  NAND4_X1 U15565 ( .A1(n15359), .A2(n13546), .A3(n13883), .A4(n13435), .ZN(
        n13436) );
  OAI211_X1 U15566 ( .C1(n6414), .C2(n13437), .A(n13436), .B(P2_B_REG_SCAN_IN), 
        .ZN(n13438) );
  MUX2_X1 U15567 ( .A(n13547), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13451), .Z(
        P2_U3562) );
  MUX2_X1 U15568 ( .A(n13592), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13451), .Z(
        P2_U3561) );
  MUX2_X1 U15569 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13439), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15570 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13594), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15571 ( .A(n13681), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13451), .Z(
        P2_U3558) );
  MUX2_X1 U15572 ( .A(n13702), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13451), .Z(
        P2_U3557) );
  MUX2_X1 U15573 ( .A(n13682), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13451), .Z(
        P2_U3556) );
  MUX2_X1 U15574 ( .A(n13701), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13451), .Z(
        P2_U3555) );
  MUX2_X1 U15575 ( .A(n13584), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13451), .Z(
        P2_U3554) );
  MUX2_X1 U15576 ( .A(n13631), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13451), .Z(
        P2_U3553) );
  MUX2_X1 U15577 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13630), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15578 ( .A(n13798), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13451), .Z(
        P2_U3551) );
  MUX2_X1 U15579 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13628), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15580 ( .A(n13797), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13451), .Z(
        P2_U3549) );
  MUX2_X1 U15581 ( .A(n13848), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13451), .Z(
        P2_U3548) );
  MUX2_X1 U15582 ( .A(n13623), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13451), .Z(
        P2_U3547) );
  MUX2_X1 U15583 ( .A(n13886), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13451), .Z(
        P2_U3546) );
  MUX2_X1 U15584 ( .A(n13568), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13451), .Z(
        P2_U3545) );
  MUX2_X1 U15585 ( .A(n13884), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13451), .Z(
        P2_U3544) );
  MUX2_X1 U15586 ( .A(n13440), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13451), .Z(
        P2_U3543) );
  MUX2_X1 U15587 ( .A(n13566), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13451), .Z(
        P2_U3542) );
  MUX2_X1 U15588 ( .A(n13441), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13451), .Z(
        P2_U3541) );
  MUX2_X1 U15589 ( .A(n13442), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13451), .Z(
        P2_U3540) );
  MUX2_X1 U15590 ( .A(n13443), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13451), .Z(
        P2_U3539) );
  MUX2_X1 U15591 ( .A(n13444), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13451), .Z(
        P2_U3538) );
  MUX2_X1 U15592 ( .A(n13445), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13451), .Z(
        P2_U3537) );
  MUX2_X1 U15593 ( .A(n13446), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13451), .Z(
        P2_U3536) );
  MUX2_X1 U15594 ( .A(n13447), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13451), .Z(
        P2_U3535) );
  MUX2_X1 U15595 ( .A(n13448), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13451), .Z(
        P2_U3534) );
  MUX2_X1 U15596 ( .A(n13449), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13451), .Z(
        P2_U3533) );
  MUX2_X1 U15597 ( .A(n13450), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13451), .Z(
        P2_U3532) );
  MUX2_X1 U15598 ( .A(n13452), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13451), .Z(
        P2_U3531) );
  MUX2_X1 U15599 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10188), .S(n13458), .Z(
        n13455) );
  INV_X1 U15600 ( .A(n13453), .ZN(n13454) );
  NAND2_X1 U15601 ( .A1(n13455), .A2(n13454), .ZN(n13456) );
  OAI211_X1 U15602 ( .C1(n13457), .C2(n13456), .A(n15315), .B(n13476), .ZN(
        n13467) );
  MUX2_X1 U15603 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11263), .S(n13458), .Z(
        n13461) );
  NAND3_X1 U15604 ( .A1(n13461), .A2(n13460), .A3(n13459), .ZN(n13462) );
  NAND3_X1 U15605 ( .A1(n15318), .A2(n13470), .A3(n13462), .ZN(n13466) );
  AOI22_X1 U15606 ( .A1(n15305), .A2(n13463), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13465) );
  NAND2_X1 U15607 ( .A1(n15273), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n13464) );
  NAND4_X1 U15608 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        P2_U3216) );
  MUX2_X1 U15609 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11430), .S(n13468), .Z(
        n13471) );
  NAND3_X1 U15610 ( .A1(n13471), .A2(n13470), .A3(n13469), .ZN(n13472) );
  NAND3_X1 U15611 ( .A1(n15318), .A2(n13473), .A3(n13472), .ZN(n13483) );
  INV_X1 U15612 ( .A(n15278), .ZN(n13478) );
  NAND3_X1 U15613 ( .A1(n13476), .A2(n13475), .A3(n13474), .ZN(n13477) );
  NAND3_X1 U15614 ( .A1(n15315), .A2(n13478), .A3(n13477), .ZN(n13482) );
  AOI22_X1 U15615 ( .A1(n15305), .A2(n13479), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13481) );
  NAND2_X1 U15616 ( .A1(n15273), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n13480) );
  NAND4_X1 U15617 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        P2_U3217) );
  INV_X1 U15618 ( .A(n13489), .ZN(n13488) );
  INV_X1 U15619 ( .A(n13484), .ZN(n13487) );
  NOR2_X1 U15620 ( .A1(n15322), .A2(n13485), .ZN(n13486) );
  AOI211_X1 U15621 ( .C1(n15305), .C2(n13488), .A(n13487), .B(n13486), .ZN(
        n13498) );
  MUX2_X1 U15622 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11275), .S(n13489), .Z(
        n13490) );
  NAND3_X1 U15623 ( .A1(n15284), .A2(n13491), .A3(n13490), .ZN(n13492) );
  NAND3_X1 U15624 ( .A1(n15318), .A2(n13501), .A3(n13492), .ZN(n13497) );
  NAND3_X1 U15625 ( .A1(n15275), .A2(n13494), .A3(n13493), .ZN(n13495) );
  NAND3_X1 U15626 ( .A1(n15315), .A2(n6636), .A3(n13495), .ZN(n13496) );
  NAND3_X1 U15627 ( .A1(n13498), .A2(n13497), .A3(n13496), .ZN(P2_U3219) );
  MUX2_X1 U15628 ( .A(n11634), .B(P2_REG2_REG_6__SCAN_IN), .S(n13509), .Z(
        n13499) );
  NAND3_X1 U15629 ( .A1(n13501), .A2(n13500), .A3(n13499), .ZN(n13502) );
  NAND3_X1 U15630 ( .A1(n15318), .A2(n13503), .A3(n13502), .ZN(n13513) );
  MUX2_X1 U15631 ( .A(n10191), .B(P2_REG1_REG_6__SCAN_IN), .S(n13509), .Z(
        n13504) );
  NAND3_X1 U15632 ( .A1(n6636), .A2(n6637), .A3(n13504), .ZN(n13505) );
  NAND3_X1 U15633 ( .A1(n15315), .A2(n13506), .A3(n13505), .ZN(n13512) );
  INV_X1 U15634 ( .A(n13507), .ZN(n13508) );
  AOI21_X1 U15635 ( .B1(n15305), .B2(n13509), .A(n13508), .ZN(n13511) );
  NAND2_X1 U15636 ( .A1(n15273), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n13510) );
  NAND4_X1 U15637 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        P2_U3220) );
  NAND2_X1 U15638 ( .A1(n13520), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U15639 ( .A1(n13515), .A2(n13514), .ZN(n13516) );
  NAND2_X1 U15640 ( .A1(n13516), .A2(n13532), .ZN(n13517) );
  NAND2_X1 U15641 ( .A1(n13536), .A2(n13517), .ZN(n13519) );
  INV_X1 U15642 ( .A(n13537), .ZN(n13518) );
  AOI21_X1 U15643 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13519), .A(n13518), 
        .ZN(n13529) );
  XNOR2_X1 U15644 ( .A(n13530), .B(n13532), .ZN(n13533) );
  XOR2_X1 U15645 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13533), .Z(n13523) );
  NAND2_X1 U15646 ( .A1(n13523), .A2(n15315), .ZN(n13528) );
  NOR2_X1 U15647 ( .A1(n15313), .A2(n13524), .ZN(n13525) );
  AOI211_X1 U15648 ( .C1(n15273), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13526), 
        .B(n13525), .ZN(n13527) );
  OAI211_X1 U15649 ( .C1(n13529), .C2(n15294), .A(n13528), .B(n13527), .ZN(
        P2_U3232) );
  INV_X1 U15650 ( .A(n13530), .ZN(n13531) );
  AOI22_X1 U15651 ( .A1(n13533), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n13532), 
        .B2(n13531), .ZN(n13535) );
  XNOR2_X1 U15652 ( .A(n13535), .B(n13534), .ZN(n13540) );
  XNOR2_X1 U15653 ( .A(n13538), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13539) );
  OR2_X2 U15654 ( .A1(n13783), .A2(n13993), .ZN(n13784) );
  NOR2_X4 U15655 ( .A1(n13784), .A2(n13988), .ZN(n13768) );
  NAND2_X1 U15656 ( .A1(n13689), .A2(n13960), .ZN(n13669) );
  INV_X1 U15657 ( .A(n13669), .ZN(n13543) );
  NAND2_X1 U15658 ( .A1(n13601), .A2(n13945), .ZN(n13550) );
  XNOR2_X1 U15659 ( .A(n13550), .B(n13942), .ZN(n13545) );
  NAND2_X1 U15660 ( .A1(n13545), .A2(n13889), .ZN(n13941) );
  AOI21_X1 U15661 ( .B1(n13546), .B2(P2_B_REG_SCAN_IN), .A(n13871), .ZN(n13593) );
  NAND2_X1 U15662 ( .A1(n13593), .A2(n13547), .ZN(n13943) );
  NOR2_X1 U15663 ( .A1(n13940), .A2(n13943), .ZN(n13552) );
  NOR2_X1 U15664 ( .A1(n13942), .A2(n13931), .ZN(n13548) );
  AOI211_X1 U15665 ( .C1(n13940), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13552), 
        .B(n13548), .ZN(n13549) );
  OAI21_X1 U15666 ( .B1(n13941), .B2(n13554), .A(n13549), .ZN(P2_U3234) );
  OAI211_X1 U15667 ( .C1(n13601), .C2(n13945), .A(n13889), .B(n13550), .ZN(
        n13944) );
  NOR2_X1 U15668 ( .A1(n13945), .A2(n13931), .ZN(n13551) );
  AOI211_X1 U15669 ( .C1(n13940), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13552), 
        .B(n13551), .ZN(n13553) );
  OAI21_X1 U15670 ( .B1(n13944), .B2(n13554), .A(n13553), .ZN(P2_U3235) );
  INV_X1 U15671 ( .A(n13555), .ZN(n13559) );
  NAND2_X1 U15672 ( .A1(n14051), .A2(n13556), .ZN(n13557) );
  NAND2_X1 U15673 ( .A1(n13559), .A2(n7841), .ZN(n13564) );
  AOI21_X1 U15674 ( .B1(n13609), .B2(n13566), .A(n13560), .ZN(n13561) );
  INV_X1 U15675 ( .A(n13565), .ZN(n13567) );
  NOR2_X1 U15676 ( .A1(n13609), .A2(n13566), .ZN(n13900) );
  NAND2_X1 U15677 ( .A1(n13882), .A2(n7844), .ZN(n13571) );
  NAND2_X1 U15678 ( .A1(n13571), .A2(n13570), .ZN(n13864) );
  NOR2_X1 U15679 ( .A1(n14008), .A2(n13573), .ZN(n13574) );
  NOR2_X1 U15680 ( .A1(n13824), .A2(n13797), .ZN(n13575) );
  NAND2_X1 U15681 ( .A1(n13824), .A2(n13797), .ZN(n13576) );
  NAND2_X1 U15682 ( .A1(n13809), .A2(n13628), .ZN(n13577) );
  INV_X1 U15683 ( .A(n13988), .ZN(n13772) );
  NAND2_X1 U15684 ( .A1(n13772), .A2(n13630), .ZN(n13580) );
  NAND2_X1 U15685 ( .A1(n13988), .A2(n13782), .ZN(n13581) );
  NAND2_X1 U15686 ( .A1(n13754), .A2(n13631), .ZN(n13582) );
  NAND2_X1 U15687 ( .A1(n13978), .A2(n13633), .ZN(n13583) );
  NAND2_X1 U15688 ( .A1(n13736), .A2(n13584), .ZN(n13585) );
  INV_X1 U15689 ( .A(n13719), .ZN(n13586) );
  NAND2_X1 U15690 ( .A1(n13972), .A2(n13741), .ZN(n13587) );
  INV_X1 U15691 ( .A(n13711), .ZN(n13700) );
  NAND2_X1 U15692 ( .A1(n13662), .A2(n13663), .ZN(n13590) );
  INV_X1 U15693 ( .A(n13674), .ZN(n13589) );
  NAND2_X1 U15694 ( .A1(n6735), .A2(n13640), .ZN(n13591) );
  AOI211_X1 U15695 ( .C1(n13656), .C2(n13594), .A(n13920), .B(n13643), .ZN(
        n13598) );
  NAND4_X1 U15696 ( .A1(n13643), .A2(n13656), .A3(n13594), .A4(n13905), .ZN(
        n13596) );
  AOI22_X1 U15697 ( .A1(n13594), .A2(n13883), .B1(n13593), .B2(n13592), .ZN(
        n13595) );
  NAND2_X1 U15698 ( .A1(n13596), .A2(n13595), .ZN(n13597) );
  AOI21_X1 U15699 ( .B1(n13650), .B2(n13598), .A(n13597), .ZN(n13599) );
  AOI211_X1 U15700 ( .C1(n13947), .C2(n13653), .A(n13926), .B(n13601), .ZN(
        n13946) );
  AOI22_X1 U15701 ( .A1(n13602), .A2(n13928), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13940), .ZN(n13603) );
  OAI21_X1 U15702 ( .B1(n13604), .B2(n13931), .A(n13603), .ZN(n13605) );
  AOI21_X1 U15703 ( .B1(n13946), .B2(n13938), .A(n13605), .ZN(n13647) );
  NAND2_X1 U15704 ( .A1(n13609), .A2(n13608), .ZN(n13606) );
  OR2_X1 U15705 ( .A1(n13609), .A2(n13608), .ZN(n13610) );
  NOR2_X1 U15706 ( .A1(n13932), .A2(n13611), .ZN(n13612) );
  OR2_X1 U15707 ( .A1(n13912), .A2(n13614), .ZN(n13615) );
  INV_X1 U15708 ( .A(n13617), .ZN(n13619) );
  AND2_X1 U15709 ( .A1(n13878), .A2(n13620), .ZN(n13621) );
  NAND2_X1 U15710 ( .A1(n14013), .A2(n13623), .ZN(n13624) );
  OR2_X1 U15711 ( .A1(n14004), .A2(n13797), .ZN(n13627) );
  INV_X1 U15712 ( .A(n13993), .ZN(n13789) );
  NAND2_X1 U15713 ( .A1(n13982), .A2(n13631), .ZN(n13730) );
  AOI21_X1 U15714 ( .B1(n13754), .B2(n13740), .A(n13633), .ZN(n13635) );
  NAND3_X1 U15715 ( .A1(n13754), .A2(n13740), .A3(n13633), .ZN(n13634) );
  NAND2_X1 U15716 ( .A1(n13720), .A2(n13719), .ZN(n13718) );
  NAND2_X1 U15717 ( .A1(n13708), .A2(n13637), .ZN(n13638) );
  NAND2_X1 U15718 ( .A1(n13962), .A2(n13702), .ZN(n13639) );
  XNOR2_X1 U15719 ( .A(n13644), .B(n13643), .ZN(n13948) );
  INV_X1 U15720 ( .A(n13948), .ZN(n13645) );
  NAND2_X1 U15721 ( .A1(n13645), .A2(n13897), .ZN(n13646) );
  OAI211_X1 U15722 ( .C1(n6464), .C2(n13940), .A(n13647), .B(n13646), .ZN(
        P2_U3236) );
  AOI21_X1 U15723 ( .B1(n13648), .B2(n13657), .A(n13920), .ZN(n13649) );
  NAND2_X1 U15724 ( .A1(n13950), .A2(n13669), .ZN(n13652) );
  AOI22_X1 U15725 ( .A1(n13654), .A2(n13928), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n13940), .ZN(n13655) );
  OAI21_X1 U15726 ( .B1(n13656), .B2(n13931), .A(n13655), .ZN(n13660) );
  NOR2_X1 U15727 ( .A1(n13952), .A2(n13935), .ZN(n13659) );
  OAI21_X1 U15728 ( .B1(n13955), .B2(n13940), .A(n13661), .ZN(P2_U3237) );
  NAND3_X1 U15729 ( .A1(n13680), .A2(n13674), .A3(n13663), .ZN(n13664) );
  NAND2_X1 U15730 ( .A1(n13956), .A2(n13880), .ZN(n13678) );
  OAI211_X1 U15731 ( .C1(n13689), .C2(n13960), .A(n13889), .B(n13669), .ZN(
        n13958) );
  INV_X1 U15732 ( .A(n13958), .ZN(n13673) );
  AOI22_X1 U15733 ( .A1(n13670), .A2(n13928), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13940), .ZN(n13671) );
  OAI21_X1 U15734 ( .B1(n13960), .B2(n13931), .A(n13671), .ZN(n13672) );
  AOI21_X1 U15735 ( .B1(n13673), .B2(n13938), .A(n13672), .ZN(n13677) );
  NAND3_X1 U15736 ( .A1(n13957), .A2(n13675), .A3(n13897), .ZN(n13676) );
  NAND3_X1 U15737 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(P2_U3238) );
  NAND2_X1 U15738 ( .A1(n13681), .A2(n13885), .ZN(n13684) );
  NAND2_X1 U15739 ( .A1(n13682), .A2(n13883), .ZN(n13683) );
  NAND2_X1 U15740 ( .A1(n13705), .A2(n13962), .ZN(n13687) );
  NAND2_X1 U15741 ( .A1(n13687), .A2(n13889), .ZN(n13688) );
  NOR2_X1 U15742 ( .A1(n13689), .A2(n13688), .ZN(n13961) );
  AOI22_X1 U15743 ( .A1(n13690), .A2(n13928), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13940), .ZN(n13691) );
  OAI21_X1 U15744 ( .B1(n13692), .B2(n13931), .A(n13691), .ZN(n13693) );
  AOI21_X1 U15745 ( .B1(n13961), .B2(n13938), .A(n13693), .ZN(n13697) );
  XNOR2_X1 U15746 ( .A(n13694), .B(n6493), .ZN(n13965) );
  INV_X1 U15747 ( .A(n13965), .ZN(n13695) );
  NAND2_X1 U15748 ( .A1(n13695), .A2(n13897), .ZN(n13696) );
  OAI211_X1 U15749 ( .C1(n13964), .C2(n13940), .A(n13697), .B(n13696), .ZN(
        P2_U3239) );
  OAI21_X1 U15750 ( .B1(n13700), .B2(n13699), .A(n13698), .ZN(n13703) );
  AOI222_X1 U15751 ( .A1(n13905), .A2(n13703), .B1(n13702), .B2(n13885), .C1(
        n13701), .C2(n13883), .ZN(n13969) );
  AOI21_X1 U15752 ( .B1(n13724), .B2(n13967), .A(n13926), .ZN(n13704) );
  AND2_X1 U15753 ( .A1(n13705), .A2(n13704), .ZN(n13966) );
  AOI22_X1 U15754 ( .A1(n13706), .A2(n13928), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13940), .ZN(n13707) );
  OAI21_X1 U15755 ( .B1(n13708), .B2(n13931), .A(n13707), .ZN(n13709) );
  AOI21_X1 U15756 ( .B1(n13966), .B2(n13938), .A(n13709), .ZN(n13714) );
  XNOR2_X1 U15757 ( .A(n13710), .B(n13711), .ZN(n13970) );
  INV_X1 U15758 ( .A(n13970), .ZN(n13712) );
  NAND2_X1 U15759 ( .A1(n13712), .A2(n13897), .ZN(n13713) );
  OAI211_X1 U15760 ( .C1(n13969), .C2(n13940), .A(n13714), .B(n13713), .ZN(
        P2_U3240) );
  XNOR2_X1 U15761 ( .A(n13719), .B(n13715), .ZN(n13717) );
  AOI21_X1 U15762 ( .B1(n13717), .B2(n13905), .A(n13716), .ZN(n13974) );
  OAI21_X1 U15763 ( .B1(n13720), .B2(n13719), .A(n13718), .ZN(n13975) );
  INV_X1 U15764 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13721) );
  OAI22_X1 U15765 ( .A1(n13722), .A2(n13837), .B1(n13721), .B2(n13880), .ZN(
        n13723) );
  AOI21_X1 U15766 ( .B1(n13972), .B2(n13853), .A(n13723), .ZN(n13727) );
  AOI21_X1 U15767 ( .B1(n13732), .B2(n13972), .A(n13926), .ZN(n13725) );
  AND2_X1 U15768 ( .A1(n13725), .A2(n13724), .ZN(n13971) );
  NAND2_X1 U15769 ( .A1(n13971), .A2(n13938), .ZN(n13726) );
  OAI211_X1 U15770 ( .C1(n13975), .C2(n13915), .A(n13727), .B(n13726), .ZN(
        n13728) );
  INV_X1 U15771 ( .A(n13728), .ZN(n13729) );
  OAI21_X1 U15772 ( .B1(n13974), .B2(n13940), .A(n13729), .ZN(P2_U3241) );
  NAND2_X1 U15773 ( .A1(n13748), .A2(n13755), .ZN(n13747) );
  NAND2_X1 U15774 ( .A1(n13747), .A2(n13730), .ZN(n13731) );
  XNOR2_X1 U15775 ( .A(n13731), .B(n13737), .ZN(n13980) );
  INV_X1 U15776 ( .A(n13749), .ZN(n13734) );
  INV_X1 U15777 ( .A(n13732), .ZN(n13733) );
  AOI211_X1 U15778 ( .C1(n13978), .C2(n13734), .A(n13926), .B(n13733), .ZN(
        n13977) );
  INV_X1 U15779 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13735) );
  OAI22_X1 U15780 ( .A1(n13736), .A2(n13931), .B1(n13735), .B2(n13880), .ZN(
        n13745) );
  XOR2_X1 U15781 ( .A(n13738), .B(n13737), .Z(n13739) );
  OAI222_X1 U15782 ( .A1(n13871), .A2(n13741), .B1(n13869), .B2(n13740), .C1(
        n13739), .C2(n13920), .ZN(n13976) );
  AOI21_X1 U15783 ( .B1(n13742), .B2(n13928), .A(n13976), .ZN(n13743) );
  NOR2_X1 U15784 ( .A1(n13743), .A2(n13940), .ZN(n13744) );
  AOI211_X1 U15785 ( .C1(n13977), .C2(n13938), .A(n13745), .B(n13744), .ZN(
        n13746) );
  OAI21_X1 U15786 ( .B1(n13915), .B2(n13980), .A(n13746), .ZN(P2_U3242) );
  OAI21_X1 U15787 ( .B1(n13748), .B2(n13755), .A(n13747), .ZN(n13985) );
  INV_X1 U15788 ( .A(n13768), .ZN(n13750) );
  AOI211_X1 U15789 ( .C1(n13982), .C2(n13750), .A(n13926), .B(n13749), .ZN(
        n13981) );
  INV_X1 U15790 ( .A(n13751), .ZN(n13752) );
  AOI22_X1 U15791 ( .A1(n13752), .A2(n13928), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13940), .ZN(n13753) );
  OAI21_X1 U15792 ( .B1(n13754), .B2(n13931), .A(n13753), .ZN(n13761) );
  AOI21_X1 U15793 ( .B1(n13756), .B2(n13755), .A(n13920), .ZN(n13759) );
  AOI21_X1 U15794 ( .B1(n13759), .B2(n13758), .A(n13757), .ZN(n13984) );
  NOR2_X1 U15795 ( .A1(n13984), .A2(n13940), .ZN(n13760) );
  AOI211_X1 U15796 ( .C1(n13981), .C2(n13938), .A(n13761), .B(n13760), .ZN(
        n13762) );
  OAI21_X1 U15797 ( .B1(n13915), .B2(n13985), .A(n13762), .ZN(P2_U3243) );
  XOR2_X1 U15798 ( .A(n13763), .B(n13764), .Z(n13990) );
  XOR2_X1 U15799 ( .A(n13765), .B(n13764), .Z(n13767) );
  OAI21_X1 U15800 ( .B1(n13767), .B2(n13920), .A(n13766), .ZN(n13986) );
  AOI211_X1 U15801 ( .C1(n13988), .C2(n13784), .A(n13926), .B(n13768), .ZN(
        n13987) );
  NAND2_X1 U15802 ( .A1(n13987), .A2(n13938), .ZN(n13771) );
  AOI22_X1 U15803 ( .A1(n13940), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13769), 
        .B2(n13928), .ZN(n13770) );
  OAI211_X1 U15804 ( .C1(n13772), .C2(n13931), .A(n13771), .B(n13770), .ZN(
        n13773) );
  AOI21_X1 U15805 ( .B1(n13986), .B2(n13880), .A(n13773), .ZN(n13774) );
  OAI21_X1 U15806 ( .B1(n13915), .B2(n13990), .A(n13774), .ZN(P2_U3244) );
  XNOR2_X1 U15807 ( .A(n13775), .B(n13779), .ZN(n13995) );
  INV_X1 U15808 ( .A(n13776), .ZN(n13777) );
  AOI21_X1 U15809 ( .B1(n13779), .B2(n13778), .A(n13777), .ZN(n13780) );
  OAI222_X1 U15810 ( .A1(n13871), .A2(n13782), .B1(n13869), .B2(n13781), .C1(
        n13920), .C2(n13780), .ZN(n13991) );
  INV_X1 U15811 ( .A(n13784), .ZN(n13785) );
  AOI211_X1 U15812 ( .C1(n13993), .C2(n13783), .A(n13926), .B(n13785), .ZN(
        n13992) );
  NAND2_X1 U15813 ( .A1(n13992), .A2(n13938), .ZN(n13788) );
  AOI22_X1 U15814 ( .A1(n13940), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13786), 
        .B2(n13928), .ZN(n13787) );
  OAI211_X1 U15815 ( .C1(n13789), .C2(n13931), .A(n13788), .B(n13787), .ZN(
        n13790) );
  AOI21_X1 U15816 ( .B1(n13991), .B2(n13880), .A(n13790), .ZN(n13791) );
  OAI21_X1 U15817 ( .B1(n13915), .B2(n13995), .A(n13791), .ZN(P2_U3245) );
  INV_X1 U15818 ( .A(n13796), .ZN(n13792) );
  XNOR2_X1 U15819 ( .A(n13793), .B(n13792), .ZN(n13810) );
  XNOR2_X1 U15820 ( .A(n13795), .B(n13796), .ZN(n13800) );
  AOI22_X1 U15821 ( .A1(n13798), .A2(n13885), .B1(n13883), .B2(n13797), .ZN(
        n13799) );
  OAI21_X1 U15822 ( .B1(n13800), .B2(n13920), .A(n13799), .ZN(n13801) );
  AOI21_X1 U15823 ( .B1(n13802), .B2(n13810), .A(n13801), .ZN(n13999) );
  INV_X1 U15824 ( .A(n13803), .ZN(n13805) );
  INV_X1 U15825 ( .A(n13783), .ZN(n13804) );
  AOI211_X1 U15826 ( .C1(n13997), .C2(n13805), .A(n13926), .B(n13804), .ZN(
        n13996) );
  INV_X1 U15827 ( .A(n13806), .ZN(n13807) );
  AOI22_X1 U15828 ( .A1(n13940), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13807), 
        .B2(n13928), .ZN(n13808) );
  OAI21_X1 U15829 ( .B1(n13809), .B2(n13931), .A(n13808), .ZN(n13813) );
  INV_X1 U15830 ( .A(n13810), .ZN(n14000) );
  NOR2_X1 U15831 ( .A1(n14000), .A2(n13811), .ZN(n13812) );
  AOI211_X1 U15832 ( .C1(n13996), .C2(n13938), .A(n13813), .B(n13812), .ZN(
        n13814) );
  OAI21_X1 U15833 ( .B1(n13999), .B2(n13940), .A(n13814), .ZN(P2_U3246) );
  XNOR2_X1 U15834 ( .A(n13815), .B(n13821), .ZN(n13817) );
  AOI21_X1 U15835 ( .B1(n13817), .B2(n13905), .A(n13816), .ZN(n14006) );
  INV_X1 U15836 ( .A(n13818), .ZN(n13819) );
  AOI21_X1 U15837 ( .B1(n13821), .B2(n13820), .A(n13819), .ZN(n14001) );
  OAI22_X1 U15838 ( .A1(n13880), .A2(n6664), .B1(n13822), .B2(n13837), .ZN(
        n13823) );
  AOI21_X1 U15839 ( .B1(n14004), .B2(n13853), .A(n13823), .ZN(n13827) );
  OAI21_X1 U15840 ( .B1(n6603), .B2(n13824), .A(n13889), .ZN(n13825) );
  NOR2_X1 U15841 ( .A1(n13825), .A2(n13803), .ZN(n14003) );
  NAND2_X1 U15842 ( .A1(n14003), .A2(n13938), .ZN(n13826) );
  OAI211_X1 U15843 ( .C1(n14001), .C2(n13935), .A(n13827), .B(n13826), .ZN(
        n13828) );
  INV_X1 U15844 ( .A(n13828), .ZN(n13829) );
  OAI21_X1 U15845 ( .B1(n14006), .B2(n13940), .A(n13829), .ZN(P2_U3247) );
  XNOR2_X1 U15846 ( .A(n13830), .B(n13835), .ZN(n13833) );
  INV_X1 U15847 ( .A(n13831), .ZN(n13832) );
  AOI21_X1 U15848 ( .B1(n13833), .B2(n13905), .A(n13832), .ZN(n14010) );
  OAI21_X1 U15849 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n14011) );
  OAI22_X1 U15850 ( .A1(n13880), .A2(n13839), .B1(n13838), .B2(n13837), .ZN(
        n13840) );
  AOI21_X1 U15851 ( .B1(n14008), .B2(n13853), .A(n13840), .ZN(n13844) );
  NAND2_X1 U15852 ( .A1(n13851), .A2(n14008), .ZN(n13841) );
  NAND2_X1 U15853 ( .A1(n13841), .A2(n13889), .ZN(n13842) );
  NOR2_X1 U15854 ( .A1(n6603), .A2(n13842), .ZN(n14007) );
  NAND2_X1 U15855 ( .A1(n14007), .A2(n13938), .ZN(n13843) );
  OAI211_X1 U15856 ( .C1(n14011), .C2(n13915), .A(n13844), .B(n13843), .ZN(
        n13845) );
  INV_X1 U15857 ( .A(n13845), .ZN(n13846) );
  OAI21_X1 U15858 ( .B1(n14010), .B2(n13940), .A(n13846), .ZN(P2_U3248) );
  XOR2_X1 U15859 ( .A(n13859), .B(n13847), .Z(n13849) );
  AOI222_X1 U15860 ( .A1(n13905), .A2(n13849), .B1(n13848), .B2(n13885), .C1(
        n13886), .C2(n13883), .ZN(n14015) );
  AOI21_X1 U15861 ( .B1(n13850), .B2(n14013), .A(n13926), .ZN(n13852) );
  AND2_X1 U15862 ( .A1(n13852), .A2(n13851), .ZN(n14012) );
  NAND2_X1 U15863 ( .A1(n14013), .A2(n13853), .ZN(n13856) );
  NAND2_X1 U15864 ( .A1(n13928), .A2(n13854), .ZN(n13855) );
  OAI211_X1 U15865 ( .C1(n13880), .C2(n13857), .A(n13856), .B(n13855), .ZN(
        n13861) );
  OAI21_X1 U15866 ( .B1(n13859), .B2(n6593), .A(n13858), .ZN(n14016) );
  NOR2_X1 U15867 ( .A1(n14016), .A2(n13915), .ZN(n13860) );
  AOI211_X1 U15868 ( .C1(n14012), .C2(n13938), .A(n13861), .B(n13860), .ZN(
        n13862) );
  OAI21_X1 U15869 ( .B1(n14015), .B2(n13940), .A(n13862), .ZN(P2_U3249) );
  XNOR2_X1 U15870 ( .A(n13863), .B(n13866), .ZN(n14021) );
  XNOR2_X1 U15871 ( .A(n13865), .B(n13866), .ZN(n13867) );
  OAI222_X1 U15872 ( .A1(n13871), .A2(n13870), .B1(n13869), .B2(n13868), .C1(
        n13867), .C2(n13920), .ZN(n14017) );
  INV_X1 U15873 ( .A(n13872), .ZN(n13890) );
  INV_X1 U15874 ( .A(n13850), .ZN(n13873) );
  AOI211_X1 U15875 ( .C1(n14019), .C2(n13890), .A(n13926), .B(n13873), .ZN(
        n14018) );
  NAND2_X1 U15876 ( .A1(n14018), .A2(n13938), .ZN(n13877) );
  INV_X1 U15877 ( .A(n13874), .ZN(n13875) );
  AOI22_X1 U15878 ( .A1(n13940), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13875), 
        .B2(n13928), .ZN(n13876) );
  OAI211_X1 U15879 ( .C1(n13878), .C2(n13931), .A(n13877), .B(n13876), .ZN(
        n13879) );
  AOI21_X1 U15880 ( .B1(n14017), .B2(n13880), .A(n13879), .ZN(n13881) );
  OAI21_X1 U15881 ( .B1(n13915), .B2(n14021), .A(n13881), .ZN(P2_U3250) );
  XOR2_X1 U15882 ( .A(n13882), .B(n13896), .Z(n13887) );
  AOI222_X1 U15883 ( .A1(n13905), .A2(n13887), .B1(n13886), .B2(n13885), .C1(
        n13884), .C2(n13883), .ZN(n14023) );
  OAI211_X1 U15884 ( .C1(n14025), .C2(n13888), .A(n13890), .B(n13889), .ZN(
        n14022) );
  INV_X1 U15885 ( .A(n14022), .ZN(n13894) );
  AOI22_X1 U15886 ( .A1(n13940), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13891), 
        .B2(n13928), .ZN(n13892) );
  OAI21_X1 U15887 ( .B1(n14025), .B2(n13931), .A(n13892), .ZN(n13893) );
  AOI21_X1 U15888 ( .B1(n13894), .B2(n13938), .A(n13893), .ZN(n13899) );
  XNOR2_X1 U15889 ( .A(n13895), .B(n13896), .ZN(n14027) );
  NAND2_X1 U15890 ( .A1(n14027), .A2(n13897), .ZN(n13898) );
  OAI211_X1 U15891 ( .C1(n14023), .C2(n13940), .A(n13899), .B(n13898), .ZN(
        P2_U3251) );
  INV_X1 U15892 ( .A(n13900), .ZN(n13901) );
  NAND2_X1 U15893 ( .A1(n13902), .A2(n13901), .ZN(n13921) );
  NOR2_X1 U15894 ( .A1(n13921), .A2(n13933), .ZN(n13919) );
  INV_X1 U15895 ( .A(n13913), .ZN(n13904) );
  NAND2_X1 U15896 ( .A1(n13904), .A2(n13903), .ZN(n13907) );
  OAI211_X1 U15897 ( .C1(n13919), .C2(n13907), .A(n13906), .B(n13905), .ZN(
        n13909) );
  AND2_X1 U15898 ( .A1(n13909), .A2(n13908), .ZN(n14033) );
  AOI211_X1 U15899 ( .C1(n14031), .C2(n13924), .A(n13926), .B(n13888), .ZN(
        n14030) );
  AOI22_X1 U15900 ( .A1(n13940), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13910), 
        .B2(n13928), .ZN(n13911) );
  OAI21_X1 U15901 ( .B1(n13912), .B2(n13931), .A(n13911), .ZN(n13917) );
  XNOR2_X1 U15902 ( .A(n13914), .B(n13913), .ZN(n14034) );
  NOR2_X1 U15903 ( .A1(n14034), .A2(n13915), .ZN(n13916) );
  AOI211_X1 U15904 ( .C1(n14030), .C2(n13938), .A(n13917), .B(n13916), .ZN(
        n13918) );
  OAI21_X1 U15905 ( .B1(n14033), .B2(n13940), .A(n13918), .ZN(P2_U3252) );
  AOI211_X1 U15906 ( .C1(n13933), .C2(n13921), .A(n13920), .B(n13919), .ZN(
        n13923) );
  NOR2_X1 U15907 ( .A1(n13923), .A2(n13922), .ZN(n14038) );
  INV_X1 U15908 ( .A(n13924), .ZN(n13925) );
  AOI211_X1 U15909 ( .C1(n14036), .C2(n13927), .A(n13926), .B(n13925), .ZN(
        n14035) );
  AOI22_X1 U15910 ( .A1(n13940), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n13929), 
        .B2(n13928), .ZN(n13930) );
  OAI21_X1 U15911 ( .B1(n13932), .B2(n13931), .A(n13930), .ZN(n13937) );
  XNOR2_X1 U15912 ( .A(n13934), .B(n13933), .ZN(n14039) );
  NOR2_X1 U15913 ( .A1(n14039), .A2(n13935), .ZN(n13936) );
  AOI211_X1 U15914 ( .C1(n14035), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        n13939) );
  OAI21_X1 U15915 ( .B1(n14038), .B2(n13940), .A(n13939), .ZN(P2_U3253) );
  OAI211_X1 U15916 ( .C1(n13942), .C2(n14024), .A(n13941), .B(n13943), .ZN(
        n14058) );
  MUX2_X1 U15917 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14058), .S(n15390), .Z(
        P2_U3530) );
  OAI211_X1 U15918 ( .C1(n13945), .C2(n14024), .A(n13944), .B(n13943), .ZN(
        n14059) );
  MUX2_X1 U15919 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14059), .S(n15390), .Z(
        P2_U3529) );
  AOI21_X1 U15920 ( .B1(n15377), .B2(n13950), .A(n13949), .ZN(n13951) );
  NAND2_X1 U15921 ( .A1(n13955), .A2(n13954), .ZN(n14060) );
  MUX2_X1 U15922 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14060), .S(n15390), .Z(
        P2_U3527) );
  NAND3_X1 U15923 ( .A1(n13957), .A2(n13675), .A3(n14028), .ZN(n13959) );
  MUX2_X1 U15924 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14061), .S(n15390), .Z(
        P2_U3526) );
  AOI21_X1 U15925 ( .B1(n15377), .B2(n13962), .A(n13961), .ZN(n13963) );
  OAI211_X1 U15926 ( .C1(n15381), .C2(n13965), .A(n13964), .B(n13963), .ZN(
        n14062) );
  MUX2_X1 U15927 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14062), .S(n15390), .Z(
        P2_U3525) );
  AOI21_X1 U15928 ( .B1(n15377), .B2(n13967), .A(n13966), .ZN(n13968) );
  OAI211_X1 U15929 ( .C1(n15381), .C2(n13970), .A(n13969), .B(n13968), .ZN(
        n14063) );
  MUX2_X1 U15930 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14063), .S(n15390), .Z(
        P2_U3524) );
  AOI21_X1 U15931 ( .B1(n15377), .B2(n13972), .A(n13971), .ZN(n13973) );
  OAI211_X1 U15932 ( .C1(n15381), .C2(n13975), .A(n13974), .B(n13973), .ZN(
        n14064) );
  MUX2_X1 U15933 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14064), .S(n15390), .Z(
        P2_U3523) );
  AOI211_X1 U15934 ( .C1(n15377), .C2(n13978), .A(n13977), .B(n13976), .ZN(
        n13979) );
  OAI21_X1 U15935 ( .B1(n15381), .B2(n13980), .A(n13979), .ZN(n14065) );
  MUX2_X1 U15936 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14065), .S(n15390), .Z(
        P2_U3522) );
  AOI21_X1 U15937 ( .B1(n15377), .B2(n13982), .A(n13981), .ZN(n13983) );
  OAI211_X1 U15938 ( .C1(n15381), .C2(n13985), .A(n13984), .B(n13983), .ZN(
        n14066) );
  MUX2_X1 U15939 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14066), .S(n15390), .Z(
        P2_U3521) );
  AOI211_X1 U15940 ( .C1(n15377), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n13989) );
  OAI21_X1 U15941 ( .B1(n15381), .B2(n13990), .A(n13989), .ZN(n14067) );
  MUX2_X1 U15942 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14067), .S(n15390), .Z(
        P2_U3520) );
  AOI211_X1 U15943 ( .C1(n15377), .C2(n13993), .A(n13992), .B(n13991), .ZN(
        n13994) );
  OAI21_X1 U15944 ( .B1(n15381), .B2(n13995), .A(n13994), .ZN(n14068) );
  MUX2_X1 U15945 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14068), .S(n15390), .Z(
        P2_U3519) );
  AOI21_X1 U15946 ( .B1(n15377), .B2(n13997), .A(n13996), .ZN(n13998) );
  OAI211_X1 U15947 ( .C1(n15371), .C2(n14000), .A(n13999), .B(n13998), .ZN(
        n14069) );
  MUX2_X1 U15948 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14069), .S(n15390), .Z(
        P2_U3518) );
  NOR2_X1 U15949 ( .A1(n14001), .A2(n15381), .ZN(n14002) );
  AOI211_X1 U15950 ( .C1(n15377), .C2(n14004), .A(n14003), .B(n14002), .ZN(
        n14005) );
  NAND2_X1 U15951 ( .A1(n14006), .A2(n14005), .ZN(n14070) );
  MUX2_X1 U15952 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14070), .S(n15390), .Z(
        P2_U3517) );
  AOI21_X1 U15953 ( .B1(n15377), .B2(n14008), .A(n14007), .ZN(n14009) );
  OAI211_X1 U15954 ( .C1(n15381), .C2(n14011), .A(n14010), .B(n14009), .ZN(
        n14071) );
  MUX2_X1 U15955 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14071), .S(n15390), .Z(
        P2_U3516) );
  AOI21_X1 U15956 ( .B1(n15377), .B2(n14013), .A(n14012), .ZN(n14014) );
  OAI211_X1 U15957 ( .C1(n15381), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        n14072) );
  MUX2_X1 U15958 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14072), .S(n15390), .Z(
        P2_U3515) );
  AOI211_X1 U15959 ( .C1(n15377), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        n14020) );
  OAI21_X1 U15960 ( .B1(n15381), .B2(n14021), .A(n14020), .ZN(n14073) );
  MUX2_X1 U15961 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14073), .S(n15390), .Z(
        P2_U3514) );
  OAI211_X1 U15962 ( .C1(n14025), .C2(n14024), .A(n14023), .B(n14022), .ZN(
        n14026) );
  AOI21_X1 U15963 ( .B1(n14028), .B2(n14027), .A(n14026), .ZN(n14075) );
  NAND2_X1 U15964 ( .A1(n15387), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n14029) );
  OAI21_X1 U15965 ( .B1(n14075), .B2(n15387), .A(n14029), .ZN(P2_U3513) );
  AOI21_X1 U15966 ( .B1(n15377), .B2(n14031), .A(n14030), .ZN(n14032) );
  OAI211_X1 U15967 ( .C1(n15381), .C2(n14034), .A(n14033), .B(n14032), .ZN(
        n14076) );
  MUX2_X1 U15968 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14076), .S(n15390), .Z(
        P2_U3512) );
  AOI21_X1 U15969 ( .B1(n15377), .B2(n14036), .A(n14035), .ZN(n14037) );
  OAI211_X1 U15970 ( .C1(n15381), .C2(n14039), .A(n14038), .B(n14037), .ZN(
        n14077) );
  MUX2_X1 U15971 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14077), .S(n15390), .Z(
        P2_U3511) );
  AOI21_X1 U15972 ( .B1(n15377), .B2(n14041), .A(n14040), .ZN(n14042) );
  OAI211_X1 U15973 ( .C1(n15381), .C2(n14044), .A(n14043), .B(n14042), .ZN(
        n14078) );
  MUX2_X1 U15974 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14078), .S(n15390), .Z(
        P2_U3510) );
  AOI21_X1 U15975 ( .B1(n15377), .B2(n14046), .A(n14045), .ZN(n14047) );
  OAI211_X1 U15976 ( .C1(n15381), .C2(n14049), .A(n14048), .B(n14047), .ZN(
        n14079) );
  MUX2_X1 U15977 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14079), .S(n15390), .Z(
        P2_U3509) );
  AOI21_X1 U15978 ( .B1(n15377), .B2(n14051), .A(n14050), .ZN(n14052) );
  OAI211_X1 U15979 ( .C1(n15381), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14080) );
  MUX2_X1 U15980 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14080), .S(n15390), .Z(
        P2_U3508) );
  OAI211_X1 U15981 ( .C1(n14057), .C2(n15371), .A(n14056), .B(n14055), .ZN(
        n14081) );
  MUX2_X1 U15982 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14081), .S(n15390), .Z(
        P2_U3499) );
  MUX2_X1 U15983 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14058), .S(n15384), .Z(
        P2_U3498) );
  MUX2_X1 U15984 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14059), .S(n15384), .Z(
        P2_U3497) );
  MUX2_X1 U15985 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14060), .S(n15384), .Z(
        P2_U3495) );
  MUX2_X1 U15986 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14062), .S(n15384), .Z(
        P2_U3493) );
  MUX2_X1 U15987 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14063), .S(n15384), .Z(
        P2_U3492) );
  MUX2_X1 U15988 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14064), .S(n15384), .Z(
        P2_U3491) );
  MUX2_X1 U15989 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14065), .S(n15384), .Z(
        P2_U3490) );
  MUX2_X1 U15990 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14066), .S(n15384), .Z(
        P2_U3489) );
  MUX2_X1 U15991 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14067), .S(n15384), .Z(
        P2_U3488) );
  MUX2_X1 U15992 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14068), .S(n15384), .Z(
        P2_U3487) );
  MUX2_X1 U15993 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14069), .S(n15384), .Z(
        P2_U3486) );
  MUX2_X1 U15994 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14070), .S(n15384), .Z(
        P2_U3484) );
  MUX2_X1 U15995 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14071), .S(n15384), .Z(
        P2_U3481) );
  MUX2_X1 U15996 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14072), .S(n15384), .Z(
        P2_U3478) );
  MUX2_X1 U15997 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14073), .S(n15384), .Z(
        P2_U3475) );
  NAND2_X1 U15998 ( .A1(n6771), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n14074) );
  OAI21_X1 U15999 ( .B1(n14075), .B2(n6771), .A(n14074), .ZN(P2_U3472) );
  MUX2_X1 U16000 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14076), .S(n15384), .Z(
        P2_U3469) );
  MUX2_X1 U16001 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14077), .S(n15384), .Z(
        P2_U3466) );
  MUX2_X1 U16002 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14078), .S(n15384), .Z(
        P2_U3463) );
  MUX2_X1 U16003 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14079), .S(n15384), .Z(
        P2_U3460) );
  MUX2_X1 U16004 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14080), .S(n15384), .Z(
        P2_U3457) );
  MUX2_X1 U16005 ( .A(P2_REG0_REG_0__SCAN_IN), .B(n14081), .S(n15384), .Z(
        P2_U3430) );
  NAND3_X1 U16006 ( .A1(n14082), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14084) );
  OAI22_X1 U16007 ( .A1(n14085), .A2(n14084), .B1(n14083), .B2(n14097), .ZN(
        n14086) );
  AOI21_X1 U16008 ( .B1(n14087), .B2(n14093), .A(n14086), .ZN(n14088) );
  INV_X1 U16009 ( .A(n14088), .ZN(P2_U3296) );
  OAI222_X1 U16010 ( .A1(n14092), .A2(n14091), .B1(n14097), .B2(n14090), .C1(
        P2_U3088), .C2(n14089), .ZN(P2_U3298) );
  NAND2_X1 U16011 ( .A1(n14094), .A2(n14093), .ZN(n14096) );
  OAI211_X1 U16012 ( .C1(n14098), .C2(n14097), .A(n14096), .B(n14095), .ZN(
        P2_U3299) );
  MUX2_X1 U16013 ( .A(n14099), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16014 ( .A(n14101), .B(n14100), .ZN(n14106) );
  AOI22_X1 U16015 ( .A1(n14480), .A2(n14239), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14103) );
  NAND2_X1 U16016 ( .A1(n14478), .A2(n14218), .ZN(n14102) );
  OAI211_X1 U16017 ( .C1(n14684), .C2(n15182), .A(n14103), .B(n14102), .ZN(
        n14104) );
  AOI21_X1 U16018 ( .B1(n14983), .B2(n14221), .A(n14104), .ZN(n14105) );
  OAI21_X1 U16019 ( .B1(n14106), .B2(n15174), .A(n14105), .ZN(P1_U3214) );
  INV_X1 U16020 ( .A(n14107), .ZN(n14108) );
  AOI21_X1 U16021 ( .B1(n14110), .B2(n14109), .A(n14108), .ZN(n14116) );
  INV_X1 U16022 ( .A(n14231), .ZN(n15171) );
  INV_X1 U16023 ( .A(n14901), .ZN(n14902) );
  NOR2_X1 U16024 ( .A1(n14902), .A2(n15259), .ZN(n15057) );
  NOR2_X1 U16025 ( .A1(n14934), .A2(n14935), .ZN(n15056) );
  NOR2_X1 U16026 ( .A1(n14236), .A2(n14862), .ZN(n14111) );
  AOI211_X1 U16027 ( .C1(n15179), .C2(n15056), .A(n14112), .B(n14111), .ZN(
        n14113) );
  OAI21_X1 U16028 ( .B1(n14903), .B2(n15182), .A(n14113), .ZN(n14114) );
  AOI21_X1 U16029 ( .B1(n15171), .B2(n15057), .A(n14114), .ZN(n14115) );
  OAI21_X1 U16030 ( .B1(n14116), .B2(n15174), .A(n14115), .ZN(P1_U3215) );
  XOR2_X1 U16031 ( .A(n14166), .B(n14117), .Z(n14121) );
  OAI22_X1 U16032 ( .A1(n14387), .A2(n14933), .B1(n14784), .B2(n14935), .ZN(
        n14754) );
  AOI22_X1 U16033 ( .A1(n14754), .A2(n15179), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14118) );
  OAI21_X1 U16034 ( .B1(n14757), .B2(n15182), .A(n14118), .ZN(n14119) );
  AOI21_X1 U16035 ( .B1(n15005), .B2(n14221), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16036 ( .B1(n14121), .B2(n15174), .A(n14120), .ZN(P1_U3216) );
  INV_X1 U16037 ( .A(n15028), .ZN(n14814) );
  OR2_X1 U16038 ( .A1(n12240), .A2(n14122), .ZN(n14214) );
  NAND2_X1 U16039 ( .A1(n14214), .A2(n14215), .ZN(n14124) );
  NAND2_X1 U16040 ( .A1(n14124), .A2(n14123), .ZN(n14126) );
  AOI21_X1 U16041 ( .B1(n14126), .B2(n14125), .A(n15174), .ZN(n14128) );
  NAND2_X1 U16042 ( .A1(n14128), .A2(n14127), .ZN(n14134) );
  INV_X1 U16043 ( .A(n14129), .ZN(n14812) );
  AND2_X1 U16044 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14639) );
  AOI21_X1 U16045 ( .B1(n14218), .B2(n14816), .A(n14639), .ZN(n14130) );
  OAI21_X1 U16046 ( .B1(n14216), .B2(n14131), .A(n14130), .ZN(n14132) );
  AOI21_X1 U16047 ( .B1(n14812), .B2(n14211), .A(n14132), .ZN(n14133) );
  OAI211_X1 U16048 ( .C1(n14814), .C2(n14242), .A(n14134), .B(n14133), .ZN(
        P1_U3219) );
  AOI21_X1 U16049 ( .B1(n14136), .B2(n14135), .A(n6506), .ZN(n14141) );
  AOI22_X1 U16050 ( .A1(n14483), .A2(n14218), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14138) );
  NAND2_X1 U16051 ( .A1(n14211), .A2(n14787), .ZN(n14137) );
  OAI211_X1 U16052 ( .C1(n14783), .C2(n14216), .A(n14138), .B(n14137), .ZN(
        n14139) );
  AOI21_X1 U16053 ( .B1(n15017), .B2(n14221), .A(n14139), .ZN(n14140) );
  OAI21_X1 U16054 ( .B1(n14141), .B2(n15174), .A(n14140), .ZN(P1_U3223) );
  INV_X1 U16055 ( .A(n14951), .ZN(n15071) );
  AOI21_X1 U16056 ( .B1(n14143), .B2(n14142), .A(n15174), .ZN(n14145) );
  NAND2_X1 U16057 ( .A1(n14145), .A2(n14144), .ZN(n14150) );
  NOR2_X1 U16058 ( .A1(n15182), .A2(n14949), .ZN(n14148) );
  OAI21_X1 U16059 ( .B1(n14236), .B2(n14934), .A(n14146), .ZN(n14147) );
  AOI211_X1 U16060 ( .C1(n14239), .C2(n14489), .A(n14148), .B(n14147), .ZN(
        n14149) );
  OAI211_X1 U16061 ( .C1(n15071), .C2(n14242), .A(n14150), .B(n14149), .ZN(
        P1_U3224) );
  OAI22_X1 U16062 ( .A1(n14679), .A2(n14933), .B1(n14387), .B2(n14935), .ZN(
        n14994) );
  OAI22_X1 U16063 ( .A1(n14722), .A2(n15182), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14153), .ZN(n14154) );
  AOI21_X1 U16064 ( .B1(n14994), .B2(n15179), .A(n14154), .ZN(n14156) );
  NAND2_X1 U16065 ( .A1(n14995), .A2(n14221), .ZN(n14155) );
  AOI21_X1 U16066 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n14165) );
  NOR2_X1 U16067 ( .A1(n15182), .A2(n14865), .ZN(n14163) );
  NAND2_X1 U16068 ( .A1(n14218), .A2(n14486), .ZN(n14161) );
  OAI211_X1 U16069 ( .C1(n14216), .C2(n14862), .A(n14161), .B(n14160), .ZN(
        n14162) );
  AOI211_X1 U16070 ( .C1(n15046), .C2(n14221), .A(n14163), .B(n14162), .ZN(
        n14164) );
  OAI21_X1 U16071 ( .B1(n14165), .B2(n15174), .A(n14164), .ZN(P1_U3226) );
  NAND2_X1 U16072 ( .A1(n14117), .A2(n14166), .ZN(n14168) );
  NAND2_X1 U16073 ( .A1(n14168), .A2(n14167), .ZN(n14169) );
  XOR2_X1 U16074 ( .A(n14170), .B(n14169), .Z(n14176) );
  NOR2_X1 U16075 ( .A1(n14171), .A2(n14935), .ZN(n14172) );
  AOI21_X1 U16076 ( .B1(n14481), .B2(n14897), .A(n14172), .ZN(n14737) );
  AOI22_X1 U16077 ( .A1(n14211), .A2(n14743), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14173) );
  OAI21_X1 U16078 ( .B1(n14737), .B2(n14198), .A(n14173), .ZN(n14174) );
  AOI21_X1 U16079 ( .B1(n14739), .B2(n14221), .A(n14174), .ZN(n14175) );
  OAI21_X1 U16080 ( .B1(n14176), .B2(n15174), .A(n14175), .ZN(P1_U3229) );
  INV_X1 U16081 ( .A(n15022), .ZN(n14186) );
  OAI211_X1 U16082 ( .C1(n14177), .C2(n14179), .A(n14178), .B(n14232), .ZN(
        n14185) );
  NAND2_X1 U16083 ( .A1(n14485), .A2(n14880), .ZN(n14181) );
  NAND2_X1 U16084 ( .A1(n14484), .A2(n14897), .ZN(n14180) );
  NAND2_X1 U16085 ( .A1(n14181), .A2(n14180), .ZN(n15021) );
  INV_X1 U16086 ( .A(n15021), .ZN(n14806) );
  OAI22_X1 U16087 ( .A1(n14806), .A2(n14198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14182), .ZN(n14183) );
  AOI21_X1 U16088 ( .B1(n14796), .B2(n14211), .A(n14183), .ZN(n14184) );
  OAI211_X1 U16089 ( .C1(n14186), .C2(n14242), .A(n14185), .B(n14184), .ZN(
        P1_U3233) );
  INV_X1 U16090 ( .A(n15065), .ZN(n14922) );
  OAI211_X1 U16091 ( .C1(n14189), .C2(n14188), .A(n14187), .B(n14232), .ZN(
        n14192) );
  OAI22_X1 U16092 ( .A1(n14301), .A2(n14935), .B1(n14333), .B2(n14933), .ZN(
        n15064) );
  AND2_X1 U16093 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14585) );
  NOR2_X1 U16094 ( .A1(n15182), .A2(n14923), .ZN(n14190) );
  AOI211_X1 U16095 ( .C1(n15179), .C2(n15064), .A(n14585), .B(n14190), .ZN(
        n14191) );
  OAI211_X1 U16096 ( .C1(n14922), .C2(n14242), .A(n14192), .B(n14191), .ZN(
        P1_U3234) );
  OAI21_X1 U16097 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n14196) );
  NAND2_X1 U16098 ( .A1(n14196), .A2(n14232), .ZN(n14201) );
  INV_X1 U16099 ( .A(n14197), .ZN(n14772) );
  AOI22_X1 U16100 ( .A1(n14482), .A2(n14897), .B1(n14880), .B2(n14484), .ZN(
        n15009) );
  NAND2_X1 U16101 ( .A1(P1_U3086), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n15454)
         );
  OAI21_X1 U16102 ( .B1(n15009), .B2(n14198), .A(n15454), .ZN(n14199) );
  AOI21_X1 U16103 ( .B1(n14772), .B2(n14211), .A(n14199), .ZN(n14200) );
  OAI211_X1 U16104 ( .C1(n14242), .C2(n9615), .A(n14201), .B(n14200), .ZN(
        P1_U3235) );
  INV_X1 U16105 ( .A(n14202), .ZN(n14203) );
  AOI21_X1 U16106 ( .B1(n14205), .B2(n14204), .A(n14203), .ZN(n14213) );
  AOI21_X1 U16107 ( .B1(n14218), .B2(n14488), .A(n14206), .ZN(n14207) );
  OAI21_X1 U16108 ( .B1(n14216), .B2(n14306), .A(n14207), .ZN(n14209) );
  NAND2_X1 U16109 ( .A1(n14303), .A2(n15255), .ZN(n15075) );
  NOR2_X1 U16110 ( .A1(n15075), .A2(n14231), .ZN(n14208) );
  AOI211_X1 U16111 ( .C1(n14211), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        n14212) );
  OAI21_X1 U16112 ( .B1(n14213), .B2(n15174), .A(n14212), .ZN(P1_U3236) );
  XOR2_X1 U16113 ( .A(n14215), .B(n14214), .Z(n14223) );
  NAND2_X1 U16114 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14617)
         );
  OAI21_X1 U16115 ( .B1(n14216), .B2(n14861), .A(n14617), .ZN(n14217) );
  AOI21_X1 U16116 ( .B1(n14218), .B2(n14485), .A(n14217), .ZN(n14219) );
  OAI21_X1 U16117 ( .B1(n14833), .B2(n15182), .A(n14219), .ZN(n14220) );
  AOI21_X1 U16118 ( .B1(n15034), .B2(n14221), .A(n14220), .ZN(n14222) );
  OAI21_X1 U16119 ( .B1(n14223), .B2(n15174), .A(n14222), .ZN(P1_U3238) );
  NAND2_X1 U16120 ( .A1(n14395), .A2(n15255), .ZN(n14988) );
  OAI22_X1 U16121 ( .A1(n14226), .A2(n14933), .B1(n14225), .B2(n14935), .ZN(
        n14705) );
  INV_X1 U16122 ( .A(n14698), .ZN(n14228) );
  OAI22_X1 U16123 ( .A1(n14228), .A2(n15182), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14227), .ZN(n14229) );
  AOI21_X1 U16124 ( .B1(n14705), .B2(n15179), .A(n14229), .ZN(n14230) );
  OAI211_X1 U16125 ( .C1(n14235), .C2(n14234), .A(n14233), .B(n14232), .ZN(
        n14241) );
  NOR2_X1 U16126 ( .A1(n15182), .A2(n14884), .ZN(n14238) );
  OAI22_X1 U16127 ( .A1(n14236), .A2(n14345), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6904), .ZN(n14237) );
  AOI211_X1 U16128 ( .C1(n14239), .C2(n14879), .A(n14238), .B(n14237), .ZN(
        n14240) );
  OAI211_X1 U16129 ( .C1(n14888), .C2(n14242), .A(n14241), .B(n14240), .ZN(
        P1_U3241) );
  NOR3_X1 U16130 ( .A1(n14243), .A2(n14935), .A3(n15106), .ZN(n14474) );
  OAI21_X1 U16131 ( .B1(n14244), .B2(n14245), .A(P1_B_REG_SCAN_IN), .ZN(n14473) );
  NAND2_X1 U16132 ( .A1(n14247), .A2(n14415), .ZN(n14249) );
  INV_X1 U16133 ( .A(n14415), .ZN(n14250) );
  NAND2_X1 U16134 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  NAND2_X2 U16135 ( .A1(n14411), .A2(n14252), .ZN(n14253) );
  INV_X4 U16136 ( .A(n14253), .ZN(n14414) );
  MUX2_X1 U16137 ( .A(n14680), .B(n14254), .S(n14414), .Z(n14407) );
  INV_X1 U16138 ( .A(n14407), .ZN(n14410) );
  NAND2_X1 U16139 ( .A1(n14438), .A2(n10741), .ZN(n14256) );
  NAND2_X1 U16140 ( .A1(n14414), .A2(n14258), .ZN(n14259) );
  INV_X1 U16141 ( .A(n14498), .ZN(n14261) );
  OR2_X1 U16142 ( .A1(n14265), .A2(n14414), .ZN(n14266) );
  AND2_X1 U16143 ( .A1(n14267), .A2(n14266), .ZN(n14271) );
  OAI21_X1 U16144 ( .B1(n14274), .B2(n14271), .A(n14270), .ZN(n14276) );
  NAND2_X1 U16145 ( .A1(n14276), .A2(n14275), .ZN(n14280) );
  MUX2_X1 U16146 ( .A(n14278), .B(n14277), .S(n14253), .Z(n14279) );
  NAND2_X1 U16147 ( .A1(n14280), .A2(n14279), .ZN(n14282) );
  MUX2_X1 U16148 ( .A(n14496), .B(n15222), .S(n14253), .Z(n14283) );
  MUX2_X1 U16149 ( .A(n15222), .B(n14496), .S(n14253), .Z(n14281) );
  INV_X1 U16150 ( .A(n14283), .ZN(n14284) );
  MUX2_X1 U16151 ( .A(n15245), .B(n14495), .S(n14427), .Z(n14286) );
  MUX2_X1 U16152 ( .A(n14495), .B(n15245), .S(n14427), .Z(n14285) );
  MUX2_X1 U16153 ( .A(n14494), .B(n15254), .S(n14427), .Z(n14288) );
  MUX2_X1 U16154 ( .A(n15254), .B(n14494), .S(n14427), .Z(n14287) );
  MUX2_X1 U16155 ( .A(n14289), .B(n14493), .S(n14427), .Z(n14292) );
  MUX2_X1 U16156 ( .A(n14493), .B(n14289), .S(n14427), .Z(n14290) );
  MUX2_X1 U16157 ( .A(n14492), .B(n14956), .S(n14427), .Z(n14294) );
  MUX2_X1 U16158 ( .A(n14956), .B(n14492), .S(n14427), .Z(n14293) );
  MUX2_X1 U16159 ( .A(n14491), .B(n14295), .S(n14414), .Z(n14298) );
  MUX2_X1 U16160 ( .A(n14491), .B(n14295), .S(n14427), .Z(n14296) );
  AOI21_X1 U16161 ( .B1(n14299), .B2(n14298), .A(n14297), .ZN(n14311) );
  NOR2_X1 U16162 ( .A1(n14299), .A2(n14298), .ZN(n14310) );
  MUX2_X1 U16163 ( .A(n14487), .B(n15065), .S(n14414), .Z(n14332) );
  NAND2_X1 U16164 ( .A1(n15065), .A2(n14427), .ZN(n14329) );
  NAND2_X1 U16165 ( .A1(n14414), .A2(n14487), .ZN(n14334) );
  NAND3_X1 U16166 ( .A1(n14332), .A2(n14329), .A3(n14334), .ZN(n14300) );
  OAI211_X1 U16167 ( .C1(n14902), .C2(n14879), .A(n14343), .B(n14300), .ZN(
        n14326) );
  MUX2_X1 U16168 ( .A(n14301), .B(n15071), .S(n14414), .Z(n14323) );
  MUX2_X1 U16169 ( .A(n14488), .B(n14951), .S(n14427), .Z(n14322) );
  MUX2_X1 U16170 ( .A(n14936), .B(n14302), .S(n14414), .Z(n14317) );
  MUX2_X1 U16171 ( .A(n14489), .B(n14303), .S(n14427), .Z(n14316) );
  OAI22_X1 U16172 ( .A1(n14323), .A2(n14322), .B1(n14317), .B2(n14316), .ZN(
        n14304) );
  OR2_X1 U16173 ( .A1(n14326), .A2(n14304), .ZN(n14319) );
  INV_X1 U16174 ( .A(n14319), .ZN(n14308) );
  MUX2_X1 U16175 ( .A(n14306), .B(n14305), .S(n14427), .Z(n14313) );
  MUX2_X1 U16176 ( .A(n14490), .B(n15079), .S(n14414), .Z(n14312) );
  NAND2_X1 U16177 ( .A1(n14313), .A2(n14312), .ZN(n14307) );
  INV_X1 U16178 ( .A(n14312), .ZN(n14315) );
  INV_X1 U16179 ( .A(n14313), .ZN(n14314) );
  AOI22_X1 U16180 ( .A1(n14317), .A2(n14316), .B1(n14315), .B2(n14314), .ZN(
        n14318) );
  NOR2_X1 U16181 ( .A1(n14319), .A2(n14318), .ZN(n14331) );
  NAND3_X1 U16182 ( .A1(n14901), .A2(n14333), .A3(n14427), .ZN(n14320) );
  OAI211_X1 U16183 ( .C1(n14343), .C2(n14414), .A(n14320), .B(n14342), .ZN(
        n14321) );
  INV_X1 U16184 ( .A(n14321), .ZN(n14328) );
  INV_X1 U16185 ( .A(n14322), .ZN(n14325) );
  INV_X1 U16186 ( .A(n14323), .ZN(n14324) );
  OR3_X1 U16187 ( .A1(n14326), .A2(n14325), .A3(n14324), .ZN(n14327) );
  OAI211_X1 U16188 ( .C1(n14329), .C2(n14332), .A(n14328), .B(n14327), .ZN(
        n14330) );
  OAI21_X1 U16189 ( .B1(n14332), .B2(n14334), .A(n14333), .ZN(n14337) );
  INV_X1 U16190 ( .A(n14332), .ZN(n14336) );
  NOR2_X1 U16191 ( .A1(n14334), .A2(n14333), .ZN(n14335) );
  AOI22_X1 U16192 ( .A1(n14337), .A2(n14902), .B1(n14336), .B2(n14335), .ZN(
        n14339) );
  INV_X1 U16193 ( .A(n14343), .ZN(n14338) );
  NAND2_X1 U16194 ( .A1(n14342), .A2(n14341), .ZN(n14344) );
  NAND3_X1 U16195 ( .A1(n14344), .A2(n14427), .A3(n14343), .ZN(n14350) );
  MUX2_X1 U16196 ( .A(n14881), .B(n15046), .S(n14414), .Z(n14360) );
  NAND2_X1 U16197 ( .A1(n14360), .A2(n14486), .ZN(n14346) );
  NAND2_X1 U16198 ( .A1(n14414), .A2(n14345), .ZN(n14355) );
  AOI21_X1 U16199 ( .B1(n14346), .B2(n14355), .A(n7717), .ZN(n14349) );
  NAND2_X1 U16200 ( .A1(n14360), .A2(n14861), .ZN(n14347) );
  OR2_X1 U16201 ( .A1(n15046), .A2(n14414), .ZN(n14351) );
  AOI21_X1 U16202 ( .B1(n14347), .B2(n14351), .A(n14844), .ZN(n14348) );
  OR2_X1 U16203 ( .A1(n14414), .A2(n14861), .ZN(n14352) );
  OAI22_X1 U16204 ( .A1(n15046), .A2(n14352), .B1(n14486), .B2(n14355), .ZN(
        n14359) );
  INV_X1 U16205 ( .A(n14351), .ZN(n14354) );
  INV_X1 U16206 ( .A(n14352), .ZN(n14353) );
  AOI21_X1 U16207 ( .B1(n14360), .B2(n14354), .A(n14353), .ZN(n14363) );
  INV_X1 U16208 ( .A(n14355), .ZN(n14356) );
  NAND2_X1 U16209 ( .A1(n14360), .A2(n14356), .ZN(n14357) );
  OAI21_X1 U16210 ( .B1(n14427), .B2(n14486), .A(n14357), .ZN(n14358) );
  NAND2_X1 U16211 ( .A1(n14358), .A2(n14844), .ZN(n14362) );
  NAND2_X1 U16212 ( .A1(n14360), .A2(n14359), .ZN(n14361) );
  OAI211_X1 U16213 ( .C1(n14363), .C2(n14844), .A(n14362), .B(n14361), .ZN(
        n14365) );
  XNOR2_X1 U16214 ( .A(n15034), .B(n14414), .ZN(n14367) );
  XNOR2_X1 U16215 ( .A(n14818), .B(n14427), .ZN(n14366) );
  MUX2_X1 U16216 ( .A(n14816), .B(n15022), .S(n14427), .Z(n14372) );
  NOR2_X1 U16217 ( .A1(n15022), .A2(n14816), .ZN(n14370) );
  OAI21_X1 U16218 ( .B1(n14372), .B2(n14370), .A(n14369), .ZN(n14374) );
  NAND2_X1 U16219 ( .A1(n14372), .A2(n14371), .ZN(n14373) );
  AND2_X1 U16220 ( .A1(n14484), .A2(n14427), .ZN(n14376) );
  OAI21_X1 U16221 ( .B1(n14484), .B2(n14427), .A(n15017), .ZN(n14375) );
  OAI21_X1 U16222 ( .B1(n14376), .B2(n15017), .A(n14375), .ZN(n14377) );
  AND2_X1 U16223 ( .A1(n14784), .A2(n14427), .ZN(n14379) );
  OAI21_X1 U16224 ( .B1(n14784), .B2(n14427), .A(n9615), .ZN(n14378) );
  OAI21_X1 U16225 ( .B1(n14379), .B2(n9615), .A(n14378), .ZN(n14380) );
  MUX2_X1 U16226 ( .A(n14482), .B(n15005), .S(n14427), .Z(n14384) );
  MUX2_X1 U16227 ( .A(n14482), .B(n15005), .S(n14414), .Z(n14381) );
  INV_X1 U16228 ( .A(n14383), .ZN(n14386) );
  INV_X1 U16229 ( .A(n14384), .ZN(n14385) );
  MUX2_X1 U16230 ( .A(n14712), .B(n14739), .S(n14414), .Z(n14389) );
  MUX2_X1 U16231 ( .A(n14387), .B(n15000), .S(n14427), .Z(n14388) );
  AOI21_X1 U16232 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n14391) );
  MUX2_X1 U16233 ( .A(n14481), .B(n14995), .S(n14427), .Z(n14393) );
  MUX2_X1 U16234 ( .A(n14481), .B(n14995), .S(n14414), .Z(n14392) );
  INV_X1 U16235 ( .A(n14393), .ZN(n14394) );
  MUX2_X1 U16236 ( .A(n14480), .B(n14395), .S(n14414), .Z(n14399) );
  MUX2_X1 U16237 ( .A(n14480), .B(n14395), .S(n14427), .Z(n14396) );
  NAND2_X1 U16238 ( .A1(n14397), .A2(n14396), .ZN(n14403) );
  INV_X1 U16239 ( .A(n14398), .ZN(n14401) );
  INV_X1 U16240 ( .A(n14399), .ZN(n14400) );
  NAND2_X1 U16241 ( .A1(n14401), .A2(n14400), .ZN(n14402) );
  MUX2_X1 U16242 ( .A(n14479), .B(n14983), .S(n14427), .Z(n14405) );
  MUX2_X1 U16243 ( .A(n14479), .B(n14983), .S(n14414), .Z(n14404) );
  INV_X1 U16244 ( .A(n14405), .ZN(n14406) );
  MUX2_X1 U16245 ( .A(n14478), .B(n14408), .S(n14427), .Z(n14409) );
  MUX2_X1 U16246 ( .A(n14477), .B(n14668), .S(n14427), .Z(n14423) );
  INV_X1 U16247 ( .A(n14411), .ZN(n14412) );
  OAI21_X1 U16248 ( .B1(n14475), .B2(n14412), .A(n14476), .ZN(n14413) );
  MUX2_X1 U16249 ( .A(n14413), .B(n14981), .S(n14414), .Z(n14425) );
  NAND2_X1 U16250 ( .A1(n14648), .A2(n14427), .ZN(n14419) );
  NAND2_X1 U16251 ( .A1(n14414), .A2(n14475), .ZN(n14428) );
  OAI21_X1 U16252 ( .B1(n14416), .B2(n14415), .A(n14428), .ZN(n14417) );
  NAND2_X1 U16253 ( .A1(n14417), .A2(n14476), .ZN(n14418) );
  NAND2_X1 U16254 ( .A1(n14419), .A2(n14418), .ZN(n14424) );
  MUX2_X1 U16255 ( .A(n14421), .B(n14420), .S(n14427), .Z(n14422) );
  INV_X1 U16256 ( .A(n14475), .ZN(n14426) );
  MUX2_X1 U16257 ( .A(n14427), .B(n14426), .S(n14643), .Z(n14430) );
  INV_X1 U16258 ( .A(n14428), .ZN(n14429) );
  NOR2_X1 U16259 ( .A1(n14430), .A2(n14429), .ZN(n14463) );
  INV_X1 U16260 ( .A(n14431), .ZN(n14433) );
  NAND2_X1 U16261 ( .A1(n14433), .A2(n14432), .ZN(n14435) );
  OR2_X1 U16262 ( .A1(n14248), .A2(n14917), .ZN(n14434) );
  NAND2_X1 U16263 ( .A1(n14435), .A2(n14434), .ZN(n14466) );
  NAND2_X1 U16264 ( .A1(n14466), .A2(n14468), .ZN(n14460) );
  NOR3_X1 U16265 ( .A1(n14459), .A2(n14463), .A3(n14460), .ZN(n14471) );
  INV_X1 U16266 ( .A(n14457), .ZN(n14462) );
  NAND4_X1 U16267 ( .A1(n14439), .A2(n14438), .A3(n14437), .A4(n14436), .ZN(
        n14441) );
  NOR4_X1 U16268 ( .A1(n15212), .A2(n14442), .A3(n14441), .A4(n14440), .ZN(
        n14445) );
  NAND3_X1 U16269 ( .A1(n14445), .A2(n9754), .A3(n14444), .ZN(n14446) );
  NOR4_X1 U16270 ( .A1(n14449), .A2(n14448), .A3(n14447), .A4(n14446), .ZN(
        n14451) );
  INV_X1 U16271 ( .A(n14856), .ZN(n14853) );
  NAND4_X1 U16272 ( .A1(n14895), .A2(n14451), .A3(n14853), .A4(n14450), .ZN(
        n14452) );
  INV_X1 U16273 ( .A(n14877), .ZN(n14874) );
  NOR4_X1 U16274 ( .A1(n14452), .A2(n14874), .A3(n14942), .A4(n14843), .ZN(
        n14453) );
  AND4_X1 U16275 ( .A1(n14804), .A2(n6411), .A3(n14453), .A4(n14824), .ZN(
        n14454) );
  NAND4_X1 U16276 ( .A1(n14752), .A2(n14768), .A3(n14454), .A4(n14780), .ZN(
        n14455) );
  XNOR2_X1 U16277 ( .A(n15000), .B(n14712), .ZN(n14732) );
  NOR4_X1 U16278 ( .A1(n14702), .A2(n14455), .A3(n14732), .A4(n14716), .ZN(
        n14456) );
  INV_X1 U16279 ( .A(n14466), .ZN(n14458) );
  INV_X1 U16280 ( .A(n14460), .ZN(n14461) );
  NAND2_X1 U16281 ( .A1(n14462), .A2(n14461), .ZN(n14465) );
  INV_X1 U16282 ( .A(n14463), .ZN(n14464) );
  MUX2_X1 U16283 ( .A(n14466), .B(n14465), .S(n14464), .Z(n14467) );
  OAI21_X1 U16284 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n14472) );
  OAI21_X1 U16285 ( .B1(n14474), .B2(n14473), .A(n14472), .ZN(P1_U3242) );
  MUX2_X1 U16286 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14475), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16287 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14476), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16288 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14477), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16289 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14478), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16290 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14479), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16291 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14480), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16292 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14481), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16293 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14712), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16294 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14482), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16295 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14483), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16296 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14484), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16297 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14816), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16298 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14485), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16299 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14818), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16300 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14486), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16301 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14881), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16302 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14896), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16303 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14879), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16304 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14487), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16305 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14488), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16306 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14489), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16307 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14490), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16308 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14491), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16309 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14492), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16310 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14493), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16311 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14494), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16312 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14495), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16313 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14496), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16314 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14497), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16315 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14265), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16316 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14498), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16317 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14499), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16318 ( .C1(n14501), .C2(n14500), .A(n15188), .B(n14517), .ZN(
        n14508) );
  OAI211_X1 U16319 ( .C1(n14510), .C2(n14502), .A(n15194), .B(n14524), .ZN(
        n14507) );
  AOI22_X1 U16320 ( .A1(n15199), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14506) );
  INV_X1 U16321 ( .A(n14503), .ZN(n14504) );
  NAND2_X1 U16322 ( .A1(n15197), .A2(n14504), .ZN(n14505) );
  NAND4_X1 U16323 ( .A1(n14508), .A2(n14507), .A3(n14506), .A4(n14505), .ZN(
        P1_U3244) );
  MUX2_X1 U16324 ( .A(n14510), .B(n14509), .S(n15106), .Z(n14512) );
  NAND2_X1 U16325 ( .A1(n14512), .A2(n14511), .ZN(n14514) );
  OAI211_X1 U16326 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14515), .A(n14514), .B(
        P1_U4016), .ZN(n15204) );
  AOI22_X1 U16327 ( .A1(n15199), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14529) );
  MUX2_X1 U16328 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10245), .S(n14522), .Z(
        n14518) );
  NAND3_X1 U16329 ( .A1(n14518), .A2(n14517), .A3(n14516), .ZN(n14519) );
  NAND2_X1 U16330 ( .A1(n14519), .A2(n14536), .ZN(n14520) );
  OAI22_X1 U16331 ( .A1(n14522), .A2(n14633), .B1(n14635), .B2(n14520), .ZN(
        n14521) );
  INV_X1 U16332 ( .A(n14521), .ZN(n14528) );
  MUX2_X1 U16333 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10262), .S(n14522), .Z(
        n14525) );
  NAND3_X1 U16334 ( .A1(n14525), .A2(n14524), .A3(n14523), .ZN(n14526) );
  NAND3_X1 U16335 ( .A1(n15194), .A2(n14541), .A3(n14526), .ZN(n14527) );
  NAND4_X1 U16336 ( .A1(n15204), .A2(n14529), .A3(n14528), .A4(n14527), .ZN(
        P1_U3245) );
  INV_X1 U16337 ( .A(n14538), .ZN(n14533) );
  OAI22_X1 U16338 ( .A1(n14583), .A2(n14531), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14530), .ZN(n14532) );
  AOI21_X1 U16339 ( .B1(n14533), .B2(n15197), .A(n14532), .ZN(n14545) );
  MUX2_X1 U16340 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10249), .S(n14538), .Z(
        n14535) );
  NAND3_X1 U16341 ( .A1(n14536), .A2(n14535), .A3(n14534), .ZN(n14537) );
  NAND3_X1 U16342 ( .A1(n15188), .A2(n15185), .A3(n14537), .ZN(n14544) );
  MUX2_X1 U16343 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10267), .S(n14538), .Z(
        n14540) );
  NAND3_X1 U16344 ( .A1(n14541), .A2(n14540), .A3(n14539), .ZN(n14542) );
  NAND3_X1 U16345 ( .A1(n15194), .A2(n15191), .A3(n14542), .ZN(n14543) );
  NAND3_X1 U16346 ( .A1(n14545), .A2(n14544), .A3(n14543), .ZN(P1_U3246) );
  OAI21_X1 U16347 ( .B1(n14583), .B2(n14547), .A(n14546), .ZN(n14548) );
  AOI21_X1 U16348 ( .B1(n14549), .B2(n15197), .A(n14548), .ZN(n14560) );
  OAI211_X1 U16349 ( .C1(n14552), .C2(n14551), .A(n15188), .B(n14550), .ZN(
        n14559) );
  NAND3_X1 U16350 ( .A1(n14555), .A2(n14554), .A3(n14553), .ZN(n14556) );
  NAND3_X1 U16351 ( .A1(n15194), .A2(n14557), .A3(n14556), .ZN(n14558) );
  NAND3_X1 U16352 ( .A1(n14560), .A2(n14559), .A3(n14558), .ZN(P1_U3249) );
  OAI21_X1 U16353 ( .B1(n14563), .B2(n14562), .A(n14561), .ZN(n14564) );
  NAND2_X1 U16354 ( .A1(n14564), .A2(n15188), .ZN(n14576) );
  OAI21_X1 U16355 ( .B1(n14583), .B2(n15548), .A(n14565), .ZN(n14566) );
  AOI21_X1 U16356 ( .B1(n14567), .B2(n15197), .A(n14566), .ZN(n14575) );
  MUX2_X1 U16357 ( .A(n11833), .B(P1_REG2_REG_9__SCAN_IN), .S(n14567), .Z(
        n14570) );
  INV_X1 U16358 ( .A(n14568), .ZN(n14569) );
  NAND2_X1 U16359 ( .A1(n14570), .A2(n14569), .ZN(n14572) );
  OAI211_X1 U16360 ( .C1(n14573), .C2(n14572), .A(n14571), .B(n15194), .ZN(
        n14574) );
  NAND3_X1 U16361 ( .A1(n14576), .A2(n14575), .A3(n14574), .ZN(P1_U3252) );
  INV_X1 U16362 ( .A(n14577), .ZN(n14582) );
  OAI21_X1 U16363 ( .B1(n14580), .B2(n14579), .A(n14578), .ZN(n14581) );
  NAND3_X1 U16364 ( .A1(n14582), .A2(n15188), .A3(n14581), .ZN(n14592) );
  INV_X1 U16365 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15116) );
  NOR2_X1 U16366 ( .A1(n14583), .A2(n15116), .ZN(n14584) );
  AOI211_X1 U16367 ( .C1(n15197), .C2(n14586), .A(n14585), .B(n14584), .ZN(
        n14591) );
  OAI211_X1 U16368 ( .C1(n14589), .C2(n14588), .A(n14587), .B(n15194), .ZN(
        n14590) );
  NAND3_X1 U16369 ( .A1(n14592), .A2(n14591), .A3(n14590), .ZN(P1_U3256) );
  AND2_X1 U16370 ( .A1(n14593), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14595) );
  MUX2_X1 U16371 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14609), .S(n14612), .Z(
        n14594) );
  OAI21_X1 U16372 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14608) );
  OR3_X1 U16373 ( .A1(n14596), .A2(n14595), .A3(n14594), .ZN(n14597) );
  NAND3_X1 U16374 ( .A1(n14608), .A2(n15194), .A3(n14597), .ZN(n14607) );
  INV_X1 U16375 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14598) );
  XNOR2_X1 U16376 ( .A(n14612), .B(n14598), .ZN(n14613) );
  XOR2_X1 U16377 ( .A(n14613), .B(n14614), .Z(n14602) );
  NAND2_X1 U16378 ( .A1(n15188), .A2(n14602), .ZN(n14603) );
  NAND2_X1 U16379 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  AOI21_X1 U16380 ( .B1(n15199), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14605), 
        .ZN(n14606) );
  OAI211_X1 U16381 ( .C1(n14633), .C2(n14610), .A(n14607), .B(n14606), .ZN(
        P1_U3260) );
  OAI21_X1 U16382 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14627) );
  XOR2_X1 U16383 ( .A(n14628), .B(n14627), .Z(n14611) );
  NAND2_X1 U16384 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14611), .ZN(n14630) );
  OAI211_X1 U16385 ( .C1(n14611), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15194), 
        .B(n14630), .ZN(n14620) );
  NAND2_X1 U16386 ( .A1(n14615), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14624) );
  OAI211_X1 U16387 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14615), .A(n15188), 
        .B(n14624), .ZN(n14616) );
  NAND2_X1 U16388 ( .A1(n14617), .A2(n14616), .ZN(n14618) );
  AOI21_X1 U16389 ( .B1(n15199), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14618), 
        .ZN(n14619) );
  OAI211_X1 U16390 ( .C1(n14633), .C2(n14621), .A(n14620), .B(n14619), .ZN(
        P1_U3261) );
  OR2_X1 U16391 ( .A1(n14622), .A2(n14621), .ZN(n14623) );
  NAND2_X1 U16392 ( .A1(n14624), .A2(n14623), .ZN(n14626) );
  NAND2_X1 U16393 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  NAND2_X1 U16394 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  XNOR2_X1 U16395 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14631), .ZN(n14638) );
  NAND2_X1 U16396 ( .A1(n14638), .A2(n15194), .ZN(n14632) );
  NAND2_X1 U16397 ( .A1(n14907), .A2(n15216), .ZN(n14966) );
  INV_X1 U16398 ( .A(n14966), .ZN(n14973) );
  NAND2_X1 U16399 ( .A1(n14640), .A2(n14973), .ZN(n14642) );
  NOR2_X1 U16400 ( .A1(n6412), .A2(n14979), .ZN(n14646) );
  AOI21_X1 U16401 ( .B1(n6412), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14646), .ZN(
        n14641) );
  OAI211_X1 U16402 ( .C1(n14643), .C2(n14921), .A(n14642), .B(n14641), .ZN(
        P1_U3263) );
  XNOR2_X1 U16403 ( .A(n9976), .B(n14981), .ZN(n14644) );
  NAND2_X1 U16404 ( .A1(n14644), .A2(n15216), .ZN(n14980) );
  NOR2_X1 U16405 ( .A1(n15220), .A2(n14645), .ZN(n14647) );
  AOI211_X1 U16406 ( .C1(n14648), .C2(n15223), .A(n14647), .B(n14646), .ZN(
        n14649) );
  OAI21_X1 U16407 ( .B1(n14980), .B2(n15225), .A(n14649), .ZN(P1_U3264) );
  NAND2_X1 U16408 ( .A1(n14651), .A2(n14650), .ZN(n14653) );
  XNOR2_X1 U16409 ( .A(n14653), .B(n14652), .ZN(n14674) );
  NAND2_X1 U16410 ( .A1(n14655), .A2(n14654), .ZN(n14657) );
  XNOR2_X1 U16411 ( .A(n14657), .B(n14656), .ZN(n14672) );
  INV_X1 U16412 ( .A(n14658), .ZN(n14661) );
  INV_X1 U16413 ( .A(n14659), .ZN(n14660) );
  AOI22_X1 U16414 ( .A1(n6412), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n14661), 
        .B2(n14660), .ZN(n14665) );
  OR3_X1 U16415 ( .A1(n14663), .A2(n14662), .A3(n15217), .ZN(n14664) );
  OAI211_X1 U16416 ( .C1(n14666), .C2(n6412), .A(n14665), .B(n14664), .ZN(
        n14667) );
  AOI21_X1 U16417 ( .B1(n14668), .B2(n15223), .A(n14667), .ZN(n14669) );
  OAI21_X1 U16418 ( .B1(n14670), .B2(n14966), .A(n14669), .ZN(n14671) );
  AOI21_X1 U16419 ( .B1(n14672), .B2(n14850), .A(n14671), .ZN(n14673) );
  OAI21_X1 U16420 ( .B1(n14674), .B2(n14910), .A(n14673), .ZN(P1_U3356) );
  INV_X1 U16421 ( .A(n14675), .ZN(n14678) );
  INV_X1 U16422 ( .A(n14676), .ZN(n14677) );
  OAI21_X1 U16423 ( .B1(n9679), .B2(n14678), .A(n14677), .ZN(n14682) );
  OAI22_X1 U16424 ( .A1(n14680), .A2(n14933), .B1(n14679), .B2(n14935), .ZN(
        n14681) );
  AOI21_X1 U16425 ( .B1(n14697), .B2(n14983), .A(n14929), .ZN(n14683) );
  INV_X1 U16426 ( .A(n14684), .ZN(n14685) );
  AOI22_X1 U16427 ( .A1(n14685), .A2(n14974), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n6412), .ZN(n14686) );
  OAI21_X1 U16428 ( .B1(n7727), .B2(n14921), .A(n14686), .ZN(n14687) );
  AOI21_X1 U16429 ( .B1(n14982), .B2(n14907), .A(n14687), .ZN(n14691) );
  XNOR2_X1 U16430 ( .A(n14688), .B(n14689), .ZN(n14985) );
  OR2_X1 U16431 ( .A1(n14985), .A2(n14910), .ZN(n14690) );
  OAI211_X1 U16432 ( .C1(n14986), .C2(n6412), .A(n14691), .B(n14690), .ZN(
        P1_U3266) );
  INV_X1 U16433 ( .A(n14749), .ZN(n14695) );
  XOR2_X1 U16434 ( .A(n14702), .B(n14696), .Z(n14991) );
  OAI211_X1 U16435 ( .C1(n14720), .C2(n14700), .A(n15216), .B(n14697), .ZN(
        n14987) );
  INV_X1 U16436 ( .A(n14987), .ZN(n14708) );
  AOI22_X1 U16437 ( .A1(n14698), .A2(n14974), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n6412), .ZN(n14699) );
  OAI21_X1 U16438 ( .B1(n14700), .B2(n14921), .A(n14699), .ZN(n14707) );
  AOI21_X1 U16439 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14704) );
  INV_X1 U16440 ( .A(n14705), .ZN(n14989) );
  AOI21_X1 U16441 ( .B1(n14990), .B2(n14989), .A(n6412), .ZN(n14706) );
  OAI21_X1 U16442 ( .B1(n14991), .B2(n14910), .A(n14709), .ZN(P1_U3267) );
  XNOR2_X1 U16443 ( .A(n14713), .B(n14716), .ZN(n14998) );
  INV_X1 U16444 ( .A(n14850), .ZN(n14873) );
  AND2_X1 U16445 ( .A1(n14732), .A2(n14733), .ZN(n14714) );
  NOR2_X1 U16446 ( .A1(n14735), .A2(n14715), .ZN(n14718) );
  INV_X1 U16447 ( .A(n14716), .ZN(n14717) );
  XNOR2_X1 U16448 ( .A(n14718), .B(n14717), .ZN(n14992) );
  NAND2_X1 U16449 ( .A1(n14992), .A2(n15227), .ZN(n14729) );
  INV_X1 U16450 ( .A(n14719), .ZN(n14721) );
  AOI211_X1 U16451 ( .C1(n14995), .C2(n14721), .A(n14929), .B(n14720), .ZN(
        n14993) );
  INV_X1 U16452 ( .A(n14722), .ZN(n14723) );
  AOI22_X1 U16453 ( .A1(n14723), .A2(n14974), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n6412), .ZN(n14725) );
  NAND2_X1 U16454 ( .A1(n14994), .A2(n15220), .ZN(n14724) );
  OAI211_X1 U16455 ( .C1(n14726), .C2(n14921), .A(n14725), .B(n14724), .ZN(
        n14727) );
  AOI21_X1 U16456 ( .B1(n14993), .B2(n14907), .A(n14727), .ZN(n14728) );
  OAI211_X1 U16457 ( .C1(n14998), .C2(n14873), .A(n14729), .B(n14728), .ZN(
        P1_U3268) );
  NAND2_X1 U16458 ( .A1(n14730), .A2(n14732), .ZN(n14731) );
  AOI21_X1 U16459 ( .B1(n14749), .B2(n14733), .A(n14732), .ZN(n14734) );
  NAND2_X1 U16460 ( .A1(n14736), .A2(n15263), .ZN(n14738) );
  NAND2_X1 U16461 ( .A1(n14740), .A2(n14739), .ZN(n14741) );
  NAND2_X1 U16462 ( .A1(n14741), .A2(n15216), .ZN(n14742) );
  OR2_X1 U16463 ( .A1(n14719), .A2(n14742), .ZN(n14999) );
  INV_X1 U16464 ( .A(n14999), .ZN(n14746) );
  AOI22_X1 U16465 ( .A1(n14743), .A2(n14974), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n6412), .ZN(n14744) );
  OAI21_X1 U16466 ( .B1(n15000), .B2(n14921), .A(n14744), .ZN(n14745) );
  AOI21_X1 U16467 ( .B1(n14746), .B2(n14907), .A(n14745), .ZN(n14747) );
  OAI21_X1 U16468 ( .B1(n6438), .B2(n6412), .A(n14747), .ZN(P1_U3269) );
  OAI21_X1 U16469 ( .B1(n14692), .B2(n14750), .A(n14749), .ZN(n15008) );
  INV_X1 U16470 ( .A(n14710), .ZN(n14753) );
  OAI21_X1 U16471 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14755) );
  AOI21_X1 U16472 ( .B1(n14755), .B2(n15251), .A(n14754), .ZN(n15007) );
  INV_X1 U16473 ( .A(n15007), .ZN(n14762) );
  XNOR2_X1 U16474 ( .A(n14771), .B(n7731), .ZN(n14756) );
  NAND2_X1 U16475 ( .A1(n15004), .A2(n14907), .ZN(n14760) );
  INV_X1 U16476 ( .A(n14757), .ZN(n14758) );
  AOI22_X1 U16477 ( .A1(n14758), .A2(n14974), .B1(n6412), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n14759) );
  OAI211_X1 U16478 ( .C1(n7731), .C2(n14921), .A(n14760), .B(n14759), .ZN(
        n14761) );
  AOI21_X1 U16479 ( .B1(n14762), .B2(n15220), .A(n14761), .ZN(n14763) );
  OAI21_X1 U16480 ( .B1(n14910), .B2(n15008), .A(n14763), .ZN(P1_U3270) );
  OAI21_X1 U16481 ( .B1(n14764), .B2(n14766), .A(n14765), .ZN(n14767) );
  INV_X1 U16482 ( .A(n14767), .ZN(n15014) );
  XNOR2_X1 U16483 ( .A(n14769), .B(n14768), .ZN(n15012) );
  OAI211_X1 U16484 ( .C1(n14770), .C2(n9615), .A(n15216), .B(n14771), .ZN(
        n15010) );
  INV_X1 U16485 ( .A(n9615), .ZN(n14775) );
  AOI22_X1 U16486 ( .A1(n6412), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14772), 
        .B2(n14974), .ZN(n14773) );
  OAI21_X1 U16487 ( .B1(n15009), .B2(n6412), .A(n14773), .ZN(n14774) );
  AOI21_X1 U16488 ( .B1(n14775), .B2(n15223), .A(n14774), .ZN(n14776) );
  OAI21_X1 U16489 ( .B1(n15010), .B2(n15225), .A(n14776), .ZN(n14777) );
  AOI21_X1 U16490 ( .B1(n15012), .B2(n14850), .A(n14777), .ZN(n14778) );
  OAI21_X1 U16491 ( .B1(n15014), .B2(n14910), .A(n14778), .ZN(P1_U3271) );
  XOR2_X1 U16492 ( .A(n14780), .B(n14779), .Z(n15019) );
  XNOR2_X1 U16493 ( .A(n14781), .B(n14780), .ZN(n14782) );
  OAI222_X1 U16494 ( .A1(n14933), .A2(n14784), .B1(n14935), .B2(n14783), .C1(
        n14782), .C2(n15050), .ZN(n15015) );
  OAI21_X1 U16495 ( .B1(n14785), .B2(n14790), .A(n15216), .ZN(n14786) );
  NOR2_X1 U16496 ( .A1(n14786), .A2(n14770), .ZN(n15016) );
  NAND2_X1 U16497 ( .A1(n15016), .A2(n14907), .ZN(n14789) );
  AOI22_X1 U16498 ( .A1(n6412), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14787), 
        .B2(n14974), .ZN(n14788) );
  OAI211_X1 U16499 ( .C1(n14790), .C2(n14921), .A(n14789), .B(n14788), .ZN(
        n14791) );
  AOI21_X1 U16500 ( .B1(n15015), .B2(n15220), .A(n14791), .ZN(n14792) );
  OAI21_X1 U16501 ( .B1(n15019), .B2(n14910), .A(n14792), .ZN(P1_U3272) );
  OAI21_X1 U16502 ( .B1(n6441), .B2(n7674), .A(n14793), .ZN(n15025) );
  NAND2_X1 U16503 ( .A1(n14811), .A2(n15022), .ZN(n14794) );
  NAND2_X1 U16504 ( .A1(n14794), .A2(n15216), .ZN(n14795) );
  NOR2_X1 U16505 ( .A1(n14785), .A2(n14795), .ZN(n15020) );
  NAND2_X1 U16506 ( .A1(n15022), .A2(n15223), .ZN(n14798) );
  AOI22_X1 U16507 ( .A1(n6412), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14796), 
        .B2(n14974), .ZN(n14797) );
  NAND2_X1 U16508 ( .A1(n14798), .A2(n14797), .ZN(n14808) );
  OR2_X1 U16509 ( .A1(n14799), .A2(n14815), .ZN(n14802) );
  AND2_X1 U16510 ( .A1(n14802), .A2(n14800), .ZN(n14805) );
  NAND2_X1 U16511 ( .A1(n14802), .A2(n14801), .ZN(n14803) );
  OAI211_X1 U16512 ( .C1(n14805), .C2(n14804), .A(n14803), .B(n15251), .ZN(
        n15023) );
  AOI21_X1 U16513 ( .B1(n15023), .B2(n14806), .A(n6412), .ZN(n14807) );
  AOI211_X1 U16514 ( .C1(n15020), .C2(n14907), .A(n14808), .B(n14807), .ZN(
        n14809) );
  OAI21_X1 U16515 ( .B1(n14910), .B2(n15025), .A(n14809), .ZN(P1_U3273) );
  XNOR2_X1 U16516 ( .A(n14810), .B(n14815), .ZN(n15031) );
  AOI211_X1 U16517 ( .C1(n15028), .C2(n14831), .A(n14929), .B(n9795), .ZN(
        n15026) );
  AOI22_X1 U16518 ( .A1(n6412), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14812), 
        .B2(n14974), .ZN(n14813) );
  OAI21_X1 U16519 ( .B1(n14814), .B2(n14921), .A(n14813), .ZN(n14821) );
  XNOR2_X1 U16520 ( .A(n14799), .B(n14815), .ZN(n14817) );
  AOI22_X1 U16521 ( .A1(n14817), .A2(n15251), .B1(n14897), .B2(n14816), .ZN(
        n15030) );
  AND2_X1 U16522 ( .A1(n14818), .A2(n14880), .ZN(n15027) );
  INV_X1 U16523 ( .A(n15027), .ZN(n14819) );
  AOI21_X1 U16524 ( .B1(n15030), .B2(n14819), .A(n6412), .ZN(n14820) );
  AOI211_X1 U16525 ( .C1(n15026), .C2(n14907), .A(n14821), .B(n14820), .ZN(
        n14822) );
  OAI21_X1 U16526 ( .B1(n14910), .B2(n15031), .A(n14822), .ZN(P1_U3274) );
  XOR2_X1 U16527 ( .A(n14823), .B(n14824), .Z(n15036) );
  XNOR2_X1 U16528 ( .A(n14825), .B(n14824), .ZN(n14826) );
  OAI222_X1 U16529 ( .A1(n14933), .A2(n14827), .B1(n14935), .B2(n14861), .C1(
        n14826), .C2(n15050), .ZN(n15032) );
  OR2_X1 U16530 ( .A1(n14828), .A2(n14829), .ZN(n14830) );
  AND3_X1 U16531 ( .A1(n14831), .A2(n15216), .A3(n14830), .ZN(n15033) );
  NAND2_X1 U16532 ( .A1(n15033), .A2(n14907), .ZN(n14836) );
  NAND2_X1 U16533 ( .A1(n6412), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14832) );
  OAI21_X1 U16534 ( .B1(n15217), .B2(n14833), .A(n14832), .ZN(n14834) );
  AOI21_X1 U16535 ( .B1(n15034), .B2(n15223), .A(n14834), .ZN(n14835) );
  NAND2_X1 U16536 ( .A1(n14836), .A2(n14835), .ZN(n14837) );
  AOI21_X1 U16537 ( .B1(n15032), .B2(n15220), .A(n14837), .ZN(n14838) );
  OAI21_X1 U16538 ( .B1(n15036), .B2(n14910), .A(n14838), .ZN(P1_U3275) );
  XOR2_X1 U16539 ( .A(n14843), .B(n14839), .Z(n15042) );
  INV_X1 U16540 ( .A(n14840), .ZN(n14841) );
  AOI21_X1 U16541 ( .B1(n14843), .B2(n14842), .A(n14841), .ZN(n15040) );
  AOI211_X1 U16542 ( .C1(n14844), .C2(n14859), .A(n14929), .B(n14828), .ZN(
        n15039) );
  NAND2_X1 U16543 ( .A1(n15039), .A2(n14907), .ZN(n14848) );
  OAI22_X1 U16544 ( .A1(n6412), .A2(n15037), .B1(n14845), .B2(n15217), .ZN(
        n14846) );
  AOI21_X1 U16545 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n6412), .A(n14846), .ZN(
        n14847) );
  OAI211_X1 U16546 ( .C1(n7717), .C2(n14921), .A(n14848), .B(n14847), .ZN(
        n14849) );
  AOI21_X1 U16547 ( .B1(n15040), .B2(n14850), .A(n14849), .ZN(n14851) );
  OAI21_X1 U16548 ( .B1(n15042), .B2(n14910), .A(n14851), .ZN(P1_U3276) );
  XNOR2_X1 U16549 ( .A(n14852), .B(n14853), .ZN(n15049) );
  OAI21_X1 U16550 ( .B1(n14857), .B2(n14856), .A(n14855), .ZN(n15043) );
  NAND2_X1 U16551 ( .A1(n15043), .A2(n15227), .ZN(n14872) );
  INV_X1 U16552 ( .A(n14859), .ZN(n14860) );
  AOI211_X1 U16553 ( .C1(n15046), .C2(n14858), .A(n14929), .B(n14860), .ZN(
        n15044) );
  INV_X1 U16554 ( .A(n15046), .ZN(n14869) );
  OR2_X1 U16555 ( .A1(n14861), .A2(n14933), .ZN(n14864) );
  OR2_X1 U16556 ( .A1(n14862), .A2(n14935), .ZN(n14863) );
  NAND2_X1 U16557 ( .A1(n14864), .A2(n14863), .ZN(n15045) );
  INV_X1 U16558 ( .A(n14865), .ZN(n14866) );
  AOI22_X1 U16559 ( .A1(n15220), .A2(n15045), .B1(n14866), .B2(n14974), .ZN(
        n14868) );
  NAND2_X1 U16560 ( .A1(n6412), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14867) );
  OAI211_X1 U16561 ( .C1(n14869), .C2(n14921), .A(n14868), .B(n14867), .ZN(
        n14870) );
  AOI21_X1 U16562 ( .B1(n15044), .B2(n14907), .A(n14870), .ZN(n14871) );
  OAI211_X1 U16563 ( .C1(n15049), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        P1_U3277) );
  XNOR2_X1 U16564 ( .A(n14875), .B(n14874), .ZN(n15055) );
  XNOR2_X1 U16565 ( .A(n14876), .B(n14877), .ZN(n14878) );
  NOR2_X1 U16566 ( .A1(n14878), .A2(n15050), .ZN(n15051) );
  OAI211_X1 U16567 ( .C1(n14900), .C2(n14888), .A(n14858), .B(n15216), .ZN(
        n14883) );
  AOI22_X1 U16568 ( .A1(n14881), .A2(n14897), .B1(n14880), .B2(n14879), .ZN(
        n14882) );
  NAND2_X1 U16569 ( .A1(n14883), .A2(n14882), .ZN(n15052) );
  NAND2_X1 U16570 ( .A1(n15052), .A2(n14907), .ZN(n14887) );
  INV_X1 U16571 ( .A(n14884), .ZN(n14885) );
  AOI22_X1 U16572 ( .A1(n6412), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14885), 
        .B2(n14974), .ZN(n14886) );
  OAI211_X1 U16573 ( .C1(n14888), .C2(n14921), .A(n14887), .B(n14886), .ZN(
        n14889) );
  AOI21_X1 U16574 ( .B1(n15051), .B2(n15220), .A(n14889), .ZN(n14890) );
  OAI21_X1 U16575 ( .B1(n14910), .B2(n15055), .A(n14890), .ZN(P1_U3278) );
  NAND2_X1 U16576 ( .A1(n14891), .A2(n14895), .ZN(n14892) );
  NAND2_X1 U16577 ( .A1(n14893), .A2(n14892), .ZN(n15061) );
  XOR2_X1 U16578 ( .A(n14894), .B(n14895), .Z(n14898) );
  AOI22_X1 U16579 ( .A1(n14898), .A2(n15251), .B1(n14897), .B2(n14896), .ZN(
        n15060) );
  INV_X1 U16580 ( .A(n15060), .ZN(n14899) );
  OAI21_X1 U16581 ( .B1(n14899), .B2(n15056), .A(n15220), .ZN(n14909) );
  AOI211_X1 U16582 ( .C1(n14901), .C2(n14912), .A(n14929), .B(n14900), .ZN(
        n15058) );
  NOR2_X1 U16583 ( .A1(n14902), .A2(n14921), .ZN(n14906) );
  OAI22_X1 U16584 ( .A1(n15220), .A2(n14904), .B1(n14903), .B2(n15217), .ZN(
        n14905) );
  AOI211_X1 U16585 ( .C1(n15058), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14908) );
  OAI211_X1 U16586 ( .C1(n15061), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        P1_U3279) );
  AOI21_X1 U16587 ( .B1(n14930), .B2(n15065), .A(n14929), .ZN(n14911) );
  AND2_X1 U16588 ( .A1(n14912), .A2(n14911), .ZN(n15063) );
  XNOR2_X1 U16589 ( .A(n14914), .B(n14919), .ZN(n14915) );
  NAND2_X1 U16590 ( .A1(n14915), .A2(n15251), .ZN(n15066) );
  INV_X1 U16591 ( .A(n15066), .ZN(n14916) );
  AOI211_X1 U16592 ( .C1(n15063), .C2(n14917), .A(n15064), .B(n14916), .ZN(
        n14928) );
  OAI21_X1 U16593 ( .B1(n14920), .B2(n14919), .A(n6642), .ZN(n15062) );
  NOR2_X1 U16594 ( .A1(n14922), .A2(n14921), .ZN(n14926) );
  OAI22_X1 U16595 ( .A1(n15220), .A2(n14924), .B1(n14923), .B2(n15217), .ZN(
        n14925) );
  AOI211_X1 U16596 ( .C1(n15062), .C2(n15227), .A(n14926), .B(n14925), .ZN(
        n14927) );
  OAI21_X1 U16597 ( .B1(n14928), .B2(n6412), .A(n14927), .ZN(P1_U3280) );
  AOI21_X1 U16598 ( .B1(n11958), .B2(n14951), .A(n14929), .ZN(n14931) );
  NAND2_X1 U16599 ( .A1(n14931), .A2(n14930), .ZN(n15069) );
  INV_X1 U16600 ( .A(n14932), .ZN(n14947) );
  OAI22_X1 U16601 ( .A1(n14936), .A2(n14935), .B1(n14934), .B2(n14933), .ZN(
        n14946) );
  NAND3_X1 U16602 ( .A1(n14939), .A2(n15263), .A3(n14938), .ZN(n14940) );
  OAI21_X1 U16603 ( .B1(n15050), .B2(n14937), .A(n14940), .ZN(n14944) );
  INV_X1 U16604 ( .A(n14937), .ZN(n14941) );
  NOR2_X1 U16605 ( .A1(n14941), .A2(n15050), .ZN(n14943) );
  MUX2_X1 U16606 ( .A(n14944), .B(n14943), .S(n14942), .Z(n14945) );
  AOI211_X1 U16607 ( .C1(n14947), .C2(n15263), .A(n14946), .B(n14945), .ZN(
        n15070) );
  OR2_X1 U16608 ( .A1(n15070), .A2(n6412), .ZN(n14953) );
  NAND2_X1 U16609 ( .A1(n6412), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n14948) );
  OAI21_X1 U16610 ( .B1(n15217), .B2(n14949), .A(n14948), .ZN(n14950) );
  AOI21_X1 U16611 ( .B1(n14951), .B2(n15223), .A(n14950), .ZN(n14952) );
  OAI211_X1 U16612 ( .C1(n15069), .C2(n15225), .A(n14953), .B(n14952), .ZN(
        P1_U3281) );
  INV_X1 U16613 ( .A(n14954), .ZN(n14955) );
  AOI22_X1 U16614 ( .A1(n15223), .A2(n14956), .B1(n14974), .B2(n14955), .ZN(
        n14957) );
  OAI21_X1 U16615 ( .B1(n14958), .B2(n14966), .A(n14957), .ZN(n14961) );
  MUX2_X1 U16616 ( .A(n14959), .B(P1_REG2_REG_8__SCAN_IN), .S(n6412), .Z(
        n14960) );
  AOI211_X1 U16617 ( .C1(n15227), .C2(n14962), .A(n14961), .B(n14960), .ZN(
        n14963) );
  INV_X1 U16618 ( .A(n14963), .ZN(P1_U3285) );
  OAI22_X1 U16619 ( .A1(n14966), .A2(n14965), .B1(n14964), .B2(n15217), .ZN(
        n14969) );
  MUX2_X1 U16620 ( .A(n14967), .B(P1_REG2_REG_1__SCAN_IN), .S(n6412), .Z(
        n14968) );
  AOI211_X1 U16621 ( .C1(n15223), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n14971) );
  INV_X1 U16622 ( .A(n14971), .ZN(P1_U3292) );
  OAI21_X1 U16623 ( .B1(n14973), .B2(n15223), .A(n14972), .ZN(n14976) );
  AOI22_X1 U16624 ( .A1(n6412), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14974), .ZN(n14975) );
  OAI211_X1 U16625 ( .C1(n6412), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        P1_U3293) );
  MUX2_X1 U16626 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14978), .S(n15272), .Z(
        P1_U3559) );
  OAI211_X1 U16627 ( .C1(n14981), .C2(n15259), .A(n14980), .B(n14979), .ZN(
        n15083) );
  MUX2_X1 U16628 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15083), .S(n15272), .Z(
        P1_U3558) );
  AOI21_X1 U16629 ( .B1(n15255), .B2(n14983), .A(n14982), .ZN(n14984) );
  MUX2_X1 U16630 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15084), .S(n15272), .Z(
        P1_U3555) );
  MUX2_X1 U16631 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15085), .S(n15272), .Z(
        P1_U3554) );
  NAND2_X1 U16632 ( .A1(n14992), .A2(n15263), .ZN(n14997) );
  AOI211_X1 U16633 ( .C1(n15255), .C2(n14995), .A(n14994), .B(n14993), .ZN(
        n14996) );
  OAI211_X1 U16634 ( .C1(n14998), .C2(n15050), .A(n14997), .B(n14996), .ZN(
        n15086) );
  MUX2_X1 U16635 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15086), .S(n15272), .Z(
        P1_U3553) );
  OAI21_X1 U16636 ( .B1(n15000), .B2(n15259), .A(n14999), .ZN(n15001) );
  INV_X1 U16637 ( .A(n15003), .ZN(P1_U3552) );
  AOI21_X1 U16638 ( .B1(n15255), .B2(n15005), .A(n15004), .ZN(n15006) );
  OAI211_X1 U16639 ( .C1(n15008), .C2(n15247), .A(n15007), .B(n15006), .ZN(
        n15089) );
  MUX2_X1 U16640 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15089), .S(n15272), .Z(
        P1_U3551) );
  OAI211_X1 U16641 ( .C1(n15259), .C2(n9615), .A(n15010), .B(n15009), .ZN(
        n15011) );
  AOI21_X1 U16642 ( .B1(n15012), .B2(n15251), .A(n15011), .ZN(n15013) );
  OAI21_X1 U16643 ( .B1(n15014), .B2(n15247), .A(n15013), .ZN(n15090) );
  MUX2_X1 U16644 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15090), .S(n15272), .Z(
        P1_U3550) );
  AOI211_X1 U16645 ( .C1(n15255), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        n15018) );
  OAI21_X1 U16646 ( .B1(n15019), .B2(n15247), .A(n15018), .ZN(n15091) );
  MUX2_X1 U16647 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15091), .S(n15272), .Z(
        P1_U3549) );
  AOI211_X1 U16648 ( .C1(n15255), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15024) );
  OAI211_X1 U16649 ( .C1(n15025), .C2(n15247), .A(n15024), .B(n15023), .ZN(
        n15092) );
  MUX2_X1 U16650 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15092), .S(n15272), .Z(
        P1_U3548) );
  AOI211_X1 U16651 ( .C1(n15255), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        n15029) );
  OAI211_X1 U16652 ( .C1(n15031), .C2(n15247), .A(n15030), .B(n15029), .ZN(
        n15093) );
  MUX2_X1 U16653 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15093), .S(n15272), .Z(
        P1_U3547) );
  AOI211_X1 U16654 ( .C1(n15255), .C2(n15034), .A(n15033), .B(n15032), .ZN(
        n15035) );
  OAI21_X1 U16655 ( .B1(n15036), .B2(n15247), .A(n15035), .ZN(n15094) );
  MUX2_X1 U16656 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15094), .S(n15272), .Z(
        P1_U3546) );
  OAI21_X1 U16657 ( .B1(n7717), .B2(n15259), .A(n15037), .ZN(n15038) );
  AOI211_X1 U16658 ( .C1(n15040), .C2(n15251), .A(n15039), .B(n15038), .ZN(
        n15041) );
  OAI21_X1 U16659 ( .B1(n15042), .B2(n15247), .A(n15041), .ZN(n15095) );
  MUX2_X1 U16660 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15095), .S(n15272), .Z(
        P1_U3545) );
  NAND2_X1 U16661 ( .A1(n15043), .A2(n15263), .ZN(n15048) );
  AOI211_X1 U16662 ( .C1(n15255), .C2(n15046), .A(n15045), .B(n15044), .ZN(
        n15047) );
  OAI211_X1 U16663 ( .C1(n15050), .C2(n15049), .A(n15048), .B(n15047), .ZN(
        n15096) );
  MUX2_X1 U16664 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15096), .S(n15272), .Z(
        P1_U3544) );
  AOI211_X1 U16665 ( .C1(n15255), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15054) );
  OAI21_X1 U16666 ( .B1(n15247), .B2(n15055), .A(n15054), .ZN(n15097) );
  MUX2_X1 U16667 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15097), .S(n15272), .Z(
        P1_U3543) );
  NOR3_X1 U16668 ( .A1(n15058), .A2(n15057), .A3(n15056), .ZN(n15059) );
  OAI211_X1 U16669 ( .C1(n15247), .C2(n15061), .A(n15060), .B(n15059), .ZN(
        n15098) );
  MUX2_X1 U16670 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15098), .S(n15272), .Z(
        P1_U3542) );
  INV_X1 U16671 ( .A(n15062), .ZN(n15068) );
  AOI211_X1 U16672 ( .C1(n15255), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        n15067) );
  OAI211_X1 U16673 ( .C1(n15068), .C2(n15247), .A(n15067), .B(n15066), .ZN(
        n15099) );
  MUX2_X1 U16674 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15099), .S(n15272), .Z(
        P1_U3541) );
  OAI211_X1 U16675 ( .C1(n15071), .C2(n15259), .A(n15070), .B(n15069), .ZN(
        n15100) );
  MUX2_X1 U16676 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15100), .S(n15272), .Z(
        P1_U3540) );
  NAND2_X1 U16677 ( .A1(n15072), .A2(n15263), .ZN(n15074) );
  NAND4_X1 U16678 ( .A1(n15076), .A2(n15075), .A3(n15074), .A4(n15073), .ZN(
        n15101) );
  MUX2_X1 U16679 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15101), .S(n15272), .Z(
        P1_U3539) );
  AOI211_X1 U16680 ( .C1(n15255), .C2(n15079), .A(n15078), .B(n15077), .ZN(
        n15080) );
  OAI21_X1 U16681 ( .B1(n15081), .B2(n15247), .A(n15080), .ZN(n15102) );
  MUX2_X1 U16682 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15102), .S(n15272), .Z(
        P1_U3538) );
  MUX2_X1 U16683 ( .A(n15082), .B(P1_REG1_REG_0__SCAN_IN), .S(n15270), .Z(
        P1_U3528) );
  MUX2_X1 U16684 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15083), .S(n15265), .Z(
        P1_U3526) );
  MUX2_X1 U16685 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15084), .S(n15265), .Z(
        P1_U3523) );
  MUX2_X1 U16686 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15085), .S(n15265), .Z(
        P1_U3522) );
  MUX2_X1 U16687 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15086), .S(n15265), .Z(
        P1_U3521) );
  INV_X1 U16688 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15088) );
  MUX2_X1 U16689 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15089), .S(n15265), .Z(
        P1_U3519) );
  MUX2_X1 U16690 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15090), .S(n15265), .Z(
        P1_U3518) );
  MUX2_X1 U16691 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15091), .S(n15265), .Z(
        P1_U3517) );
  MUX2_X1 U16692 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15092), .S(n15265), .Z(
        P1_U3516) );
  MUX2_X1 U16693 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15093), .S(n15265), .Z(
        P1_U3515) );
  MUX2_X1 U16694 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15094), .S(n15265), .Z(
        P1_U3513) );
  MUX2_X1 U16695 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15095), .S(n15265), .Z(
        P1_U3510) );
  MUX2_X1 U16696 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15096), .S(n15265), .Z(
        P1_U3507) );
  MUX2_X1 U16697 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15097), .S(n15265), .Z(
        P1_U3504) );
  MUX2_X1 U16698 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15098), .S(n15265), .Z(
        P1_U3501) );
  MUX2_X1 U16699 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15099), .S(n15265), .Z(
        P1_U3498) );
  MUX2_X1 U16700 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15100), .S(n15265), .Z(
        P1_U3495) );
  MUX2_X1 U16701 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15101), .S(n15265), .Z(
        P1_U3492) );
  MUX2_X1 U16702 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n15102), .S(n15265), .Z(
        P1_U3489) );
  OAI222_X1 U16703 ( .A1(n15105), .A2(n15104), .B1(P1_U3086), .B2(n9333), .C1(
        n10976), .C2(n15103), .ZN(P1_U3325) );
  OAI222_X1 U16704 ( .A1(n15105), .A2(n15108), .B1(n10976), .B2(n15107), .C1(
        n15106), .C2(P1_U3086), .ZN(P1_U3328) );
  MUX2_X1 U16705 ( .A(n14245), .B(n15109), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16706 ( .A(n6639), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NAND2_X1 U16707 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15113), .ZN(n15114) );
  NAND2_X1 U16708 ( .A1(n15115), .A2(n15114), .ZN(n15118) );
  NAND2_X1 U16709 ( .A1(n15116), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15117) );
  NAND2_X1 U16710 ( .A1(n15118), .A2(n15117), .ZN(n15127) );
  INV_X1 U16711 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15472) );
  NAND2_X1 U16712 ( .A1(n15472), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15128) );
  OAI21_X1 U16713 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n15472), .A(n15128), 
        .ZN(n15119) );
  XNOR2_X1 U16714 ( .A(n15127), .B(n15119), .ZN(n15120) );
  OAI21_X1 U16715 ( .B1(n15122), .B2(n15124), .A(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n15123) );
  OAI21_X1 U16716 ( .B1(n7304), .B2(n15124), .A(n15123), .ZN(SUB_1596_U66) );
  AND2_X1 U16717 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15125), .ZN(n15126) );
  NAND2_X1 U16718 ( .A1(n15129), .A2(n15128), .ZN(n15134) );
  INV_X1 U16719 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U16720 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15130), .ZN(n15137) );
  INV_X1 U16721 ( .A(n15137), .ZN(n15131) );
  AOI21_X1 U16722 ( .B1(n15132), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15131), 
        .ZN(n15133) );
  NAND2_X1 U16723 ( .A1(n15134), .A2(n15133), .ZN(n15138) );
  OR2_X1 U16724 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  NAND2_X1 U16725 ( .A1(n15138), .A2(n15135), .ZN(n15142) );
  XOR2_X1 U16726 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15142), .Z(n15136) );
  XNOR2_X1 U16727 ( .A(n15140), .B(n15136), .ZN(SUB_1596_U65) );
  NAND2_X1 U16728 ( .A1(n15138), .A2(n15137), .ZN(n15146) );
  XNOR2_X1 U16729 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n15139) );
  XNOR2_X1 U16730 ( .A(n15146), .B(n15139), .ZN(n15141) );
  NAND2_X1 U16731 ( .A1(n6923), .A2(n15144), .ZN(n15143) );
  XNOR2_X1 U16732 ( .A(n15143), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OR2_X1 U16733 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15147), .ZN(n15145) );
  NAND2_X1 U16734 ( .A1(n15146), .A2(n15145), .ZN(n15149) );
  NAND2_X1 U16735 ( .A1(n15147), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15148) );
  NAND2_X1 U16736 ( .A1(n15149), .A2(n15148), .ZN(n15156) );
  XNOR2_X1 U16737 ( .A(n15156), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15155) );
  XNOR2_X1 U16738 ( .A(n15155), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U16739 ( .A1(n15152), .A2(n15154), .ZN(n15153) );
  XNOR2_X1 U16740 ( .A(n15153), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U16741 ( .A(n15155), .ZN(n15158) );
  NOR2_X1 U16742 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15156), .ZN(n15157) );
  AOI21_X1 U16743 ( .B1(n15158), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15157), 
        .ZN(n15164) );
  XNOR2_X1 U16744 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15159) );
  XNOR2_X1 U16745 ( .A(n15160), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  INV_X1 U16746 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U16747 ( .A1(n15448), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15163) );
  INV_X1 U16748 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15162) );
  AOI22_X1 U16749 ( .A1(n15164), .A2(n15163), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15162), .ZN(n15167) );
  XNOR2_X1 U16750 ( .A(n15165), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15166) );
  AOI21_X1 U16751 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15168) );
  OAI21_X1 U16752 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n15168), 
        .ZN(U28) );
  AOI21_X1 U16753 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15169) );
  OAI21_X1 U16754 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15169), 
        .ZN(U29) );
  AND2_X1 U16755 ( .A1(n15255), .A2(n15170), .ZN(n15232) );
  AOI22_X1 U16756 ( .A1(n15171), .A2(n15232), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15181) );
  INV_X1 U16757 ( .A(n15172), .ZN(n15178) );
  AOI211_X1 U16758 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15177) );
  AOI21_X1 U16759 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n15180) );
  OAI211_X1 U16760 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n15182), .A(n15181), .B(
        n15180), .ZN(P1_U3218) );
  MUX2_X1 U16761 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10252), .S(n15195), .Z(
        n15183) );
  NAND3_X1 U16762 ( .A1(n15185), .A2(n15184), .A3(n15183), .ZN(n15186) );
  NAND3_X1 U16763 ( .A1(n15188), .A2(n15187), .A3(n15186), .ZN(n15203) );
  NAND3_X1 U16764 ( .A1(n15191), .A2(n15190), .A3(n15189), .ZN(n15192) );
  NAND3_X1 U16765 ( .A1(n15194), .A2(n15193), .A3(n15192), .ZN(n15202) );
  INV_X1 U16766 ( .A(n15195), .ZN(n15196) );
  NAND2_X1 U16767 ( .A1(n15197), .A2(n15196), .ZN(n15201) );
  AND2_X1 U16768 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15198) );
  AOI21_X1 U16769 ( .B1(n15199), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n15198), .ZN(
        n15200) );
  AND4_X1 U16770 ( .A1(n15203), .A2(n15202), .A3(n15201), .A4(n15200), .ZN(
        n15205) );
  NAND2_X1 U16771 ( .A1(n15205), .A2(n15204), .ZN(P1_U3247) );
  XNOR2_X1 U16772 ( .A(n15207), .B(n15206), .ZN(n15210) );
  INV_X1 U16773 ( .A(n15208), .ZN(n15209) );
  AOI21_X1 U16774 ( .B1(n15210), .B2(n15251), .A(n15209), .ZN(n15238) );
  OAI21_X1 U16775 ( .B1(n15213), .B2(n15212), .A(n15211), .ZN(n15241) );
  OAI211_X1 U16776 ( .C1(n9794), .C2(n15237), .A(n15216), .B(n15215), .ZN(
        n15236) );
  OAI22_X1 U16777 ( .A1(n15220), .A2(n15219), .B1(n15218), .B2(n15217), .ZN(
        n15221) );
  AOI21_X1 U16778 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15224) );
  OAI21_X1 U16779 ( .B1(n15225), .B2(n15236), .A(n15224), .ZN(n15226) );
  AOI21_X1 U16780 ( .B1(n15227), .B2(n15241), .A(n15226), .ZN(n15228) );
  OAI21_X1 U16781 ( .B1(n6412), .B2(n15238), .A(n15228), .ZN(P1_U3289) );
  AND2_X1 U16782 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15230), .ZN(P1_U3294) );
  AND2_X1 U16783 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15230), .ZN(P1_U3295) );
  AND2_X1 U16784 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15230), .ZN(P1_U3296) );
  AND2_X1 U16785 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15230), .ZN(P1_U3297) );
  AND2_X1 U16786 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15230), .ZN(P1_U3298) );
  AND2_X1 U16787 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15230), .ZN(P1_U3299) );
  AND2_X1 U16788 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15230), .ZN(P1_U3300) );
  AND2_X1 U16789 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15230), .ZN(P1_U3301) );
  AND2_X1 U16790 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15230), .ZN(P1_U3302) );
  AND2_X1 U16791 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15230), .ZN(P1_U3303) );
  AND2_X1 U16792 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15230), .ZN(P1_U3304) );
  AND2_X1 U16793 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15230), .ZN(P1_U3305) );
  INV_X1 U16794 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15469) );
  NOR2_X1 U16795 ( .A1(n15229), .A2(n15469), .ZN(P1_U3306) );
  AND2_X1 U16796 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15230), .ZN(P1_U3307) );
  AND2_X1 U16797 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15230), .ZN(P1_U3308) );
  AND2_X1 U16798 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15230), .ZN(P1_U3309) );
  INV_X1 U16799 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15511) );
  NOR2_X1 U16800 ( .A1(n15229), .A2(n15511), .ZN(P1_U3310) );
  AND2_X1 U16801 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15230), .ZN(P1_U3311) );
  AND2_X1 U16802 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15230), .ZN(P1_U3312) );
  AND2_X1 U16803 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15230), .ZN(P1_U3313) );
  AND2_X1 U16804 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15230), .ZN(P1_U3314) );
  AND2_X1 U16805 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15230), .ZN(P1_U3315) );
  AND2_X1 U16806 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15230), .ZN(P1_U3316) );
  AND2_X1 U16807 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15230), .ZN(P1_U3317) );
  AND2_X1 U16808 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15230), .ZN(P1_U3318) );
  AND2_X1 U16809 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15230), .ZN(P1_U3319) );
  AND2_X1 U16810 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15230), .ZN(P1_U3320) );
  AND2_X1 U16811 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15230), .ZN(P1_U3321) );
  AND2_X1 U16812 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15230), .ZN(P1_U3322) );
  AND2_X1 U16813 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15230), .ZN(P1_U3323) );
  INV_X1 U16814 ( .A(n15231), .ZN(n15233) );
  NOR3_X1 U16815 ( .A1(n15234), .A2(n15233), .A3(n15232), .ZN(n15266) );
  INV_X1 U16816 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U16817 ( .A1(n15265), .A2(n15266), .B1(n15235), .B2(n15264), .ZN(
        P1_U3468) );
  OAI21_X1 U16818 ( .B1(n15237), .B2(n15259), .A(n15236), .ZN(n15240) );
  INV_X1 U16819 ( .A(n15238), .ZN(n15239) );
  AOI211_X1 U16820 ( .C1(n15263), .C2(n15241), .A(n15240), .B(n15239), .ZN(
        n15267) );
  INV_X1 U16821 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U16822 ( .A1(n15265), .A2(n15267), .B1(n15242), .B2(n15264), .ZN(
        P1_U3471) );
  AOI211_X1 U16823 ( .C1(n15255), .C2(n15245), .A(n15244), .B(n15243), .ZN(
        n15246) );
  OAI21_X1 U16824 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15249) );
  AOI21_X1 U16825 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15268) );
  AOI22_X1 U16826 ( .A1(n15265), .A2(n15268), .B1(n9388), .B2(n15264), .ZN(
        P1_U3474) );
  AOI211_X1 U16827 ( .C1(n15255), .C2(n15254), .A(n15253), .B(n15252), .ZN(
        n15269) );
  INV_X1 U16828 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15256) );
  AOI22_X1 U16829 ( .A1(n15265), .A2(n15269), .B1(n15256), .B2(n15264), .ZN(
        P1_U3477) );
  OAI211_X1 U16830 ( .C1(n15260), .C2(n15259), .A(n15258), .B(n15257), .ZN(
        n15261) );
  AOI21_X1 U16831 ( .B1(n15263), .B2(n15262), .A(n15261), .ZN(n15271) );
  AOI22_X1 U16832 ( .A1(n15265), .A2(n15271), .B1(n9421), .B2(n15264), .ZN(
        P1_U3480) );
  AOI22_X1 U16833 ( .A1(n15272), .A2(n15266), .B1(n10249), .B2(n15270), .ZN(
        P1_U3531) );
  AOI22_X1 U16834 ( .A1(n15272), .A2(n15267), .B1(n10252), .B2(n15270), .ZN(
        P1_U3532) );
  AOI22_X1 U16835 ( .A1(n15272), .A2(n15268), .B1(n10244), .B2(n15270), .ZN(
        P1_U3533) );
  AOI22_X1 U16836 ( .A1(n15272), .A2(n15269), .B1(n10314), .B2(n15270), .ZN(
        P1_U3534) );
  AOI22_X1 U16837 ( .A1(n15272), .A2(n15271), .B1(n9425), .B2(n15270), .ZN(
        P1_U3535) );
  NOR2_X1 U16838 ( .A1(n15273), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16839 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15289) );
  INV_X1 U16840 ( .A(n15274), .ZN(n15282) );
  INV_X1 U16841 ( .A(n15275), .ZN(n15280) );
  NOR3_X1 U16842 ( .A1(n15278), .A2(n15277), .A3(n15276), .ZN(n15279) );
  NOR3_X1 U16843 ( .A1(n15300), .A2(n15280), .A3(n15279), .ZN(n15281) );
  AOI211_X1 U16844 ( .C1(n15305), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        n15288) );
  OAI211_X1 U16845 ( .C1(n15286), .C2(n15285), .A(n15318), .B(n15284), .ZN(
        n15287) );
  OAI211_X1 U16846 ( .C1(n15322), .C2(n15289), .A(n15288), .B(n15287), .ZN(
        P2_U3218) );
  INV_X1 U16847 ( .A(n15290), .ZN(n15292) );
  NAND3_X1 U16848 ( .A1(n15293), .A2(n15292), .A3(n15291), .ZN(n15295) );
  AOI21_X1 U16849 ( .B1(n15296), .B2(n15295), .A(n15294), .ZN(n15303) );
  AOI21_X1 U16850 ( .B1(n15299), .B2(n15298), .A(n15297), .ZN(n15301) );
  NOR2_X1 U16851 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  AOI211_X1 U16852 ( .C1(n15305), .C2(n15304), .A(n15303), .B(n15302), .ZN(
        n15307) );
  NAND2_X1 U16853 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15306)
         );
  OAI211_X1 U16854 ( .C1(n15308), .C2(n15322), .A(n15307), .B(n15306), .ZN(
        P2_U3226) );
  XOR2_X1 U16855 ( .A(n15310), .B(n15309), .Z(n15316) );
  OAI21_X1 U16856 ( .B1(n15313), .B2(n15312), .A(n15311), .ZN(n15314) );
  AOI21_X1 U16857 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(n15321) );
  XOR2_X1 U16858 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n15317), .Z(n15319) );
  NAND2_X1 U16859 ( .A1(n15319), .A2(n15318), .ZN(n15320) );
  OAI211_X1 U16860 ( .C1(n15322), .C2(n7086), .A(n15321), .B(n15320), .ZN(
        P2_U3228) );
  INV_X1 U16861 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15324) );
  NOR2_X1 U16862 ( .A1(n15354), .A2(n15324), .ZN(P2_U3266) );
  INV_X1 U16863 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15325) );
  NOR2_X1 U16864 ( .A1(n15354), .A2(n15325), .ZN(P2_U3267) );
  INV_X1 U16865 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15326) );
  NOR2_X1 U16866 ( .A1(n15354), .A2(n15326), .ZN(P2_U3268) );
  INV_X1 U16867 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15327) );
  NOR2_X1 U16868 ( .A1(n15354), .A2(n15327), .ZN(P2_U3269) );
  INV_X1 U16869 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15328) );
  NOR2_X1 U16870 ( .A1(n15338), .A2(n15328), .ZN(P2_U3270) );
  INV_X1 U16871 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15329) );
  NOR2_X1 U16872 ( .A1(n15338), .A2(n15329), .ZN(P2_U3271) );
  INV_X1 U16873 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15330) );
  NOR2_X1 U16874 ( .A1(n15338), .A2(n15330), .ZN(P2_U3272) );
  INV_X1 U16875 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U16876 ( .A1(n15338), .A2(n15331), .ZN(P2_U3273) );
  INV_X1 U16877 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U16878 ( .A1(n15338), .A2(n15332), .ZN(P2_U3274) );
  INV_X1 U16879 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15333) );
  NOR2_X1 U16880 ( .A1(n15338), .A2(n15333), .ZN(P2_U3275) );
  INV_X1 U16881 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U16882 ( .A1(n15338), .A2(n15334), .ZN(P2_U3276) );
  INV_X1 U16883 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16884 ( .A1(n15338), .A2(n15335), .ZN(P2_U3277) );
  INV_X1 U16885 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U16886 ( .A1(n15338), .A2(n15336), .ZN(P2_U3278) );
  INV_X1 U16887 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U16888 ( .A1(n15338), .A2(n15337), .ZN(P2_U3279) );
  INV_X1 U16889 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15339) );
  NOR2_X1 U16890 ( .A1(n15354), .A2(n15339), .ZN(P2_U3280) );
  INV_X1 U16891 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U16892 ( .A1(n15354), .A2(n15340), .ZN(P2_U3281) );
  INV_X1 U16893 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U16894 ( .A1(n15354), .A2(n15341), .ZN(P2_U3282) );
  INV_X1 U16895 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U16896 ( .A1(n15354), .A2(n15342), .ZN(P2_U3283) );
  INV_X1 U16897 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U16898 ( .A1(n15354), .A2(n15343), .ZN(P2_U3284) );
  INV_X1 U16899 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15344) );
  NOR2_X1 U16900 ( .A1(n15354), .A2(n15344), .ZN(P2_U3285) );
  INV_X1 U16901 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15508) );
  NOR2_X1 U16902 ( .A1(n15354), .A2(n15508), .ZN(P2_U3286) );
  INV_X1 U16903 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15345) );
  NOR2_X1 U16904 ( .A1(n15354), .A2(n15345), .ZN(P2_U3287) );
  INV_X1 U16905 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15346) );
  NOR2_X1 U16906 ( .A1(n15354), .A2(n15346), .ZN(P2_U3288) );
  INV_X1 U16907 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U16908 ( .A1(n15354), .A2(n15347), .ZN(P2_U3289) );
  INV_X1 U16909 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15557) );
  NOR2_X1 U16910 ( .A1(n15354), .A2(n15557), .ZN(P2_U3290) );
  INV_X1 U16911 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U16912 ( .A1(n15354), .A2(n15348), .ZN(P2_U3291) );
  INV_X1 U16913 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U16914 ( .A1(n15354), .A2(n15349), .ZN(P2_U3292) );
  INV_X1 U16915 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15350) );
  NOR2_X1 U16916 ( .A1(n15354), .A2(n15350), .ZN(P2_U3293) );
  INV_X1 U16917 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15351) );
  NOR2_X1 U16918 ( .A1(n15354), .A2(n15351), .ZN(P2_U3294) );
  INV_X1 U16919 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15352) );
  NOR2_X1 U16920 ( .A1(n15354), .A2(n15352), .ZN(P2_U3295) );
  OAI22_X1 U16921 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n15354), .B1(n15356), .B2(
        n15353), .ZN(n15355) );
  INV_X1 U16922 ( .A(n15355), .ZN(P2_U3416) );
  AOI22_X1 U16923 ( .A1(n15359), .A2(n15358), .B1(n15357), .B2(n15356), .ZN(
        P2_U3417) );
  AOI21_X1 U16924 ( .B1(n15377), .B2(n15361), .A(n15360), .ZN(n15362) );
  OAI211_X1 U16925 ( .C1(n15381), .C2(n15364), .A(n15363), .B(n15362), .ZN(
        n15365) );
  INV_X1 U16926 ( .A(n15365), .ZN(n15385) );
  INV_X1 U16927 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U16928 ( .A1(n15384), .A2(n15385), .B1(n15366), .B2(n6771), .ZN(
        P2_U3436) );
  AOI21_X1 U16929 ( .B1(n15377), .B2(n15368), .A(n15367), .ZN(n15369) );
  OAI211_X1 U16930 ( .C1(n15372), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        n15373) );
  INV_X1 U16931 ( .A(n15373), .ZN(n15386) );
  INV_X1 U16932 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15374) );
  AOI22_X1 U16933 ( .A1(n15384), .A2(n15386), .B1(n15374), .B2(n6771), .ZN(
        P2_U3442) );
  AOI21_X1 U16934 ( .B1(n15377), .B2(n15376), .A(n15375), .ZN(n15378) );
  OAI211_X1 U16935 ( .C1(n15381), .C2(n15380), .A(n15379), .B(n15378), .ZN(
        n15382) );
  INV_X1 U16936 ( .A(n15382), .ZN(n15389) );
  INV_X1 U16937 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15383) );
  AOI22_X1 U16938 ( .A1(n15384), .A2(n15389), .B1(n15383), .B2(n6771), .ZN(
        P2_U3451) );
  AOI22_X1 U16939 ( .A1(n15390), .A2(n15385), .B1(n10188), .B2(n15387), .ZN(
        P2_U3501) );
  AOI22_X1 U16940 ( .A1(n15390), .A2(n15386), .B1(n10190), .B2(n15387), .ZN(
        P2_U3503) );
  AOI22_X1 U16941 ( .A1(n15390), .A2(n15389), .B1(n15388), .B2(n15387), .ZN(
        P2_U3506) );
  NOR2_X1 U16942 ( .A1(P3_U3897), .A2(n15391), .ZN(P3_U3150) );
  AOI211_X1 U16943 ( .C1(n15395), .C2(n15394), .A(n15393), .B(n15392), .ZN(
        n15432) );
  INV_X1 U16944 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U16945 ( .A1(n15431), .A2(n15432), .B1(n15396), .B2(n15429), .ZN(
        P3_U3393) );
  INV_X1 U16946 ( .A(n15425), .ZN(n15398) );
  OAI21_X1 U16947 ( .B1(n15399), .B2(n15398), .A(n15397), .ZN(n15400) );
  NOR2_X1 U16948 ( .A1(n15401), .A2(n15400), .ZN(n15433) );
  INV_X1 U16949 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U16950 ( .A1(n15431), .A2(n15433), .B1(n15402), .B2(n15429), .ZN(
        P3_U3396) );
  AOI22_X1 U16951 ( .A1(n15404), .A2(n15425), .B1(n15423), .B2(n15403), .ZN(
        n15405) );
  AND2_X1 U16952 ( .A1(n15406), .A2(n15405), .ZN(n15434) );
  INV_X1 U16953 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U16954 ( .A1(n15431), .A2(n15434), .B1(n15407), .B2(n15429), .ZN(
        P3_U3402) );
  AOI22_X1 U16955 ( .A1(n15409), .A2(n15425), .B1(n15423), .B2(n15408), .ZN(
        n15410) );
  AND2_X1 U16956 ( .A1(n15411), .A2(n15410), .ZN(n15436) );
  INV_X1 U16957 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15412) );
  AOI22_X1 U16958 ( .A1(n15431), .A2(n15436), .B1(n15412), .B2(n15429), .ZN(
        P3_U3405) );
  AOI22_X1 U16959 ( .A1(n15414), .A2(n15425), .B1(n15423), .B2(n15413), .ZN(
        n15415) );
  AND2_X1 U16960 ( .A1(n15416), .A2(n15415), .ZN(n15437) );
  INV_X1 U16961 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U16962 ( .A1(n15431), .A2(n15437), .B1(n15417), .B2(n15429), .ZN(
        P3_U3408) );
  NOR2_X1 U16963 ( .A1(n15419), .A2(n15418), .ZN(n15421) );
  AOI211_X1 U16964 ( .C1(n15425), .C2(n15422), .A(n15421), .B(n15420), .ZN(
        n15439) );
  INV_X1 U16965 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U16966 ( .A1(n15431), .A2(n15439), .B1(n15513), .B2(n15429), .ZN(
        P3_U3411) );
  AOI22_X1 U16967 ( .A1(n15426), .A2(n15425), .B1(n15424), .B2(n15423), .ZN(
        n15427) );
  AND2_X1 U16968 ( .A1(n15428), .A2(n15427), .ZN(n15441) );
  INV_X1 U16969 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U16970 ( .A1(n15431), .A2(n15441), .B1(n15430), .B2(n15429), .ZN(
        P3_U3414) );
  AOI22_X1 U16971 ( .A1(n15589), .A2(n15432), .B1(n10518), .B2(n15440), .ZN(
        P3_U3460) );
  AOI22_X1 U16972 ( .A1(n15589), .A2(n15433), .B1(n10517), .B2(n15440), .ZN(
        P3_U3461) );
  AOI22_X1 U16973 ( .A1(n15589), .A2(n15434), .B1(n10610), .B2(n15440), .ZN(
        P3_U3463) );
  INV_X1 U16974 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15435) );
  AOI22_X1 U16975 ( .A1(n15589), .A2(n15436), .B1(n15435), .B2(n15440), .ZN(
        P3_U3464) );
  AOI22_X1 U16976 ( .A1(n15589), .A2(n15437), .B1(n10629), .B2(n15440), .ZN(
        P3_U3465) );
  INV_X1 U16977 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U16978 ( .A1(n15589), .A2(n15439), .B1(n15438), .B2(n15440), .ZN(
        P3_U3466) );
  AOI22_X1 U16979 ( .A1(n15589), .A2(n15441), .B1(n10869), .B2(n15440), .ZN(
        P3_U3467) );
  NOR4_X1 U16980 ( .A1(P3_REG0_REG_7__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(P1_WR_REG_SCAN_IN), .A4(n15508), .ZN(n15445) );
  NOR4_X1 U16981 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P1_REG1_REG_27__SCAN_IN), 
        .A3(P1_REG2_REG_7__SCAN_IN), .A4(n15545), .ZN(n15444) );
  NOR4_X1 U16982 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .A3(P2_ADDR_REG_11__SCAN_IN), .A4(P3_DATAO_REG_10__SCAN_IN), .ZN(
        n15443) );
  INV_X1 U16983 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15533) );
  INV_X1 U16984 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n15535) );
  INV_X1 U16985 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15526) );
  NOR4_X1 U16986 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n15533), .A3(n15535), .A4(
        n15526), .ZN(n15442) );
  NAND4_X1 U16987 ( .A1(n15445), .A2(n15444), .A3(n15443), .A4(n15442), .ZN(
        n15467) );
  NAND4_X1 U16988 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(P3_REG1_REG_16__SCAN_IN), 
        .A3(P1_IR_REG_4__SCAN_IN), .A4(n15569), .ZN(n15466) );
  NAND4_X1 U16989 ( .A1(n15448), .A2(n15447), .A3(n15446), .A4(
        P3_REG1_REG_25__SCAN_IN), .ZN(n15451) );
  NOR3_X1 U16990 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .A3(P1_REG2_REG_28__SCAN_IN), .ZN(n15449) );
  NAND4_X1 U16991 ( .A1(n15532), .A2(P1_DATAO_REG_10__SCAN_IN), .A3(
        P1_DATAO_REG_11__SCAN_IN), .A4(n15449), .ZN(n15450) );
  INV_X1 U16992 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15570) );
  OR4_X1 U16993 ( .A1(n15451), .A2(n15450), .A3(n15570), .A4(n15557), .ZN(
        n15465) );
  NOR4_X1 U16994 ( .A1(P3_REG2_REG_7__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), 
        .A3(n15542), .A4(n15475), .ZN(n15463) );
  NOR4_X1 U16995 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        n7417), .A4(n15472), .ZN(n15462) );
  NAND4_X1 U16996 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), 
        .A3(P1_D_REG_1__SCAN_IN), .A4(n15452), .ZN(n15453) );
  NOR4_X1 U16997 ( .A1(n15454), .A2(n15498), .A3(n10031), .A4(n15453), .ZN(
        n15461) );
  NAND4_X1 U16998 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_ADDR_REG_12__SCAN_IN), .A4(n15512), .ZN(n15459) );
  INV_X1 U16999 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n15457) );
  NAND4_X1 U17000 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), 
        .A3(P3_ADDR_REG_17__SCAN_IN), .A4(n7526), .ZN(n15456) );
  NAND4_X1 U17001 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(SI_11_), .A3(
        P2_REG2_REG_7__SCAN_IN), .A4(P1_IR_REG_3__SCAN_IN), .ZN(n15455) );
  OR4_X1 U17002 ( .A1(n15457), .A2(P2_REG3_REG_9__SCAN_IN), .A3(n15456), .A4(
        n15455), .ZN(n15458) );
  INV_X1 U17003 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15485) );
  NOR4_X1 U17004 ( .A1(n15459), .A2(n15458), .A3(P1_REG0_REG_16__SCAN_IN), 
        .A4(n15485), .ZN(n15460) );
  NAND4_X1 U17005 ( .A1(n15463), .A2(n15462), .A3(n15461), .A4(n15460), .ZN(
        n15464) );
  NOR4_X1 U17006 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15586) );
  AOI22_X1 U17007 ( .A1(P1_U3086), .A2(keyinput5), .B1(keyinput34), .B2(n15469), .ZN(n15468) );
  OAI221_X1 U17008 ( .B1(P1_U3086), .B2(keyinput5), .C1(n15469), .C2(
        keyinput34), .A(n15468), .ZN(n15481) );
  AOI22_X1 U17009 ( .A1(n15472), .A2(keyinput26), .B1(n15471), .B2(keyinput47), 
        .ZN(n15470) );
  OAI221_X1 U17010 ( .B1(n15472), .B2(keyinput26), .C1(n15471), .C2(keyinput47), .A(n15470), .ZN(n15480) );
  AOI22_X1 U17011 ( .A1(n15475), .A2(keyinput62), .B1(n15474), .B2(keyinput8), 
        .ZN(n15473) );
  OAI221_X1 U17012 ( .B1(n15475), .B2(keyinput62), .C1(n15474), .C2(keyinput8), 
        .A(n15473), .ZN(n15479) );
  XNOR2_X1 U17013 ( .A(P3_REG2_REG_9__SCAN_IN), .B(keyinput1), .ZN(n15477) );
  XNOR2_X1 U17014 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput49), .ZN(n15476) );
  NAND2_X1 U17015 ( .A1(n15477), .A2(n15476), .ZN(n15478) );
  NOR4_X1 U17016 ( .A1(n15481), .A2(n15480), .A3(n15479), .A4(n15478), .ZN(
        n15524) );
  AOI22_X1 U17017 ( .A1(n15483), .A2(keyinput56), .B1(keyinput33), .B2(n10119), 
        .ZN(n15482) );
  OAI221_X1 U17018 ( .B1(n15483), .B2(keyinput56), .C1(n10119), .C2(keyinput33), .A(n15482), .ZN(n15493) );
  AOI22_X1 U17019 ( .A1(n15486), .A2(keyinput16), .B1(n15485), .B2(keyinput31), 
        .ZN(n15484) );
  OAI221_X1 U17020 ( .B1(n15486), .B2(keyinput16), .C1(n15485), .C2(keyinput31), .A(n15484), .ZN(n15492) );
  XOR2_X1 U17021 ( .A(n15457), .B(keyinput58), .Z(n15490) );
  XNOR2_X1 U17022 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput40), .ZN(n15489) );
  XNOR2_X1 U17023 ( .A(P3_REG1_REG_12__SCAN_IN), .B(keyinput17), .ZN(n15488)
         );
  XNOR2_X1 U17024 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput15), .ZN(n15487) );
  NAND4_X1 U17025 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15491) );
  NOR3_X1 U17026 ( .A1(n15493), .A2(n15492), .A3(n15491), .ZN(n15523) );
  AOI22_X1 U17027 ( .A1(n15495), .A2(keyinput48), .B1(n7526), .B2(keyinput28), 
        .ZN(n15494) );
  OAI221_X1 U17028 ( .B1(n15495), .B2(keyinput48), .C1(n7526), .C2(keyinput28), 
        .A(n15494), .ZN(n15505) );
  AOI22_X1 U17029 ( .A1(n15498), .A2(keyinput19), .B1(n15497), .B2(keyinput11), 
        .ZN(n15496) );
  OAI221_X1 U17030 ( .B1(n15498), .B2(keyinput19), .C1(n15497), .C2(keyinput11), .A(n15496), .ZN(n15504) );
  XNOR2_X1 U17031 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput29), .ZN(n15502) );
  XNOR2_X1 U17032 ( .A(P3_IR_REG_25__SCAN_IN), .B(keyinput52), .ZN(n15501) );
  XNOR2_X1 U17033 ( .A(SI_11_), .B(keyinput44), .ZN(n15500) );
  XNOR2_X1 U17034 ( .A(keyinput45), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n15499) );
  NAND4_X1 U17035 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15503) );
  NOR3_X1 U17036 ( .A1(n15505), .A2(n15504), .A3(n15503), .ZN(n15522) );
  INV_X1 U17037 ( .A(P1_WR_REG_SCAN_IN), .ZN(n15507) );
  AOI22_X1 U17038 ( .A1(n15508), .A2(keyinput55), .B1(keyinput9), .B2(n15507), 
        .ZN(n15506) );
  OAI221_X1 U17039 ( .B1(n15508), .B2(keyinput55), .C1(n15507), .C2(keyinput9), 
        .A(n15506), .ZN(n15520) );
  AOI22_X1 U17040 ( .A1(n15511), .A2(keyinput18), .B1(keyinput10), .B2(n15510), 
        .ZN(n15509) );
  OAI221_X1 U17041 ( .B1(n15511), .B2(keyinput18), .C1(n15510), .C2(keyinput10), .A(n15509), .ZN(n15519) );
  XNOR2_X1 U17042 ( .A(n15512), .B(keyinput20), .ZN(n15518) );
  XOR2_X1 U17043 ( .A(n15513), .B(keyinput41), .Z(n15516) );
  XNOR2_X1 U17044 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput38), .ZN(n15515) );
  XNOR2_X1 U17045 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput54), .ZN(n15514) );
  NAND3_X1 U17046 ( .A1(n15516), .A2(n15515), .A3(n15514), .ZN(n15517) );
  NOR4_X1 U17047 ( .A1(n15520), .A2(n15519), .A3(n15518), .A4(n15517), .ZN(
        n15521) );
  NAND4_X1 U17048 ( .A1(n15524), .A2(n15523), .A3(n15522), .A4(n15521), .ZN(
        n15585) );
  AOI22_X1 U17049 ( .A1(n15527), .A2(keyinput63), .B1(keyinput46), .B2(n15526), 
        .ZN(n15525) );
  OAI221_X1 U17050 ( .B1(n15527), .B2(keyinput63), .C1(n15526), .C2(keyinput46), .A(n15525), .ZN(n15540) );
  AOI22_X1 U17051 ( .A1(n15530), .A2(keyinput7), .B1(n15529), .B2(keyinput6), 
        .ZN(n15528) );
  OAI221_X1 U17052 ( .B1(n15530), .B2(keyinput7), .C1(n15529), .C2(keyinput6), 
        .A(n15528), .ZN(n15539) );
  AOI22_X1 U17053 ( .A1(n15533), .A2(keyinput42), .B1(n15532), .B2(keyinput4), 
        .ZN(n15531) );
  OAI221_X1 U17054 ( .B1(n15533), .B2(keyinput42), .C1(n15532), .C2(keyinput4), 
        .A(n15531), .ZN(n15538) );
  INV_X1 U17055 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U17056 ( .A1(n15536), .A2(keyinput3), .B1(keyinput53), .B2(n15535), 
        .ZN(n15534) );
  OAI221_X1 U17057 ( .B1(n15536), .B2(keyinput3), .C1(n15535), .C2(keyinput53), 
        .A(n15534), .ZN(n15537) );
  NOR4_X1 U17058 ( .A1(n15540), .A2(n15539), .A3(n15538), .A4(n15537), .ZN(
        n15583) );
  AOI22_X1 U17059 ( .A1(n15543), .A2(keyinput43), .B1(keyinput0), .B2(n15542), 
        .ZN(n15541) );
  OAI221_X1 U17060 ( .B1(n15543), .B2(keyinput43), .C1(n15542), .C2(keyinput0), 
        .A(n15541), .ZN(n15555) );
  INV_X1 U17061 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U17062 ( .A1(n15546), .A2(keyinput21), .B1(n15545), .B2(keyinput57), 
        .ZN(n15544) );
  OAI221_X1 U17063 ( .B1(n15546), .B2(keyinput21), .C1(n15545), .C2(keyinput57), .A(n15544), .ZN(n15554) );
  AOI22_X1 U17064 ( .A1(n15549), .A2(keyinput12), .B1(n15548), .B2(keyinput23), 
        .ZN(n15547) );
  OAI221_X1 U17065 ( .B1(n15549), .B2(keyinput12), .C1(n15548), .C2(keyinput23), .A(n15547), .ZN(n15553) );
  AOI22_X1 U17066 ( .A1(n10322), .A2(keyinput60), .B1(n15551), .B2(keyinput36), 
        .ZN(n15550) );
  OAI221_X1 U17067 ( .B1(n10322), .B2(keyinput60), .C1(n15551), .C2(keyinput36), .A(n15550), .ZN(n15552) );
  NOR4_X1 U17068 ( .A1(n15555), .A2(n15554), .A3(n15553), .A4(n15552), .ZN(
        n15582) );
  AOI22_X1 U17069 ( .A1(n10031), .A2(keyinput32), .B1(n15557), .B2(keyinput25), 
        .ZN(n15556) );
  OAI221_X1 U17070 ( .B1(n10031), .B2(keyinput32), .C1(n15557), .C2(keyinput25), .A(n15556), .ZN(n15567) );
  INV_X1 U17071 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15560) );
  AOI22_X1 U17072 ( .A1(n15560), .A2(keyinput37), .B1(n15559), .B2(keyinput2), 
        .ZN(n15558) );
  OAI221_X1 U17073 ( .B1(n15560), .B2(keyinput37), .C1(n15559), .C2(keyinput2), 
        .A(n15558), .ZN(n15566) );
  XNOR2_X1 U17074 ( .A(SI_20_), .B(keyinput50), .ZN(n15564) );
  XNOR2_X1 U17075 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput39), .ZN(n15563)
         );
  XNOR2_X1 U17076 ( .A(P3_REG1_REG_25__SCAN_IN), .B(keyinput30), .ZN(n15562)
         );
  XNOR2_X1 U17077 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput51), .ZN(n15561) );
  NAND4_X1 U17078 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15565) );
  NOR3_X1 U17079 ( .A1(n15567), .A2(n15566), .A3(n15565), .ZN(n15581) );
  AOI22_X1 U17080 ( .A1(n15570), .A2(keyinput61), .B1(n15569), .B2(keyinput24), 
        .ZN(n15568) );
  OAI221_X1 U17081 ( .B1(n15570), .B2(keyinput61), .C1(n15569), .C2(keyinput24), .A(n15568), .ZN(n15579) );
  XNOR2_X1 U17082 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput22), .ZN(n15574)
         );
  XNOR2_X1 U17083 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(keyinput13), .ZN(n15573)
         );
  XNOR2_X1 U17084 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput14), .ZN(n15572) );
  XNOR2_X1 U17085 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput59), .ZN(n15571) );
  NAND4_X1 U17086 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15578) );
  XNOR2_X1 U17087 ( .A(n15575), .B(keyinput27), .ZN(n15577) );
  XNOR2_X1 U17088 ( .A(keyinput35), .B(n9180), .ZN(n15576) );
  NOR4_X1 U17089 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15580) );
  NAND4_X1 U17090 ( .A1(n15583), .A2(n15582), .A3(n15581), .A4(n15580), .ZN(
        n15584) );
  NOR3_X1 U17091 ( .A1(n15586), .A2(n15585), .A3(n15584), .ZN(n15591) );
  NAND2_X1 U17092 ( .A1(n15587), .A2(n15589), .ZN(n15588) );
  OAI21_X1 U17093 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n15589), .A(n15588), .ZN(
        n15590) );
  XNOR2_X1 U17094 ( .A(n15591), .B(n15590), .ZN(P3_U3462) );
  CLKBUF_X2 U7168 ( .A(n13215), .Z(n13372) );
  CLKBUF_X2 U7163 ( .A(n12298), .Z(n6401) );
  INV_X1 U7149 ( .A(n15429), .ZN(n15431) );
  OR2_X1 U7198 ( .A1(n12569), .A2(n6620), .ZN(n6999) );
  AND3_X1 U7212 ( .A1(n6400), .A2(n7734), .A3(n6531), .ZN(n7218) );
  CLKBUF_X1 U7216 ( .A(n8062), .Z(n8389) );
  CLKBUF_X2 U7228 ( .A(n8029), .Z(n10431) );
  CLKBUF_X1 U7248 ( .A(n8816), .Z(n6418) );
  CLKBUF_X2 U7269 ( .A(n9970), .Z(n6406) );
  CLKBUF_X1 U7592 ( .A(n12055), .Z(n12056) );
  CLKBUF_X1 U9995 ( .A(n11722), .Z(n6403) );
  AOI211_X1 U14447 ( .C1(n14907), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14709) );
endmodule

