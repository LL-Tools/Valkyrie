

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4265, n4266, n4267, n4268, n4271, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054;

  INV_X4 U4771 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4772 ( .A(n6241), .ZN(n8529) );
  INV_X1 U4773 ( .A(n5160), .ZN(n7739) );
  INV_X2 U4774 ( .A(n9264), .ZN(n9045) );
  AND2_X1 U4775 ( .A1(n7930), .A2(n7747), .ZN(n7865) );
  CLKBUF_X1 U4776 ( .A(n5089), .Z(n5408) );
  INV_X1 U4777 ( .A(n7952), .ZN(n5744) );
  INV_X2 U4778 ( .A(n6094), .ZN(n5775) );
  INV_X4 U4779 ( .A(n4483), .ZN(n5759) );
  NAND2_X1 U4780 ( .A1(n4451), .A2(n5065), .ZN(n5075) );
  CLKBUF_X1 U4781 ( .A(n9536), .Z(n4265) );
  NOR2_X1 U4782 ( .A1(n6826), .A2(n9045), .ZN(n9536) );
  INV_X1 U4783 ( .A(n8919), .ZN(n8760) );
  INV_X1 U4784 ( .A(n5735), .ZN(n6239) );
  OR2_X1 U4785 ( .A1(n5999), .A2(n7659), .ZN(n6020) );
  CLKBUF_X2 U4786 ( .A(n5090), .Z(n5164) );
  OR2_X1 U4787 ( .A1(n5939), .A2(n5938), .ZN(n5944) );
  INV_X1 U4788 ( .A(n6897), .ZN(n9560) );
  INV_X1 U4789 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  BUF_X1 U4790 ( .A(n5048), .Z(n6337) );
  INV_X1 U4791 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5091) );
  OAI211_X1 U4792 ( .C1(n8497), .C2(n4314), .A(n4809), .B(n4807), .ZN(n8583)
         );
  NAND2_X1 U4793 ( .A1(n7959), .A2(n4530), .ZN(n5751) );
  OR2_X1 U4794 ( .A1(n5656), .A2(n5992), .ZN(n5658) );
  INV_X1 U4795 ( .A(n6328), .ZN(n8130) );
  NAND2_X2 U4797 ( .A1(n5487), .A2(n7062), .ZN(n7742) );
  INV_X2 U4798 ( .A(n4434), .ZN(n8236) );
  NOR2_X2 U4799 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5731) );
  XNOR2_X2 U4800 ( .A(n5706), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7934) );
  NAND2_X2 U4801 ( .A1(n9444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5706) );
  AOI21_X2 U4802 ( .B1(n5534), .B2(n7917), .A(n4855), .ZN(n5535) );
  AOI21_X2 U4803 ( .B1(n5469), .B2(n6494), .A(n4852), .ZN(n5534) );
  OAI211_X2 U4804 ( .C1(n4482), .C2(n6476), .A(n5764), .B(n5763), .ZN(n6897)
         );
  XNOR2_X2 U4805 ( .A(n5658), .B(n5657), .ZN(n8959) );
  NAND3_X1 U4806 ( .A1(n4792), .A2(n8054), .A3(n8299), .ZN(n8017) );
  OAI21_X1 U4807 ( .B1(n8764), .B2(n8815), .A(n8763), .ZN(n8775) );
  OAI21_X1 U4808 ( .B1(n8623), .B2(n6101), .A(n4396), .ZN(n4395) );
  INV_X1 U4809 ( .A(n8497), .ZN(n8498) );
  NAND2_X1 U4810 ( .A1(n7748), .A2(n7745), .ZN(n7881) );
  NAND2_X2 U4811 ( .A1(n5074), .A2(n5536), .ZN(n7748) );
  NAND2_X1 U4812 ( .A1(n8671), .A2(n8821), .ZN(n8784) );
  INV_X1 U4813 ( .A(n9566), .ZN(n8664) );
  INV_X1 U4814 ( .A(n6854), .ZN(n6941) );
  OR2_X1 U4815 ( .A1(n5965), .A2(n5964), .ZN(n5999) );
  INV_X1 U4816 ( .A(n5835), .ZN(n5780) );
  BUF_X1 U4817 ( .A(n5019), .Z(n4986) );
  AND4_X1 U4818 ( .A1(n4341), .A2(n4580), .A3(n4578), .A4(n4579), .ZN(n5454)
         );
  INV_X2 U4819 ( .A(n4877), .ZN(n4266) );
  OAI21_X1 U4820 ( .B1(n7705), .B2(n7704), .A(n7720), .ZN(n4639) );
  NOR2_X1 U4821 ( .A1(n6302), .A2(n6301), .ZN(n6311) );
  NAND2_X1 U4822 ( .A1(n8777), .A2(n4302), .ZN(n8922) );
  NAND2_X1 U4823 ( .A1(n4640), .A2(n7838), .ZN(n7982) );
  OAI21_X1 U4824 ( .B1(n8775), .B2(n9051), .A(n4398), .ZN(n4397) );
  NAND3_X1 U4825 ( .A1(n6153), .A2(n6154), .A3(n8513), .ZN(n8511) );
  NOR2_X1 U4826 ( .A1(n4385), .A2(n8592), .ZN(n4384) );
  NAND2_X1 U4827 ( .A1(n4572), .A2(n4571), .ZN(n9174) );
  NAND2_X1 U4828 ( .A1(n4393), .A2(n4799), .ZN(n6152) );
  AOI21_X1 U4829 ( .B1(n5507), .B2(n4630), .A(n4628), .ZN(n4627) );
  NAND2_X1 U4830 ( .A1(n4395), .A2(n4394), .ZN(n8523) );
  NAND2_X1 U4831 ( .A1(n8623), .A2(n6101), .ZN(n4394) );
  AND2_X1 U4832 ( .A1(n4382), .A2(n8591), .ZN(n4381) );
  INV_X1 U4833 ( .A(n8104), .ZN(n4787) );
  NAND2_X1 U4834 ( .A1(n6174), .A2(n8512), .ZN(n4382) );
  OAI22_X1 U4835 ( .A1(n7595), .A2(n4375), .B1(n4377), .B2(n6012), .ZN(n6048)
         );
  OAI21_X1 U4836 ( .B1(n5508), .B2(n4629), .A(n7822), .ZN(n4628) );
  NOR2_X1 U4837 ( .A1(n5508), .A2(n4631), .ZN(n4630) );
  INV_X1 U4838 ( .A(n8620), .ZN(n4396) );
  OR2_X1 U4839 ( .A1(n9233), .A2(n8939), .ZN(n6365) );
  OR2_X1 U4840 ( .A1(n6157), .A2(n8515), .ZN(n6177) );
  NAND2_X1 U4841 ( .A1(n5882), .A2(n5881), .ZN(n7206) );
  NAND2_X2 U4842 ( .A1(n6826), .A2(n9309), .ZN(n9287) );
  NAND2_X2 U4843 ( .A1(n8146), .A2(n9778), .ZN(n7758) );
  INV_X1 U4844 ( .A(n6687), .ZN(n8144) );
  INV_X1 U4845 ( .A(n6634), .ZN(n4267) );
  NAND2_X1 U4846 ( .A1(n8945), .A2(n8664), .ZN(n8826) );
  AND4_X1 U4847 ( .A1(n5096), .A2(n5095), .A3(n5094), .A4(n5093), .ZN(n5104)
         );
  OAI211_X1 U4848 ( .C1(n5853), .C2(n6475), .A(n5784), .B(n5783), .ZN(n6854)
         );
  OAI211_X1 U4849 ( .C1(n6337), .C2(n6597), .A(n5103), .B(n5102), .ZN(n6724)
         );
  NOR2_X1 U4850 ( .A1(n6351), .A2(n6922), .ZN(n6924) );
  AND2_X1 U4851 ( .A1(n5025), .A2(n8495), .ZN(n5090) );
  NAND4_X1 U4852 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(n5757)
         );
  AND2_X2 U4853 ( .A1(n8491), .A2(n8495), .ZN(n7721) );
  AND4_X1 U4854 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n6886)
         );
  OAI22_X1 U4855 ( .A1(n7737), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n5160), .B2(
        n6474), .ZN(n4450) );
  OR2_X1 U4856 ( .A1(n6389), .A2(n5687), .ZN(n6818) );
  AND2_X1 U4857 ( .A1(n5025), .A2(n5026), .ZN(n5092) );
  AND2_X1 U4858 ( .A1(n5670), .A2(n6261), .ZN(n8921) );
  XNOR2_X1 U4859 ( .A(n5055), .B(n5054), .ZN(n5487) );
  INV_X2 U4860 ( .A(n4482), .ZN(n5758) );
  NAND2_X1 U4861 ( .A1(n5683), .A2(n6260), .ZN(n6441) );
  OR2_X1 U4862 ( .A1(n5751), .A2(n5736), .ZN(n5738) );
  INV_X2 U4863 ( .A(n5751), .ZN(n5773) );
  OR2_X1 U4864 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U4865 ( .A1(n6265), .A2(n8893), .ZN(n6389) );
  CLKBUF_X2 U4866 ( .A(n5780), .Z(n4271) );
  CLKBUF_X1 U4867 ( .A(n4482), .Z(n5853) );
  INV_X1 U4868 ( .A(n5025), .ZN(n8491) );
  AND2_X1 U4869 ( .A1(n5439), .A2(n5438), .ZN(n7747) );
  NAND2_X2 U4870 ( .A1(n4530), .A2(n5707), .ZN(n8771) );
  XNOR2_X1 U4871 ( .A(n5435), .B(n5441), .ZN(n7062) );
  NAND2_X1 U4872 ( .A1(n5459), .A2(n5460), .ZN(n7513) );
  MUX2_X1 U4873 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5461), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5462) );
  NAND2_X1 U4874 ( .A1(n5677), .A2(n5681), .ZN(n7591) );
  XNOR2_X1 U4875 ( .A(n5675), .B(n5674), .ZN(n8893) );
  NAND2_X2 U4876 ( .A1(n4987), .A2(n4986), .ZN(n7928) );
  NAND2_X1 U4877 ( .A1(n5655), .A2(n5701), .ZN(n6280) );
  MUX2_X1 U4878 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5676), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5677) );
  NOR2_X1 U4879 ( .A1(n5221), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5235) );
  INV_X2 U4880 ( .A(n8487), .ZN(n8494) );
  NAND2_X1 U4881 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NAND2_X2 U4882 ( .A1(n7731), .A2(P1_U3086), .ZN(n7960) );
  NAND2_X1 U4883 ( .A1(n5701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5702) );
  OR2_X1 U4884 ( .A1(n5678), .A2(n4830), .ZN(n5681) );
  NAND2_X1 U4885 ( .A1(n5454), .A2(n4992), .ZN(n5463) );
  AND2_X1 U4886 ( .A1(n5661), .A2(n4573), .ZN(n5705) );
  NAND2_X1 U4887 ( .A1(n4670), .A2(n4669), .ZN(n4877) );
  AND4_X1 U4888 ( .A1(n4317), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n5650)
         );
  AND2_X1 U4889 ( .A1(n5434), .A2(n4976), .ZN(n5432) );
  AND4_X1 U4890 ( .A1(n5644), .A2(n5643), .A3(n4828), .A4(n4827), .ZN(n4826)
         );
  AND4_X1 U4891 ( .A1(n5993), .A2(n5990), .A3(n5645), .A4(n6031), .ZN(n5646)
         );
  NOR2_X1 U4892 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4827) );
  INV_X2 U4893 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U4894 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4828) );
  INV_X1 U4895 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5990) );
  INV_X1 U4896 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9050) );
  INV_X1 U4897 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10005) );
  INV_X1 U4898 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U4899 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4966) );
  NOR2_X1 U4900 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4967) );
  NAND2_X1 U4901 ( .A1(n8511), .A2(n4384), .ZN(n4383) );
  AND2_X2 U4902 ( .A1(n7934), .A2(n7959), .ZN(n6094) );
  NAND2_X2 U4903 ( .A1(n5734), .A2(n4479), .ZN(n7952) );
  AND2_X1 U4904 ( .A1(n8491), .A2(n8495), .ZN(n4268) );
  NAND2_X2 U4905 ( .A1(n9145), .A2(n9144), .ZN(n9130) );
  OAI22_X2 U4906 ( .A1(n9180), .A2(n4334), .B1(n4528), .B2(n4281), .ZN(n9145)
         );
  OR2_X2 U4907 ( .A1(n8321), .A2(n4715), .ZN(n4714) );
  OAI222_X1 U4908 ( .A1(n7964), .A2(n10020), .B1(P1_U3086), .B2(n8959), .C1(
        n7960), .C2(n7667), .ZN(P1_U3328) );
  OAI21_X2 U4909 ( .B1(n8436), .B2(n8133), .A(n5363), .ZN(n8264) );
  XNOR2_X1 U4910 ( .A(n5743), .B(n5744), .ZN(n6397) );
  NAND2_X1 U4911 ( .A1(n4526), .A2(n4524), .ZN(n4898) );
  AND2_X1 U4912 ( .A1(n4654), .A2(n4525), .ZN(n4524) );
  INV_X1 U4913 ( .A(n5173), .ZN(n4525) );
  OR2_X1 U4914 ( .A1(n8648), .A2(n9171), .ZN(n4400) );
  NAND2_X1 U4915 ( .A1(n8651), .A2(n9171), .ZN(n4401) );
  NAND2_X1 U4916 ( .A1(n8015), .A2(n8122), .ZN(n4747) );
  NAND2_X1 U4917 ( .A1(n8531), .A2(n6241), .ZN(n4796) );
  AOI21_X1 U4918 ( .B1(n4543), .B2(n4545), .A(n4315), .ZN(n4542) );
  INV_X1 U4919 ( .A(n4547), .ZN(n4543) );
  NAND2_X1 U4920 ( .A1(n6051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U4921 ( .A(n4911), .B(SI_12_), .ZN(n5219) );
  NOR2_X1 U4922 ( .A1(n4656), .A2(n4653), .ZN(n4527) );
  INV_X1 U4923 ( .A(n5140), .ZN(n4653) );
  INV_X1 U4924 ( .A(n5159), .ZN(n4656) );
  INV_X1 U4925 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U4926 ( .A1(n5835), .A2(n4266), .ZN(n4483) );
  NAND2_X1 U4927 ( .A1(n4727), .A2(n4305), .ZN(n4419) );
  OR2_X1 U4928 ( .A1(n7808), .A2(n8347), .ZN(n4418) );
  NAND2_X1 U4929 ( .A1(n4598), .A2(n4412), .ZN(n4411) );
  AND2_X1 U4930 ( .A1(n4596), .A2(n4295), .ZN(n4412) );
  OR2_X1 U4931 ( .A1(n7789), .A2(n7865), .ZN(n4598) );
  AOI21_X1 U4932 ( .B1(n4597), .B2(n7865), .A(n7897), .ZN(n4596) );
  NAND2_X1 U4933 ( .A1(n4295), .A2(n4594), .ZN(n4410) );
  NAND2_X1 U4934 ( .A1(n4595), .A2(n4705), .ZN(n4594) );
  INV_X1 U4935 ( .A(n7795), .ZN(n4595) );
  INV_X1 U4936 ( .A(n4505), .ZN(n4504) );
  OAI21_X1 U4937 ( .B1(n9142), .B2(n4304), .A(n8748), .ZN(n4505) );
  INV_X1 U4938 ( .A(n5280), .ZN(n4926) );
  NAND2_X1 U4939 ( .A1(n4747), .A2(n4300), .ZN(n4743) );
  INV_X1 U4940 ( .A(n7866), .ZN(n4440) );
  NAND2_X1 U4941 ( .A1(n7855), .A2(n7854), .ZN(n4439) );
  AND2_X1 U4942 ( .A1(n4638), .A2(n4637), .ZN(n7926) );
  OAI21_X1 U4943 ( .B1(n4639), .B2(n7727), .A(n8374), .ZN(n4638) );
  NAND2_X1 U4944 ( .A1(n4639), .A2(n7913), .ZN(n4637) );
  NAND2_X1 U4945 ( .A1(n4981), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4983) );
  OR2_X1 U4946 ( .A1(n8442), .A2(n7694), .ZN(n7828) );
  OR2_X1 U4947 ( .A1(n5133), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U4948 ( .A1(n5075), .A2(n5538), .ZN(n7745) );
  OR2_X1 U4949 ( .A1(n8448), .A2(n8301), .ZN(n7822) );
  OR2_X1 U4950 ( .A1(n7351), .A2(n7464), .ZN(n7797) );
  INV_X1 U4951 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5053) );
  INV_X1 U4952 ( .A(n4969), .ZN(n4580) );
  AND2_X1 U4953 ( .A1(n6389), .A2(n6441), .ZN(n5689) );
  OR2_X1 U4954 ( .A1(n9337), .A2(n9134), .ZN(n8880) );
  AND2_X1 U4955 ( .A1(n4568), .A2(n4331), .ZN(n4567) );
  AND2_X1 U4956 ( .A1(n9379), .A2(n8940), .ZN(n6364) );
  OR2_X1 U4957 ( .A1(n7605), .A2(n7632), .ZN(n8709) );
  NAND2_X1 U4958 ( .A1(n7711), .A2(n7710), .ZN(n7730) );
  OR2_X1 U4959 ( .A1(n7707), .A2(n7706), .ZN(n7711) );
  NAND2_X1 U4960 ( .A1(n5385), .A2(n5384), .ZN(n5398) );
  INV_X1 U4961 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4833) );
  INV_X1 U4962 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5651) );
  AOI21_X1 U4963 ( .B1(n5342), .B2(n4695), .A(n4692), .ZN(n4691) );
  NAND2_X1 U4964 ( .A1(n4693), .A2(n4960), .ZN(n4692) );
  NAND2_X1 U4965 ( .A1(n4695), .A2(n4697), .ZN(n4693) );
  NOR2_X1 U4966 ( .A1(n5673), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U4967 ( .A1(n4928), .A2(n4927), .ZN(n5301) );
  INV_X1 U4968 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5993) );
  OAI21_X1 U4969 ( .B1(n4372), .B2(n4368), .A(n4367), .ZN(n5234) );
  AOI21_X1 U4970 ( .B1(n4366), .B2(n4898), .A(n4321), .ZN(n4367) );
  INV_X1 U4971 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U4972 ( .A1(n5556), .A2(n5557), .ZN(n4762) );
  INV_X1 U4973 ( .A(n5538), .ZN(n5074) );
  AND2_X1 U4974 ( .A1(n8079), .A2(n8080), .ZN(n5582) );
  NAND2_X1 U4975 ( .A1(n6685), .A2(n4276), .ZN(n4768) );
  OAI21_X1 U4976 ( .B1(n9616), .B2(n4454), .A(n4452), .ZN(n9631) );
  AOI21_X1 U4977 ( .B1(n7244), .B2(n7268), .A(n4453), .ZN(n4452) );
  INV_X1 U4978 ( .A(n9633), .ZN(n4453) );
  XNOR2_X1 U4979 ( .A(n7550), .B(n7556), .ZN(n9731) );
  NOR2_X1 U4980 ( .A1(n8177), .A2(n4457), .ZN(n8198) );
  NOR2_X1 U4981 ( .A1(n8181), .A2(n8154), .ZN(n4457) );
  AND2_X1 U4982 ( .A1(n6326), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U4983 ( .A1(n4718), .A2(n4717), .ZN(n7692) );
  OR2_X1 U4984 ( .A1(n8442), .A2(n8312), .ZN(n4717) );
  AND2_X1 U4985 ( .A1(n4713), .A2(n4712), .ZN(n4711) );
  OR2_X1 U4986 ( .A1(n8458), .A2(n8085), .ZN(n8324) );
  INV_X1 U4987 ( .A(n5487), .ZN(n8243) );
  OR2_X1 U4988 ( .A1(n5232), .A2(n4710), .ZN(n4709) );
  INV_X1 U4989 ( .A(n5218), .ZN(n4710) );
  INV_X1 U4990 ( .A(n6724), .ZN(n9778) );
  BUF_X1 U4991 ( .A(n5454), .Z(n5474) );
  AND2_X1 U4992 ( .A1(n6238), .A2(n6237), .ZN(n8540) );
  AOI21_X1 U4993 ( .B1(n4542), .B2(n4544), .A(n4316), .ZN(n4540) );
  INV_X1 U4994 ( .A(n4545), .ZN(n4544) );
  OR2_X1 U4995 ( .A1(n9108), .A2(n6375), .ZN(n6377) );
  NAND2_X1 U4996 ( .A1(n9130), .A2(n8867), .ZN(n4510) );
  INV_X1 U4997 ( .A(n9116), .ZN(n9147) );
  INV_X1 U4998 ( .A(n8940), .ZN(n9262) );
  NAND2_X1 U4999 ( .A1(n4327), .A2(n4280), .ZN(n4556) );
  AND2_X1 U5000 ( .A1(n8905), .A2(n6280), .ZN(n9299) );
  INV_X1 U5001 ( .A(n9553), .ZN(n9295) );
  NAND2_X1 U5002 ( .A1(n8770), .A2(n8769), .ZN(n9052) );
  AND2_X1 U5003 ( .A1(n4960), .A2(n4959), .ZN(n5032) );
  NAND2_X1 U5004 ( .A1(n5661), .A2(n5662), .ZN(n6051) );
  NAND2_X1 U5005 ( .A1(n4371), .A2(n4910), .ZN(n5220) );
  NAND2_X1 U5006 ( .A1(n4887), .A2(n4886), .ZN(n5139) );
  XNOR2_X1 U5007 ( .A(n7542), .B(n7556), .ZN(n9729) );
  NOR2_X1 U5008 ( .A1(n7544), .A2(n7545), .ZN(n8152) );
  XNOR2_X1 U5009 ( .A(n7705), .B(n7915), .ZN(n7995) );
  NAND2_X1 U5010 ( .A1(n4449), .A2(n4602), .ZN(n4448) );
  NOR2_X1 U5011 ( .A1(n7762), .A2(n7763), .ZN(n4602) );
  NOR2_X1 U5012 ( .A1(n4619), .A2(n4600), .ZN(n4599) );
  INV_X1 U5013 ( .A(n4601), .ZN(n4600) );
  AOI21_X1 U5014 ( .B1(n7766), .B2(n7767), .A(n7857), .ZN(n4601) );
  AND2_X1 U5015 ( .A1(n7777), .A2(n4422), .ZN(n7787) );
  INV_X1 U5016 ( .A(n7783), .ZN(n4422) );
  AND2_X1 U5017 ( .A1(n4416), .A2(n4414), .ZN(n7816) );
  INV_X1 U5018 ( .A(n4415), .ZN(n4414) );
  OAI21_X1 U5019 ( .B1(n4418), .B2(n4417), .A(n4275), .ZN(n4415) );
  OAI21_X1 U5020 ( .B1(n4278), .B2(n4320), .A(n4585), .ZN(n4589) );
  AOI21_X1 U5021 ( .B1(n4591), .B2(n4587), .A(n4586), .ZN(n4585) );
  OR2_X1 U5022 ( .A1(n4405), .A2(n4404), .ZN(n7834) );
  NAND2_X1 U5023 ( .A1(n7829), .A2(n7832), .ZN(n4404) );
  AOI21_X1 U5024 ( .B1(n4408), .B2(n4407), .A(n4406), .ZN(n4405) );
  MUX2_X1 U5025 ( .A(n7828), .B(n7827), .S(n7857), .Z(n7829) );
  OR3_X1 U5026 ( .A1(n8868), .A2(n8760), .A3(n8654), .ZN(n8658) );
  OR2_X1 U5027 ( .A1(n8650), .A2(n8649), .ZN(n4402) );
  AND2_X1 U5028 ( .A1(n4504), .A2(n8779), .ZN(n4503) );
  AND2_X1 U5029 ( .A1(n4501), .A2(n4500), .ZN(n8751) );
  NAND2_X1 U5030 ( .A1(n4504), .A2(n4284), .ZN(n4500) );
  AND2_X1 U5031 ( .A1(n6318), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U5032 ( .A1(n4675), .A2(n5416), .ZN(n4674) );
  INV_X1 U5033 ( .A(n5397), .ZN(n4675) );
  INV_X1 U5034 ( .A(n5416), .ZN(n4676) );
  OR2_X1 U5035 ( .A1(n7852), .A2(n4333), .ZN(n7855) );
  AND2_X1 U5036 ( .A1(n7852), .A2(n7853), .ZN(n7866) );
  NAND2_X1 U5037 ( .A1(n4660), .A2(n4658), .ZN(n7856) );
  AND2_X1 U5038 ( .A1(n4659), .A2(n6324), .ZN(n4658) );
  NOR2_X1 U5039 ( .A1(n9379), .A2(n9233), .ZN(n4497) );
  AND2_X1 U5040 ( .A1(n4289), .A2(n4390), .ZN(n4389) );
  NAND2_X1 U5041 ( .A1(n4683), .A2(n4391), .ZN(n4390) );
  INV_X1 U5042 ( .A(n4927), .ZN(n4391) );
  INV_X1 U5043 ( .A(n4910), .ZN(n4370) );
  INV_X1 U5044 ( .A(n5219), .ZN(n4913) );
  INV_X1 U5045 ( .A(SI_1_), .ZN(n4666) );
  AOI21_X1 U5046 ( .B1(n4670), .B2(n4669), .A(n4484), .ZN(n4668) );
  NAND3_X1 U5047 ( .A1(n9050), .A2(n4523), .A3(n4522), .ZN(n4670) );
  INV_X1 U5048 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4522) );
  NAND3_X1 U5049 ( .A1(n4403), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4669) );
  INV_X1 U5050 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4403) );
  INV_X1 U5051 ( .A(n8025), .ZN(n4778) );
  AOI21_X1 U5052 ( .B1(n8025), .B2(n8026), .A(n4777), .ZN(n4776) );
  OR2_X1 U5053 ( .A1(n5599), .A2(n4749), .ZN(n5600) );
  NOR2_X1 U5054 ( .A1(n7861), .A2(n7860), .ZN(n7862) );
  INV_X1 U5055 ( .A(n7855), .ZN(n7868) );
  NOR3_X1 U5056 ( .A1(n7866), .A2(n7865), .A3(n7864), .ZN(n7867) );
  NAND2_X1 U5057 ( .A1(n6525), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U5058 ( .A1(n4477), .A2(n4311), .ZN(n4476) );
  OR2_X1 U5059 ( .A1(n6523), .A2(n6522), .ZN(n4477) );
  NAND2_X1 U5060 ( .A1(n4651), .A2(n4309), .ZN(n7243) );
  INV_X1 U5061 ( .A(n4743), .ZN(n4742) );
  NOR2_X1 U5062 ( .A1(n4742), .A2(n4738), .ZN(n4737) );
  INV_X1 U5063 ( .A(n4746), .ZN(n4738) );
  OAI21_X1 U5064 ( .B1(n7890), .B2(n4617), .A(n7769), .ZN(n4616) );
  NAND2_X1 U5065 ( .A1(n6766), .A2(n7760), .ZN(n4617) );
  NAND2_X1 U5066 ( .A1(n4739), .A2(n4743), .ZN(n6313) );
  NAND2_X1 U5067 ( .A1(n4745), .A2(n4294), .ZN(n4739) );
  OR2_X1 U5068 ( .A1(n7978), .A2(n8122), .ZN(n7847) );
  OR2_X1 U5069 ( .A1(n8268), .A2(n8279), .ZN(n7837) );
  AOI21_X1 U5070 ( .B1(n4726), .B2(n4725), .A(n4308), .ZN(n4724) );
  INV_X1 U5071 ( .A(n4728), .ZN(n4725) );
  NAND4_X1 U5072 ( .A1(n4577), .A2(n4992), .A3(n4579), .A4(n4297), .ZN(n4991)
         );
  NOR2_X1 U5073 ( .A1(n4969), .A2(n4975), .ZN(n4577) );
  INV_X1 U5074 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5476) );
  INV_X1 U5075 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4977) );
  INV_X1 U5076 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U5077 ( .A1(n4788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5314) );
  AND2_X1 U5078 ( .A1(n4791), .A2(n4790), .ZN(n4789) );
  NOR2_X1 U5079 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5084) );
  AOI21_X1 U5080 ( .B1(n4796), .B2(n9556), .A(n4318), .ZN(n5728) );
  AOI21_X1 U5081 ( .B1(n4800), .B2(n4801), .A(n4348), .ZN(n4799) );
  NAND2_X1 U5082 ( .A1(n8523), .A2(n4801), .ZN(n4393) );
  OR2_X1 U5083 ( .A1(n6396), .A2(n8543), .ZN(n8860) );
  OR2_X1 U5084 ( .A1(n9327), .A2(n9094), .ZN(n8859) );
  NAND2_X1 U5085 ( .A1(n4509), .A2(n4507), .ZN(n9092) );
  AOI21_X1 U5086 ( .B1(n4292), .B2(n4513), .A(n4508), .ZN(n4507) );
  INV_X1 U5087 ( .A(n8881), .ZN(n4508) );
  OR2_X1 U5088 ( .A1(n9368), .A2(n9221), .ZN(n9189) );
  INV_X1 U5089 ( .A(n9237), .ZN(n4520) );
  OR2_X1 U5090 ( .A1(n9389), .A2(n9260), .ZN(n8723) );
  NOR2_X1 U5091 ( .A1(n7674), .A2(n7637), .ZN(n4490) );
  NOR2_X1 U5092 ( .A1(n4831), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4576) );
  AND2_X1 U5093 ( .A1(n5366), .A2(n4964), .ZN(n5364) );
  NAND2_X1 U5094 ( .A1(n4701), .A2(n4948), .ZN(n4700) );
  INV_X1 U5095 ( .A(n5352), .ZN(n4701) );
  INV_X1 U5096 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5671) );
  AND2_X1 U5097 ( .A1(n4685), .A2(n4373), .ZN(n4372) );
  AOI21_X1 U5098 ( .B1(n4837), .B2(n4689), .A(n4688), .ZN(n4687) );
  INV_X1 U5099 ( .A(n4903), .ZN(n4688) );
  INV_X1 U5100 ( .A(n4897), .ZN(n4689) );
  OR2_X1 U5101 ( .A1(n5900), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5920) );
  AOI21_X1 U5102 ( .B1(n5159), .B2(n4655), .A(n4322), .ZN(n4654) );
  INV_X1 U5103 ( .A(n4890), .ZN(n4655) );
  INV_X1 U5104 ( .A(n5540), .ZN(n5597) );
  NAND2_X1 U5105 ( .A1(n5558), .A2(n4764), .ZN(n4763) );
  INV_X1 U5106 ( .A(n5553), .ZN(n4764) );
  AND2_X1 U5107 ( .A1(n4783), .A2(n4781), .ZN(n8066) );
  AOI21_X1 U5108 ( .B1(n6914), .B2(n4782), .A(n5551), .ZN(n4781) );
  OR2_X1 U5109 ( .A1(n6793), .A2(n4779), .ZN(n4783) );
  AND2_X1 U5110 ( .A1(n5550), .A2(n6978), .ZN(n5551) );
  XNOR2_X1 U5111 ( .A(n5603), .B(n5601), .ZN(n8116) );
  NAND2_X1 U5112 ( .A1(n5561), .A2(n7457), .ZN(n7460) );
  AND2_X1 U5113 ( .A1(n5521), .A2(n5520), .ZN(n5629) );
  AND2_X1 U5114 ( .A1(n5430), .A2(n5429), .ZN(n6328) );
  AND4_X1 U5115 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n8110)
         );
  AND4_X1 U5116 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n5297)
         );
  AND4_X1 U5117 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n6687)
         );
  NAND4_X1 U5118 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n5538)
         );
  OAI21_X1 U5119 ( .B1(n6525), .B2(P2_REG2_REG_2__SCAN_IN), .A(n4470), .ZN(
        n6464) );
  OR2_X1 U5120 ( .A1(n6463), .A2(n6464), .ZN(n4469) );
  XNOR2_X1 U5121 ( .A(n6525), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6522) );
  OR2_X1 U5122 ( .A1(n6599), .A2(n6600), .ZN(n4651) );
  XNOR2_X1 U5123 ( .A(n7243), .B(n9627), .ZN(n9616) );
  NAND2_X1 U5124 ( .A1(n9616), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U5125 ( .A1(n9648), .A2(n7247), .ZN(n9666) );
  NAND2_X1 U5126 ( .A1(n9666), .A2(n9667), .ZN(n9665) );
  NAND2_X1 U5127 ( .A1(n4983), .A2(n4982), .ZN(n4987) );
  NAND2_X1 U5128 ( .A1(n4984), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5129 ( .A1(n4472), .A2(n4351), .ZN(n7550) );
  NAND2_X1 U5130 ( .A1(n7546), .A2(n4473), .ZN(n4472) );
  INV_X1 U5131 ( .A(n7549), .ZN(n4473) );
  NAND2_X1 U5132 ( .A1(n8158), .A2(n8159), .ZN(n8160) );
  NAND2_X1 U5133 ( .A1(n8160), .A2(n8161), .ZN(n8180) );
  OR2_X1 U5134 ( .A1(n5390), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5406) );
  AND3_X1 U5135 ( .A1(n5361), .A2(n5360), .A3(n5359), .ZN(n7694) );
  NAND2_X1 U5136 ( .A1(n4328), .A2(n4273), .ZN(n4713) );
  NAND2_X1 U5137 ( .A1(n8326), .A2(n5341), .ZN(n4716) );
  NAND2_X1 U5138 ( .A1(n4273), .A2(n5341), .ZN(n4715) );
  AOI21_X1 U5139 ( .B1(n8340), .B2(n8458), .A(n7682), .ZN(n8321) );
  OR2_X1 U5140 ( .A1(n5323), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5335) );
  OR2_X1 U5141 ( .A1(n5305), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5321) );
  OR2_X1 U5142 ( .A1(n5270), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5289) );
  OR2_X1 U5143 ( .A1(n5200), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5225) );
  AND2_X1 U5144 ( .A1(n4647), .A2(n7778), .ZN(n4645) );
  INV_X1 U5145 ( .A(n7785), .ZN(n4647) );
  OR2_X1 U5146 ( .A1(n6974), .A2(n6973), .ZN(n4648) );
  AND2_X1 U5147 ( .A1(n5498), .A2(n7756), .ZN(n4649) );
  NAND2_X1 U5148 ( .A1(n6711), .A2(n7761), .ZN(n4650) );
  INV_X1 U5149 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4999) );
  AND4_X1 U5150 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n6874)
         );
  NAND2_X1 U5151 ( .A1(n6730), .A2(n6731), .ZN(n6720) );
  INV_X1 U5152 ( .A(n7847), .ZN(n4626) );
  NAND2_X1 U5153 ( .A1(n4324), .A2(n4750), .ZN(n4744) );
  NAND2_X1 U5154 ( .A1(n5512), .A2(n7842), .ZN(n7966) );
  INV_X1 U5155 ( .A(n8360), .ZN(n8302) );
  INV_X1 U5156 ( .A(n8362), .ZN(n8300) );
  NAND2_X1 U5157 ( .A1(n8321), .A2(n8320), .ZN(n8319) );
  INV_X1 U5158 ( .A(n7814), .ZN(n4634) );
  AOI21_X1 U5159 ( .B1(n7814), .B2(n4635), .A(n4633), .ZN(n4632) );
  NAND2_X1 U5160 ( .A1(n7813), .A2(n7878), .ZN(n4635) );
  NAND2_X1 U5161 ( .A1(n5334), .A2(n5333), .ZN(n8399) );
  NOR2_X1 U5162 ( .A1(n5311), .A2(n4729), .ZN(n4728) );
  INV_X1 U5163 ( .A(n5298), .ZN(n4729) );
  NAND2_X1 U5164 ( .A1(n8357), .A2(n5296), .ZN(n5299) );
  NAND2_X1 U5165 ( .A1(n4608), .A2(n4606), .ZN(n8346) );
  AOI21_X1 U5166 ( .B1(n4610), .B2(n4613), .A(n4607), .ZN(n4606) );
  INV_X1 U5167 ( .A(n7804), .ZN(n4613) );
  AND2_X1 U5168 ( .A1(n7809), .A2(n7812), .ZN(n8359) );
  AOI21_X1 U5169 ( .B1(n4707), .B2(n4709), .A(n4705), .ZN(n4704) );
  AND2_X1 U5170 ( .A1(n5619), .A2(n7865), .ZN(n8362) );
  AND3_X1 U5171 ( .A1(n5131), .A2(n5130), .A3(n5129), .ZN(n9788) );
  AND3_X1 U5172 ( .A1(n4307), .A2(n5088), .A3(n5087), .ZN(n9773) );
  NAND2_X1 U5173 ( .A1(n7381), .A2(n7174), .ZN(n9816) );
  OR2_X1 U5174 ( .A1(n5523), .A2(n7918), .ZN(n5626) );
  NAND2_X1 U5175 ( .A1(n8484), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5018) );
  AND2_X1 U5176 ( .A1(n5024), .A2(n8484), .ZN(n5026) );
  INV_X1 U5177 ( .A(n4975), .ZN(n4578) );
  AND2_X1 U5178 ( .A1(n5432), .A2(n4702), .ZN(n5453) );
  AND2_X1 U5179 ( .A1(n4977), .A2(n5476), .ZN(n4702) );
  NAND2_X1 U5180 ( .A1(n5235), .A2(n5052), .ZN(n5283) );
  INV_X1 U5181 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5248) );
  INV_X1 U5182 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5049) );
  CLKBUF_X1 U5183 ( .A(n5084), .Z(n5085) );
  NAND2_X1 U5184 ( .A1(n5691), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U5185 ( .A1(n5692), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5885) );
  INV_X1 U5186 ( .A(n5859), .ZN(n5692) );
  NAND2_X1 U5187 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U5188 ( .A1(n5866), .A2(n6168), .ZN(n5867) );
  AND2_X1 U5189 ( .A1(n5852), .A2(n5877), .ZN(n4824) );
  INV_X1 U5190 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5928) );
  AND2_X1 U5191 ( .A1(n6247), .A2(n6248), .ZN(n6246) );
  NOR2_X1 U5192 ( .A1(n4845), .A2(n6115), .ZN(n4802) );
  NAND2_X1 U5193 ( .A1(n6196), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U5194 ( .A1(n5989), .A2(n4380), .ZN(n4375) );
  AOI21_X1 U5195 ( .B1(n4379), .B2(n5989), .A(n4378), .ZN(n4377) );
  NOR2_X1 U5196 ( .A1(n4854), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5197 ( .A1(n6066), .A2(n4813), .ZN(n4812) );
  NOR2_X1 U5198 ( .A1(n6064), .A2(n4854), .ZN(n4810) );
  AND2_X1 U5199 ( .A1(n4811), .A2(n6047), .ZN(n4808) );
  NAND2_X1 U5200 ( .A1(n5693), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5929) );
  INV_X1 U5201 ( .A(n5904), .ZN(n5693) );
  AND2_X1 U5202 ( .A1(n4803), .A2(n4298), .ZN(n8602) );
  NAND2_X1 U5203 ( .A1(n4804), .A2(n4806), .ZN(n4803) );
  INV_X1 U5204 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U5205 ( .A1(n5699), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6140) );
  INV_X1 U5206 ( .A(n6121), .ZN(n5699) );
  OAI22_X1 U5207 ( .A1(n6822), .A2(n8532), .B1(n9560), .B2(n5735), .ZN(n5765)
         );
  XNOR2_X1 U5208 ( .A(n4794), .B(n8529), .ZN(n5749) );
  NAND2_X1 U5209 ( .A1(n7952), .A2(n4796), .ZN(n4795) );
  INV_X1 U5210 ( .A(n8563), .ZN(n4821) );
  AND2_X1 U5211 ( .A1(n6227), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U5212 ( .A1(n8563), .A2(n4820), .ZN(n4819) );
  INV_X1 U5213 ( .A(n6193), .ZN(n4820) );
  NAND2_X1 U5214 ( .A1(n5667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  INV_X1 U5215 ( .A(n8771), .ZN(n6413) );
  NOR2_X1 U5216 ( .A1(n4493), .A2(n9051), .ZN(n4491) );
  NAND2_X1 U5217 ( .A1(n4540), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5218 ( .A1(n4538), .A2(n8815), .ZN(n4537) );
  INV_X1 U5219 ( .A(n4542), .ZN(n4538) );
  NAND2_X1 U5220 ( .A1(n4550), .A2(n4546), .ZN(n4545) );
  AND2_X1 U5221 ( .A1(n8859), .A2(n8759), .ZN(n9078) );
  NOR2_X1 U5222 ( .A1(n6378), .A2(n4548), .ZN(n4547) );
  INV_X1 U5223 ( .A(n6376), .ZN(n4548) );
  NOR2_X1 U5224 ( .A1(n9123), .A2(n9337), .ZN(n9098) );
  NAND2_X1 U5225 ( .A1(n4566), .A2(n4564), .ZN(n9108) );
  AOI21_X1 U5226 ( .B1(n4567), .B2(n4569), .A(n4565), .ZN(n4564) );
  NOR2_X1 U5227 ( .A1(n9127), .A2(n9147), .ZN(n4565) );
  NAND2_X1 U5228 ( .A1(n4279), .A2(n4312), .ZN(n4568) );
  NOR2_X1 U5229 ( .A1(n9139), .A2(n6374), .ZN(n4858) );
  NAND2_X1 U5230 ( .A1(n4279), .A2(n4570), .ZN(n4569) );
  INV_X1 U5231 ( .A(n6369), .ZN(n4570) );
  INV_X1 U5232 ( .A(n9194), .ZN(n9156) );
  AND2_X1 U5233 ( .A1(n8864), .A2(n8861), .ZN(n9164) );
  OR2_X1 U5234 ( .A1(n9180), .A2(n9179), .ZN(n9183) );
  OR2_X1 U5235 ( .A1(n6119), .A2(n6118), .ZN(n6121) );
  NAND2_X1 U5236 ( .A1(n4552), .A2(n4551), .ZN(n9225) );
  NAND2_X1 U5237 ( .A1(n4349), .A2(n6363), .ZN(n4551) );
  AND4_X1 U5238 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n9240)
         );
  NAND2_X1 U5239 ( .A1(n9258), .A2(n9257), .ZN(n4521) );
  OR2_X1 U5240 ( .A1(n9384), .A2(n9240), .ZN(n8737) );
  NAND2_X1 U5241 ( .A1(n9252), .A2(n9251), .ZN(n9250) );
  NOR2_X1 U5242 ( .A1(n9305), .A2(n9389), .ZN(n9273) );
  NOR2_X1 U5243 ( .A1(n4562), .A2(n6362), .ZN(n4561) );
  AOI21_X1 U5244 ( .B1(n4347), .B2(n4560), .A(n4287), .ZN(n4559) );
  INV_X1 U5245 ( .A(n6362), .ZN(n4560) );
  INV_X1 U5246 ( .A(n8942), .ZN(n7616) );
  NOR2_X1 U5247 ( .A1(n7534), .A2(n7637), .ZN(n7619) );
  OR2_X1 U5248 ( .A1(n7477), .A2(n7605), .ZN(n7534) );
  NAND2_X1 U5249 ( .A1(n8797), .A2(n6402), .ZN(n8834) );
  OR3_X1 U5250 ( .A1(n8793), .A2(n8791), .A3(n6401), .ZN(n6402) );
  OAI21_X1 U5251 ( .B1(n7096), .B2(n4533), .A(n4531), .ZN(n7040) );
  AOI21_X1 U5252 ( .B1(n8790), .B2(n4532), .A(n4313), .ZN(n4531) );
  NAND2_X1 U5253 ( .A1(n7097), .A2(n8789), .ZN(n7096) );
  OR2_X1 U5254 ( .A1(n6893), .A2(n6854), .ZN(n6952) );
  INV_X1 U5255 ( .A(n6959), .ZN(n7073) );
  OAI21_X1 U5256 ( .B1(n5743), .B2(n7952), .A(n6812), .ZN(n6885) );
  INV_X1 U5257 ( .A(n9299), .ZN(n9263) );
  INV_X1 U5258 ( .A(n9298), .ZN(n9261) );
  NOR2_X1 U5259 ( .A1(n7952), .A2(n9556), .ZN(n6894) );
  INV_X1 U5260 ( .A(n9229), .ZN(n9306) );
  INV_X1 U5261 ( .A(n9112), .ZN(n9337) );
  INV_X1 U5262 ( .A(n9152), .ZN(n9348) );
  NAND2_X1 U5263 ( .A1(n6017), .A2(n6016), .ZN(n7650) );
  AND2_X1 U5264 ( .A1(n9557), .A2(n6266), .ZN(n9567) );
  AND2_X1 U5265 ( .A1(n6409), .A2(n8923), .ZN(n9553) );
  AND2_X1 U5266 ( .A1(n6532), .A2(n6264), .ZN(n6531) );
  NAND2_X1 U5267 ( .A1(n6259), .A2(n6260), .ZN(n6421) );
  XNOR2_X1 U5268 ( .A(n7735), .B(n7734), .ZN(n8768) );
  OAI21_X1 U5269 ( .B1(n7730), .B2(n7729), .A(n7728), .ZN(n7735) );
  XNOR2_X1 U5270 ( .A(n7730), .B(n7729), .ZN(n8765) );
  INV_X1 U5271 ( .A(n4831), .ZN(n4575) );
  XNOR2_X1 U5272 ( .A(n5403), .B(n5402), .ZN(n7640) );
  XNOR2_X1 U5273 ( .A(n5682), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5274 ( .A1(n5681), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5682) );
  XNOR2_X1 U5275 ( .A(n5398), .B(n5397), .ZN(n7608) );
  INV_X1 U5276 ( .A(n4700), .ZN(n4699) );
  OAI21_X1 U5277 ( .B1(n4700), .B2(n4698), .A(n4954), .ZN(n4697) );
  INV_X1 U5278 ( .A(n4949), .ZN(n4698) );
  NAND2_X1 U5279 ( .A1(n5329), .A2(n5330), .ZN(n4945) );
  OAI21_X1 U5280 ( .B1(n5329), .B2(n5330), .A(n4944), .ZN(n4946) );
  OR2_X1 U5281 ( .A1(n5685), .A2(n5992), .ZN(n5686) );
  NAND2_X1 U5282 ( .A1(n6089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5283 ( .A1(n4678), .A2(n4680), .ZN(n5047) );
  NAND2_X1 U5284 ( .A1(n5301), .A2(n4683), .ZN(n4678) );
  NAND2_X1 U5285 ( .A1(n4679), .A2(n4933), .ZN(n5313) );
  INV_X1 U5286 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5645) );
  XNOR2_X1 U5287 ( .A(n5282), .B(n5281), .ZN(n6786) );
  NAND2_X1 U5288 ( .A1(n4921), .A2(n4920), .ZN(n5265) );
  XNOR2_X1 U5289 ( .A(n5179), .B(n4837), .ZN(n6534) );
  NAND2_X1 U5290 ( .A1(n4882), .A2(n4881), .ZN(n4364) );
  AND4_X1 U5291 ( .A1(n5243), .A2(n5242), .A3(n5241), .A4(n5240), .ZN(n7464)
         );
  NAND2_X1 U5292 ( .A1(n5035), .A2(n5034), .ZN(n8021) );
  NAND2_X1 U5293 ( .A1(n4787), .A2(n4303), .ZN(n8081) );
  NAND2_X1 U5294 ( .A1(n8115), .A2(n4282), .ZN(n8006) );
  AOI21_X1 U5295 ( .B1(n5597), .B2(n6640), .A(n4267), .ZN(n6701) );
  AND4_X1 U5296 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7217)
         );
  AND2_X1 U5297 ( .A1(n5031), .A2(n5030), .ZN(n8266) );
  NAND2_X1 U5298 ( .A1(n5543), .A2(n8146), .ZN(n4772) );
  XNOR2_X1 U5299 ( .A(n5544), .B(n6759), .ZN(n6686) );
  CLKBUF_X1 U5300 ( .A(n5074), .Z(n7703) );
  AND4_X1 U5301 ( .A1(n5045), .A2(n5044), .A3(n5043), .A4(n5042), .ZN(n8085)
         );
  AND3_X1 U5302 ( .A1(n5146), .A2(n5145), .A3(n5144), .ZN(n9794) );
  XNOR2_X1 U5303 ( .A(n5433), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U5304 ( .A1(n4428), .A2(n7871), .ZN(n4427) );
  INV_X1 U5305 ( .A(n7927), .ZN(n4432) );
  AOI21_X1 U5306 ( .B1(n4430), .B2(n7872), .A(n4851), .ZN(n4429) );
  INV_X1 U5307 ( .A(n7694), .ZN(n8312) );
  INV_X1 U5308 ( .A(n8029), .ZN(n8313) );
  INV_X1 U5309 ( .A(n8085), .ZN(n8340) );
  INV_X1 U5310 ( .A(n5297), .ZN(n8349) );
  INV_X1 U5311 ( .A(n7464), .ZN(n8136) );
  INV_X1 U5312 ( .A(n6874), .ZN(n8143) );
  NAND2_X1 U5313 ( .A1(n9729), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9728) );
  OR2_X1 U5314 ( .A1(n8152), .A2(n8153), .ZN(n4459) );
  AND2_X1 U5315 ( .A1(n4459), .A2(n4458), .ZN(n8177) );
  INV_X1 U5316 ( .A(n8155), .ZN(n4458) );
  AOI21_X1 U5317 ( .B1(n6341), .B2(n8365), .A(n6340), .ZN(n7994) );
  AND2_X1 U5318 ( .A1(n5420), .A2(n5419), .ZN(n7854) );
  NAND2_X1 U5319 ( .A1(n5224), .A2(n5223), .ZN(n7790) );
  INV_X1 U5320 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8485) );
  NAND2_X1 U5321 ( .A1(n5925), .A2(n5924), .ZN(n7523) );
  AND2_X1 U5322 ( .A1(n8547), .A2(n8603), .ZN(n8535) );
  INV_X1 U5323 ( .A(n8937), .ZN(n9181) );
  AND4_X1 U5324 ( .A1(n5954), .A2(n5953), .A3(n5952), .A4(n5951), .ZN(n7632)
         );
  AND2_X1 U5325 ( .A1(n6380), .A2(n6379), .ZN(n9085) );
  NAND2_X1 U5326 ( .A1(n4510), .A2(n8779), .ZN(n9114) );
  OAI21_X1 U5327 ( .B1(n9130), .B2(n4513), .A(n4292), .ZN(n9113) );
  NAND2_X1 U5328 ( .A1(n6156), .A2(n6155), .ZN(n9171) );
  INV_X1 U5329 ( .A(n7746), .ZN(n4443) );
  AND2_X1 U5330 ( .A1(n7748), .A2(n7865), .ZN(n4442) );
  NAND2_X1 U5331 ( .A1(n4582), .A2(n7857), .ZN(n4581) );
  NAND2_X1 U5332 ( .A1(n4583), .A2(n7748), .ZN(n4582) );
  NAND2_X1 U5333 ( .A1(n6634), .A2(n7174), .ZN(n4584) );
  NAND2_X1 U5334 ( .A1(n8826), .A2(n8760), .ZN(n8666) );
  INV_X1 U5335 ( .A(n8666), .ZN(n8665) );
  AND2_X1 U5336 ( .A1(n4447), .A2(n4444), .ZN(n7776) );
  AOI21_X1 U5337 ( .B1(n4599), .B2(n4448), .A(n7890), .ZN(n4447) );
  OAI21_X1 U5338 ( .B1(n4446), .B2(n7762), .A(n7760), .ZN(n4445) );
  OAI21_X1 U5339 ( .B1(n7787), .B2(n4285), .A(n7788), .ZN(n4597) );
  AND2_X1 U5340 ( .A1(n4421), .A2(n7784), .ZN(n7789) );
  OR2_X1 U5341 ( .A1(n7787), .A2(n4335), .ZN(n4421) );
  INV_X1 U5342 ( .A(n7812), .ZN(n4417) );
  NAND2_X1 U5343 ( .A1(n7879), .A2(n8324), .ZN(n4590) );
  INV_X1 U5344 ( .A(n4590), .ZN(n4587) );
  NAND2_X1 U5345 ( .A1(n7878), .A2(n7810), .ZN(n4591) );
  OR2_X1 U5346 ( .A1(n4420), .A2(n4419), .ZN(n4413) );
  NAND2_X1 U5347 ( .A1(n4411), .A2(n4410), .ZN(n4420) );
  NAND2_X1 U5348 ( .A1(n4592), .A2(n4409), .ZN(n4408) );
  AND2_X1 U5349 ( .A1(n4588), .A2(n7818), .ZN(n4409) );
  NAND2_X1 U5350 ( .A1(n8304), .A2(n7824), .ZN(n4406) );
  INV_X1 U5351 ( .A(n7825), .ZN(n4407) );
  OAI21_X1 U5352 ( .B1(n7840), .B2(n8271), .A(n7839), .ZN(n7846) );
  AOI21_X1 U5353 ( .B1(n4605), .B2(n4604), .A(n4603), .ZN(n7852) );
  NOR2_X1 U5354 ( .A1(n7967), .A2(n7845), .ZN(n4604) );
  NAND2_X1 U5355 ( .A1(n7846), .A2(n7983), .ZN(n4605) );
  OR2_X1 U5356 ( .A1(n7851), .A2(n7850), .ZN(n4603) );
  NAND2_X1 U5357 ( .A1(n4503), .A2(n4299), .ZN(n4499) );
  AOI21_X1 U5358 ( .B1(n4503), .B2(n4284), .A(n4325), .ZN(n4502) );
  INV_X1 U5359 ( .A(n5046), .ZN(n4677) );
  AND2_X1 U5360 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4993) );
  AND2_X1 U5361 ( .A1(n5052), .A2(n4970), .ZN(n4791) );
  INV_X1 U5362 ( .A(n4802), .ZN(n4800) );
  OAI21_X1 U5363 ( .B1(n8690), .B2(n8793), .A(n8702), .ZN(n6400) );
  AOI21_X1 U5364 ( .B1(n4673), .B2(n4676), .A(n4358), .ZN(n4672) );
  INV_X1 U5365 ( .A(n4696), .ZN(n4695) );
  OAI21_X1 U5366 ( .B1(n4697), .B2(n4699), .A(n5032), .ZN(n4696) );
  INV_X1 U5367 ( .A(n5343), .ZN(n4947) );
  INV_X1 U5368 ( .A(n4683), .ZN(n4392) );
  AND2_X1 U5369 ( .A1(n4924), .A2(n5278), .ZN(n4925) );
  INV_X1 U5370 ( .A(n5263), .ZN(n4923) );
  INV_X1 U5371 ( .A(SI_15_), .ZN(n4922) );
  AND2_X1 U5372 ( .A1(n4277), .A2(n4369), .ZN(n4366) );
  INV_X1 U5373 ( .A(n4784), .ZN(n4780) );
  INV_X1 U5374 ( .A(n5549), .ZN(n4782) );
  NOR2_X1 U5375 ( .A1(n5558), .A2(n4753), .ZN(n4752) );
  NAND2_X1 U5376 ( .A1(n4760), .A2(n4762), .ZN(n4753) );
  INV_X1 U5377 ( .A(n7110), .ZN(n4758) );
  NOR2_X1 U5378 ( .A1(n4759), .A2(n4756), .ZN(n4755) );
  INV_X1 U5379 ( .A(n4762), .ZN(n4756) );
  AND2_X1 U5380 ( .A1(n8420), .A2(n7741), .ZN(n7919) );
  INV_X1 U5381 ( .A(n7919), .ZN(n7875) );
  AND2_X1 U5382 ( .A1(n4469), .A2(n4470), .ZN(n6595) );
  NAND2_X1 U5383 ( .A1(n9634), .A2(n7227), .ZN(n7228) );
  NAND2_X1 U5384 ( .A1(n8180), .A2(n4471), .ZN(n8203) );
  NAND2_X1 U5385 ( .A1(n8178), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5386 ( .A1(n7847), .A2(n4625), .ZN(n4624) );
  INV_X1 U5387 ( .A(n7848), .ZN(n4625) );
  NOR2_X1 U5388 ( .A1(n4626), .A2(n7843), .ZN(n4621) );
  INV_X1 U5389 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7112) );
  NAND2_X1 U5390 ( .A1(n6759), .A2(n4735), .ZN(n4734) );
  AND2_X1 U5391 ( .A1(n5470), .A2(n6490), .ZN(n5519) );
  NAND2_X1 U5392 ( .A1(n7958), .A2(n7739), .ZN(n4660) );
  AND2_X1 U5393 ( .A1(n4750), .A2(n8271), .ZN(n4746) );
  OR2_X1 U5394 ( .A1(n8021), .A2(n8299), .ZN(n7832) );
  NAND2_X1 U5395 ( .A1(n4632), .A2(n4634), .ZN(n4629) );
  INV_X1 U5396 ( .A(n4632), .ZN(n4631) );
  AND2_X1 U5397 ( .A1(n4611), .A2(n7812), .ZN(n4610) );
  NAND2_X1 U5398 ( .A1(n4612), .A2(n7804), .ZN(n4611) );
  INV_X1 U5399 ( .A(n7803), .ZN(n4612) );
  NAND2_X1 U5400 ( .A1(n4994), .A2(n4995), .ZN(n4434) );
  AND2_X1 U5401 ( .A1(n4991), .A2(n4990), .ZN(n4995) );
  NAND2_X1 U5402 ( .A1(n5463), .A2(n4993), .ZN(n4994) );
  INV_X1 U5403 ( .A(n4989), .ZN(n4990) );
  AND2_X1 U5404 ( .A1(n4978), .A2(n5457), .ZN(n4979) );
  INV_X1 U5405 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4978) );
  INV_X1 U5406 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4973) );
  INV_X1 U5407 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5457) );
  INV_X1 U5408 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5251) );
  INV_X1 U5409 ( .A(n5980), .ZN(n4379) );
  INV_X1 U5410 ( .A(n7658), .ZN(n4378) );
  INV_X1 U5411 ( .A(n8513), .ZN(n4385) );
  INV_X1 U5412 ( .A(n8499), .ZN(n4813) );
  NOR2_X1 U5413 ( .A1(n9327), .A2(n9101), .ZN(n4494) );
  OR2_X1 U5414 ( .A1(n9101), .A2(n8540), .ZN(n8886) );
  NAND2_X1 U5415 ( .A1(n9424), .A2(n9212), .ZN(n4571) );
  OR2_X1 U5416 ( .A1(n9201), .A2(n9212), .ZN(n8782) );
  INV_X1 U5417 ( .A(n4840), .ZN(n4554) );
  AND2_X1 U5418 ( .A1(n6363), .A2(n9251), .ZN(n4553) );
  AND2_X1 U5419 ( .A1(n4280), .A2(n4561), .ZN(n4557) );
  NAND2_X1 U5420 ( .A1(n4490), .A2(n9441), .ZN(n4489) );
  NAND2_X1 U5421 ( .A1(n8701), .A2(n8692), .ZN(n8793) );
  NAND2_X1 U5422 ( .A1(n4515), .A2(n4514), .ZN(n8701) );
  INV_X1 U5423 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5884) );
  INV_X1 U5424 ( .A(n4853), .ZN(n4532) );
  NAND2_X1 U5425 ( .A1(n9167), .A2(n6393), .ZN(n9168) );
  NAND2_X1 U5426 ( .A1(n9255), .A2(n4497), .ZN(n9228) );
  AND2_X1 U5427 ( .A1(n9273), .A2(n6392), .ZN(n9255) );
  OR2_X1 U5428 ( .A1(n8919), .A2(n8907), .ZN(n6861) );
  XNOR2_X1 U5429 ( .A(n7709), .B(n7708), .ZN(n7707) );
  INV_X1 U5430 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4832) );
  AND2_X1 U5431 ( .A1(n5415), .A2(n5389), .ZN(n5397) );
  AND2_X1 U5432 ( .A1(n5384), .A2(n5370), .ZN(n5382) );
  INV_X1 U5433 ( .A(SI_20_), .ZN(n5330) );
  NAND2_X1 U5434 ( .A1(n4388), .A2(n4386), .ZN(n5329) );
  AOI21_X1 U5435 ( .B1(n4389), .B2(n4392), .A(n4387), .ZN(n4386) );
  NAND2_X1 U5436 ( .A1(n4928), .A2(n4389), .ZN(n4388) );
  INV_X1 U5437 ( .A(n4943), .ZN(n4387) );
  INV_X1 U5438 ( .A(n4681), .ZN(n4680) );
  OAI21_X1 U5439 ( .B1(n4938), .B2(n4682), .A(n4937), .ZN(n4681) );
  NAND2_X1 U5440 ( .A1(n5300), .A2(n4933), .ZN(n4682) );
  NOR2_X1 U5441 ( .A1(n4938), .A2(n4684), .ZN(n4683) );
  INV_X1 U5442 ( .A(n4933), .ZN(n4684) );
  NAND2_X1 U5443 ( .A1(n4907), .A2(n4906), .ZN(n4910) );
  AOI21_X1 U5444 ( .B1(n4277), .B2(n4690), .A(n4323), .ZN(n4685) );
  OAI21_X1 U5445 ( .B1(n7731), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4878), .ZN(
        n4879) );
  NAND2_X1 U5446 ( .A1(n7731), .A2(n6480), .ZN(n4878) );
  OAI211_X1 U5447 ( .C1(n4665), .C2(n4668), .A(n4663), .B(n4662), .ZN(n5062)
         );
  NAND2_X1 U5448 ( .A1(n4664), .A2(SI_1_), .ZN(n4663) );
  AND2_X1 U5449 ( .A1(n5546), .A2(n8143), .ZN(n4786) );
  NAND2_X1 U5450 ( .A1(n6836), .A2(n4785), .ZN(n4784) );
  INV_X1 U5451 ( .A(n4786), .ZN(n4785) );
  AND2_X1 U5452 ( .A1(n8035), .A2(n5595), .ZN(n8055) );
  OR2_X1 U5453 ( .A1(n6685), .A2(n6686), .ZN(n4769) );
  OAI21_X1 U5454 ( .B1(n4757), .B2(n4754), .A(n4751), .ZN(n7337) );
  NAND2_X1 U5455 ( .A1(n4763), .A2(n4755), .ZN(n4754) );
  AOI21_X1 U5456 ( .B1(n4752), .B2(n4763), .A(n4286), .ZN(n4751) );
  INV_X1 U5457 ( .A(n8064), .ZN(n4757) );
  NAND2_X1 U5458 ( .A1(n4774), .A2(n4301), .ZN(n8091) );
  NAND2_X1 U5459 ( .A1(n4776), .A2(n4778), .ZN(n4773) );
  NAND2_X1 U5460 ( .A1(n8064), .A2(n5553), .ZN(n7312) );
  NAND2_X1 U5461 ( .A1(n4431), .A2(n4344), .ZN(n4430) );
  NAND2_X1 U5462 ( .A1(n7870), .A2(n7869), .ZN(n4431) );
  INV_X1 U5463 ( .A(n4430), .ZN(n4428) );
  XNOR2_X1 U5464 ( .A(n4476), .B(n4475), .ZN(n6592) );
  AOI21_X1 U5465 ( .B1(n6592), .B2(P2_REG1_REG_3__SCAN_IN), .A(n4474), .ZN(
        n6593) );
  AND2_X1 U5466 ( .A1(n4476), .A2(n6597), .ZN(n4474) );
  NOR2_X1 U5467 ( .A1(n5127), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U5468 ( .A1(n9617), .A2(n7226), .ZN(n9635) );
  NAND2_X1 U5469 ( .A1(n9635), .A2(n9636), .ZN(n9634) );
  NAND2_X1 U5470 ( .A1(n9631), .A2(n7245), .ZN(n7246) );
  OR2_X1 U5471 ( .A1(n5156), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5171) );
  XNOR2_X1 U5472 ( .A(n7228), .B(n9660), .ZN(n9651) );
  INV_X1 U5473 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U5474 ( .A1(n9665), .A2(n7248), .ZN(n7249) );
  NAND2_X1 U5475 ( .A1(n9744), .A2(n4478), .ZN(n8157) );
  NAND2_X1 U5476 ( .A1(n9765), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4478) );
  AOI21_X1 U5477 ( .B1(n9729), .B2(n4353), .A(n4455), .ZN(n8150) );
  OAI21_X1 U5478 ( .B1(n7543), .B2(n4456), .A(n4359), .ZN(n4455) );
  INV_X1 U5479 ( .A(n9752), .ZN(n4456) );
  XNOR2_X1 U5480 ( .A(n8203), .B(n8210), .ZN(n8182) );
  OR2_X1 U5481 ( .A1(n4467), .A2(n4361), .ZN(n4466) );
  INV_X1 U5482 ( .A(n4741), .ZN(n4740) );
  NAND2_X1 U5483 ( .A1(n8264), .A2(n4737), .ZN(n4736) );
  OAI21_X1 U5484 ( .B1(n4294), .B2(n4742), .A(n6312), .ZN(n4741) );
  NAND2_X1 U5485 ( .A1(n5374), .A2(n5373), .ZN(n5390) );
  INV_X1 U5486 ( .A(n5375), .ZN(n5374) );
  INV_X1 U5487 ( .A(n5356), .ZN(n5016) );
  NAND2_X1 U5488 ( .A1(n5014), .A2(n5013), .ZN(n5347) );
  INV_X1 U5489 ( .A(n5335), .ZN(n5014) );
  NAND2_X1 U5490 ( .A1(n5012), .A2(n5011), .ZN(n5323) );
  NAND2_X1 U5491 ( .A1(n5010), .A2(n5009), .ZN(n5305) );
  INV_X1 U5492 ( .A(n5289), .ZN(n5010) );
  INV_X1 U5493 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5007) );
  INV_X1 U5494 ( .A(n5256), .ZN(n5008) );
  NAND2_X1 U5495 ( .A1(n5006), .A2(n5005), .ZN(n5256) );
  INV_X1 U5496 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5005) );
  INV_X1 U5497 ( .A(n5238), .ZN(n5006) );
  INV_X1 U5498 ( .A(n5185), .ZN(n5003) );
  AND4_X1 U5499 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n6978)
         );
  NAND2_X1 U5500 ( .A1(n4618), .A2(n4615), .ZN(n6902) );
  INV_X1 U5501 ( .A(n4616), .ZN(n4615) );
  NOR2_X1 U5502 ( .A1(n7890), .A2(n4619), .ZN(n4614) );
  INV_X1 U5503 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5001) );
  INV_X1 U5504 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U5505 ( .A1(n5077), .A2(n5076), .ZN(n6730) );
  AND2_X1 U5506 ( .A1(n5526), .A2(n5488), .ZN(n6631) );
  NOR2_X1 U5507 ( .A1(n9818), .A2(n7747), .ZN(n5615) );
  AND2_X1 U5508 ( .A1(n8250), .A2(n8249), .ZN(n8421) );
  NOR2_X1 U5509 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NOR2_X1 U5510 ( .A1(n7009), .A2(n8300), .ZN(n5450) );
  NAND2_X1 U5511 ( .A1(n8264), .A2(n4746), .ZN(n4745) );
  NOR2_X1 U5512 ( .A1(n4642), .A2(n7830), .ZN(n4641) );
  INV_X1 U5513 ( .A(n7837), .ZN(n4642) );
  AND2_X1 U5514 ( .A1(n7841), .A2(n7842), .ZN(n7983) );
  AND2_X1 U5515 ( .A1(n5396), .A2(n5395), .ZN(n8267) );
  AOI21_X1 U5516 ( .B1(n8021), .B2(n8134), .A(n5362), .ZN(n8277) );
  OAI22_X1 U5517 ( .A1(n5299), .A2(n4721), .B1(n4724), .B2(n5328), .ZN(n7681)
         );
  AND2_X1 U5518 ( .A1(n7903), .A2(n4730), .ZN(n4719) );
  OR2_X1 U5519 ( .A1(n7485), .A2(n7484), .ZN(n7899) );
  INV_X1 U5520 ( .A(n4708), .ZN(n4707) );
  OAI21_X1 U5521 ( .B1(n4709), .B2(n7012), .A(n5231), .ZN(n4708) );
  NAND2_X1 U5522 ( .A1(n4644), .A2(n4643), .ZN(n4646) );
  AOI21_X1 U5523 ( .B1(n4645), .B2(n6973), .A(n4335), .ZN(n4643) );
  NAND2_X1 U5524 ( .A1(n5463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5465) );
  AND2_X1 U5525 ( .A1(n5432), .A2(n4977), .ZN(n5475) );
  CLKBUF_X1 U5526 ( .A(n5434), .Z(n5435) );
  OR2_X1 U5527 ( .A1(n5171), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5180) );
  OR2_X1 U5528 ( .A1(n5097), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5127) );
  AOI22_X1 U5529 ( .A1(n5851), .A2(n5850), .B1(n7067), .B2(n5849), .ZN(n5852)
         );
  NAND2_X1 U5530 ( .A1(n6998), .A2(n5846), .ZN(n4825) );
  NAND2_X1 U5531 ( .A1(n6988), .A2(n5878), .ZN(n5899) );
  AND2_X1 U5532 ( .A1(n6648), .A2(n5729), .ZN(n7948) );
  INV_X1 U5533 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5964) );
  AND2_X1 U5534 ( .A1(n6193), .A2(n6192), .ZN(n8591) );
  OR2_X1 U5535 ( .A1(n5885), .A2(n5884), .ZN(n5904) );
  NAND2_X1 U5536 ( .A1(n4793), .A2(n6649), .ZN(n6648) );
  NAND2_X1 U5537 ( .A1(n5694), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5965) );
  OR2_X1 U5538 ( .A1(n6822), .A2(n8531), .ZN(n5767) );
  NAND2_X1 U5539 ( .A1(n8562), .A2(n8563), .ZN(n6299) );
  NAND2_X1 U5540 ( .A1(n5695), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6036) );
  AND2_X1 U5541 ( .A1(n4814), .A2(n4813), .ZN(n8572) );
  NOR2_X1 U5542 ( .A1(n8778), .A2(n4399), .ZN(n4398) );
  AND2_X1 U5543 ( .A1(n9051), .A2(n8919), .ZN(n4399) );
  AND2_X1 U5544 ( .A1(n6387), .A2(n6386), .ZN(n8543) );
  AND4_X1 U5545 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9260)
         );
  AND2_X1 U5546 ( .A1(n6271), .A2(n6231), .ZN(n9102) );
  AND2_X1 U5547 ( .A1(n6277), .A2(n6276), .ZN(n9094) );
  NAND2_X1 U5548 ( .A1(n4512), .A2(n8779), .ZN(n4511) );
  INV_X1 U5549 ( .A(n8867), .ZN(n4512) );
  OR2_X1 U5550 ( .A1(n9348), .A2(n9157), .ZN(n9129) );
  AND2_X1 U5551 ( .A1(n6218), .A2(n6217), .ZN(n9134) );
  NOR2_X1 U5552 ( .A1(n9348), .A2(n9168), .ZN(n9148) );
  OR2_X1 U5553 ( .A1(n6177), .A2(n8595), .ZN(n6197) );
  AND2_X1 U5554 ( .A1(n9129), .A2(n8862), .ZN(n9144) );
  INV_X1 U5555 ( .A(n8861), .ZN(n4528) );
  OR2_X1 U5556 ( .A1(n6371), .A2(n6370), .ZN(n9140) );
  INV_X1 U5557 ( .A(n6140), .ZN(n6139) );
  NAND2_X1 U5558 ( .A1(n9255), .A2(n4495), .ZN(n9199) );
  AND2_X1 U5559 ( .A1(n4283), .A2(n9424), .ZN(n4495) );
  AND3_X1 U5560 ( .A1(n6124), .A2(n6123), .A3(n6122), .ZN(n9221) );
  AOI21_X1 U5561 ( .B1(n4518), .B2(n9251), .A(n4517), .ZN(n4516) );
  INV_X1 U5562 ( .A(n8736), .ZN(n4517) );
  NAND2_X1 U5563 ( .A1(n5698), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6119) );
  INV_X1 U5564 ( .A(n6105), .ZN(n5698) );
  AND2_X1 U5565 ( .A1(n8660), .A2(n8872), .ZN(n9224) );
  NAND2_X1 U5566 ( .A1(n5697), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6092) );
  INV_X1 U5567 ( .A(n6074), .ZN(n5697) );
  NAND2_X1 U5568 ( .A1(n5696), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6056) );
  INV_X1 U5569 ( .A(n6036), .ZN(n5696) );
  OR2_X1 U5570 ( .A1(n6056), .A2(n6055), .ZN(n6074) );
  NOR2_X1 U5571 ( .A1(n7534), .A2(n4488), .ZN(n7648) );
  INV_X1 U5572 ( .A(n4490), .ZN(n4488) );
  AND2_X1 U5573 ( .A1(n8710), .A2(n8841), .ZN(n8801) );
  AND3_X1 U5574 ( .A1(n7099), .A2(n4274), .A3(n4485), .ZN(n7402) );
  NOR2_X1 U5575 ( .A1(n7206), .A2(n7307), .ZN(n4485) );
  OR2_X1 U5576 ( .A1(n7307), .A2(n4514), .ZN(n6355) );
  NAND2_X1 U5577 ( .A1(n7099), .A2(n9575), .ZN(n7052) );
  AND4_X1 U5578 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n7085)
         );
  AND4_X2 U5579 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n8663)
         );
  OR2_X1 U5580 ( .A1(n6817), .A2(n6816), .ZN(n6826) );
  NAND2_X1 U5581 ( .A1(n6195), .A2(n6194), .ZN(n9343) );
  INV_X1 U5582 ( .A(n7523), .ZN(n6356) );
  OR2_X1 U5583 ( .A1(n6817), .A2(n6428), .ZN(n6432) );
  INV_X1 U5584 ( .A(n9595), .ZN(n9571) );
  XNOR2_X1 U5585 ( .A(n7707), .B(SI_29_), .ZN(n7958) );
  NAND2_X1 U5586 ( .A1(n5651), .A2(n4833), .ZN(n4830) );
  AND2_X1 U5587 ( .A1(n4317), .A2(n5663), .ZN(n5664) );
  NAND2_X1 U5588 ( .A1(n5672), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  INV_X1 U5589 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U5590 ( .A1(n6087), .A2(n6086), .ZN(n6089) );
  NAND2_X1 U5591 ( .A1(n4686), .A2(n4687), .ZN(n5194) );
  OR2_X1 U5592 ( .A1(n4898), .A2(n4690), .ZN(n4686) );
  OR2_X1 U5593 ( .A1(n5879), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U5594 ( .A1(n4526), .A2(n4654), .ZN(n5174) );
  OR2_X1 U5595 ( .A1(n6793), .A2(n4784), .ZN(n6835) );
  INV_X1 U5596 ( .A(n8004), .ZN(n5605) );
  NAND2_X1 U5597 ( .A1(n6835), .A2(n5549), .ZN(n6915) );
  NAND2_X1 U5598 ( .A1(n8024), .A2(n5583), .ZN(n4775) );
  NAND2_X1 U5599 ( .A1(n4763), .A2(n4762), .ZN(n4761) );
  NOR2_X1 U5600 ( .A1(n8064), .A2(n4766), .ZN(n4765) );
  AND2_X1 U5601 ( .A1(n4769), .A2(n4276), .ZN(n6757) );
  INV_X1 U5602 ( .A(n4769), .ZN(n6684) );
  NAND2_X1 U5603 ( .A1(n5616), .A2(n7996), .ZN(n8072) );
  OAI22_X1 U5604 ( .A1(n6700), .A2(n6701), .B1(n5539), .B2(n8148), .ZN(n6693)
         );
  CLKBUF_X1 U5605 ( .A(n5104), .Z(n6732) );
  OR2_X1 U5606 ( .A1(n5545), .A2(n8144), .ZN(n4770) );
  AOI21_X1 U5607 ( .B1(n4276), .B2(n6686), .A(n6758), .ZN(n4767) );
  NAND2_X1 U5608 ( .A1(n7460), .A2(n5563), .ZN(n7500) );
  NAND2_X1 U5609 ( .A1(n5631), .A2(n5630), .ZN(n8124) );
  INV_X1 U5610 ( .A(n7933), .ZN(n4425) );
  INV_X1 U5611 ( .A(n8267), .ZN(n8132) );
  NAND4_X1 U5612 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), .ZN(n8147)
         );
  CLKBUF_X1 U5613 ( .A(n5538), .Z(n8148) );
  INV_X1 U5614 ( .A(P2_U3893), .ZN(n8215) );
  INV_X1 U5615 ( .A(n4469), .ZN(n6524) );
  INV_X1 U5616 ( .A(n4651), .ZN(n7239) );
  NAND2_X1 U5617 ( .A1(n9615), .A2(n7244), .ZN(n9632) );
  XNOR2_X1 U5618 ( .A(n7246), .B(n9660), .ZN(n9649) );
  NAND2_X1 U5619 ( .A1(n9649), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U5620 ( .A1(n9716), .A2(n7235), .ZN(n7546) );
  NAND2_X1 U5621 ( .A1(n9730), .A2(n7551), .ZN(n9746) );
  NAND2_X1 U5622 ( .A1(n9746), .A2(n9745), .ZN(n9744) );
  NAND2_X1 U5623 ( .A1(n9728), .A2(n7543), .ZN(n9758) );
  XNOR2_X1 U5624 ( .A(n8150), .B(n8151), .ZN(n7544) );
  XNOR2_X1 U5625 ( .A(n8157), .B(n8151), .ZN(n7552) );
  NAND2_X1 U5626 ( .A1(n4467), .A2(n4361), .ZN(n4465) );
  NOR2_X1 U5627 ( .A1(n8202), .A2(n8237), .ZN(n4462) );
  NOR2_X1 U5628 ( .A1(n8199), .A2(n8200), .ZN(n8201) );
  INV_X1 U5629 ( .A(n7854), .ZN(n8260) );
  NAND2_X1 U5630 ( .A1(n5510), .A2(n7877), .ZN(n8272) );
  NAND2_X1 U5631 ( .A1(n4714), .A2(n4713), .ZN(n8297) );
  NAND2_X1 U5632 ( .A1(n4648), .A2(n4645), .ZN(n7011) );
  AND2_X1 U5633 ( .A1(n5184), .A2(n5183), .ZN(n9810) );
  OAI21_X1 U5634 ( .B1(n6767), .B2(n6766), .A(n7760), .ZN(n6880) );
  NAND2_X1 U5635 ( .A1(n6489), .A2(n5615), .ZN(n7996) );
  NAND2_X1 U5636 ( .A1(n4650), .A2(n7756), .ZN(n6751) );
  OR2_X1 U5637 ( .A1(n7737), .A2(n9974), .ZN(n5103) );
  INV_X1 U5638 ( .A(n8330), .ZN(n8369) );
  INV_X2 U5639 ( .A(n8336), .ZN(n8366) );
  AOI21_X1 U5640 ( .B1(n8768), .B2(n7739), .A(n7738), .ZN(n8374) );
  AOI21_X1 U5641 ( .B1(n7608), .B2(n7739), .A(n4356), .ZN(n8379) );
  AND2_X1 U5642 ( .A1(n4997), .A2(n4996), .ZN(n8387) );
  NAND2_X1 U5643 ( .A1(n7718), .A2(n7717), .ZN(n8424) );
  OR2_X1 U5644 ( .A1(n7995), .A2(n9818), .ZN(n6342) );
  INV_X1 U5645 ( .A(n4622), .ZN(n6327) );
  AOI21_X1 U5646 ( .B1(n7966), .B2(n7848), .A(n4626), .ZN(n4622) );
  NAND2_X1 U5647 ( .A1(n5405), .A2(n5404), .ZN(n7978) );
  INV_X1 U5648 ( .A(n8379), .ZN(n7991) );
  INV_X1 U5649 ( .A(n8387), .ZN(n8436) );
  NAND2_X1 U5650 ( .A1(n5355), .A2(n5354), .ZN(n8442) );
  NAND2_X1 U5651 ( .A1(n8319), .A2(n5341), .ZN(n8311) );
  OAI21_X1 U5652 ( .B1(n5507), .B2(n4634), .A(n4632), .ZN(n8309) );
  NAND2_X1 U5653 ( .A1(n5057), .A2(n5056), .ZN(n8458) );
  NAND2_X1 U5654 ( .A1(n5320), .A2(n5319), .ZN(n8465) );
  NAND2_X1 U5655 ( .A1(n4723), .A2(n4726), .ZN(n8339) );
  NAND2_X1 U5656 ( .A1(n5299), .A2(n4728), .ZN(n4723) );
  NAND2_X1 U5657 ( .A1(n5304), .A2(n5303), .ZN(n8471) );
  NAND2_X1 U5658 ( .A1(n5299), .A2(n5298), .ZN(n8348) );
  NAND2_X1 U5659 ( .A1(n5288), .A2(n5287), .ZN(n8478) );
  NAND2_X1 U5660 ( .A1(n4609), .A2(n7804), .ZN(n8355) );
  NAND2_X1 U5661 ( .A1(n7483), .A2(n7803), .ZN(n4609) );
  NAND2_X1 U5662 ( .A1(n5269), .A2(n5268), .ZN(n7498) );
  NAND2_X1 U5663 ( .A1(n5237), .A2(n5236), .ZN(n7351) );
  NAND2_X1 U5664 ( .A1(n4706), .A2(n5218), .ZN(n7118) );
  NAND2_X1 U5665 ( .A1(n7017), .A2(n7012), .ZN(n4706) );
  INV_X1 U5666 ( .A(n8428), .ZN(n8477) );
  NAND2_X1 U5667 ( .A1(n6489), .A2(n6488), .ZN(n6498) );
  NOR2_X1 U5668 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4593) );
  INV_X1 U5669 ( .A(n5026), .ZN(n8495) );
  INV_X1 U5670 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7515) );
  MUX2_X1 U5671 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5456), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5459) );
  NAND2_X1 U5672 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  INV_X1 U5673 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7383) );
  INV_X1 U5674 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7176) );
  INV_X1 U5675 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U5676 ( .A1(n5316), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  INV_X1 U5677 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6870) );
  INV_X1 U5678 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6792) );
  INV_X1 U5679 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9963) );
  INV_X1 U5680 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6540) );
  INV_X1 U5681 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6497) );
  INV_X1 U5682 ( .A(n9643), .ZN(n7275) );
  OR2_X1 U5683 ( .A1(n5085), .A2(n8485), .ZN(n4652) );
  XNOR2_X1 U5684 ( .A(n6263), .B(n6262), .ZN(n6532) );
  AOI21_X1 U5685 ( .B1(n6303), .B2(n6248), .A(n6247), .ZN(n6268) );
  INV_X1 U5686 ( .A(n4814), .ZN(n8500) );
  AOI21_X1 U5687 ( .B1(n8511), .B2(n8513), .A(n8512), .ZN(n8510) );
  INV_X1 U5688 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U5689 ( .A1(n5944), .A2(n5940), .ZN(n7516) );
  XNOR2_X1 U5690 ( .A(n5790), .B(n5788), .ZN(n6779) );
  NAND2_X1 U5691 ( .A1(n4817), .A2(n4815), .ZN(n8539) );
  AND2_X1 U5692 ( .A1(n6246), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U5693 ( .A1(n4818), .A2(n4821), .ZN(n4816) );
  INV_X1 U5694 ( .A(n9085), .ZN(n9327) );
  INV_X1 U5695 ( .A(n4480), .ZN(n4479) );
  OAI22_X1 U5696 ( .A1(n4484), .A2(n4483), .B1(n4482), .B2(n4481), .ZN(n4480)
         );
  NAND2_X1 U5697 ( .A1(n4804), .A2(n4802), .ZN(n4798) );
  NAND2_X1 U5698 ( .A1(n6054), .A2(n6053), .ZN(n9389) );
  AND4_X1 U5699 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n7050)
         );
  NOR2_X1 U5700 ( .A1(n4810), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U5701 ( .A1(n6048), .A2(n4811), .ZN(n4809) );
  OAI211_X2 U5702 ( .C1(n5853), .C2(n6481), .A(n5801), .B(n5800), .ZN(n9566)
         );
  AND2_X1 U5703 ( .A1(n6283), .A2(n6281), .ZN(n8627) );
  NAND2_X1 U5704 ( .A1(n7595), .A2(n5980), .ZN(n4376) );
  NAND2_X1 U5705 ( .A1(n6153), .A2(n8513), .ZN(n8612) );
  NAND2_X1 U5706 ( .A1(n4365), .A2(n6138), .ZN(n9357) );
  NAND2_X1 U5707 ( .A1(n7379), .A2(n5758), .ZN(n4365) );
  AND2_X1 U5708 ( .A1(n6293), .A2(n6267), .ZN(n8603) );
  INV_X1 U5709 ( .A(n8607), .ZN(n8635) );
  NAND2_X1 U5710 ( .A1(n6034), .A2(n6033), .ZN(n9308) );
  INV_X1 U5711 ( .A(n8610), .ZN(n8641) );
  INV_X1 U5712 ( .A(n8540), .ZN(n9117) );
  NAND2_X1 U5713 ( .A1(n6203), .A2(n6202), .ZN(n9116) );
  NAND2_X1 U5714 ( .A1(n6163), .A2(n6162), .ZN(n8937) );
  OR2_X1 U5715 ( .A1(n6099), .A2(n6098), .ZN(n8940) );
  INV_X1 U5716 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6624) );
  INV_X1 U5717 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6622) );
  INV_X1 U5718 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6620) );
  AND4_X1 U5719 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n6959)
         );
  INV_X1 U5720 ( .A(n8663), .ZN(n8945) );
  OR2_X1 U5721 ( .A1(n5751), .A2(n5752), .ZN(n5756) );
  OR2_X1 U5722 ( .A1(n8771), .A2(n5739), .ZN(n5741) );
  NAND2_X1 U5723 ( .A1(n5773), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5718) );
  AND2_X1 U5724 ( .A1(n5923), .A2(n5945), .ZN(n9458) );
  INV_X1 U5725 ( .A(n7358), .ZN(n9516) );
  AND2_X1 U5726 ( .A1(n6611), .A2(n6578), .ZN(n9885) );
  NOR2_X1 U5727 ( .A1(n9053), .A2(n9306), .ZN(n9319) );
  NAND2_X1 U5728 ( .A1(n4540), .A2(n8815), .ZN(n4539) );
  OAI21_X1 U5729 ( .B1(n4540), .B2(n4549), .A(n4536), .ZN(n4535) );
  NAND2_X1 U5730 ( .A1(n4541), .A2(n4545), .ZN(n9075) );
  AND2_X1 U5731 ( .A1(n6208), .A2(n6207), .ZN(n9112) );
  NAND2_X1 U5732 ( .A1(n4563), .A2(n4568), .ZN(n9122) );
  OR2_X1 U5733 ( .A1(n9197), .A2(n4569), .ZN(n4563) );
  AND2_X1 U5734 ( .A1(n6176), .A2(n6175), .ZN(n9152) );
  NAND2_X1 U5735 ( .A1(n9183), .A2(n4281), .ZN(n9155) );
  INV_X1 U5736 ( .A(n9357), .ZN(n9178) );
  NAND2_X1 U5737 ( .A1(n6103), .A2(n6102), .ZN(n9233) );
  NAND2_X1 U5738 ( .A1(n4521), .A2(n8737), .ZN(n9238) );
  NAND2_X1 U5739 ( .A1(n9250), .A2(n4840), .ZN(n9236) );
  NAND2_X1 U5740 ( .A1(n6072), .A2(n6071), .ZN(n9384) );
  NAND2_X1 U5741 ( .A1(n4558), .A2(n4559), .ZN(n9304) );
  NAND2_X1 U5742 ( .A1(n7618), .A2(n4561), .ZN(n4558) );
  AOI21_X1 U5743 ( .B1(n7618), .B2(n8803), .A(n4347), .ZN(n7641) );
  NAND2_X1 U5744 ( .A1(n6403), .A2(n8710), .ZN(n7614) );
  NAND2_X1 U5745 ( .A1(n5948), .A2(n5947), .ZN(n7605) );
  NAND2_X1 U5746 ( .A1(n4529), .A2(n8834), .ZN(n7399) );
  NAND2_X1 U5747 ( .A1(n6964), .A2(n8790), .ZN(n6963) );
  NAND2_X1 U5748 ( .A1(n7096), .A2(n4853), .ZN(n6964) );
  AND2_X1 U5749 ( .A1(n8914), .A2(n8819), .ZN(n9557) );
  NAND2_X1 U5750 ( .A1(n5963), .A2(n5962), .ZN(n7637) );
  INV_X1 U5751 ( .A(n9171), .ZN(n6393) );
  INV_X1 U5752 ( .A(n9233), .ZN(n9429) );
  INV_X1 U5753 ( .A(n7650), .ZN(n9441) );
  OAI211_X1 U5754 ( .C1(n5853), .C2(n6484), .A(n5822), .B(n5821), .ZN(n7107)
         );
  NAND2_X1 U5755 ( .A1(n9598), .A2(n9567), .ZN(n9440) );
  XNOR2_X1 U5756 ( .A(n5418), .B(n6317), .ZN(n7961) );
  NAND2_X1 U5757 ( .A1(n5417), .A2(n5416), .ZN(n6319) );
  NAND2_X1 U5758 ( .A1(n5652), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5653) );
  AND2_X1 U5759 ( .A1(n5661), .A2(n4574), .ZN(n5656) );
  NAND2_X1 U5760 ( .A1(n5680), .A2(n4291), .ZN(n7512) );
  XNOR2_X1 U5761 ( .A(n5033), .B(n5032), .ZN(n7421) );
  INV_X1 U5762 ( .A(n4694), .ZN(n5033) );
  INV_X1 U5763 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7380) );
  INV_X1 U5764 ( .A(n8921), .ZN(n8914) );
  INV_X1 U5765 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7173) );
  INV_X1 U5766 ( .A(n6265), .ZN(n8819) );
  INV_X1 U5767 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6972) );
  INV_X1 U5769 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9948) );
  INV_X1 U5770 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6788) );
  INV_X1 U5771 ( .A(n5661), .ZN(n6049) );
  AND2_X1 U5772 ( .A1(n6015), .A2(n6030), .ZN(n9532) );
  INV_X1 U5773 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6627) );
  INV_X1 U5774 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9945) );
  INV_X1 U5775 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6538) );
  INV_X1 U5776 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6535) );
  INV_X1 U5777 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U5778 ( .A1(n4657), .A2(n4890), .ZN(n5158) );
  OR2_X1 U5779 ( .A1(n5840), .A2(n5839), .ZN(n6570) );
  NAND2_X1 U5780 ( .A1(n4424), .A2(n4423), .ZN(P2_U3296) );
  OR2_X1 U5781 ( .A1(n7932), .A2(n7931), .ZN(n4423) );
  NAND2_X1 U5782 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  INV_X1 U5783 ( .A(n4459), .ZN(n8156) );
  OAI21_X1 U5784 ( .B1(n7667), .B2(n8492), .A(n4436), .ZN(P2_U3268) );
  AND2_X1 U5785 ( .A1(n4438), .A2(n4437), .ZN(n4436) );
  OR2_X1 U5786 ( .A1(n8494), .A2(n9972), .ZN(n4438) );
  INV_X1 U5787 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6478) );
  OR2_X1 U5788 ( .A1(n8448), .A2(n5351), .ZN(n4273) );
  AND2_X1 U5789 ( .A1(n9575), .A2(n7198), .ZN(n4274) );
  AND2_X1 U5790 ( .A1(n7879), .A2(n7811), .ZN(n4275) );
  NAND2_X1 U5791 ( .A1(n5544), .A2(n6759), .ZN(n4276) );
  AND2_X1 U5792 ( .A1(n4687), .A2(n5195), .ZN(n4277) );
  INV_X1 U5793 ( .A(n8779), .ZN(n4513) );
  AND2_X1 U5794 ( .A1(n4413), .A2(n4418), .ZN(n4278) );
  OR2_X1 U5795 ( .A1(n6374), .A2(n6373), .ZN(n4279) );
  NAND2_X1 U5796 ( .A1(n9436), .A2(n8505), .ZN(n4280) );
  AND2_X1 U5797 ( .A1(n9164), .A2(n8863), .ZN(n4281) );
  AND2_X1 U5798 ( .A1(n5604), .A2(n5605), .ZN(n4282) );
  INV_X1 U5799 ( .A(n8347), .ZN(n4727) );
  INV_X1 U5800 ( .A(n9556), .ZN(n6922) );
  AND2_X1 U5801 ( .A1(n4497), .A2(n4496), .ZN(n4283) );
  INV_X1 U5802 ( .A(n9051), .ZN(n9408) );
  NAND2_X1 U5803 ( .A1(n8767), .A2(n8766), .ZN(n9051) );
  INV_X1 U5804 ( .A(n4845), .ZN(n4805) );
  NOR2_X1 U5805 ( .A1(n6134), .A2(n8552), .ZN(n4845) );
  NAND2_X1 U5806 ( .A1(n8747), .A2(n9144), .ZN(n4284) );
  NAND2_X1 U5807 ( .A1(n4326), .A2(n4805), .ZN(n4801) );
  OR2_X1 U5808 ( .A1(n8471), .A2(n8110), .ZN(n7811) );
  OR2_X1 U5809 ( .A1(n7785), .A2(n7786), .ZN(n4285) );
  NAND2_X1 U5810 ( .A1(n6048), .A2(n6047), .ZN(n8497) );
  AND2_X1 U5811 ( .A1(n4758), .A2(n7792), .ZN(n4286) );
  NOR2_X1 U5812 ( .A1(n9441), .A2(n7660), .ZN(n4287) );
  INV_X1 U5813 ( .A(n7609), .ZN(n5473) );
  NAND2_X1 U5814 ( .A1(n5467), .A2(n5466), .ZN(n7609) );
  OR2_X1 U5815 ( .A1(n6759), .A2(n4735), .ZN(n4288) );
  AND2_X1 U5816 ( .A1(n4680), .A2(n4677), .ZN(n4289) );
  AND2_X1 U5817 ( .A1(n5381), .A2(n5380), .ZN(n8279) );
  INV_X1 U5818 ( .A(n8279), .ZN(n4749) );
  AND4_X1 U5819 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n7401)
         );
  INV_X1 U5820 ( .A(n7401), .ZN(n4514) );
  NOR2_X1 U5821 ( .A1(n4355), .A2(n5107), .ZN(n6712) );
  INV_X1 U5822 ( .A(n7813), .ZN(n4586) );
  INV_X1 U5823 ( .A(n8202), .ZN(n4468) );
  AND2_X1 U5824 ( .A1(n5266), .A2(n5253), .ZN(n9754) );
  NAND2_X2 U5825 ( .A1(n5707), .A2(n7934), .ZN(n5774) );
  INV_X1 U5826 ( .A(n6715), .ZN(n4735) );
  NOR2_X1 U5827 ( .A1(n8103), .A2(n4841), .ZN(n4290) );
  INV_X1 U5828 ( .A(n8523), .ZN(n4804) );
  INV_X1 U5829 ( .A(n4796), .ZN(n5735) );
  OR2_X1 U5830 ( .A1(n6048), .A2(n6047), .ZN(n4814) );
  OR2_X1 U5831 ( .A1(n5678), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4291) );
  NAND2_X1 U5833 ( .A1(n5835), .A2(n7731), .ZN(n4482) );
  AND2_X1 U5834 ( .A1(n9115), .A2(n4511), .ZN(n4292) );
  NAND2_X1 U5835 ( .A1(n4898), .A2(n4277), .ZN(n4374) );
  INV_X1 U5836 ( .A(n8815), .ZN(n4549) );
  NAND2_X1 U5837 ( .A1(n8860), .A2(n8888), .ZN(n8815) );
  AND2_X1 U5838 ( .A1(n9098), .A2(n4492), .ZN(n4293) );
  AND2_X1 U5839 ( .A1(n4744), .A2(n4747), .ZN(n4294) );
  INV_X1 U5840 ( .A(n7760), .ZN(n4619) );
  AND2_X1 U5841 ( .A1(n7800), .A2(n7801), .ZN(n7900) );
  INV_X1 U5842 ( .A(n8803), .ZN(n4562) );
  INV_X1 U5843 ( .A(n7934), .ZN(n4530) );
  INV_X1 U5844 ( .A(n7898), .ZN(n4705) );
  AND2_X1 U5845 ( .A1(n7900), .A2(n7799), .ZN(n4295) );
  AND2_X1 U5846 ( .A1(n8379), .A2(n8267), .ZN(n4296) );
  INV_X1 U5847 ( .A(n9089), .ZN(n4546) );
  AND3_X1 U5848 ( .A1(n4972), .A2(n4971), .A3(n4980), .ZN(n4297) );
  NAND2_X1 U5849 ( .A1(n8116), .A2(n8267), .ZN(n8115) );
  NAND2_X1 U5850 ( .A1(n4792), .A2(n8054), .ZN(n8016) );
  INV_X1 U5851 ( .A(n5558), .ZN(n4766) );
  NAND2_X1 U5852 ( .A1(n4798), .A2(n4801), .ZN(n8553) );
  NAND2_X1 U5853 ( .A1(n6114), .A2(n6113), .ZN(n4298) );
  AND3_X1 U5854 ( .A1(n8745), .A2(n8744), .A3(n8746), .ZN(n4299) );
  AND2_X1 U5855 ( .A1(n7978), .A2(n8131), .ZN(n4300) );
  NAND2_X1 U5856 ( .A1(n5661), .A2(n5650), .ZN(n5678) );
  OR2_X1 U5857 ( .A1(n8436), .A2(n8266), .ZN(n7877) );
  INV_X1 U5858 ( .A(n9379), .ZN(n9247) );
  NAND2_X1 U5859 ( .A1(n6091), .A2(n6090), .ZN(n9379) );
  AND2_X1 U5860 ( .A1(n4773), .A2(n8090), .ZN(n4301) );
  INV_X1 U5861 ( .A(n7747), .ZN(n7174) );
  NAND2_X1 U5862 ( .A1(n5998), .A2(n5997), .ZN(n7674) );
  AND2_X1 U5863 ( .A1(n4397), .A2(n8920), .ZN(n4302) );
  NAND2_X1 U5864 ( .A1(n5346), .A2(n5345), .ZN(n8448) );
  INV_X1 U5865 ( .A(n6378), .ZN(n4550) );
  AND2_X1 U5866 ( .A1(n4290), .A2(n5578), .ZN(n4303) );
  AND2_X1 U5867 ( .A1(n7991), .A2(n8267), .ZN(n7844) );
  AND3_X1 U5868 ( .A1(n4402), .A2(n4401), .A3(n4400), .ZN(n4304) );
  AND2_X1 U5869 ( .A1(n7899), .A2(n7802), .ZN(n4305) );
  INV_X1 U5870 ( .A(n9101), .ZN(n6394) );
  NAND2_X1 U5871 ( .A1(n6229), .A2(n6228), .ZN(n9101) );
  INV_X1 U5872 ( .A(n5761), .ZN(n4829) );
  AND2_X1 U5873 ( .A1(n5805), .A2(n5791), .ZN(n4306) );
  NAND2_X1 U5874 ( .A1(n4727), .A2(n4731), .ZN(n4726) );
  NAND2_X1 U5875 ( .A1(n6382), .A2(n6381), .ZN(n6396) );
  OR2_X1 U5876 ( .A1(n7737), .A2(n6477), .ZN(n4307) );
  AND2_X1 U5877 ( .A1(n8465), .A2(n8350), .ZN(n4308) );
  OR2_X1 U5878 ( .A1(n7241), .A2(n7240), .ZN(n4309) );
  NAND2_X1 U5879 ( .A1(n9308), .A2(n9282), .ZN(n4310) );
  OR2_X1 U5880 ( .A1(n6521), .A2(n9834), .ZN(n4311) );
  NAND2_X1 U5881 ( .A1(n4858), .A2(n4571), .ZN(n4312) );
  OR2_X1 U5882 ( .A1(n8399), .A2(n8313), .ZN(n5341) );
  NOR2_X1 U5883 ( .A1(n8944), .A2(n7074), .ZN(n4313) );
  INV_X1 U5884 ( .A(n5311), .ZN(n4731) );
  OR2_X1 U5885 ( .A1(n8478), .A2(n5297), .ZN(n7809) );
  INV_X1 U5886 ( .A(n7809), .ZN(n4607) );
  INV_X1 U5887 ( .A(n4493), .ZN(n4492) );
  NAND2_X1 U5888 ( .A1(n4494), .A2(n9068), .ZN(n4493) );
  OR2_X1 U5889 ( .A1(n4854), .A2(n6065), .ZN(n4314) );
  AND2_X1 U5890 ( .A1(n9085), .A2(n9094), .ZN(n4315) );
  AND2_X1 U5891 ( .A1(n8934), .A2(n9327), .ZN(n4316) );
  AND2_X1 U5892 ( .A1(n6086), .A2(n5671), .ZN(n4317) );
  INV_X1 U5893 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5021) );
  AND2_X1 U5894 ( .A1(n6351), .A2(n6168), .ZN(n4318) );
  INV_X1 U5895 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5657) );
  AND2_X1 U5896 ( .A1(n5611), .A2(n8117), .ZN(n4319) );
  OR2_X1 U5897 ( .A1(n4590), .A2(n4607), .ZN(n4320) );
  AND2_X1 U5898 ( .A1(n4912), .A2(SI_12_), .ZN(n4321) );
  AND2_X1 U5899 ( .A1(n4892), .A2(SI_7_), .ZN(n4322) );
  AND2_X1 U5900 ( .A1(n4905), .A2(SI_10_), .ZN(n4323) );
  OR2_X1 U5901 ( .A1(n4748), .A2(n4296), .ZN(n4324) );
  OR2_X1 U5902 ( .A1(n8465), .A2(n5577), .ZN(n7879) );
  NAND2_X1 U5903 ( .A1(n8880), .A2(n8780), .ZN(n4325) );
  NAND2_X1 U5904 ( .A1(n6135), .A2(n4298), .ZN(n4326) );
  INV_X1 U5905 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U5906 ( .A1(n7110), .A2(n8137), .ZN(n4760) );
  NAND2_X1 U5907 ( .A1(n4559), .A2(n4310), .ZN(n4327) );
  NAND2_X1 U5908 ( .A1(n8310), .A2(n4716), .ZN(n4328) );
  OR2_X1 U5909 ( .A1(n7767), .A2(n7757), .ZN(n4329) );
  OR2_X1 U5910 ( .A1(n7991), .A2(n8267), .ZN(n7842) );
  AND2_X1 U5911 ( .A1(n4542), .A2(n4549), .ZN(n4330) );
  OR2_X1 U5912 ( .A1(n9343), .A2(n9116), .ZN(n4331) );
  AND3_X1 U5913 ( .A1(n5650), .A2(n5652), .A3(n4576), .ZN(n4332) );
  AND2_X1 U5914 ( .A1(n7915), .A2(n7853), .ZN(n4333) );
  OR2_X1 U5915 ( .A1(n9179), .A2(n4528), .ZN(n4334) );
  INV_X1 U5916 ( .A(n7818), .ZN(n4633) );
  NAND2_X1 U5917 ( .A1(n7788), .A2(n7780), .ZN(n4335) );
  NOR2_X1 U5918 ( .A1(n4419), .A2(n4417), .ZN(n4336) );
  NOR2_X1 U5919 ( .A1(n8201), .A2(n8202), .ZN(n4337) );
  AND2_X1 U5920 ( .A1(n4562), .A2(n8710), .ZN(n4338) );
  INV_X1 U5921 ( .A(n4369), .ZN(n4368) );
  NOR2_X1 U5922 ( .A1(n4913), .A2(n4370), .ZN(n4369) );
  OR2_X1 U5923 ( .A1(n9827), .A2(n7217), .ZN(n7784) );
  AND2_X1 U5924 ( .A1(n5565), .A2(n5563), .ZN(n4339) );
  AND2_X1 U5925 ( .A1(n9183), .A2(n8863), .ZN(n4340) );
  AND2_X1 U5926 ( .A1(n4972), .A2(n4971), .ZN(n4341) );
  INV_X1 U5927 ( .A(n4519), .ZN(n4518) );
  NAND2_X1 U5928 ( .A1(n4520), .A2(n8737), .ZN(n4519) );
  INV_X1 U5929 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U5930 ( .A1(n5944), .A2(n4823), .ZN(n7595) );
  AND2_X1 U5931 ( .A1(n4775), .A2(n8025), .ZN(n4342) );
  AND2_X1 U5932 ( .A1(n9255), .A2(n9247), .ZN(n4343) );
  NOR2_X1 U5933 ( .A1(n9199), .A2(n9357), .ZN(n9167) );
  NAND2_X1 U5934 ( .A1(n5235), .A2(n4791), .ZN(n5285) );
  AND2_X1 U5935 ( .A1(n5712), .A2(n5711), .ZN(n9212) );
  INV_X1 U5936 ( .A(n9660), .ZN(n7265) );
  NAND2_X1 U5937 ( .A1(n4376), .A2(n5989), .ZN(n7657) );
  XNOR2_X1 U5938 ( .A(n5686), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6265) );
  AND2_X1 U5939 ( .A1(n7828), .A2(n7826), .ZN(n8304) );
  INV_X1 U5940 ( .A(n8304), .ZN(n4712) );
  AND3_X1 U5941 ( .A1(n4826), .A2(n4829), .A3(n4834), .ZN(n5960) );
  NAND2_X1 U5942 ( .A1(n5856), .A2(n5855), .ZN(n7051) );
  NAND2_X1 U5943 ( .A1(n4787), .A2(n4290), .ZN(n7936) );
  AND4_X1 U5944 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n7027)
         );
  AND3_X1 U5945 ( .A1(n5040), .A2(n5039), .A3(n5038), .ZN(n8299) );
  AND4_X1 U5946 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7600)
         );
  AND4_X1 U5947 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n7331)
         );
  INV_X1 U5948 ( .A(n7504), .ZN(n8135) );
  AND4_X1 U5949 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n7504)
         );
  NAND2_X1 U5950 ( .A1(n5372), .A2(n5371), .ZN(n8268) );
  NAND2_X1 U5951 ( .A1(n9255), .A2(n4283), .ZN(n4498) );
  NAND2_X1 U5952 ( .A1(n8374), .A2(n8250), .ZN(n4344) );
  AND2_X1 U5953 ( .A1(n7726), .A2(n5447), .ZN(n7009) );
  INV_X1 U5954 ( .A(n7009), .ZN(n4659) );
  AND2_X1 U5955 ( .A1(n4521), .A2(n4518), .ZN(n4345) );
  AND2_X1 U5956 ( .A1(n4822), .A2(n5944), .ZN(n4346) );
  AND2_X1 U5957 ( .A1(n7674), .A2(n8941), .ZN(n4347) );
  NOR2_X1 U5958 ( .A1(n6137), .A2(n6136), .ZN(n4348) );
  INV_X1 U5959 ( .A(n6012), .ZN(n4380) );
  INV_X1 U5960 ( .A(n6115), .ZN(n4806) );
  AND2_X1 U5961 ( .A1(n8521), .A2(n8520), .ZN(n6115) );
  NOR2_X1 U5962 ( .A1(n8268), .A2(n4749), .ZN(n4748) );
  OR2_X1 U5963 ( .A1(n6364), .A2(n4554), .ZN(n4349) );
  AND2_X1 U5964 ( .A1(n4839), .A2(n4920), .ZN(n4350) );
  AND2_X1 U5965 ( .A1(n5660), .A2(n5659), .ZN(n9424) );
  INV_X1 U5966 ( .A(n9424), .ZN(n9201) );
  NAND2_X1 U5967 ( .A1(n5687), .A2(n8893), .ZN(n6266) );
  NAND2_X1 U5968 ( .A1(n5903), .A2(n5902), .ZN(n7307) );
  INV_X1 U5969 ( .A(n7307), .ZN(n4515) );
  NAND2_X1 U5970 ( .A1(n6117), .A2(n6116), .ZN(n9368) );
  INV_X1 U5971 ( .A(n9368), .ZN(n4496) );
  OR2_X1 U5972 ( .A1(n7548), .A2(n7547), .ZN(n4351) );
  INV_X1 U5973 ( .A(n7865), .ZN(n7857) );
  NAND2_X1 U5974 ( .A1(n4646), .A2(n7784), .ZN(n7121) );
  NAND2_X1 U5975 ( .A1(n4648), .A2(n7778), .ZN(n7023) );
  NAND2_X1 U5976 ( .A1(n8921), .A2(n5687), .ZN(n6278) );
  INV_X1 U5977 ( .A(n8089), .ZN(n4777) );
  NAND2_X1 U5978 ( .A1(n4825), .A2(n5852), .ZN(n6987) );
  NAND2_X1 U5979 ( .A1(n5792), .A2(n4306), .ZN(n6803) );
  NAND2_X1 U5980 ( .A1(n5792), .A2(n5791), .ZN(n6801) );
  NAND2_X1 U5981 ( .A1(n7099), .A2(n4274), .ZN(n4352) );
  NOR3_X1 U5982 ( .A1(n7534), .A2(n9308), .A3(n4489), .ZN(n4486) );
  AND2_X1 U5983 ( .A1(n9752), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4353) );
  XNOR2_X1 U5984 ( .A(n5899), .B(n5897), .ZN(n7202) );
  NOR2_X1 U5985 ( .A1(n6793), .A2(n4786), .ZN(n4354) );
  INV_X1 U5986 ( .A(n4487), .ZN(n9307) );
  NOR2_X1 U5987 ( .A1(n7534), .A2(n4489), .ZN(n4487) );
  AND2_X1 U5988 ( .A1(n6720), .A2(n5108), .ZN(n4355) );
  NOR2_X1 U5989 ( .A1(n7737), .A2(n7610), .ZN(n4356) );
  NAND2_X1 U5990 ( .A1(n5475), .A2(n5474), .ZN(n4357) );
  AND2_X1 U5991 ( .A1(n6321), .A2(n6320), .ZN(n4358) );
  NAND2_X1 U5992 ( .A1(n9765), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4359) );
  NOR2_X1 U5993 ( .A1(n4765), .A2(n4761), .ZN(n4360) );
  INV_X1 U5994 ( .A(n5757), .ZN(n6822) );
  NAND4_X1 U5995 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n8149)
         );
  AND2_X1 U5996 ( .A1(n8230), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4361) );
  INV_X1 U5997 ( .A(n8181), .ZN(n8178) );
  INV_X1 U5998 ( .A(n4464), .ZN(n4463) );
  OAI21_X1 U5999 ( .B1(n4466), .B2(n4468), .A(n4465), .ZN(n4464) );
  INV_X1 U6000 ( .A(n8237), .ZN(n4467) );
  AND2_X1 U6001 ( .A1(n4463), .A2(n4466), .ZN(n4362) );
  OR2_X1 U6002 ( .A1(n4464), .A2(n4462), .ZN(n4363) );
  INV_X1 U6003 ( .A(n6597), .ZN(n4475) );
  INV_X1 U6004 ( .A(n6474), .ZN(n4481) );
  INV_X1 U6005 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4484) );
  INV_X1 U6006 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4523) );
  OR2_X2 U6007 ( .A1(n7411), .A2(n7900), .ZN(n7413) );
  NAND2_X1 U6008 ( .A1(n5245), .A2(n5244), .ZN(n7411) );
  NAND2_X1 U6009 ( .A1(n4714), .A2(n4711), .ZN(n4718) );
  NAND2_X1 U6010 ( .A1(n4364), .A2(n5126), .ZN(n4887) );
  XNOR2_X1 U6011 ( .A(n5126), .B(n4364), .ZN(n6484) );
  XNOR2_X1 U6012 ( .A(n5353), .B(n5352), .ZN(n7379) );
  NAND2_X1 U6013 ( .A1(n4372), .A2(n4374), .ZN(n4371) );
  NAND2_X1 U6014 ( .A1(n4374), .A2(n4685), .ZN(n5207) );
  INV_X1 U6015 ( .A(n5208), .ZN(n4373) );
  NAND2_X2 U6016 ( .A1(n4383), .A2(n4381), .ZN(n8590) );
  OAI21_X2 U6017 ( .B1(n8590), .B2(n4821), .A(n4818), .ZN(n6303) );
  NAND2_X1 U6018 ( .A1(n6803), .A2(n5808), .ZN(n6998) );
  NAND3_X1 U6019 ( .A1(n4670), .A2(n4669), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4667) );
  NAND3_X1 U6020 ( .A1(n4411), .A2(n4410), .A3(n4336), .ZN(n4416) );
  NAND3_X1 U6021 ( .A1(n4432), .A2(n4429), .A3(n4427), .ZN(n4426) );
  NAND2_X2 U6022 ( .A1(n7928), .A2(n4434), .ZN(n5048) );
  CLKBUF_X1 U6023 ( .A(n8236), .Z(n4433) );
  AND2_X1 U6024 ( .A1(n4433), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6447) );
  XNOR2_X1 U6025 ( .A(n4435), .B(n4433), .ZN(n5619) );
  INV_X1 U6026 ( .A(n7928), .ZN(n4435) );
  MUX2_X1 U6027 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n8236), .Z(n6443) );
  MUX2_X1 U6028 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n8236), .Z(n9609) );
  MUX2_X1 U6029 ( .A(P2_REG1_REG_2__SCAN_IN), .B(P2_REG2_REG_2__SCAN_IN), .S(
        n8236), .Z(n6517) );
  MUX2_X1 U6030 ( .A(P2_REG1_REG_3__SCAN_IN), .B(P2_REG2_REG_3__SCAN_IN), .S(
        n8236), .Z(n6588) );
  MUX2_X1 U6031 ( .A(P2_REG1_REG_4__SCAN_IN), .B(P2_REG2_REG_4__SCAN_IN), .S(
        n8236), .Z(n7271) );
  MUX2_X1 U6032 ( .A(n7267), .B(n7268), .S(n8236), .Z(n7272) );
  MUX2_X1 U6033 ( .A(P2_REG1_REG_6__SCAN_IN), .B(P2_REG2_REG_6__SCAN_IN), .S(
        n4433), .Z(n7276) );
  MUX2_X1 U6034 ( .A(P2_REG1_REG_7__SCAN_IN), .B(P2_REG2_REG_7__SCAN_IN), .S(
        n4433), .Z(n7266) );
  MUX2_X1 U6035 ( .A(P2_REG1_REG_8__SCAN_IN), .B(P2_REG2_REG_8__SCAN_IN), .S(
        n4433), .Z(n7264) );
  MUX2_X1 U6036 ( .A(P2_REG1_REG_9__SCAN_IN), .B(P2_REG2_REG_9__SCAN_IN), .S(
        n4433), .Z(n7262) );
  MUX2_X1 U6037 ( .A(P2_REG1_REG_10__SCAN_IN), .B(P2_REG2_REG_10__SCAN_IN), 
        .S(n4433), .Z(n7260) );
  MUX2_X1 U6038 ( .A(P2_REG1_REG_11__SCAN_IN), .B(P2_REG2_REG_11__SCAN_IN), 
        .S(n4433), .Z(n7258) );
  MUX2_X1 U6039 ( .A(P2_REG1_REG_12__SCAN_IN), .B(P2_REG2_REG_12__SCAN_IN), 
        .S(n4433), .Z(n7559) );
  MUX2_X1 U6040 ( .A(P2_REG1_REG_13__SCAN_IN), .B(P2_REG2_REG_13__SCAN_IN), 
        .S(n4433), .Z(n7557) );
  MUX2_X1 U6041 ( .A(P2_REG1_REG_14__SCAN_IN), .B(P2_REG2_REG_14__SCAN_IN), 
        .S(n4433), .Z(n7555) );
  MUX2_X1 U6042 ( .A(P2_REG1_REG_15__SCAN_IN), .B(P2_REG2_REG_15__SCAN_IN), 
        .S(n4433), .Z(n8167) );
  MUX2_X1 U6043 ( .A(P2_REG1_REG_16__SCAN_IN), .B(P2_REG2_REG_16__SCAN_IN), 
        .S(n4433), .Z(n8163) );
  MUX2_X1 U6044 ( .A(P2_REG1_REG_17__SCAN_IN), .B(P2_REG2_REG_17__SCAN_IN), 
        .S(n4433), .Z(n8207) );
  MUX2_X1 U6045 ( .A(P2_REG1_REG_18__SCAN_IN), .B(P2_REG2_REG_18__SCAN_IN), 
        .S(n4433), .Z(n8212) );
  NAND2_X1 U6046 ( .A1(n4433), .A2(P2_STATE_REG_SCAN_IN), .ZN(n4437) );
  NAND4_X1 U6047 ( .A1(n4440), .A2(n7913), .A3(n7856), .A4(n4439), .ZN(n7863)
         );
  INV_X1 U6048 ( .A(n7881), .ZN(n7744) );
  NAND2_X1 U6049 ( .A1(n4581), .A2(n4441), .ZN(n7754) );
  OAI21_X1 U6050 ( .B1(n7881), .B2(n4443), .A(n4442), .ZN(n4441) );
  NAND2_X1 U6051 ( .A1(n4580), .A2(n4579), .ZN(n5209) );
  NAND2_X1 U6052 ( .A1(n4445), .A2(n7857), .ZN(n4444) );
  AOI21_X1 U6053 ( .B1(n7765), .B2(n7758), .A(n4329), .ZN(n4446) );
  NAND2_X1 U6054 ( .A1(n7765), .A2(n7764), .ZN(n4449) );
  INV_X1 U6055 ( .A(n4450), .ZN(n4451) );
  INV_X2 U6056 ( .A(n5075), .ZN(n5536) );
  INV_X1 U6057 ( .A(n7244), .ZN(n4454) );
  NAND2_X1 U6058 ( .A1(n8201), .A2(n4362), .ZN(n4460) );
  OAI211_X1 U6059 ( .C1(n8201), .C2(n4363), .A(n4460), .B(n9737), .ZN(n4461)
         );
  NAND2_X1 U6060 ( .A1(n4461), .A2(n8248), .ZN(P2_U3201) );
  NAND3_X1 U6061 ( .A1(n7099), .A2(n4274), .A3(n6391), .ZN(n7293) );
  INV_X1 U6062 ( .A(n4486), .ZN(n9305) );
  AND2_X1 U6063 ( .A1(n9098), .A2(n4494), .ZN(n9081) );
  NAND2_X1 U6064 ( .A1(n9098), .A2(n4491), .ZN(n9059) );
  NAND2_X1 U6065 ( .A1(n9098), .A2(n6394), .ZN(n9099) );
  INV_X1 U6066 ( .A(n4498), .ZN(n9213) );
  NAND2_X1 U6067 ( .A1(n4499), .A2(n4502), .ZN(n8752) );
  NAND4_X1 U6068 ( .A1(n8745), .A2(n8744), .A3(n8746), .A4(n4504), .ZN(n4501)
         );
  XNOR2_X1 U6069 ( .A(n4506), .B(n5663), .ZN(n5687) );
  NAND2_X2 U6070 ( .A1(n9045), .A2(n8914), .ZN(n8919) );
  NAND2_X1 U6071 ( .A1(n9130), .A2(n4292), .ZN(n4509) );
  OAI21_X1 U6072 ( .B1(n9258), .B2(n4519), .A(n4516), .ZN(n9220) );
  NAND2_X1 U6073 ( .A1(n5139), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U6074 ( .A1(n6403), .A2(n4338), .ZN(n7642) );
  NAND2_X1 U6075 ( .A1(n7642), .A2(n6404), .ZN(n6405) );
  NAND3_X1 U6076 ( .A1(n4529), .A2(n8834), .A3(n8796), .ZN(n7397) );
  NAND2_X1 U6077 ( .A1(n8833), .A2(n6957), .ZN(n4529) );
  INV_X1 U6078 ( .A(n5707), .ZN(n7959) );
  INV_X1 U6079 ( .A(n8790), .ZN(n4533) );
  NAND2_X1 U6080 ( .A1(n6377), .A2(n4330), .ZN(n4534) );
  OAI211_X1 U6081 ( .C1(n6377), .C2(n4539), .A(n4535), .B(n4534), .ZN(n9064)
         );
  NAND2_X1 U6082 ( .A1(n6377), .A2(n4547), .ZN(n4541) );
  NAND2_X1 U6083 ( .A1(n6377), .A2(n6376), .ZN(n9090) );
  NAND2_X1 U6084 ( .A1(n9252), .A2(n4553), .ZN(n4552) );
  NAND2_X1 U6085 ( .A1(n7618), .A2(n4557), .ZN(n4555) );
  NAND2_X1 U6086 ( .A1(n4555), .A2(n4556), .ZN(n9272) );
  NAND2_X1 U6087 ( .A1(n9197), .A2(n4567), .ZN(n4566) );
  OR2_X1 U6088 ( .A1(n9197), .A2(n6369), .ZN(n4572) );
  NAND2_X1 U6089 ( .A1(n5661), .A2(n4332), .ZN(n5701) );
  AND2_X1 U6090 ( .A1(n5650), .A2(n4576), .ZN(n4573) );
  AND2_X1 U6091 ( .A1(n5650), .A2(n4575), .ZN(n4574) );
  NOR2_X2 U6092 ( .A1(n5097), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4579) );
  NAND3_X1 U6093 ( .A1(n4584), .A2(n7746), .A3(n7745), .ZN(n4583) );
  NAND2_X1 U6094 ( .A1(n4589), .A2(n7865), .ZN(n4588) );
  NAND2_X1 U6095 ( .A1(n7817), .A2(n7857), .ZN(n4592) );
  NAND2_X1 U6096 ( .A1(n4985), .A2(n4984), .ZN(n5019) );
  NAND2_X1 U6097 ( .A1(n4985), .A2(n4593), .ZN(n8484) );
  NOR2_X1 U6098 ( .A1(n7755), .A2(n7882), .ZN(n7765) );
  AOI21_X1 U6099 ( .B1(n7754), .B2(n7885), .A(n7753), .ZN(n7755) );
  MUX2_X1 U6100 ( .A(n7836), .B(n7835), .S(n7857), .Z(n7840) );
  XNOR2_X1 U6101 ( .A(n5018), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5025) );
  OAI211_X1 U6102 ( .C1(n7776), .C2(n7775), .A(n7892), .B(n7774), .ZN(n7777)
         );
  NAND2_X1 U6103 ( .A1(n6948), .A2(n6949), .ZN(n7102) );
  NAND2_X1 U6104 ( .A1(n9279), .A2(n8723), .ZN(n9258) );
  NAND2_X1 U6105 ( .A1(n7471), .A2(n8709), .ZN(n7526) );
  NAND2_X1 U6106 ( .A1(n6821), .A2(n6924), .ZN(n6820) );
  NAND2_X1 U6107 ( .A1(n9219), .A2(n8872), .ZN(n8897) );
  INV_X8 U6108 ( .A(n4266), .ZN(n7731) );
  NAND2_X1 U6109 ( .A1(n5139), .A2(n5140), .ZN(n4657) );
  NAND2_X1 U6110 ( .A1(n7483), .A2(n4610), .ZN(n4608) );
  NAND2_X1 U6111 ( .A1(n6767), .A2(n4614), .ZN(n4618) );
  NAND2_X1 U6112 ( .A1(n4620), .A2(n4623), .ZN(n6330) );
  NAND2_X1 U6113 ( .A1(n5512), .A2(n4621), .ZN(n4620) );
  INV_X1 U6114 ( .A(n4627), .ZN(n8305) );
  NAND2_X1 U6115 ( .A1(n5507), .A2(n7878), .ZN(n8323) );
  INV_X1 U6116 ( .A(n8149), .ZN(n4636) );
  NAND3_X1 U6117 ( .A1(n4267), .A2(n7745), .A3(n7748), .ZN(n6655) );
  NAND2_X1 U6118 ( .A1(n4636), .A2(n9771), .ZN(n6634) );
  NAND2_X1 U6119 ( .A1(n5510), .A2(n4641), .ZN(n4640) );
  NAND2_X1 U6120 ( .A1(n6974), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6121 ( .A1(n4650), .A2(n4649), .ZN(n5499) );
  XNOR2_X2 U6122 ( .A(n4652), .B(n5086), .ZN(n6525) );
  NAND2_X1 U6123 ( .A1(n4660), .A2(n6324), .ZN(n6345) );
  NAND2_X1 U6124 ( .A1(n4661), .A2(n4667), .ZN(n4864) );
  INV_X1 U6125 ( .A(n4668), .ZN(n4661) );
  NAND2_X1 U6126 ( .A1(n4668), .A2(SI_1_), .ZN(n4662) );
  INV_X1 U6127 ( .A(n4667), .ZN(n4664) );
  NAND2_X1 U6128 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U6129 ( .A1(n5279), .A2(n4925), .ZN(n4928) );
  NAND2_X1 U6130 ( .A1(n4921), .A2(n4350), .ZN(n5279) );
  NAND2_X1 U6131 ( .A1(n5398), .A2(n4673), .ZN(n4671) );
  NAND2_X1 U6132 ( .A1(n4671), .A2(n4672), .ZN(n7709) );
  NAND2_X1 U6133 ( .A1(n5398), .A2(n5397), .ZN(n5417) );
  OR2_X1 U6134 ( .A1(n5301), .A2(n5300), .ZN(n4679) );
  NAND2_X1 U6135 ( .A1(n4898), .A2(n4897), .ZN(n5179) );
  INV_X1 U6136 ( .A(n4837), .ZN(n4690) );
  INV_X1 U6137 ( .A(n4691), .ZN(n5365) );
  AOI21_X1 U6138 ( .B1(n5342), .B2(n4699), .A(n4697), .ZN(n4694) );
  OAI21_X1 U6139 ( .B1(n5342), .B2(n4949), .A(n4948), .ZN(n5353) );
  AND2_X2 U6140 ( .A1(n5453), .A2(n4979), .ZN(n4992) );
  NAND2_X1 U6141 ( .A1(n4704), .A2(n4703), .ZN(n5245) );
  NAND2_X1 U6142 ( .A1(n7017), .A2(n4707), .ZN(n4703) );
  OAI21_X1 U6143 ( .B1(n7017), .B2(n4709), .A(n4707), .ZN(n7344) );
  NAND2_X1 U6144 ( .A1(n4726), .A2(n4719), .ZN(n4720) );
  OAI22_X2 U6145 ( .A1(n4720), .A2(n5299), .B1(n4722), .B2(n4724), .ZN(n7682)
         );
  NAND2_X1 U6146 ( .A1(n4726), .A2(n4730), .ZN(n4721) );
  NAND2_X1 U6147 ( .A1(n7903), .A2(n4730), .ZN(n4722) );
  INV_X1 U6148 ( .A(n5328), .ZN(n4730) );
  NAND2_X1 U6149 ( .A1(n5107), .A2(n4734), .ZN(n4732) );
  NAND3_X1 U6150 ( .A1(n4733), .A2(n4732), .A3(n4288), .ZN(n6752) );
  NAND3_X1 U6151 ( .A1(n6720), .A2(n5108), .A3(n4734), .ZN(n4733) );
  NAND2_X1 U6152 ( .A1(n6752), .A2(n6750), .ZN(n5132) );
  NAND2_X1 U6153 ( .A1(n4736), .A2(n4740), .ZN(n6315) );
  NAND2_X1 U6154 ( .A1(n4745), .A2(n4744), .ZN(n7968) );
  AOI21_X1 U6155 ( .B1(n8264), .B2(n8271), .A(n4748), .ZN(n7984) );
  NAND2_X1 U6156 ( .A1(n7991), .A2(n8132), .ZN(n4750) );
  NAND2_X1 U6157 ( .A1(n4768), .A2(n4767), .ZN(n4771) );
  NAND2_X1 U6158 ( .A1(n4771), .A2(n4770), .ZN(n6794) );
  NAND2_X1 U6159 ( .A1(n6641), .A2(n4772), .ZN(n6685) );
  NAND2_X1 U6160 ( .A1(n8024), .A2(n4776), .ZN(n4774) );
  NAND2_X1 U6161 ( .A1(n4780), .A2(n6914), .ZN(n4779) );
  NAND2_X1 U6162 ( .A1(n5235), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U6163 ( .A1(n7460), .A2(n4339), .ZN(n7501) );
  NOR2_X1 U6164 ( .A1(n4969), .A2(n5097), .ZN(n5196) );
  INV_X1 U6165 ( .A(n5209), .ZN(n5050) );
  NAND2_X1 U6166 ( .A1(n8115), .A2(n5604), .ZN(n8005) );
  NAND3_X1 U6167 ( .A1(n8115), .A2(n4282), .A3(n4319), .ZN(n5640) );
  NAND2_X1 U6168 ( .A1(n5592), .A2(n5591), .ZN(n8054) );
  NAND2_X1 U6169 ( .A1(n5590), .A2(n5589), .ZN(n4792) );
  OAI21_X1 U6170 ( .B1(n6649), .B2(n4793), .A(n6648), .ZN(n8961) );
  NAND2_X1 U6171 ( .A1(n5728), .A2(n5724), .ZN(n4793) );
  XNOR2_X2 U6172 ( .A(n5702), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6173 ( .A1(n5743), .A2(n6168), .ZN(n4797) );
  NAND2_X1 U6174 ( .A1(n4797), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6175 ( .A1(n8590), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U6176 ( .A1(n8590), .A2(n6193), .ZN(n8562) );
  NAND2_X1 U6177 ( .A1(n5940), .A2(n5943), .ZN(n4823) );
  NAND2_X1 U6178 ( .A1(n4825), .A2(n4824), .ZN(n6988) );
  AND4_X2 U6179 ( .A1(n4826), .A2(n4829), .A3(n4834), .A4(n5646), .ZN(n5661)
         );
  NAND2_X1 U6180 ( .A1(n4829), .A2(n4834), .ZN(n5817) );
  NAND3_X1 U6181 ( .A1(n5651), .A2(n4833), .A3(n4832), .ZN(n4831) );
  NAND2_X1 U6182 ( .A1(n6361), .A2(n4838), .ZN(n7618) );
  AND2_X1 U6183 ( .A1(n6319), .A2(n6316), .ZN(n5418) );
  OR2_X1 U6184 ( .A1(n8670), .A2(n6399), .ZN(n8661) );
  NAND2_X1 U6185 ( .A1(n4917), .A2(n4916), .ZN(n5247) );
  XNOR2_X1 U6186 ( .A(n5101), .B(n5100), .ZN(n6475) );
  NAND2_X1 U6187 ( .A1(n5050), .A2(n5049), .ZN(n5221) );
  AOI21_X1 U6188 ( .B1(n5019), .B2(P2_IR_REG_31__SCAN_IN), .A(n5021), .ZN(
        n5020) );
  INV_X1 U6189 ( .A(n7721), .ZN(n6333) );
  XNOR2_X1 U6190 ( .A(n5536), .B(n5540), .ZN(n5537) );
  NAND4_X2 U6191 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .ZN(n6351)
         );
  INV_X2 U6192 ( .A(n9589), .ZN(n9598) );
  INV_X2 U6193 ( .A(n9605), .ZN(n9608) );
  AND2_X1 U6194 ( .A1(n10005), .A2(n5642), .ZN(n4834) );
  OR2_X1 U6195 ( .A1(n9598), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n4835) );
  OR2_X1 U6196 ( .A1(n9608), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4836) );
  AND2_X1 U6197 ( .A1(n4903), .A2(n4902), .ZN(n4837) );
  INV_X1 U6198 ( .A(n8613), .ZN(n6154) );
  OR2_X1 U6199 ( .A1(n7577), .A2(n7616), .ZN(n4838) );
  OR2_X1 U6200 ( .A1(n4923), .A2(n4922), .ZN(n4839) );
  OR2_X1 U6201 ( .A1(n6392), .A2(n9240), .ZN(n4840) );
  AND2_X1 U6202 ( .A1(n5576), .A2(n5577), .ZN(n4841) );
  OR2_X1 U6203 ( .A1(n7999), .A2(n8386), .ZN(n4842) );
  OR2_X1 U6204 ( .A1(n9068), .A2(n9401), .ZN(n4843) );
  AND2_X1 U6205 ( .A1(n8859), .A2(n4859), .ZN(n4844) );
  NAND2_X1 U6206 ( .A1(n4946), .A2(n4945), .ZN(n5342) );
  OR2_X1 U6207 ( .A1(n6394), .A2(n8610), .ZN(n4846) );
  OR2_X1 U6208 ( .A1(n9068), .A2(n9440), .ZN(n4847) );
  OR2_X1 U6209 ( .A1(n7999), .A2(n8428), .ZN(n4848) );
  OR2_X1 U6210 ( .A1(n9274), .A2(n9260), .ZN(n4849) );
  OAI21_X1 U6211 ( .B1(n8346), .B2(n5506), .A(n7810), .ZN(n8337) );
  OR2_X1 U6212 ( .A1(n9429), .A2(n9241), .ZN(n4850) );
  INV_X1 U6213 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5703) );
  INV_X1 U6214 ( .A(n9098), .ZN(n9109) );
  AND3_X1 U6215 ( .A1(n7926), .A2(n8243), .A3(n7740), .ZN(n4851) );
  INV_X1 U6216 ( .A(n5092), .ZN(n5443) );
  AND2_X1 U6217 ( .A1(n7609), .A2(n7513), .ZN(n4852) );
  AND2_X1 U6218 ( .A1(n5350), .A2(n5349), .ZN(n8301) );
  INV_X1 U6219 ( .A(n8301), .ZN(n5351) );
  OR2_X1 U6220 ( .A1(n7073), .A2(n7107), .ZN(n4853) );
  AND2_X1 U6221 ( .A1(n6069), .A2(n6068), .ZN(n4854) );
  AND2_X1 U6222 ( .A1(n7747), .A2(n7062), .ZN(n4855) );
  INV_X1 U6223 ( .A(n8365), .ZN(n9768) );
  NAND2_X1 U6224 ( .A1(n5523), .A2(n7873), .ZN(n8365) );
  INV_X1 U6225 ( .A(n7911), .ZN(n5431) );
  OR2_X1 U6226 ( .A1(n8946), .A2(n6854), .ZN(n4856) );
  NOR3_X1 U6227 ( .A1(n7898), .A2(n7897), .A3(n7896), .ZN(n4857) );
  NAND2_X1 U6228 ( .A1(n5367), .A2(n5366), .ZN(n5383) );
  OR2_X1 U6229 ( .A1(n8757), .A2(n8760), .ZN(n4859) );
  AND2_X1 U6230 ( .A1(n5529), .A2(n5528), .ZN(n9831) );
  AND2_X2 U6231 ( .A1(n6631), .A2(n5493), .ZN(n9851) );
  AND2_X1 U6232 ( .A1(n7877), .A2(n7832), .ZN(n4860) );
  INV_X1 U6233 ( .A(n7206), .ZN(n6391) );
  INV_X1 U6234 ( .A(n7085), .ZN(n5866) );
  XNOR2_X1 U6235 ( .A(n5749), .B(n5747), .ZN(n7946) );
  INV_X1 U6236 ( .A(n7876), .ZN(n7833) );
  AOI21_X1 U6237 ( .B1(n7834), .B2(n4860), .A(n7833), .ZN(n7835) );
  INV_X1 U6238 ( .A(n8350), .ZN(n5577) );
  INV_X1 U6239 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4970) );
  AND2_X1 U6240 ( .A1(n4970), .A2(n4790), .ZN(n4971) );
  AND2_X1 U6241 ( .A1(n8758), .A2(n4844), .ZN(n8762) );
  INV_X1 U6242 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5643) );
  INV_X1 U6243 ( .A(n7484), .ZN(n5276) );
  INV_X1 U6244 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5652) );
  OR2_X1 U6245 ( .A1(n4926), .A2(SI_16_), .ZN(n4924) );
  NAND2_X1 U6246 ( .A1(n8260), .A2(n8130), .ZN(n6314) );
  INV_X1 U6247 ( .A(n5150), .ZN(n5002) );
  NOR2_X1 U6248 ( .A1(n8122), .A2(n8302), .ZN(n5449) );
  AND2_X1 U6249 ( .A1(n6187), .A2(n6186), .ZN(n6189) );
  NAND2_X1 U6250 ( .A1(n6209), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6230) );
  INV_X1 U6251 ( .A(n6020), .ZN(n5695) );
  OR2_X1 U6252 ( .A1(n6230), .A2(n9906), .ZN(n6271) );
  INV_X1 U6253 ( .A(n6197), .ZN(n6196) );
  NAND2_X1 U6254 ( .A1(n9247), .A2(n9262), .ZN(n6363) );
  INV_X1 U6255 ( .A(n5949), .ZN(n5694) );
  OR2_X1 U6256 ( .A1(n5757), .A2(n6897), .ZN(n6352) );
  INV_X1 U6257 ( .A(SI_17_), .ZN(n4929) );
  INV_X1 U6258 ( .A(n8142), .ZN(n5548) );
  NAND2_X1 U6259 ( .A1(n5552), .A2(n8140), .ZN(n5553) );
  NAND2_X1 U6260 ( .A1(n8038), .A2(n5600), .ZN(n5603) );
  INV_X1 U6261 ( .A(n9695), .ZN(n7261) );
  INV_X1 U6262 ( .A(n7850), .ZN(n7915) );
  OR2_X1 U6263 ( .A1(n5358), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5037) );
  INV_X1 U6264 ( .A(n5321), .ZN(n5012) );
  NAND2_X1 U6265 ( .A1(n5500), .A2(n7773), .ZN(n5501) );
  NAND2_X1 U6266 ( .A1(n5002), .A2(n5001), .ZN(n5165) );
  INV_X1 U6267 ( .A(n7737), .ZN(n5318) );
  OR2_X1 U6268 ( .A1(n7742), .A2(n7857), .ZN(n5628) );
  NAND2_X1 U6269 ( .A1(n5021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5022) );
  XNOR2_X1 U6270 ( .A(n5869), .B(n8529), .ZN(n5872) );
  OR2_X1 U6271 ( .A1(n5929), .A2(n5928), .ZN(n5949) );
  INV_X1 U6272 ( .A(n9384), .ZN(n6392) );
  AND2_X1 U6273 ( .A1(n6301), .A2(n6300), .ZN(n6227) );
  NAND2_X1 U6274 ( .A1(n6139), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6157) );
  OR2_X1 U6275 ( .A1(n6092), .A2(n7431), .ZN(n6105) );
  OR2_X1 U6276 ( .A1(n5775), .A2(n6892), .ZN(n5755) );
  OR2_X1 U6277 ( .A1(n7389), .A2(n7388), .ZN(n7386) );
  NAND2_X1 U6278 ( .A1(n9294), .A2(n6406), .ZN(n9279) );
  NOR2_X1 U6279 ( .A1(n7605), .A2(n6358), .ZN(n6359) );
  OR2_X1 U6280 ( .A1(n8945), .A2(n9566), .ZN(n6353) );
  OR2_X1 U6281 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  INV_X1 U6282 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6283 ( .A1(n4930), .A2(n4929), .ZN(n4933) );
  NAND2_X1 U6284 ( .A1(n5234), .A2(n4914), .ZN(n4917) );
  NAND2_X1 U6285 ( .A1(n5003), .A2(n8067), .ZN(n5200) );
  NAND2_X1 U6286 ( .A1(n8081), .A2(n5582), .ZN(n8024) );
  INV_X1 U6287 ( .A(n7499), .ZN(n5565) );
  INV_X1 U6288 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8067) );
  INV_X1 U6289 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7317) );
  OR2_X1 U6290 ( .A1(n5406), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6291 ( .A1(n5016), .A2(n5015), .ZN(n5358) );
  OR3_X1 U6292 ( .A1(n7683), .A2(n7682), .A3(n9768), .ZN(n7685) );
  NAND2_X1 U6293 ( .A1(n5008), .A2(n5007), .ZN(n5270) );
  OR2_X1 U6294 ( .A1(n5165), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6295 ( .A1(n5000), .A2(n4999), .ZN(n5133) );
  INV_X1 U6296 ( .A(n8131), .ZN(n8122) );
  INV_X1 U6297 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6347) );
  OR2_X1 U6298 ( .A1(n7743), .A2(n7930), .ZN(n9818) );
  OR2_X1 U6299 ( .A1(n6304), .A2(n5774), .ZN(n6218) );
  AND2_X1 U6300 ( .A1(n9521), .A2(n9520), .ZN(n9523) );
  AND2_X1 U6301 ( .A1(n7386), .A2(n7370), .ZN(n7371) );
  AND2_X1 U6302 ( .A1(n8921), .A2(n6265), .ZN(n8905) );
  INV_X1 U6303 ( .A(n6396), .ZN(n9068) );
  AND2_X1 U6304 ( .A1(n6441), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6264) );
  INV_X1 U6305 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5662) );
  INV_X1 U6306 ( .A(n8121), .ZN(n8107) );
  AOI22_X1 U6307 ( .A1(n6693), .A2(n6694), .B1(n6703), .B2(n5542), .ZN(n6643)
         );
  NAND2_X1 U6308 ( .A1(n7501), .A2(n5568), .ZN(n7583) );
  INV_X1 U6309 ( .A(n8052), .ZN(n8117) );
  OR2_X1 U6310 ( .A1(n7997), .A2(n5443), .ZN(n7726) );
  AND4_X1 U6311 ( .A1(n5340), .A2(n5339), .A3(n5338), .A4(n5337), .ZN(n8029)
         );
  INV_X1 U6312 ( .A(n9622), .ZN(n9750) );
  INV_X1 U6313 ( .A(n9664), .ZN(n9743) );
  AND2_X1 U6314 ( .A1(n5448), .A2(n7865), .ZN(n8360) );
  INV_X1 U6315 ( .A(n8372), .ZN(n8333) );
  INV_X1 U6316 ( .A(n8386), .ZN(n8413) );
  AND2_X1 U6317 ( .A1(n5492), .A2(n5491), .ZN(n5493) );
  INV_X1 U6318 ( .A(n9816), .ZN(n9828) );
  AND2_X1 U6319 ( .A1(n6437), .A2(n6493), .ZN(n6489) );
  INV_X1 U6320 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5086) );
  OR2_X1 U6321 ( .A1(n6295), .A2(n6427), .ZN(n9309) );
  OAI21_X1 U6322 ( .B1(n9112), .B2(n8610), .A(n6307), .ZN(n6308) );
  OR2_X1 U6323 ( .A1(n9135), .A2(n5774), .ZN(n6203) );
  AND4_X1 U6324 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n7529)
         );
  INV_X1 U6325 ( .A(n9522), .ZN(n9879) );
  AND2_X1 U6326 ( .A1(n6543), .A2(n6542), .ZN(n6611) );
  AND2_X1 U6327 ( .A1(n7442), .A2(n7441), .ZN(n7446) );
  AND2_X1 U6328 ( .A1(n9557), .A2(n8893), .ZN(n9229) );
  AND2_X1 U6329 ( .A1(n8880), .A2(n8881), .ZN(n9115) );
  INV_X1 U6330 ( .A(n9144), .ZN(n9142) );
  NOR2_X1 U6331 ( .A1(n6280), .A2(n6411), .ZN(n9298) );
  NAND2_X1 U6332 ( .A1(n6900), .A2(n6849), .ZN(n9545) );
  OAI21_X1 U6333 ( .B1(n6421), .B2(P1_D_REG_0__SCAN_IN), .A(n9443), .ZN(n6814)
         );
  NAND2_X1 U6334 ( .A1(n6848), .A2(n6861), .ZN(n9595) );
  MUX2_X1 U6335 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9449), .S(n5835), .Z(n9556) );
  INV_X1 U6336 ( .A(n6337), .ZN(n6440) );
  INV_X1 U6337 ( .A(n8268), .ZN(n8429) );
  AND2_X1 U6338 ( .A1(n5610), .A2(n5609), .ZN(n8052) );
  INV_X1 U6339 ( .A(n8072), .ZN(n8128) );
  INV_X1 U6340 ( .A(n6978), .ZN(n8141) );
  INV_X1 U6341 ( .A(n5104), .ZN(n8146) );
  OR2_X1 U6342 ( .A1(P2_U3150), .A2(n6450), .ZN(n9664) );
  INV_X1 U6343 ( .A(n9696), .ZN(n9766) );
  AND2_X2 U6344 ( .A1(n6636), .A2(n7996), .ZN(n8336) );
  NAND2_X1 U6345 ( .A1(n8366), .A2(n6710), .ZN(n8372) );
  NAND2_X1 U6346 ( .A1(n9851), .A2(n9828), .ZN(n8386) );
  NAND2_X1 U6347 ( .A1(n9851), .A2(n9808), .ZN(n8416) );
  INV_X1 U6348 ( .A(n9851), .ZN(n9848) );
  INV_X1 U6349 ( .A(n8021), .ZN(n8292) );
  NAND2_X1 U6350 ( .A1(n9829), .A2(n9808), .ZN(n8481) );
  INV_X2 U6351 ( .A(n9831), .ZN(n9829) );
  AND2_X1 U6352 ( .A1(n7422), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6493) );
  INV_X1 U6353 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7424) );
  INV_X1 U6354 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6787) );
  INV_X1 U6355 ( .A(n9668), .ZN(n7263) );
  NAND2_X1 U6356 ( .A1(n8536), .A2(n8535), .ZN(n8551) );
  INV_X1 U6357 ( .A(n9343), .ZN(n9127) );
  INV_X1 U6358 ( .A(n7107), .ZN(n9543) );
  AND2_X1 U6359 ( .A1(n6296), .A2(n9309), .ZN(n8610) );
  INV_X1 U6360 ( .A(n6308), .ZN(n6309) );
  INV_X1 U6361 ( .A(n9094), .ZN(n8934) );
  NAND2_X1 U6362 ( .A1(n6147), .A2(n6146), .ZN(n9194) );
  INV_X1 U6363 ( .A(n7050), .ZN(n8944) );
  NAND2_X1 U6364 ( .A1(n6543), .A2(n6541), .ZN(n9892) );
  INV_X1 U6365 ( .A(n9545), .ZN(n9290) );
  NAND2_X1 U6366 ( .A1(n9608), .A2(n9567), .ZN(n9401) );
  OR2_X1 U6367 ( .A1(n6432), .A2(n6814), .ZN(n9605) );
  INV_X1 U6368 ( .A(n9052), .ZN(n9405) );
  INV_X1 U6369 ( .A(n9308), .ZN(n9436) );
  OR2_X1 U6370 ( .A1(n6432), .A2(n6431), .ZN(n9589) );
  NAND2_X1 U6371 ( .A1(n6531), .A2(n6421), .ZN(n9550) );
  OR2_X1 U6372 ( .A1(n5996), .A2(n5995), .ZN(n7358) );
  INV_X1 U6373 ( .A(n5062), .ZN(n4863) );
  AND2_X1 U6374 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U6375 ( .A1(n4877), .A2(n4861), .ZN(n5721) );
  AND2_X1 U6376 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U6377 ( .A1(n4266), .A2(n4862), .ZN(n5072) );
  NAND2_X1 U6378 ( .A1(n5721), .A2(n5072), .ZN(n5063) );
  NAND2_X1 U6379 ( .A1(n4863), .A2(n5063), .ZN(n4866) );
  NAND2_X1 U6380 ( .A1(n4864), .A2(SI_1_), .ZN(n4865) );
  NAND2_X1 U6381 ( .A1(n4866), .A2(n4865), .ZN(n5082) );
  INV_X1 U6382 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6477) );
  INV_X1 U6383 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4867) );
  MUX2_X1 U6384 ( .A(n6477), .B(n4867), .S(n4877), .Z(n4868) );
  XNOR2_X1 U6385 ( .A(n4868), .B(SI_2_), .ZN(n5083) );
  NAND2_X1 U6386 ( .A1(n5082), .A2(n5083), .ZN(n4871) );
  INV_X1 U6387 ( .A(n4868), .ZN(n4869) );
  NAND2_X1 U6388 ( .A1(n4869), .A2(SI_2_), .ZN(n4870) );
  NAND2_X1 U6389 ( .A1(n4871), .A2(n4870), .ZN(n5101) );
  INV_X1 U6390 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9974) );
  INV_X1 U6391 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4872) );
  MUX2_X1 U6392 ( .A(n9974), .B(n4872), .S(n4877), .Z(n4873) );
  XNOR2_X1 U6393 ( .A(n4873), .B(SI_3_), .ZN(n5100) );
  NAND2_X1 U6394 ( .A1(n5101), .A2(n5100), .ZN(n4876) );
  INV_X1 U6395 ( .A(n4873), .ZN(n4874) );
  NAND2_X1 U6396 ( .A1(n4874), .A2(SI_3_), .ZN(n4875) );
  NAND2_X1 U6397 ( .A1(n4876), .A2(n4875), .ZN(n5116) );
  INV_X1 U6398 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6482) );
  INV_X1 U6399 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6480) );
  XNOR2_X1 U6400 ( .A(n4879), .B(SI_4_), .ZN(n5117) );
  NAND2_X1 U6401 ( .A1(n5116), .A2(n5117), .ZN(n4882) );
  INV_X1 U6402 ( .A(n4879), .ZN(n4880) );
  NAND2_X1 U6403 ( .A1(n4880), .A2(SI_4_), .ZN(n4881) );
  INV_X1 U6404 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6618) );
  INV_X1 U6405 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4883) );
  MUX2_X1 U6406 ( .A(n6618), .B(n4883), .S(n7731), .Z(n4884) );
  XNOR2_X1 U6407 ( .A(n4884), .B(SI_5_), .ZN(n5126) );
  INV_X1 U6408 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6409 ( .A1(n4885), .A2(SI_5_), .ZN(n4886) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6485) );
  INV_X1 U6411 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U6412 ( .A(n6485), .B(n6487), .S(n7731), .Z(n4888) );
  XNOR2_X1 U6413 ( .A(n4888), .B(SI_6_), .ZN(n5140) );
  INV_X1 U6414 ( .A(n4888), .ZN(n4889) );
  NAND2_X1 U6415 ( .A1(n4889), .A2(SI_6_), .ZN(n4890) );
  INV_X1 U6416 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U6417 ( .A(n6497), .B(n6495), .S(n7731), .Z(n4891) );
  XNOR2_X1 U6418 ( .A(n4891), .B(SI_7_), .ZN(n5159) );
  INV_X1 U6419 ( .A(n4891), .ZN(n4892) );
  MUX2_X1 U6420 ( .A(n6620), .B(n9991), .S(n7731), .Z(n4894) );
  INV_X1 U6421 ( .A(SI_8_), .ZN(n4893) );
  NAND2_X1 U6422 ( .A1(n4894), .A2(n4893), .ZN(n4897) );
  INV_X1 U6423 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6424 ( .A1(n4895), .A2(SI_8_), .ZN(n4896) );
  NAND2_X1 U6425 ( .A1(n4897), .A2(n4896), .ZN(n5173) );
  MUX2_X1 U6426 ( .A(n6622), .B(n6535), .S(n7731), .Z(n4900) );
  INV_X1 U6427 ( .A(SI_9_), .ZN(n4899) );
  NAND2_X1 U6428 ( .A1(n4900), .A2(n4899), .ZN(n4903) );
  INV_X1 U6429 ( .A(n4900), .ZN(n4901) );
  NAND2_X1 U6430 ( .A1(n4901), .A2(SI_9_), .ZN(n4902) );
  MUX2_X1 U6431 ( .A(n6540), .B(n6538), .S(n7731), .Z(n4904) );
  XNOR2_X1 U6432 ( .A(n4904), .B(SI_10_), .ZN(n5195) );
  INV_X1 U6433 ( .A(n4904), .ZN(n4905) );
  MUX2_X1 U6434 ( .A(n6624), .B(n9945), .S(n7731), .Z(n4907) );
  INV_X1 U6435 ( .A(SI_11_), .ZN(n4906) );
  INV_X1 U6436 ( .A(n4907), .ZN(n4908) );
  NAND2_X1 U6437 ( .A1(n4908), .A2(SI_11_), .ZN(n4909) );
  NAND2_X1 U6438 ( .A1(n4910), .A2(n4909), .ZN(n5208) );
  MUX2_X1 U6439 ( .A(n9963), .B(n6627), .S(n7731), .Z(n4911) );
  INV_X1 U6440 ( .A(n4911), .ZN(n4912) );
  MUX2_X1 U6441 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7731), .Z(n4915) );
  XNOR2_X1 U6442 ( .A(n4915), .B(SI_13_), .ZN(n5233) );
  INV_X1 U6443 ( .A(n5233), .ZN(n4914) );
  NAND2_X1 U6444 ( .A1(n4915), .A2(SI_13_), .ZN(n4916) );
  MUX2_X1 U6445 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7731), .Z(n4919) );
  XNOR2_X1 U6446 ( .A(n4919), .B(SI_14_), .ZN(n5246) );
  INV_X1 U6447 ( .A(n5246), .ZN(n4918) );
  NAND2_X1 U6448 ( .A1(n5247), .A2(n4918), .ZN(n4921) );
  NAND2_X1 U6449 ( .A1(n4919), .A2(SI_14_), .ZN(n4920) );
  MUX2_X1 U6450 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7731), .Z(n5263) );
  MUX2_X1 U6451 ( .A(n6787), .B(n6788), .S(n7731), .Z(n5280) );
  NAND2_X1 U6452 ( .A1(n4923), .A2(n4922), .ZN(n5278) );
  NAND2_X1 U6453 ( .A1(n4926), .A2(SI_16_), .ZN(n4927) );
  MUX2_X1 U6454 ( .A(n6792), .B(n9948), .S(n7731), .Z(n4930) );
  INV_X1 U6455 ( .A(n4930), .ZN(n4931) );
  NAND2_X1 U6456 ( .A1(n4931), .A2(SI_17_), .ZN(n4932) );
  NAND2_X1 U6457 ( .A1(n4933), .A2(n4932), .ZN(n5300) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n4934) );
  MUX2_X1 U6459 ( .A(n6870), .B(n4934), .S(n7731), .Z(n4935) );
  XNOR2_X1 U6460 ( .A(n4935), .B(SI_18_), .ZN(n5312) );
  INV_X1 U6461 ( .A(n5312), .ZN(n4938) );
  INV_X1 U6462 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6463 ( .A1(n4936), .A2(SI_18_), .ZN(n4937) );
  MUX2_X1 U6464 ( .A(n7957), .B(n6972), .S(n7731), .Z(n4940) );
  INV_X1 U6465 ( .A(SI_19_), .ZN(n4939) );
  NAND2_X1 U6466 ( .A1(n4940), .A2(n4939), .ZN(n4943) );
  INV_X1 U6467 ( .A(n4940), .ZN(n4941) );
  NAND2_X1 U6468 ( .A1(n4941), .A2(SI_19_), .ZN(n4942) );
  NAND2_X1 U6469 ( .A1(n4943), .A2(n4942), .ZN(n5046) );
  MUX2_X1 U6470 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7731), .Z(n5331) );
  INV_X1 U6471 ( .A(n5331), .ZN(n4944) );
  MUX2_X1 U6472 ( .A(n7176), .B(n7173), .S(n7731), .Z(n5343) );
  NOR2_X1 U6473 ( .A1(n4947), .A2(SI_21_), .ZN(n4949) );
  NAND2_X1 U6474 ( .A1(n4947), .A2(SI_21_), .ZN(n4948) );
  MUX2_X1 U6475 ( .A(n7383), .B(n7380), .S(n7731), .Z(n4951) );
  INV_X1 U6476 ( .A(SI_22_), .ZN(n4950) );
  NAND2_X1 U6477 ( .A1(n4951), .A2(n4950), .ZN(n4954) );
  INV_X1 U6478 ( .A(n4951), .ZN(n4952) );
  NAND2_X1 U6479 ( .A1(n4952), .A2(SI_22_), .ZN(n4953) );
  NAND2_X1 U6480 ( .A1(n4954), .A2(n4953), .ZN(n5352) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4955) );
  MUX2_X1 U6482 ( .A(n7424), .B(n4955), .S(n7731), .Z(n4957) );
  INV_X1 U6483 ( .A(SI_23_), .ZN(n4956) );
  NAND2_X1 U6484 ( .A1(n4957), .A2(n4956), .ZN(n4960) );
  INV_X1 U6485 ( .A(n4957), .ZN(n4958) );
  NAND2_X1 U6486 ( .A1(n4958), .A2(SI_23_), .ZN(n4959) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7511) );
  MUX2_X1 U6488 ( .A(n7515), .B(n7511), .S(n7731), .Z(n4962) );
  INV_X1 U6489 ( .A(SI_24_), .ZN(n4961) );
  NAND2_X1 U6490 ( .A1(n4962), .A2(n4961), .ZN(n5366) );
  INV_X1 U6491 ( .A(n4962), .ZN(n4963) );
  NAND2_X1 U6492 ( .A1(n4963), .A2(SI_24_), .ZN(n4964) );
  XNOR2_X1 U6493 ( .A(n5365), .B(n5364), .ZN(n7510) );
  NOR2_X1 U6494 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4968) );
  NAND4_X1 U6495 ( .A1(n4968), .A2(n4967), .A3(n4966), .A4(n4965), .ZN(n4969)
         );
  NAND2_X1 U6496 ( .A1(n5084), .A2(n5086), .ZN(n5097) );
  NAND2_X1 U6497 ( .A1(n5251), .A2(n5248), .ZN(n5051) );
  INV_X1 U6498 ( .A(n5051), .ZN(n4972) );
  NOR2_X1 U6499 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4974) );
  NAND4_X1 U6500 ( .A1(n4974), .A2(n4973), .A3(n5049), .A4(n5053), .ZN(n4975)
         );
  NOR2_X1 U6501 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4980) );
  INV_X1 U6502 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6503 ( .A1(n4991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4981) );
  INV_X1 U6504 ( .A(n4991), .ZN(n4985) );
  INV_X1 U6505 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6506 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4988) );
  AOI22_X1 U6507 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n8485), .B1(n4988), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6509 ( .A1(n7510), .A2(n7739), .ZN(n4997) );
  NAND2_X4 U6510 ( .A1(n5048), .A2(n7731), .ZN(n7737) );
  OR2_X1 U6511 ( .A1(n7737), .A2(n7515), .ZN(n4996) );
  NAND2_X1 U6512 ( .A1(n5091), .A2(n4998), .ZN(n5120) );
  INV_X1 U6513 ( .A(n5120), .ZN(n5000) );
  NAND2_X1 U6514 ( .A1(n7317), .A2(n7112), .ZN(n5004) );
  OR2_X2 U6515 ( .A1(n5225), .A2(n5004), .ZN(n5238) );
  INV_X1 U6516 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5009) );
  INV_X1 U6517 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5011) );
  INV_X1 U6518 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5013) );
  OR2_X2 U6519 ( .A1(n5347), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5356) );
  INV_X1 U6520 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5015) );
  OR2_X2 U6521 ( .A1(n5037), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6522 ( .A1(n5037), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6523 ( .A1(n5375), .A2(n5017), .ZN(n8281) );
  INV_X1 U6524 ( .A(n5020), .ZN(n5023) );
  NAND2_X1 U6525 ( .A1(n5023), .A2(n5022), .ZN(n5024) );
  NAND2_X1 U6526 ( .A1(n8281), .A2(n5213), .ZN(n5031) );
  INV_X1 U6527 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8435) );
  AND2_X2 U6528 ( .A1(n8491), .A2(n5026), .ZN(n5089) );
  NAND2_X1 U6529 ( .A1(n5408), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6530 ( .A1(n5164), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5027) );
  OAI211_X1 U6531 ( .C1(n6333), .C2(n8435), .A(n5028), .B(n5027), .ZN(n5029)
         );
  INV_X1 U6532 ( .A(n5029), .ZN(n5030) );
  INV_X1 U6533 ( .A(n8266), .ZN(n8133) );
  NAND2_X1 U6534 ( .A1(n7421), .A2(n7739), .ZN(n5035) );
  OR2_X1 U6535 ( .A1(n7737), .A2(n7424), .ZN(n5034) );
  NAND2_X1 U6536 ( .A1(n5358), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U6537 ( .A1(n5037), .A2(n5036), .ZN(n8290) );
  NAND2_X1 U6538 ( .A1(n8290), .A2(n5213), .ZN(n5040) );
  AOI22_X1 U6539 ( .A1(n5164), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5089), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6540 ( .A1(n4268), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5038) );
  INV_X1 U6541 ( .A(n8299), .ZN(n8134) );
  NAND2_X1 U6542 ( .A1(n5408), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6543 ( .A1(n4268), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U6544 ( .A1(n5323), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6545 ( .A1(n5335), .A2(n5041), .ZN(n7941) );
  NAND2_X1 U6546 ( .A1(n5213), .A2(n7941), .ZN(n5043) );
  NAND2_X1 U6547 ( .A1(n5164), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5042) );
  XNOR2_X1 U6548 ( .A(n5047), .B(n5046), .ZN(n6971) );
  NAND2_X1 U6549 ( .A1(n6971), .A2(n7739), .ZN(n5057) );
  NOR2_X1 U6550 ( .A1(n5051), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6551 ( .A1(n5314), .A2(n5053), .ZN(n5316) );
  INV_X1 U6552 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U6553 ( .A1(n5318), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6440), .B2(
        n8243), .ZN(n5056) );
  NAND2_X1 U6554 ( .A1(n4268), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6555 ( .A1(n5092), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6556 ( .A1(n5090), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6557 ( .A1(n5089), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5058) );
  XNOR2_X1 U6558 ( .A(n5062), .B(n5063), .ZN(n6474) );
  NAND2_X1 U6559 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5064) );
  XNOR2_X1 U6560 ( .A(n5064), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6510) );
  OR2_X1 U6561 ( .A1(n6337), .A2(n6510), .ZN(n5065) );
  NAND2_X1 U6562 ( .A1(n7721), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6563 ( .A1(n5089), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6564 ( .A1(n5092), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6565 ( .A1(n5090), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6566 ( .A1(n4266), .A2(SI_0_), .ZN(n5071) );
  INV_X1 U6567 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6568 ( .A1(n5071), .A2(n5070), .ZN(n5073) );
  AND2_X1 U6569 ( .A1(n5073), .A2(n5072), .ZN(n8496) );
  MUX2_X1 U6570 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8496), .S(n6337), .Z(n9771) );
  NAND2_X1 U6571 ( .A1(n8149), .A2(n9771), .ZN(n6656) );
  NAND2_X1 U6572 ( .A1(n7881), .A2(n6656), .ZN(n5077) );
  NAND2_X1 U6573 ( .A1(n7703), .A2(n5075), .ZN(n5076) );
  NAND2_X1 U6574 ( .A1(n5089), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6575 ( .A1(n7721), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6576 ( .A1(n5092), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6577 ( .A1(n5090), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U6578 ( .A(n5082), .B(n5083), .ZN(n6476) );
  OR2_X1 U6579 ( .A1(n5160), .A2(n6476), .ZN(n5088) );
  OR2_X1 U6580 ( .A1(n6337), .A2(n6525), .ZN(n5087) );
  XNOR2_X1 U6581 ( .A(n8147), .B(n9773), .ZN(n6731) );
  INV_X1 U6582 ( .A(n8147), .ZN(n6703) );
  NAND2_X1 U6583 ( .A1(n6703), .A2(n9773), .ZN(n6719) );
  NAND2_X1 U6584 ( .A1(n5089), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6585 ( .A1(n5090), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6586 ( .A1(n7721), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6587 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND2_X1 U6588 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5099) );
  INV_X1 U6589 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5098) );
  XNOR2_X1 U6590 ( .A(n5099), .B(n5098), .ZN(n6597) );
  OR2_X1 U6591 ( .A1(n5160), .A2(n6475), .ZN(n5102) );
  NAND2_X1 U6592 ( .A1(n6732), .A2(n9778), .ZN(n5105) );
  AND2_X1 U6593 ( .A1(n6719), .A2(n5105), .ZN(n5108) );
  NAND2_X1 U6594 ( .A1(n5104), .A2(n6724), .ZN(n7764) );
  INV_X1 U6596 ( .A(n5105), .ZN(n5106) );
  NOR2_X1 U6597 ( .A1(n7880), .A2(n5106), .ZN(n5107) );
  NAND2_X1 U6598 ( .A1(n5164), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6599 ( .A1(n5089), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5112) );
  INV_X2 U6600 ( .A(n5443), .ZN(n5213) );
  NAND2_X1 U6601 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5109) );
  NAND2_X1 U6602 ( .A1(n5120), .A2(n5109), .ZN(n6714) );
  NAND2_X1 U6603 ( .A1(n5213), .A2(n6714), .ZN(n5111) );
  NAND2_X1 U6604 ( .A1(n7721), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5110) );
  AND4_X2 U6605 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n6759)
         );
  NAND2_X1 U6606 ( .A1(n5127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5115) );
  INV_X1 U6607 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6608 ( .A(n5115), .B(n5114), .ZN(n7270) );
  XNOR2_X1 U6609 ( .A(n5116), .B(n5117), .ZN(n6481) );
  OR2_X1 U6610 ( .A1(n5160), .A2(n6481), .ZN(n5119) );
  OR2_X1 U6611 ( .A1(n7737), .A2(n6482), .ZN(n5118) );
  OAI211_X1 U6612 ( .C1(n6337), .C2(n7270), .A(n5119), .B(n5118), .ZN(n6715)
         );
  NAND2_X1 U6613 ( .A1(n5089), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6614 ( .A1(n5164), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6615 ( .A1(n5120), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6616 ( .A1(n5133), .A2(n5121), .ZN(n6762) );
  NAND2_X1 U6617 ( .A1(n5213), .A2(n6762), .ZN(n5123) );
  NAND2_X1 U6618 ( .A1(n7721), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5122) );
  OR2_X1 U6619 ( .A1(n5160), .A2(n6484), .ZN(n5131) );
  OR2_X1 U6620 ( .A1(n7737), .A2(n6618), .ZN(n5130) );
  OR2_X1 U6621 ( .A1(n5142), .A2(n8485), .ZN(n5128) );
  XNOR2_X1 U6622 ( .A(n5128), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9627) );
  INV_X1 U6623 ( .A(n9627), .ZN(n7242) );
  OR2_X1 U6624 ( .A1(n6337), .A2(n7242), .ZN(n5129) );
  NAND2_X1 U6625 ( .A1(n6687), .A2(n9788), .ZN(n6750) );
  INV_X1 U6626 ( .A(n9788), .ZN(n6761) );
  NAND2_X1 U6627 ( .A1(n8144), .A2(n6761), .ZN(n6749) );
  NAND2_X1 U6628 ( .A1(n5132), .A2(n6749), .ZN(n6772) );
  NAND2_X1 U6629 ( .A1(n5089), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6630 ( .A1(n5164), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6631 ( .A1(n5133), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6632 ( .A1(n5150), .A2(n5134), .ZN(n6768) );
  NAND2_X1 U6633 ( .A1(n5213), .A2(n6768), .ZN(n5136) );
  NAND2_X1 U6634 ( .A1(n7721), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5135) );
  XNOR2_X1 U6635 ( .A(n5139), .B(n5140), .ZN(n6486) );
  OR2_X1 U6636 ( .A1(n5160), .A2(n6486), .ZN(n5146) );
  OR2_X1 U6637 ( .A1(n7737), .A2(n6485), .ZN(n5145) );
  INV_X1 U6638 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6639 ( .A1(n5142), .A2(n5141), .ZN(n5156) );
  NAND2_X1 U6640 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5143) );
  XNOR2_X1 U6641 ( .A(n5143), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9643) );
  OR2_X1 U6642 ( .A1(n6337), .A2(n7275), .ZN(n5144) );
  NAND2_X1 U6643 ( .A1(n6874), .A2(n9794), .ZN(n5147) );
  NAND2_X1 U6644 ( .A1(n6772), .A2(n5147), .ZN(n5149) );
  INV_X1 U6645 ( .A(n9794), .ZN(n6770) );
  NAND2_X1 U6646 ( .A1(n8143), .A2(n6770), .ZN(n5148) );
  NAND2_X1 U6647 ( .A1(n5149), .A2(n5148), .ZN(n6872) );
  INV_X1 U6648 ( .A(n6872), .ZN(n5163) );
  NAND2_X1 U6649 ( .A1(n5408), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U6650 ( .A1(n5150), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6651 ( .A1(n5165), .A2(n5151), .ZN(n6877) );
  NAND2_X1 U6652 ( .A1(n5213), .A2(n6877), .ZN(n5154) );
  NAND2_X1 U6653 ( .A1(n5164), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6654 ( .A1(n7721), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6655 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n8142)
         );
  NAND2_X1 U6656 ( .A1(n5171), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  XNOR2_X1 U6657 ( .A(n5157), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9660) );
  XNOR2_X1 U6658 ( .A(n5158), .B(n5159), .ZN(n6496) );
  OR2_X1 U6659 ( .A1(n5160), .A2(n6496), .ZN(n5162) );
  OR2_X1 U6660 ( .A1(n7737), .A2(n6497), .ZN(n5161) );
  OAI211_X1 U6661 ( .C1(n6337), .C2(n7265), .A(n5162), .B(n5161), .ZN(n6881)
         );
  XNOR2_X1 U6662 ( .A(n8142), .B(n6881), .ZN(n7768) );
  NAND2_X1 U6663 ( .A1(n5163), .A2(n7890), .ZN(n6905) );
  NAND2_X1 U6664 ( .A1(n5164), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6665 ( .A1(n5408), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6666 ( .A1(n5165), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6667 ( .A1(n5185), .A2(n5166), .ZN(n6919) );
  NAND2_X1 U6668 ( .A1(n5213), .A2(n6919), .ZN(n5168) );
  NAND2_X1 U6669 ( .A1(n7721), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6670 ( .A1(n5180), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  XNOR2_X1 U6671 ( .A(n5172), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9668) );
  XNOR2_X1 U6672 ( .A(n5174), .B(n5173), .ZN(n6500) );
  NAND2_X1 U6673 ( .A1(n6500), .A2(n7739), .ZN(n5176) );
  OR2_X1 U6674 ( .A1(n7737), .A2(n6620), .ZN(n5175) );
  OAI211_X1 U6675 ( .C1(n6337), .C2(n7263), .A(n5176), .B(n5175), .ZN(n6911)
         );
  NAND2_X1 U6676 ( .A1(n6978), .A2(n6911), .ZN(n7772) );
  INV_X1 U6677 ( .A(n6911), .ZN(n9805) );
  NAND2_X1 U6678 ( .A1(n8141), .A2(n9805), .ZN(n7773) );
  NAND2_X1 U6679 ( .A1(n7772), .A2(n7773), .ZN(n7889) );
  INV_X1 U6680 ( .A(n6881), .ZN(n9798) );
  NAND2_X1 U6681 ( .A1(n5548), .A2(n9798), .ZN(n6904) );
  AND2_X1 U6682 ( .A1(n7889), .A2(n6904), .ZN(n5177) );
  NAND2_X1 U6683 ( .A1(n6905), .A2(n5177), .ZN(n6903) );
  NAND2_X1 U6684 ( .A1(n8141), .A2(n6911), .ZN(n5178) );
  NAND2_X1 U6685 ( .A1(n6903), .A2(n5178), .ZN(n6976) );
  NAND2_X1 U6686 ( .A1(n6534), .A2(n7739), .ZN(n5184) );
  OAI21_X1 U6687 ( .B1(n5180), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5182) );
  INV_X1 U6688 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U6689 ( .A(n5182), .B(n5181), .ZN(n9695) );
  AOI22_X1 U6690 ( .A1(n5318), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6440), .B2(
        n7261), .ZN(n5183) );
  NAND2_X1 U6691 ( .A1(n5164), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6692 ( .A1(n5408), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6693 ( .A1(n5185), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6694 ( .A1(n5200), .A2(n5186), .ZN(n8074) );
  NAND2_X1 U6695 ( .A1(n5213), .A2(n8074), .ZN(n5188) );
  NAND2_X1 U6696 ( .A1(n7721), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6697 ( .A1(n9810), .A2(n7027), .ZN(n5191) );
  NAND2_X1 U6698 ( .A1(n6976), .A2(n5191), .ZN(n5193) );
  INV_X1 U6699 ( .A(n9810), .ZN(n8073) );
  INV_X1 U6700 ( .A(n7027), .ZN(n8140) );
  NAND2_X1 U6701 ( .A1(n8073), .A2(n8140), .ZN(n5192) );
  NAND2_X1 U6702 ( .A1(n5193), .A2(n5192), .ZN(n7026) );
  XNOR2_X1 U6703 ( .A(n5194), .B(n5195), .ZN(n6537) );
  NAND2_X1 U6704 ( .A1(n6537), .A2(n7739), .ZN(n5199) );
  OR2_X1 U6705 ( .A1(n5196), .A2(n8485), .ZN(n5197) );
  XNOR2_X1 U6706 ( .A(n5197), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9697) );
  AOI22_X1 U6707 ( .A1(n5318), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6440), .B2(
        n9697), .ZN(n5198) );
  NAND2_X1 U6708 ( .A1(n5199), .A2(n5198), .ZN(n7035) );
  NAND2_X1 U6709 ( .A1(n5408), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6710 ( .A1(n5200), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6711 ( .A1(n5225), .A2(n5201), .ZN(n7220) );
  NAND2_X1 U6712 ( .A1(n5213), .A2(n7220), .ZN(n5204) );
  NAND2_X1 U6713 ( .A1(n7721), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6714 ( .A1(n5164), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5202) );
  NAND4_X1 U6715 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n8139)
         );
  OR2_X1 U6716 ( .A1(n7035), .A2(n8139), .ZN(n7025) );
  NAND2_X1 U6717 ( .A1(n7026), .A2(n7025), .ZN(n5206) );
  NAND2_X1 U6718 ( .A1(n7035), .A2(n8139), .ZN(n7024) );
  NAND2_X1 U6719 ( .A1(n5206), .A2(n7024), .ZN(n7017) );
  XNOR2_X1 U6720 ( .A(n5207), .B(n5208), .ZN(n6606) );
  NAND2_X1 U6721 ( .A1(n6606), .A2(n7739), .ZN(n5212) );
  NAND2_X1 U6722 ( .A1(n5209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U6723 ( .A(n5210), .B(n5049), .ZN(n9726) );
  INV_X1 U6724 ( .A(n9726), .ZN(n7257) );
  AOI22_X1 U6725 ( .A1(n5318), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6440), .B2(
        n7257), .ZN(n5211) );
  NAND2_X1 U6726 ( .A1(n5212), .A2(n5211), .ZN(n9827) );
  NAND2_X1 U6727 ( .A1(n5408), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6728 ( .A1(n5164), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6729 ( .A(n5225), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U6730 ( .A1(n5213), .A2(n7318), .ZN(n5215) );
  NAND2_X1 U6731 ( .A1(n7721), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6732 ( .A1(n9827), .A2(n7217), .ZN(n7788) );
  NAND2_X1 U6733 ( .A1(n7784), .A2(n7788), .ZN(n7012) );
  INV_X1 U6734 ( .A(n7217), .ZN(n8138) );
  NAND2_X1 U6735 ( .A1(n9827), .A2(n8138), .ZN(n5218) );
  XNOR2_X1 U6736 ( .A(n5220), .B(n5219), .ZN(n6626) );
  NAND2_X1 U6737 ( .A1(n6626), .A2(n7739), .ZN(n5224) );
  NAND2_X1 U6738 ( .A1(n5221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5222) );
  XNOR2_X1 U6739 ( .A(n5222), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7548) );
  AOI22_X1 U6740 ( .A1(n5318), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6440), .B2(
        n7548), .ZN(n5223) );
  NAND2_X1 U6741 ( .A1(n5164), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6742 ( .A1(n5408), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5229) );
  OAI21_X1 U6743 ( .B1(n5225), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6744 ( .A1(n5226), .A2(n5238), .ZN(n7179) );
  NAND2_X1 U6745 ( .A1(n5213), .A2(n7179), .ZN(n5228) );
  NAND2_X1 U6746 ( .A1(n7721), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5227) );
  NAND4_X1 U6747 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n8137)
         );
  AND2_X1 U6748 ( .A1(n7790), .A2(n8137), .ZN(n5232) );
  OR2_X1 U6749 ( .A1(n7790), .A2(n8137), .ZN(n5231) );
  XNOR2_X1 U6750 ( .A(n5234), .B(n5233), .ZN(n6652) );
  NAND2_X1 U6751 ( .A1(n6652), .A2(n7739), .ZN(n5237) );
  OR2_X1 U6752 ( .A1(n5235), .A2(n8485), .ZN(n5249) );
  XNOR2_X1 U6753 ( .A(n5249), .B(n5248), .ZN(n9741) );
  INV_X1 U6754 ( .A(n9741), .ZN(n7556) );
  AOI22_X1 U6755 ( .A1(n5318), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6440), .B2(
        n7556), .ZN(n5236) );
  NAND2_X1 U6756 ( .A1(n5164), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6757 ( .A1(n5408), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6758 ( .A1(n5238), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6759 ( .A1(n5256), .A2(n5239), .ZN(n7453) );
  NAND2_X1 U6760 ( .A1(n5213), .A2(n7453), .ZN(n5241) );
  NAND2_X1 U6761 ( .A1(n7721), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6762 ( .A1(n7351), .A2(n7464), .ZN(n7798) );
  NAND2_X1 U6763 ( .A1(n7797), .A2(n7798), .ZN(n7898) );
  OR2_X1 U6764 ( .A1(n7351), .A2(n8136), .ZN(n5244) );
  XNOR2_X1 U6765 ( .A(n5247), .B(n5246), .ZN(n6707) );
  NAND2_X1 U6766 ( .A1(n6707), .A2(n7739), .ZN(n5255) );
  NAND2_X1 U6767 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NAND2_X1 U6768 ( .A1(n5250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6769 ( .A1(n5252), .A2(n5251), .ZN(n5266) );
  OR2_X1 U6770 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  AOI22_X1 U6771 ( .A1(n5318), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6440), .B2(
        n9754), .ZN(n5254) );
  NAND2_X1 U6772 ( .A1(n5255), .A2(n5254), .ZN(n7410) );
  NAND2_X1 U6773 ( .A1(n5164), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6774 ( .A1(n5408), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6775 ( .A1(n5256), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6776 ( .A1(n5270), .A2(n5257), .ZN(n7466) );
  NAND2_X1 U6777 ( .A1(n5092), .A2(n7466), .ZN(n5259) );
  NAND2_X1 U6778 ( .A1(n4268), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6779 ( .A1(n7410), .A2(n7504), .ZN(n7800) );
  NAND2_X1 U6780 ( .A1(n7410), .A2(n7504), .ZN(n7801) );
  NAND2_X1 U6781 ( .A1(n7410), .A2(n8135), .ZN(n5262) );
  NAND2_X1 U6782 ( .A1(n7413), .A2(n5262), .ZN(n7486) );
  INV_X1 U6783 ( .A(n7486), .ZN(n5277) );
  XNOR2_X1 U6784 ( .A(n5263), .B(SI_15_), .ZN(n5264) );
  XNOR2_X1 U6785 ( .A(n5265), .B(n5264), .ZN(n6745) );
  NAND2_X1 U6786 ( .A1(n6745), .A2(n7739), .ZN(n5269) );
  NAND2_X1 U6787 ( .A1(n5266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5267) );
  XNOR2_X1 U6788 ( .A(n5267), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8151) );
  AOI22_X1 U6789 ( .A1(n5318), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6440), .B2(
        n8151), .ZN(n5268) );
  NAND2_X1 U6790 ( .A1(n5408), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6791 ( .A1(n5270), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6792 ( .A1(n5289), .A2(n5271), .ZN(n7506) );
  NAND2_X1 U6793 ( .A1(n5213), .A2(n7506), .ZN(n5274) );
  NAND2_X1 U6794 ( .A1(n5164), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5273) );
  NAND2_X1 U6795 ( .A1(n7721), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5272) );
  NAND4_X1 U6796 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n8361)
         );
  AND2_X1 U6797 ( .A1(n7498), .A2(n8361), .ZN(n7484) );
  NAND2_X1 U6798 ( .A1(n5277), .A2(n5276), .ZN(n8357) );
  NAND2_X1 U6799 ( .A1(n5279), .A2(n5278), .ZN(n5282) );
  XNOR2_X1 U6800 ( .A(n5280), .B(SI_16_), .ZN(n5281) );
  NAND2_X1 U6801 ( .A1(n6786), .A2(n7739), .ZN(n5288) );
  NAND2_X1 U6802 ( .A1(n5283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5284) );
  MUX2_X1 U6803 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5284), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5286) );
  AND2_X1 U6804 ( .A1(n5286), .A2(n5285), .ZN(n8181) );
  AOI22_X1 U6805 ( .A1(n5318), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6440), .B2(
        n8181), .ZN(n5287) );
  NAND2_X1 U6806 ( .A1(n5164), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6807 ( .A1(n5408), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6808 ( .A1(n5289), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6809 ( .A1(n5305), .A2(n5290), .ZN(n8367) );
  NAND2_X1 U6810 ( .A1(n5213), .A2(n8367), .ZN(n5292) );
  NAND2_X1 U6811 ( .A1(n4268), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6812 ( .A1(n8478), .A2(n5297), .ZN(n7812) );
  INV_X1 U6813 ( .A(n8359), .ZN(n5295) );
  OR2_X1 U6814 ( .A1(n7498), .A2(n8361), .ZN(n8356) );
  AND2_X1 U6815 ( .A1(n5295), .A2(n8356), .ZN(n5296) );
  NAND2_X1 U6816 ( .A1(n8478), .A2(n8349), .ZN(n5298) );
  XNOR2_X1 U6817 ( .A(n5301), .B(n5300), .ZN(n6790) );
  NAND2_X1 U6818 ( .A1(n6790), .A2(n7739), .ZN(n5304) );
  NAND2_X1 U6819 ( .A1(n5285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6820 ( .A(n5302), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8210) );
  AOI22_X1 U6821 ( .A1(n5318), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6440), .B2(
        n8210), .ZN(n5303) );
  NAND2_X1 U6822 ( .A1(n5408), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6823 ( .A1(n7721), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6824 ( .A1(n5305), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6825 ( .A1(n5321), .A2(n5306), .ZN(n8352) );
  NAND2_X1 U6826 ( .A1(n5213), .A2(n8352), .ZN(n5308) );
  NAND2_X1 U6827 ( .A1(n5164), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6828 ( .A1(n8471), .A2(n8110), .ZN(n7810) );
  NAND2_X1 U6829 ( .A1(n7811), .A2(n7810), .ZN(n8347) );
  INV_X1 U6830 ( .A(n8110), .ZN(n8363) );
  AND2_X1 U6831 ( .A1(n8471), .A2(n8363), .ZN(n5311) );
  XNOR2_X1 U6832 ( .A(n5313), .B(n5312), .ZN(n6810) );
  NAND2_X1 U6833 ( .A1(n6810), .A2(n7739), .ZN(n5320) );
  INV_X1 U6834 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6835 ( .A1(n5315), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5317) );
  AND2_X1 U6836 ( .A1(n5317), .A2(n5316), .ZN(n8220) );
  AOI22_X1 U6837 ( .A1(n5318), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6440), .B2(
        n8220), .ZN(n5319) );
  NAND2_X1 U6838 ( .A1(n5408), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6839 ( .A1(n5321), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6840 ( .A1(n5323), .A2(n5322), .ZN(n8343) );
  NAND2_X1 U6841 ( .A1(n5213), .A2(n8343), .ZN(n5326) );
  NAND2_X1 U6842 ( .A1(n5164), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6843 ( .A1(n7721), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5324) );
  NAND4_X1 U6844 ( .A1(n5327), .A2(n5326), .A3(n5325), .A4(n5324), .ZN(n8350)
         );
  NOR2_X1 U6845 ( .A1(n8465), .A2(n8350), .ZN(n5328) );
  NAND2_X1 U6846 ( .A1(n8458), .A2(n8085), .ZN(n7813) );
  NAND2_X1 U6847 ( .A1(n8324), .A2(n7813), .ZN(n7903) );
  XNOR2_X1 U6848 ( .A(n5331), .B(n5330), .ZN(n5332) );
  XNOR2_X1 U6849 ( .A(n5329), .B(n5332), .ZN(n7061) );
  NAND2_X1 U6850 ( .A1(n7061), .A2(n7739), .ZN(n5334) );
  INV_X1 U6851 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7063) );
  OR2_X1 U6852 ( .A1(n7737), .A2(n7063), .ZN(n5333) );
  NAND2_X1 U6853 ( .A1(n5164), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6854 ( .A1(n5408), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6855 ( .A1(n5335), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6856 ( .A1(n5347), .A2(n5336), .ZN(n8328) );
  NAND2_X1 U6857 ( .A1(n5213), .A2(n8328), .ZN(n5338) );
  NAND2_X1 U6858 ( .A1(n7721), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5337) );
  OR2_X1 U6859 ( .A1(n8399), .A2(n8029), .ZN(n7819) );
  NAND2_X1 U6860 ( .A1(n8399), .A2(n8029), .ZN(n7818) );
  NAND2_X1 U6861 ( .A1(n7819), .A2(n7818), .ZN(n8320) );
  XNOR2_X1 U6862 ( .A(n5343), .B(SI_21_), .ZN(n5344) );
  XNOR2_X1 U6863 ( .A(n5342), .B(n5344), .ZN(n7172) );
  NAND2_X1 U6864 ( .A1(n7172), .A2(n7739), .ZN(n5346) );
  OR2_X1 U6865 ( .A1(n7737), .A2(n7176), .ZN(n5345) );
  NAND2_X1 U6866 ( .A1(n5347), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6867 ( .A1(n5356), .A2(n5348), .ZN(n8316) );
  AOI22_X1 U6868 ( .A1(n8316), .A2(n5213), .B1(n4268), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5350) );
  AOI22_X1 U6869 ( .A1(n5164), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5089), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6870 ( .A1(n8448), .A2(n8301), .ZN(n7823) );
  NAND2_X1 U6871 ( .A1(n7822), .A2(n7823), .ZN(n8310) );
  INV_X1 U6872 ( .A(n8448), .ZN(n8033) );
  NAND2_X1 U6873 ( .A1(n7379), .A2(n7739), .ZN(n5355) );
  OR2_X1 U6874 ( .A1(n7737), .A2(n7383), .ZN(n5354) );
  NAND2_X1 U6875 ( .A1(n5356), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6876 ( .A1(n5358), .A2(n5357), .ZN(n8303) );
  NAND2_X1 U6877 ( .A1(n8303), .A2(n5213), .ZN(n5361) );
  AOI22_X1 U6878 ( .A1(n5164), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n5089), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6879 ( .A1(n7721), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6880 ( .A1(n8442), .A2(n7694), .ZN(n7826) );
  AOI21_X1 U6881 ( .B1(n8292), .B2(n8299), .A(n7692), .ZN(n5362) );
  OAI21_X1 U6882 ( .B1(n8266), .B2(n8387), .A(n8277), .ZN(n5363) );
  NAND2_X1 U6883 ( .A1(n5365), .A2(n5364), .ZN(n5367) );
  INV_X1 U6884 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7594) );
  INV_X1 U6885 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7590) );
  MUX2_X1 U6886 ( .A(n7594), .B(n7590), .S(n7731), .Z(n5368) );
  INV_X1 U6887 ( .A(SI_25_), .ZN(n10012) );
  NAND2_X1 U6888 ( .A1(n5368), .A2(n10012), .ZN(n5384) );
  INV_X1 U6889 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6890 ( .A1(n5369), .A2(SI_25_), .ZN(n5370) );
  XNOR2_X1 U6891 ( .A(n5383), .B(n5382), .ZN(n7589) );
  NAND2_X1 U6892 ( .A1(n7589), .A2(n7739), .ZN(n5372) );
  OR2_X1 U6893 ( .A1(n7737), .A2(n7594), .ZN(n5371) );
  INV_X1 U6894 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6895 ( .A1(n5375), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6896 ( .A1(n5390), .A2(n5376), .ZN(n8270) );
  NAND2_X1 U6897 ( .A1(n8270), .A2(n5213), .ZN(n5381) );
  INV_X1 U6898 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10010) );
  NAND2_X1 U6899 ( .A1(n5164), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6900 ( .A1(n5408), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5377) );
  OAI211_X1 U6901 ( .C1(n10010), .C2(n6333), .A(n5378), .B(n5377), .ZN(n5379)
         );
  INV_X1 U6902 ( .A(n5379), .ZN(n5380) );
  NAND2_X1 U6903 ( .A1(n8268), .A2(n8279), .ZN(n7838) );
  NAND2_X1 U6904 ( .A1(n7837), .A2(n7838), .ZN(n8271) );
  NAND2_X1 U6905 ( .A1(n5383), .A2(n5382), .ZN(n5385) );
  INV_X1 U6906 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7610) );
  INV_X1 U6907 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9964) );
  MUX2_X1 U6908 ( .A(n7610), .B(n9964), .S(n7731), .Z(n5387) );
  INV_X1 U6909 ( .A(SI_26_), .ZN(n5386) );
  NAND2_X1 U6910 ( .A1(n5387), .A2(n5386), .ZN(n5415) );
  INV_X1 U6911 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U6912 ( .A1(n5388), .A2(SI_26_), .ZN(n5389) );
  NAND2_X1 U6913 ( .A1(n5390), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6914 ( .A1(n5406), .A2(n5391), .ZN(n8125) );
  NAND2_X1 U6915 ( .A1(n8125), .A2(n5213), .ZN(n5396) );
  INV_X1 U6916 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U6917 ( .A1(n5164), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6918 ( .A1(n5408), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5392) );
  OAI211_X1 U6919 ( .C1(n7986), .C2(n6333), .A(n5393), .B(n5392), .ZN(n5394)
         );
  INV_X1 U6920 ( .A(n5394), .ZN(n5395) );
  NAND2_X1 U6921 ( .A1(n5417), .A2(n5415), .ZN(n5403) );
  INV_X1 U6922 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9972) );
  INV_X1 U6923 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10020) );
  MUX2_X1 U6924 ( .A(n9972), .B(n10020), .S(n7731), .Z(n5400) );
  INV_X1 U6925 ( .A(SI_27_), .ZN(n5399) );
  NAND2_X1 U6926 ( .A1(n5400), .A2(n5399), .ZN(n5414) );
  INV_X1 U6927 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6928 ( .A1(n5401), .A2(SI_27_), .ZN(n6316) );
  AND2_X1 U6929 ( .A1(n5414), .A2(n6316), .ZN(n5402) );
  NAND2_X1 U6930 ( .A1(n7640), .A2(n7739), .ZN(n5405) );
  OR2_X1 U6931 ( .A1(n7737), .A2(n9972), .ZN(n5404) );
  NAND2_X1 U6932 ( .A1(n5406), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6933 ( .A1(n5423), .A2(n5407), .ZN(n8008) );
  NAND2_X1 U6934 ( .A1(n8008), .A2(n5213), .ZN(n5413) );
  INV_X1 U6935 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U6936 ( .A1(n5164), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6937 ( .A1(n5408), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U6938 ( .C1(n7970), .C2(n6333), .A(n5410), .B(n5409), .ZN(n5411)
         );
  INV_X1 U6939 ( .A(n5411), .ZN(n5412) );
  NAND2_X2 U6940 ( .A1(n5413), .A2(n5412), .ZN(n8131) );
  INV_X1 U6941 ( .A(n7978), .ZN(n8015) );
  AND2_X1 U6942 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7680) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7963) );
  MUX2_X1 U6945 ( .A(n7680), .B(n7963), .S(n7731), .Z(n6321) );
  XNOR2_X1 U6946 ( .A(n6321), .B(SI_28_), .ZN(n6317) );
  NAND2_X1 U6947 ( .A1(n7961), .A2(n7739), .ZN(n5420) );
  OR2_X1 U6948 ( .A1(n7737), .A2(n7680), .ZN(n5419) );
  INV_X1 U6949 ( .A(n5423), .ZN(n5422) );
  INV_X1 U6950 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6951 ( .A1(n5422), .A2(n5421), .ZN(n7997) );
  NAND2_X1 U6952 ( .A1(n5423), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6953 ( .A1(n7997), .A2(n5424), .ZN(n8259) );
  NAND2_X1 U6954 ( .A1(n8259), .A2(n5213), .ZN(n5430) );
  INV_X1 U6955 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6956 ( .A1(n5164), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6957 ( .A1(n5408), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5425) );
  OAI211_X1 U6958 ( .C1(n5427), .C2(n6333), .A(n5426), .B(n5425), .ZN(n5428)
         );
  INV_X1 U6959 ( .A(n5428), .ZN(n5429) );
  XNOR2_X1 U6960 ( .A(n7854), .B(n8130), .ZN(n7911) );
  XNOR2_X1 U6961 ( .A(n6313), .B(n5431), .ZN(n5442) );
  NAND2_X1 U6962 ( .A1(n5474), .A2(n5432), .ZN(n5438) );
  NAND2_X1 U6963 ( .A1(n5438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6964 ( .A1(n8243), .A2(n7930), .ZN(n5523) );
  NAND2_X1 U6965 ( .A1(n5474), .A2(n5435), .ZN(n5436) );
  NAND2_X1 U6966 ( .A1(n5436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5437) );
  MUX2_X1 U6967 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5437), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5439) );
  INV_X1 U6968 ( .A(n5474), .ZN(n5440) );
  NAND2_X1 U6969 ( .A1(n5440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5441) );
  INV_X1 U6970 ( .A(n7062), .ZN(n5522) );
  NAND2_X1 U6971 ( .A1(n7747), .A2(n5522), .ZN(n7873) );
  NAND2_X1 U6972 ( .A1(n5442), .A2(n8365), .ZN(n5452) );
  NAND2_X1 U6973 ( .A1(n5164), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6974 ( .A1(n5408), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5444) );
  OAI211_X1 U6975 ( .C1(n6347), .C2(n6333), .A(n5445), .B(n5444), .ZN(n5446)
         );
  INV_X1 U6976 ( .A(n5446), .ZN(n5447) );
  INV_X1 U6977 ( .A(n5619), .ZN(n5448) );
  NAND2_X1 U6978 ( .A1(n5452), .A2(n5451), .ZN(n8255) );
  NAND2_X1 U6979 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  AND2_X1 U6980 ( .A1(n5453), .A2(n5457), .ZN(n5458) );
  NAND2_X1 U6981 ( .A1(n5474), .A2(n5458), .ZN(n5460) );
  XNOR2_X1 U6982 ( .A(n7513), .B(P2_B_REG_SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6983 ( .A1(n5460), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6984 ( .A1(n5462), .A2(n5463), .ZN(n7592) );
  INV_X1 U6985 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5464) );
  OR2_X1 U6986 ( .A1(n5465), .A2(n5464), .ZN(n5467) );
  NAND2_X1 U6987 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  AOI21_X2 U6988 ( .B1(n5468), .B2(n7592), .A(n7609), .ZN(n5469) );
  INV_X1 U6989 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6494) );
  INV_X1 U6990 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U6991 ( .A1(n5469), .A2(n6492), .ZN(n5470) );
  NAND2_X1 U6992 ( .A1(n7609), .A2(n7592), .ZN(n6490) );
  NAND2_X1 U6993 ( .A1(n5534), .A2(n5519), .ZN(n5526) );
  INV_X1 U6994 ( .A(n7513), .ZN(n5472) );
  INV_X1 U6995 ( .A(n7592), .ZN(n5471) );
  NAND3_X1 U6996 ( .A1(n5473), .A2(n5472), .A3(n5471), .ZN(n6437) );
  NAND2_X1 U6997 ( .A1(n4357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U6998 ( .A(n5477), .B(n5476), .ZN(n7422) );
  NOR4_X1 U6999 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U7000 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5480) );
  NOR4_X1 U7001 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5479) );
  NOR4_X1 U7002 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5478) );
  NAND4_X1 U7003 ( .A1(n10008), .A2(n5480), .A3(n5479), .A4(n5478), .ZN(n5486)
         );
  NOR4_X1 U7004 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5484) );
  NOR4_X1 U7005 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5483) );
  NOR4_X1 U7006 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5482) );
  NOR4_X1 U7007 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5481) );
  NAND4_X1 U7008 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n5485)
         );
  OAI21_X1 U7009 ( .B1(n5486), .B2(n5485), .A(n5469), .ZN(n5518) );
  NAND2_X1 U7010 ( .A1(n7742), .A2(n7865), .ZN(n5623) );
  AND3_X1 U7011 ( .A1(n6489), .A2(n5518), .A3(n5623), .ZN(n5488) );
  INV_X1 U7012 ( .A(n5534), .ZN(n5520) );
  NAND2_X1 U7013 ( .A1(n8243), .A2(n7062), .ZN(n7743) );
  NAND2_X1 U7014 ( .A1(n5487), .A2(n7930), .ZN(n5513) );
  OR2_X1 U7015 ( .A1(n5513), .A2(n7062), .ZN(n5489) );
  AND2_X1 U7016 ( .A1(n5489), .A2(n7857), .ZN(n6632) );
  OAI21_X1 U7017 ( .B1(n5520), .B2(n5615), .A(n6632), .ZN(n5492) );
  INV_X1 U7018 ( .A(n5519), .ZN(n6629) );
  INV_X1 U7019 ( .A(n6632), .ZN(n5490) );
  NAND2_X1 U7020 ( .A1(n6629), .A2(n5490), .ZN(n5491) );
  MUX2_X1 U7021 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8255), .S(n9851), .Z(n5494)
         );
  INV_X1 U7022 ( .A(n5494), .ZN(n5517) );
  NAND2_X1 U7023 ( .A1(n6655), .A2(n7748), .ZN(n6729) );
  INV_X1 U7024 ( .A(n6731), .ZN(n7885) );
  NAND2_X1 U7025 ( .A1(n6729), .A2(n7885), .ZN(n5495) );
  INV_X1 U7026 ( .A(n9773), .ZN(n6695) );
  NAND2_X1 U7027 ( .A1(n6703), .A2(n6695), .ZN(n7749) );
  NAND2_X1 U7028 ( .A1(n5495), .A2(n7749), .ZN(n6718) );
  INV_X1 U7029 ( .A(n7880), .ZN(n5496) );
  NAND2_X1 U7030 ( .A1(n6718), .A2(n5496), .ZN(n5497) );
  NAND2_X1 U7031 ( .A1(n5497), .A2(n7764), .ZN(n6711) );
  INV_X1 U7032 ( .A(n6759), .ZN(n8145) );
  NAND2_X1 U7033 ( .A1(n8145), .A2(n4735), .ZN(n7761) );
  NAND2_X1 U7034 ( .A1(n6759), .A2(n6715), .ZN(n7756) );
  NOR2_X1 U7035 ( .A1(n8144), .A2(n9788), .ZN(n7767) );
  INV_X1 U7036 ( .A(n7767), .ZN(n5498) );
  NAND2_X1 U7037 ( .A1(n8144), .A2(n9788), .ZN(n7759) );
  NAND2_X1 U7038 ( .A1(n5499), .A2(n7759), .ZN(n6767) );
  AND2_X1 U7039 ( .A1(n8143), .A2(n9794), .ZN(n6766) );
  NAND2_X1 U7040 ( .A1(n6874), .A2(n6770), .ZN(n7760) );
  NAND2_X1 U7041 ( .A1(n8142), .A2(n9798), .ZN(n7769) );
  INV_X1 U7042 ( .A(n6902), .ZN(n5500) );
  NAND2_X1 U7043 ( .A1(n5501), .A2(n7772), .ZN(n6974) );
  XNOR2_X1 U7044 ( .A(n7027), .B(n8073), .ZN(n6973) );
  NAND2_X1 U7045 ( .A1(n9810), .A2(n8140), .ZN(n7778) );
  INV_X1 U7046 ( .A(n7035), .ZN(n9817) );
  AND2_X1 U7047 ( .A1(n9817), .A2(n8139), .ZN(n7785) );
  INV_X1 U7048 ( .A(n8139), .ZN(n8070) );
  NAND2_X1 U7049 ( .A1(n7035), .A2(n8070), .ZN(n7780) );
  XNOR2_X1 U7050 ( .A(n7790), .B(n8137), .ZN(n7796) );
  NAND2_X1 U7051 ( .A1(n7121), .A2(n7796), .ZN(n5503) );
  INV_X1 U7052 ( .A(n8137), .ZN(n7792) );
  OR2_X1 U7053 ( .A1(n7790), .A2(n7792), .ZN(n5502) );
  NAND2_X1 U7054 ( .A1(n5503), .A2(n5502), .ZN(n7347) );
  NAND2_X1 U7055 ( .A1(n7347), .A2(n7798), .ZN(n5504) );
  NAND2_X1 U7056 ( .A1(n5504), .A2(n7797), .ZN(n7417) );
  NAND2_X1 U7057 ( .A1(n7417), .A2(n7801), .ZN(n5505) );
  NAND2_X1 U7058 ( .A1(n5505), .A2(n7800), .ZN(n7483) );
  INV_X1 U7059 ( .A(n8361), .ZN(n5564) );
  NAND2_X1 U7060 ( .A1(n7498), .A2(n5564), .ZN(n7803) );
  OR2_X1 U7061 ( .A1(n7498), .A2(n5564), .ZN(n7804) );
  INV_X1 U7062 ( .A(n7811), .ZN(n5506) );
  NAND2_X1 U7063 ( .A1(n8337), .A2(n7879), .ZN(n5507) );
  NAND2_X1 U7064 ( .A1(n8465), .A2(n5577), .ZN(n7878) );
  AND2_X1 U7065 ( .A1(n7819), .A2(n8324), .ZN(n7814) );
  INV_X1 U7066 ( .A(n7823), .ZN(n5508) );
  INV_X1 U7067 ( .A(n7828), .ZN(n5509) );
  AOI21_X1 U7068 ( .B1(n8305), .B2(n7826), .A(n5509), .ZN(n7691) );
  NAND2_X1 U7069 ( .A1(n7691), .A2(n7832), .ZN(n8283) );
  NAND2_X1 U7070 ( .A1(n8436), .A2(n8266), .ZN(n7876) );
  NAND2_X1 U7071 ( .A1(n8021), .A2(n8299), .ZN(n8282) );
  AND2_X1 U7072 ( .A1(n7876), .A2(n8282), .ZN(n7831) );
  NAND2_X1 U7073 ( .A1(n8283), .A2(n7831), .ZN(n5510) );
  INV_X1 U7074 ( .A(n7982), .ZN(n5511) );
  NAND2_X1 U7075 ( .A1(n5511), .A2(n7841), .ZN(n5512) );
  NAND2_X1 U7076 ( .A1(n7978), .A2(n8122), .ZN(n7848) );
  XNOR2_X1 U7077 ( .A(n6327), .B(n5431), .ZN(n8263) );
  INV_X1 U7078 ( .A(n7930), .ZN(n7381) );
  NAND2_X1 U7079 ( .A1(n7742), .A2(n5513), .ZN(n5514) );
  NAND3_X1 U7080 ( .A1(n5628), .A2(n9816), .A3(n5514), .ZN(n7031) );
  NAND2_X1 U7081 ( .A1(n7031), .A2(n9818), .ZN(n9808) );
  OAI22_X1 U7082 ( .A1(n8263), .A2(n8416), .B1(n7854), .B2(n8386), .ZN(n5515)
         );
  INV_X1 U7083 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U7084 ( .A1(n5517), .A2(n5516), .ZN(P2_U3487) );
  INV_X1 U7085 ( .A(n5518), .ZN(n5525) );
  NOR2_X1 U7086 ( .A1(n5519), .A2(n5525), .ZN(n5521) );
  NAND2_X1 U7087 ( .A1(n5629), .A2(n6489), .ZN(n5617) );
  NAND2_X1 U7088 ( .A1(n7174), .A2(n5522), .ZN(n7918) );
  NOR2_X1 U7089 ( .A1(n9828), .A2(n7865), .ZN(n5524) );
  NAND2_X1 U7090 ( .A1(n5626), .A2(n5524), .ZN(n5608) );
  NAND2_X1 U7091 ( .A1(n7743), .A2(n9828), .ZN(n8276) );
  AND2_X1 U7092 ( .A1(n5608), .A2(n8276), .ZN(n5621) );
  OR2_X1 U7093 ( .A1(n5617), .A2(n5621), .ZN(n5529) );
  NOR2_X1 U7094 ( .A1(n5526), .A2(n5525), .ZN(n5622) );
  NAND2_X1 U7095 ( .A1(n5622), .A2(n6489), .ZN(n5614) );
  AND2_X1 U7096 ( .A1(n5628), .A2(n5626), .ZN(n5527) );
  OR2_X1 U7097 ( .A1(n5614), .A2(n5527), .ZN(n5528) );
  MUX2_X1 U7098 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8255), .S(n9829), .Z(n5530)
         );
  INV_X1 U7099 ( .A(n5530), .ZN(n5533) );
  NAND2_X1 U7100 ( .A1(n9829), .A2(n9828), .ZN(n8428) );
  OAI22_X1 U7101 ( .A1(n8263), .A2(n8481), .B1(n7854), .B2(n8428), .ZN(n5531)
         );
  INV_X1 U7102 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U7103 ( .A1(n5533), .A2(n5532), .ZN(P2_U3455) );
  INV_X1 U7104 ( .A(n7918), .ZN(n7917) );
  NAND2_X2 U7105 ( .A1(n5535), .A2(n7742), .ZN(n5540) );
  CLKBUF_X3 U7106 ( .A(n5540), .Z(n5606) );
  XNOR2_X1 U7107 ( .A(n9794), .B(n5606), .ZN(n5546) );
  XNOR2_X1 U7108 ( .A(n9778), .B(n5540), .ZN(n5543) );
  XNOR2_X1 U7109 ( .A(n5537), .B(n7703), .ZN(n6700) );
  INV_X1 U7110 ( .A(n9771), .ZN(n6640) );
  INV_X1 U7111 ( .A(n5537), .ZN(n5539) );
  XNOR2_X1 U7112 ( .A(n5540), .B(n9773), .ZN(n5541) );
  XNOR2_X1 U7113 ( .A(n5541), .B(n6703), .ZN(n6694) );
  INV_X1 U7114 ( .A(n5541), .ZN(n5542) );
  XNOR2_X1 U7115 ( .A(n5543), .B(n6732), .ZN(n6642) );
  NAND2_X1 U7116 ( .A1(n6643), .A2(n6642), .ZN(n6641) );
  XNOR2_X1 U7117 ( .A(n6715), .B(n5606), .ZN(n5544) );
  XNOR2_X1 U7118 ( .A(n9788), .B(n5606), .ZN(n5545) );
  XNOR2_X1 U7119 ( .A(n8144), .B(n5545), .ZN(n6758) );
  XNOR2_X1 U7120 ( .A(n8143), .B(n5546), .ZN(n6795) );
  NOR2_X1 U7121 ( .A1(n6794), .A2(n6795), .ZN(n6793) );
  XNOR2_X1 U7122 ( .A(n6881), .B(n5606), .ZN(n5547) );
  XNOR2_X1 U7123 ( .A(n5547), .B(n8142), .ZN(n6836) );
  NAND2_X1 U7124 ( .A1(n5547), .A2(n5548), .ZN(n5549) );
  XNOR2_X1 U7125 ( .A(n6911), .B(n5606), .ZN(n5550) );
  XNOR2_X1 U7126 ( .A(n8141), .B(n5550), .ZN(n6914) );
  XNOR2_X1 U7127 ( .A(n9810), .B(n5606), .ZN(n5552) );
  XNOR2_X1 U7128 ( .A(n5552), .B(n7027), .ZN(n8065) );
  NAND2_X1 U7129 ( .A1(n8066), .A2(n8065), .ZN(n8064) );
  XNOR2_X1 U7130 ( .A(n7035), .B(n5606), .ZN(n7311) );
  XNOR2_X1 U7131 ( .A(n7012), .B(n5606), .ZN(n7315) );
  AOI21_X1 U7132 ( .B1(n8070), .B2(n7311), .A(n7315), .ZN(n5558) );
  NAND3_X1 U7133 ( .A1(n7035), .A2(n5597), .A3(n8139), .ZN(n5554) );
  OAI211_X1 U7134 ( .C1(n5597), .C2(n7217), .A(n7012), .B(n5554), .ZN(n5557)
         );
  INV_X1 U7135 ( .A(n7012), .ZN(n7894) );
  NAND2_X1 U7136 ( .A1(n7785), .A2(n5606), .ZN(n5555) );
  OAI211_X1 U7137 ( .C1(n7217), .C2(n5606), .A(n7894), .B(n5555), .ZN(n5556)
         );
  INV_X1 U7138 ( .A(n7790), .ZN(n7791) );
  XNOR2_X1 U7139 ( .A(n7791), .B(n5606), .ZN(n7110) );
  XNOR2_X1 U7140 ( .A(n7351), .B(n5597), .ZN(n5559) );
  NOR2_X1 U7141 ( .A1(n5559), .A2(n8136), .ZN(n7458) );
  AOI21_X1 U7142 ( .B1(n5559), .B2(n8136), .A(n7458), .ZN(n7338) );
  NAND2_X1 U7143 ( .A1(n7337), .A2(n7338), .ZN(n7336) );
  INV_X1 U7144 ( .A(n7458), .ZN(n5560) );
  NAND2_X1 U7145 ( .A1(n7336), .A2(n5560), .ZN(n5561) );
  XNOR2_X1 U7146 ( .A(n7410), .B(n5606), .ZN(n5562) );
  XNOR2_X1 U7147 ( .A(n5562), .B(n8135), .ZN(n7457) );
  NAND2_X1 U7148 ( .A1(n5562), .A2(n7504), .ZN(n5563) );
  XNOR2_X1 U7149 ( .A(n7498), .B(n5606), .ZN(n5566) );
  XNOR2_X1 U7150 ( .A(n5566), .B(n5564), .ZN(n7499) );
  INV_X1 U7151 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7152 ( .A1(n5567), .A2(n8361), .ZN(n5568) );
  XNOR2_X1 U7153 ( .A(n8478), .B(n5606), .ZN(n5569) );
  XNOR2_X1 U7154 ( .A(n5569), .B(n8349), .ZN(n7582) );
  NAND2_X1 U7155 ( .A1(n7583), .A2(n7582), .ZN(n5572) );
  INV_X1 U7156 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7157 ( .A1(n5570), .A2(n8349), .ZN(n5571) );
  NAND2_X1 U7158 ( .A1(n5572), .A2(n5571), .ZN(n8045) );
  XNOR2_X1 U7159 ( .A(n8471), .B(n5606), .ZN(n5573) );
  NAND2_X1 U7160 ( .A1(n5573), .A2(n8110), .ZN(n8099) );
  OAI21_X1 U7161 ( .B1(n5573), .B2(n8110), .A(n8099), .ZN(n8047) );
  XNOR2_X1 U7162 ( .A(n8465), .B(n5606), .ZN(n5576) );
  XNOR2_X1 U7163 ( .A(n5576), .B(n8350), .ZN(n8100) );
  INV_X1 U7164 ( .A(n8100), .ZN(n5575) );
  OR2_X1 U7165 ( .A1(n8047), .A2(n5575), .ZN(n5574) );
  NOR2_X1 U7166 ( .A1(n8045), .A2(n5574), .ZN(n8104) );
  NOR2_X1 U7167 ( .A1(n5575), .A2(n8099), .ZN(n8103) );
  XNOR2_X1 U7168 ( .A(n8458), .B(n5606), .ZN(n5580) );
  XNOR2_X1 U7169 ( .A(n5580), .B(n8085), .ZN(n7937) );
  INV_X1 U7170 ( .A(n7937), .ZN(n5578) );
  XNOR2_X1 U7171 ( .A(n8399), .B(n5597), .ZN(n5579) );
  NOR2_X1 U7172 ( .A1(n5579), .A2(n8313), .ZN(n8026) );
  AOI21_X1 U7173 ( .B1(n5579), .B2(n8313), .A(n8026), .ZN(n8079) );
  INV_X1 U7174 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7175 ( .A1(n5581), .A2(n8340), .ZN(n8080) );
  INV_X1 U7176 ( .A(n8026), .ZN(n5583) );
  XNOR2_X1 U7177 ( .A(n8448), .B(n5606), .ZN(n5584) );
  NAND2_X1 U7178 ( .A1(n5584), .A2(n8301), .ZN(n8089) );
  INV_X1 U7179 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7180 ( .A1(n5585), .A2(n5351), .ZN(n5586) );
  AND2_X1 U7181 ( .A1(n8089), .A2(n5586), .ZN(n8025) );
  XNOR2_X1 U7182 ( .A(n8442), .B(n5606), .ZN(n5587) );
  XNOR2_X1 U7183 ( .A(n5587), .B(n8312), .ZN(n8090) );
  NAND2_X1 U7184 ( .A1(n5587), .A2(n7694), .ZN(n5588) );
  NAND2_X1 U7185 ( .A1(n8091), .A2(n5588), .ZN(n5592) );
  INV_X1 U7186 ( .A(n5592), .ZN(n5590) );
  XNOR2_X1 U7187 ( .A(n8021), .B(n5606), .ZN(n5591) );
  INV_X1 U7188 ( .A(n5591), .ZN(n5589) );
  NAND2_X1 U7189 ( .A1(n8017), .A2(n8054), .ZN(n5596) );
  XNOR2_X1 U7190 ( .A(n8387), .B(n5597), .ZN(n5593) );
  NAND2_X1 U7191 ( .A1(n5593), .A2(n8266), .ZN(n8035) );
  INV_X1 U7192 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7193 ( .A1(n5594), .A2(n8133), .ZN(n5595) );
  NAND2_X1 U7194 ( .A1(n5596), .A2(n8055), .ZN(n8034) );
  NAND2_X1 U7195 ( .A1(n8034), .A2(n8035), .ZN(n5598) );
  XNOR2_X1 U7196 ( .A(n8268), .B(n5597), .ZN(n5599) );
  XNOR2_X1 U7197 ( .A(n5599), .B(n8279), .ZN(n8036) );
  NAND2_X1 U7198 ( .A1(n5598), .A2(n8036), .ZN(n8038) );
  XNOR2_X1 U7199 ( .A(n8379), .B(n5606), .ZN(n5601) );
  INV_X1 U7200 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7201 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  XNOR2_X1 U7202 ( .A(n7978), .B(n5606), .ZN(n5634) );
  XNOR2_X1 U7203 ( .A(n5634), .B(n8122), .ZN(n8004) );
  XNOR2_X1 U7204 ( .A(n6328), .B(n5606), .ZN(n5607) );
  XNOR2_X1 U7205 ( .A(n7854), .B(n5607), .ZN(n5635) );
  INV_X1 U7206 ( .A(n5635), .ZN(n5611) );
  OR2_X1 U7207 ( .A1(n5617), .A2(n5626), .ZN(n5610) );
  OR2_X1 U7208 ( .A1(n5614), .A2(n5608), .ZN(n5609) );
  INV_X1 U7209 ( .A(n5634), .ZN(n5612) );
  AOI21_X1 U7210 ( .B1(n5612), .B2(n8131), .A(n8052), .ZN(n5613) );
  NAND3_X1 U7211 ( .A1(n8006), .A2(n5613), .A3(n5635), .ZN(n5639) );
  OR2_X1 U7212 ( .A1(n5614), .A2(n9816), .ZN(n5616) );
  OR2_X1 U7213 ( .A1(n5617), .A2(n5628), .ZN(n5620) );
  INV_X1 U7214 ( .A(n5620), .ZN(n5618) );
  NAND2_X1 U7215 ( .A1(n5618), .A2(n5619), .ZN(n8121) );
  NOR2_X2 U7216 ( .A1(n5620), .A2(n5619), .ZN(n8119) );
  AOI22_X1 U7217 ( .A1(n8131), .A2(n8119), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n5633) );
  OR2_X1 U7218 ( .A1(n5622), .A2(n5621), .ZN(n5625) );
  AND3_X1 U7219 ( .A1(n6437), .A2(n7422), .A3(n5623), .ZN(n5624) );
  OAI211_X1 U7220 ( .C1(n5629), .C2(n5626), .A(n5625), .B(n5624), .ZN(n5627)
         );
  NAND2_X1 U7221 ( .A1(n5627), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5631) );
  INV_X1 U7222 ( .A(n5628), .ZN(n6635) );
  NAND2_X1 U7223 ( .A1(n6489), .A2(n6635), .ZN(n7929) );
  OR2_X1 U7224 ( .A1(n5629), .A2(n7929), .ZN(n5630) );
  NAND2_X1 U7225 ( .A1(n8259), .A2(n8124), .ZN(n5632) );
  OAI211_X1 U7226 ( .C1(n7009), .C2(n8121), .A(n5633), .B(n5632), .ZN(n5637)
         );
  NOR4_X1 U7227 ( .A1(n5635), .A2(n8122), .A3(n5634), .A4(n8052), .ZN(n5636)
         );
  AOI211_X1 U7228 ( .C1(n8260), .C2(n8072), .A(n5637), .B(n5636), .ZN(n5638)
         );
  NAND3_X1 U7229 ( .A1(n5640), .A2(n5639), .A3(n5638), .ZN(P2_U3160) );
  NAND2_X1 U7230 ( .A1(n5731), .A2(n5641), .ZN(n5761) );
  NOR2_X1 U7231 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5644) );
  NOR2_X1 U7232 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5649) );
  NOR2_X1 U7233 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5648) );
  NOR2_X1 U7234 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5647) );
  OAI21_X1 U7235 ( .B1(n5705), .B2(n5992), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5654) );
  NAND2_X2 U7236 ( .A1(n6280), .A2(n8959), .ZN(n5835) );
  NAND2_X1 U7237 ( .A1(n7172), .A2(n5758), .ZN(n5660) );
  NAND2_X1 U7238 ( .A1(n5759), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5659) );
  INV_X1 U7239 ( .A(n6051), .ZN(n5665) );
  INV_X1 U7240 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7241 ( .A1(n5665), .A2(n5664), .ZN(n5673) );
  INV_X1 U7242 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7243 ( .A1(n5685), .A2(n5666), .ZN(n5667) );
  NAND2_X1 U7244 ( .A1(n5669), .A2(n5668), .ZN(n6261) );
  NAND2_X1 U7245 ( .A1(n6070), .A2(n5671), .ZN(n5672) );
  NAND2_X1 U7246 ( .A1(n5673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5675) );
  INV_X1 U7247 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7248 ( .A1(n4291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7249 ( .A1(n5678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5679) );
  MUX2_X1 U7250 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5679), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5680) );
  NOR2_X1 U7251 ( .A1(n7591), .A2(n7512), .ZN(n5683) );
  OAI21_X1 U7252 ( .B1(n8921), .B2(n6266), .A(n6441), .ZN(n5684) );
  INV_X1 U7253 ( .A(n5684), .ZN(n5688) );
  NAND2_X4 U7254 ( .A1(n5688), .A2(n6818), .ZN(n8531) );
  NAND2_X4 U7255 ( .A1(n5689), .A2(n6278), .ZN(n6241) );
  NAND2_X1 U7256 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5811) );
  INV_X1 U7257 ( .A(n5811), .ZN(n5690) );
  NAND2_X1 U7258 ( .A1(n5690), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5828) );
  INV_X1 U7259 ( .A(n5828), .ZN(n5691) );
  INV_X1 U7260 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6055) );
  INV_X1 U7261 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7431) );
  INV_X1 U7262 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6118) );
  INV_X1 U7263 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U7264 ( .A1(n6121), .A2(n8557), .ZN(n5700) );
  NAND2_X1 U7265 ( .A1(n6140), .A2(n5700), .ZN(n9203) );
  AND2_X1 U7266 ( .A1(n5652), .A2(n5703), .ZN(n5704) );
  NAND2_X1 U7267 ( .A1(n5705), .A2(n5704), .ZN(n9444) );
  OR2_X1 U7268 ( .A1(n9203), .A2(n5774), .ZN(n5712) );
  INV_X1 U7269 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U7270 ( .A1(n6413), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7271 ( .A1(n5773), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5708) );
  OAI211_X1 U7272 ( .C1(n9202), .C2(n5775), .A(n5709), .B(n5708), .ZN(n5710)
         );
  INV_X1 U7273 ( .A(n5710), .ZN(n5711) );
  INV_X1 U7274 ( .A(n6389), .ZN(n6929) );
  AND2_X4 U7275 ( .A1(n6929), .A2(n6441), .ZN(n6168) );
  INV_X2 U7276 ( .A(n6168), .ZN(n8532) );
  OAI22_X1 U7277 ( .A1(n9424), .A2(n5735), .B1(n9212), .B2(n8532), .ZN(n5713)
         );
  XNOR2_X1 U7278 ( .A(n5713), .B(n6241), .ZN(n6137) );
  OAI22_X1 U7279 ( .A1(n9424), .A2(n8532), .B1(n9212), .B2(n8531), .ZN(n6136)
         );
  INV_X1 U7280 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6928) );
  OR2_X1 U7281 ( .A1(n5774), .A2(n6928), .ZN(n5717) );
  INV_X1 U7282 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5714) );
  OR2_X1 U7283 ( .A1(n5775), .A2(n5714), .ZN(n5716) );
  INV_X1 U7284 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5723) );
  OR2_X1 U7285 ( .A1(n8771), .A2(n5723), .ZN(n5715) );
  NAND2_X1 U7286 ( .A1(n7731), .A2(SI_0_), .ZN(n5720) );
  INV_X1 U7287 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7288 ( .A1(n5720), .A2(n5719), .ZN(n5722) );
  AND2_X1 U7289 ( .A1(n5722), .A2(n5721), .ZN(n9449) );
  OR2_X1 U7290 ( .A1(n6441), .A2(n5723), .ZN(n5724) );
  INV_X1 U7291 ( .A(n8531), .ZN(n6219) );
  NAND2_X1 U7292 ( .A1(n6351), .A2(n6219), .ZN(n5727) );
  INV_X1 U7293 ( .A(n6441), .ZN(n5725) );
  AOI22_X1 U7294 ( .A1(n9556), .A2(n6168), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5725), .ZN(n5726) );
  NAND2_X1 U7295 ( .A1(n5727), .A2(n5726), .ZN(n6649) );
  NAND2_X1 U7296 ( .A1(n5728), .A2(n8529), .ZN(n5729) );
  NAND2_X1 U7297 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5730) );
  MUX2_X1 U7298 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5730), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5733) );
  INV_X1 U7299 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7300 ( .A1(n5733), .A2(n5732), .ZN(n6561) );
  INV_X1 U7301 ( .A(n6561), .ZN(n8949) );
  NAND2_X1 U7302 ( .A1(n5780), .A2(n8949), .ZN(n5734) );
  INV_X1 U7303 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U7304 ( .A1(n6094), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5737) );
  AND2_X1 U7305 ( .A1(n5738), .A2(n5737), .ZN(n5742) );
  INV_X1 U7306 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5739) );
  INV_X1 U7307 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8947) );
  OR2_X1 U7308 ( .A1(n5774), .A2(n8947), .ZN(n5740) );
  NAND2_X1 U7309 ( .A1(n5743), .A2(n6219), .ZN(n5746) );
  OR2_X1 U7310 ( .A1(n5744), .A2(n8532), .ZN(n5745) );
  NAND2_X1 U7311 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  NAND2_X1 U7312 ( .A1(n7948), .A2(n7946), .ZN(n7947) );
  INV_X1 U7313 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7314 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7315 ( .A1(n7947), .A2(n5750), .ZN(n6740) );
  INV_X1 U7316 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5752) );
  INV_X1 U7317 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6892) );
  INV_X1 U7318 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6544) );
  OR2_X1 U7319 ( .A1(n8771), .A2(n6544), .ZN(n5754) );
  INV_X1 U7320 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8968) );
  OR2_X1 U7321 ( .A1(n5774), .A2(n8968), .ZN(n5753) );
  NAND2_X1 U7322 ( .A1(n5759), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5764) );
  NOR2_X1 U7323 ( .A1(n5731), .A2(n5992), .ZN(n5760) );
  MUX2_X1 U7324 ( .A(n5992), .B(n5760), .S(P1_IR_REG_2__SCAN_IN), .Z(n5762) );
  NOR2_X1 U7325 ( .A1(n5762), .A2(n4829), .ZN(n8971) );
  NAND2_X1 U7326 ( .A1(n4271), .A2(n8971), .ZN(n5763) );
  XNOR2_X1 U7327 ( .A(n5765), .B(n8529), .ZN(n5770) );
  NAND2_X1 U7328 ( .A1(n6897), .A2(n6168), .ZN(n5766) );
  NAND2_X1 U7329 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  XNOR2_X1 U7330 ( .A(n5770), .B(n5768), .ZN(n6739) );
  NAND2_X1 U7331 ( .A1(n6740), .A2(n6739), .ZN(n5772) );
  INV_X1 U7332 ( .A(n5768), .ZN(n5769) );
  NAND2_X1 U7333 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  NAND2_X1 U7334 ( .A1(n5772), .A2(n5771), .ZN(n6778) );
  NAND2_X1 U7335 ( .A1(n5773), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5779) );
  OR2_X1 U7336 ( .A1(n5774), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5778) );
  INV_X1 U7337 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6564) );
  OR2_X1 U7338 ( .A1(n5775), .A2(n6564), .ZN(n5777) );
  INV_X1 U7339 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6547) );
  OR2_X1 U7340 ( .A1(n8771), .A2(n6547), .ZN(n5776) );
  NAND2_X1 U7341 ( .A1(n5759), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7342 ( .A1(n5761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7343 ( .A1(n5781), .A2(n10005), .ZN(n5798) );
  OR2_X1 U7344 ( .A1(n5781), .A2(n10005), .ZN(n5782) );
  AND2_X1 U7345 ( .A1(n5798), .A2(n5782), .ZN(n8984) );
  NAND2_X1 U7346 ( .A1(n4271), .A2(n8984), .ZN(n5783) );
  OAI22_X1 U7347 ( .A1(n6886), .A2(n8532), .B1(n6941), .B2(n5735), .ZN(n5785)
         );
  XNOR2_X1 U7348 ( .A(n5785), .B(n8529), .ZN(n5790) );
  OR2_X1 U7349 ( .A1(n6886), .A2(n8531), .ZN(n5787) );
  NAND2_X1 U7350 ( .A1(n6854), .A2(n6168), .ZN(n5786) );
  NAND2_X1 U7351 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  NAND2_X1 U7352 ( .A1(n6778), .A2(n6779), .ZN(n5792) );
  INV_X1 U7353 ( .A(n5788), .ZN(n5789) );
  NAND2_X1 U7354 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  INV_X1 U7355 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6951) );
  OR2_X1 U7356 ( .A1(n5775), .A2(n6951), .ZN(n5797) );
  OAI21_X1 U7357 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5811), .ZN(n6953) );
  OR2_X1 U7358 ( .A1(n5774), .A2(n6953), .ZN(n5796) );
  NAND2_X1 U7359 ( .A1(n5773), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5795) );
  INV_X1 U7360 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5793) );
  OR2_X1 U7361 ( .A1(n8771), .A2(n5793), .ZN(n5794) );
  NAND2_X1 U7362 ( .A1(n5759), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7363 ( .A1(n5798), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U7364 ( .A(n5799), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U7365 ( .A1(n5780), .A2(n6566), .ZN(n5800) );
  OAI22_X1 U7366 ( .A1(n8663), .A2(n8532), .B1(n8664), .B2(n5735), .ZN(n5802)
         );
  XNOR2_X1 U7367 ( .A(n5802), .B(n6241), .ZN(n5807) );
  OR2_X1 U7368 ( .A1(n8663), .A2(n8531), .ZN(n5804) );
  NAND2_X1 U7369 ( .A1(n9566), .A2(n6168), .ZN(n5803) );
  NAND2_X1 U7370 ( .A1(n5804), .A2(n5803), .ZN(n5806) );
  XNOR2_X1 U7371 ( .A(n5807), .B(n5806), .ZN(n6802) );
  INV_X1 U7372 ( .A(n6802), .ZN(n5805) );
  NAND2_X1 U7373 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  NAND2_X1 U7374 ( .A1(n6413), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5816) );
  INV_X1 U7375 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5809) );
  OR2_X1 U7376 ( .A1(n5751), .A2(n5809), .ZN(n5815) );
  INV_X1 U7377 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7378 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U7379 ( .A1(n5828), .A2(n5812), .ZN(n7003) );
  OR2_X1 U7380 ( .A1(n5774), .A2(n7003), .ZN(n5814) );
  INV_X1 U7381 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7382 ( .A1(n5775), .A2(n6568), .ZN(n5813) );
  NAND2_X1 U7383 ( .A1(n5759), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7384 ( .A1(n5817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5818) );
  MUX2_X1 U7385 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5818), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5820) );
  NOR2_X1 U7386 ( .A1(n5817), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5838) );
  INV_X1 U7387 ( .A(n5838), .ZN(n5819) );
  AND2_X1 U7388 ( .A1(n5820), .A2(n5819), .ZN(n9011) );
  NAND2_X1 U7389 ( .A1(n4271), .A2(n9011), .ZN(n5821) );
  OAI22_X1 U7390 ( .A1(n6959), .A2(n8532), .B1(n9543), .B2(n5735), .ZN(n5823)
         );
  XNOR2_X1 U7391 ( .A(n5823), .B(n8529), .ZN(n6999) );
  OR2_X1 U7392 ( .A1(n6959), .A2(n8531), .ZN(n5825) );
  NAND2_X1 U7393 ( .A1(n7107), .A2(n6168), .ZN(n5824) );
  AND2_X1 U7394 ( .A1(n5825), .A2(n5824), .ZN(n7001) );
  NAND2_X1 U7395 ( .A1(n5773), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5834) );
  INV_X1 U7396 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5826) );
  OR2_X1 U7397 ( .A1(n5775), .A2(n5826), .ZN(n5833) );
  INV_X1 U7398 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U7399 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  NAND2_X1 U7400 ( .A1(n5859), .A2(n5829), .ZN(n6965) );
  OR2_X1 U7401 ( .A1(n5774), .A2(n6965), .ZN(n5832) );
  INV_X1 U7402 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5830) );
  OR2_X1 U7403 ( .A1(n8771), .A2(n5830), .ZN(n5831) );
  NOR2_X1 U7404 ( .A1(n5838), .A2(n5992), .ZN(n5836) );
  MUX2_X1 U7405 ( .A(n5992), .B(n5836), .S(P1_IR_REG_6__SCAN_IN), .Z(n5840) );
  INV_X1 U7406 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7407 ( .A1(n5838), .A2(n5837), .ZN(n5879) );
  INV_X1 U7408 ( .A(n5879), .ZN(n5839) );
  OR2_X1 U7409 ( .A1(n6486), .A2(n5853), .ZN(n5842) );
  NAND2_X1 U7410 ( .A1(n5759), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U7411 ( .C1(n5835), .C2(n6570), .A(n5842), .B(n5841), .ZN(n7074)
         );
  INV_X1 U7412 ( .A(n7074), .ZN(n9575) );
  OAI22_X1 U7413 ( .A1(n7050), .A2(n8532), .B1(n9575), .B2(n5735), .ZN(n5843)
         );
  XNOR2_X1 U7414 ( .A(n5843), .B(n8529), .ZN(n7069) );
  OR2_X1 U7415 ( .A1(n7050), .A2(n8531), .ZN(n5845) );
  NAND2_X1 U7416 ( .A1(n7074), .A2(n6168), .ZN(n5844) );
  AND2_X1 U7417 ( .A1(n5845), .A2(n5844), .ZN(n5847) );
  AOI22_X1 U7418 ( .A1(n6999), .A2(n7001), .B1(n7069), .B2(n5847), .ZN(n5846)
         );
  OAI21_X1 U7419 ( .B1(n6999), .B2(n7001), .A(n5847), .ZN(n5851) );
  INV_X1 U7420 ( .A(n7069), .ZN(n5850) );
  INV_X1 U7421 ( .A(n6999), .ZN(n7067) );
  INV_X1 U7422 ( .A(n7001), .ZN(n5848) );
  INV_X1 U7423 ( .A(n5847), .ZN(n7068) );
  AND2_X1 U7424 ( .A1(n5848), .A2(n7068), .ZN(n5849) );
  OR2_X1 U7425 ( .A1(n6496), .A2(n5853), .ZN(n5856) );
  NAND2_X1 U7426 ( .A1(n5879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7427 ( .A(n5854), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U7428 ( .A1(n5759), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4271), .B2(
        n6574), .ZN(n5855) );
  NAND2_X1 U7429 ( .A1(n7051), .A2(n6239), .ZN(n5868) );
  NAND2_X1 U7430 ( .A1(n5773), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5865) );
  INV_X1 U7431 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7432 ( .A1(n5775), .A2(n5857), .ZN(n5864) );
  INV_X1 U7433 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7434 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  NAND2_X1 U7435 ( .A1(n5885), .A2(n5860), .ZN(n7054) );
  OR2_X1 U7436 ( .A1(n5774), .A2(n7054), .ZN(n5863) );
  INV_X1 U7437 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5861) );
  OR2_X1 U7438 ( .A1(n8771), .A2(n5861), .ZN(n5862) );
  OR2_X1 U7439 ( .A1(n7085), .A2(n8531), .ZN(n5871) );
  NAND2_X1 U7440 ( .A1(n7051), .A2(n6168), .ZN(n5870) );
  AND2_X1 U7441 ( .A1(n5871), .A2(n5870), .ZN(n5873) );
  NAND2_X1 U7442 ( .A1(n5872), .A2(n5873), .ZN(n5878) );
  INV_X1 U7443 ( .A(n5872), .ZN(n5875) );
  INV_X1 U7444 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7445 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  NAND2_X1 U7446 ( .A1(n5878), .A2(n5876), .ZN(n6990) );
  INV_X1 U7447 ( .A(n6990), .ZN(n5877) );
  NAND2_X1 U7448 ( .A1(n6500), .A2(n5758), .ZN(n5882) );
  NAND2_X1 U7449 ( .A1(n5900), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7450 ( .A(n5880), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9480) );
  AOI22_X1 U7451 ( .A1(n5759), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4271), .B2(
        n9480), .ZN(n5881) );
  NAND2_X1 U7452 ( .A1(n7206), .A2(n6239), .ZN(n5893) );
  NAND2_X1 U7453 ( .A1(n5773), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5891) );
  INV_X1 U7454 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5883) );
  OR2_X1 U7455 ( .A1(n8771), .A2(n5883), .ZN(n5890) );
  NAND2_X1 U7456 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7457 ( .A1(n5904), .A2(n5886), .ZN(n7207) );
  OR2_X1 U7458 ( .A1(n5774), .A2(n7207), .ZN(n5889) );
  INV_X1 U7459 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7460 ( .A1(n5775), .A2(n5887), .ZN(n5888) );
  OR2_X1 U7461 ( .A1(n7331), .A2(n8532), .ZN(n5892) );
  NAND2_X1 U7462 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  XNOR2_X1 U7463 ( .A(n5894), .B(n6241), .ZN(n5897) );
  NAND2_X1 U7464 ( .A1(n7206), .A2(n6168), .ZN(n5896) );
  OR2_X1 U7465 ( .A1(n7331), .A2(n8531), .ZN(n5895) );
  AND2_X1 U7466 ( .A1(n5896), .A2(n5895), .ZN(n7204) );
  NAND2_X1 U7467 ( .A1(n7202), .A2(n7204), .ZN(n7203) );
  INV_X1 U7468 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U7469 ( .A1(n5899), .A2(n5898), .ZN(n7324) );
  NAND2_X1 U7470 ( .A1(n6534), .A2(n5758), .ZN(n5903) );
  NAND2_X1 U7471 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5901) );
  XNOR2_X1 U7472 ( .A(n5901), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6673) );
  AOI22_X1 U7473 ( .A1(n5759), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4271), .B2(
        n6673), .ZN(n5902) );
  NAND2_X1 U7474 ( .A1(n7307), .A2(n6239), .ZN(n5912) );
  NAND2_X1 U7475 ( .A1(n5773), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7476 ( .A1(n8771), .A2(n9603), .ZN(n5909) );
  INV_X1 U7477 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U7478 ( .A1(n5904), .A2(n6580), .ZN(n5905) );
  NAND2_X1 U7479 ( .A1(n5929), .A2(n5905), .ZN(n7328) );
  OR2_X1 U7480 ( .A1(n5774), .A2(n7328), .ZN(n5908) );
  INV_X1 U7481 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5906) );
  OR2_X1 U7482 ( .A1(n5775), .A2(n5906), .ZN(n5907) );
  OR2_X1 U7483 ( .A1(n7401), .A2(n8532), .ZN(n5911) );
  NAND2_X1 U7484 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  XNOR2_X1 U7485 ( .A(n5913), .B(n6241), .ZN(n5916) );
  NOR2_X1 U7486 ( .A1(n7401), .A2(n8531), .ZN(n5914) );
  AOI21_X1 U7487 ( .B1(n7307), .B2(n6168), .A(n5914), .ZN(n5917) );
  XNOR2_X1 U7488 ( .A(n5916), .B(n5917), .ZN(n7326) );
  AND2_X1 U7489 ( .A1(n7324), .A2(n7326), .ZN(n5915) );
  NAND2_X1 U7490 ( .A1(n7203), .A2(n5915), .ZN(n7325) );
  INV_X1 U7491 ( .A(n5916), .ZN(n5918) );
  OR2_X1 U7492 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  NAND2_X1 U7493 ( .A1(n7325), .A2(n5919), .ZN(n5939) );
  NAND2_X1 U7494 ( .A1(n6537), .A2(n5758), .ZN(n5925) );
  OAI21_X1 U7495 ( .B1(n5920), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5922) );
  INV_X1 U7496 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5921) );
  OR2_X1 U7497 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  NAND2_X1 U7498 ( .A1(n5922), .A2(n5921), .ZN(n5945) );
  AOI22_X1 U7499 ( .A1(n5759), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4271), .B2(
        n9458), .ZN(n5924) );
  NAND2_X1 U7500 ( .A1(n7523), .A2(n6239), .ZN(n5936) );
  NAND2_X1 U7501 ( .A1(n6413), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5934) );
  INV_X1 U7502 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7503 ( .A1(n5751), .A2(n5926), .ZN(n5933) );
  INV_X1 U7504 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5927) );
  OR2_X1 U7505 ( .A1(n5775), .A2(n5927), .ZN(n5932) );
  NAND2_X1 U7506 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  NAND2_X1 U7507 ( .A1(n5949), .A2(n5930), .ZN(n7521) );
  OR2_X1 U7508 ( .A1(n5774), .A2(n7521), .ZN(n5931) );
  OR2_X1 U7509 ( .A1(n7600), .A2(n8532), .ZN(n5935) );
  NAND2_X1 U7510 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  XNOR2_X1 U7511 ( .A(n5937), .B(n6241), .ZN(n5938) );
  NAND2_X1 U7512 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U7513 ( .A1(n7523), .A2(n6168), .ZN(n5942) );
  OR2_X1 U7514 ( .A1(n7600), .A2(n8531), .ZN(n5941) );
  NAND2_X1 U7515 ( .A1(n5942), .A2(n5941), .ZN(n7517) );
  INV_X1 U7516 ( .A(n7517), .ZN(n5943) );
  NAND2_X1 U7517 ( .A1(n6606), .A2(n5758), .ZN(n5948) );
  NAND2_X1 U7518 ( .A1(n5945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7519 ( .A(n5946), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U7520 ( .A1(n5759), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5780), .B2(
        n6675), .ZN(n5947) );
  NAND2_X1 U7521 ( .A1(n7605), .A2(n6239), .ZN(n5956) );
  NAND2_X1 U7522 ( .A1(n5773), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5954) );
  INV_X1 U7523 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6674) );
  OR2_X1 U7524 ( .A1(n8771), .A2(n6674), .ZN(n5953) );
  INV_X1 U7525 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U7526 ( .A1(n5949), .A2(n7599), .ZN(n5950) );
  NAND2_X1 U7527 ( .A1(n5965), .A2(n5950), .ZN(n7603) );
  OR2_X1 U7528 ( .A1(n5774), .A2(n7603), .ZN(n5952) );
  INV_X1 U7529 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7476) );
  OR2_X1 U7530 ( .A1(n5775), .A2(n7476), .ZN(n5951) );
  OR2_X1 U7531 ( .A1(n7632), .A2(n8532), .ZN(n5955) );
  NAND2_X1 U7532 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  XNOR2_X1 U7533 ( .A(n5957), .B(n6241), .ZN(n5982) );
  NAND2_X1 U7534 ( .A1(n7605), .A2(n6168), .ZN(n5959) );
  OR2_X1 U7535 ( .A1(n7632), .A2(n8531), .ZN(n5958) );
  NAND2_X1 U7536 ( .A1(n5959), .A2(n5958), .ZN(n5983) );
  NAND2_X1 U7537 ( .A1(n5982), .A2(n5983), .ZN(n7596) );
  NAND2_X1 U7538 ( .A1(n6626), .A2(n5758), .ZN(n5963) );
  OR2_X1 U7539 ( .A1(n5960), .A2(n5992), .ZN(n5961) );
  XNOR2_X1 U7540 ( .A(n5961), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7365) );
  AOI22_X1 U7541 ( .A1(n5759), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5780), .B2(
        n7365), .ZN(n5962) );
  NAND2_X1 U7542 ( .A1(n7637), .A2(n6239), .ZN(n5973) );
  NAND2_X1 U7543 ( .A1(n5773), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5971) );
  INV_X1 U7544 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7535) );
  OR2_X1 U7545 ( .A1(n5775), .A2(n7535), .ZN(n5970) );
  NAND2_X1 U7546 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  NAND2_X1 U7547 ( .A1(n5999), .A2(n5966), .ZN(n7635) );
  OR2_X1 U7548 ( .A1(n5774), .A2(n7635), .ZN(n5969) );
  INV_X1 U7549 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5967) );
  OR2_X1 U7550 ( .A1(n8771), .A2(n5967), .ZN(n5968) );
  NAND4_X1 U7551 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n8942)
         );
  NAND2_X1 U7552 ( .A1(n8942), .A2(n6168), .ZN(n5972) );
  NAND2_X1 U7553 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  XNOR2_X1 U7554 ( .A(n5974), .B(n6241), .ZN(n5978) );
  INV_X1 U7555 ( .A(n5978), .ZN(n5976) );
  AND2_X1 U7556 ( .A1(n8942), .A2(n6219), .ZN(n5975) );
  AOI21_X1 U7557 ( .B1(n7637), .B2(n6168), .A(n5975), .ZN(n5977) );
  NAND2_X1 U7558 ( .A1(n5976), .A2(n5977), .ZN(n5986) );
  INV_X1 U7559 ( .A(n5986), .ZN(n5979) );
  XNOR2_X1 U7560 ( .A(n5978), .B(n5977), .ZN(n7630) );
  OR2_X1 U7561 ( .A1(n5979), .A2(n7630), .ZN(n5981) );
  AND2_X1 U7562 ( .A1(n7596), .A2(n5981), .ZN(n5980) );
  INV_X1 U7563 ( .A(n5981), .ZN(n5988) );
  INV_X1 U7564 ( .A(n5982), .ZN(n5985) );
  INV_X1 U7565 ( .A(n5983), .ZN(n5984) );
  NAND2_X1 U7566 ( .A1(n5985), .A2(n5984), .ZN(n7627) );
  AND2_X1 U7567 ( .A1(n7627), .A2(n5986), .ZN(n5987) );
  OR2_X1 U7568 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7569 ( .A1(n6652), .A2(n5758), .ZN(n5998) );
  AND2_X1 U7570 ( .A1(n5960), .A2(n5990), .ZN(n5994) );
  NOR2_X1 U7571 ( .A1(n5994), .A2(n5992), .ZN(n5991) );
  MUX2_X1 U7572 ( .A(n5992), .B(n5991), .S(P1_IR_REG_13__SCAN_IN), .Z(n5996)
         );
  NAND2_X1 U7573 ( .A1(n5994), .A2(n5993), .ZN(n6014) );
  INV_X1 U7574 ( .A(n6014), .ZN(n5995) );
  AOI22_X1 U7575 ( .A1(n5759), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4271), .B2(
        n9516), .ZN(n5997) );
  NAND2_X1 U7576 ( .A1(n7674), .A2(n6239), .ZN(n6006) );
  NAND2_X1 U7577 ( .A1(n5773), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6004) );
  INV_X1 U7578 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7621) );
  OR2_X1 U7579 ( .A1(n5775), .A2(n7621), .ZN(n6003) );
  NAND2_X1 U7580 ( .A1(n5999), .A2(n7659), .ZN(n6000) );
  NAND2_X1 U7581 ( .A1(n6020), .A2(n6000), .ZN(n7663) );
  OR2_X1 U7582 ( .A1(n5774), .A2(n7663), .ZN(n6002) );
  INV_X1 U7583 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7357) );
  OR2_X1 U7584 ( .A1(n8771), .A2(n7357), .ZN(n6001) );
  OR2_X1 U7585 ( .A1(n7529), .A2(n8532), .ZN(n6005) );
  NAND2_X1 U7586 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  XNOR2_X1 U7587 ( .A(n6007), .B(n6241), .ZN(n6009) );
  NOR2_X1 U7588 ( .A1(n7529), .A2(n8531), .ZN(n6008) );
  AOI21_X1 U7589 ( .B1(n7674), .B2(n6168), .A(n6008), .ZN(n6010) );
  XNOR2_X1 U7590 ( .A(n6009), .B(n6010), .ZN(n7658) );
  INV_X1 U7591 ( .A(n6009), .ZN(n6011) );
  AND2_X1 U7592 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  NAND2_X1 U7593 ( .A1(n6707), .A2(n5758), .ZN(n6017) );
  NAND2_X1 U7594 ( .A1(n6014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6013) );
  MUX2_X1 U7595 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6013), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6015) );
  OR2_X1 U7596 ( .A1(n6014), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6030) );
  AOI22_X1 U7597 ( .A1(n5759), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4271), .B2(
        n9532), .ZN(n6016) );
  NAND2_X1 U7598 ( .A1(n7650), .A2(n6239), .ZN(n6027) );
  NAND2_X1 U7599 ( .A1(n5773), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6025) );
  INV_X1 U7600 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6018) );
  OR2_X1 U7601 ( .A1(n5775), .A2(n6018), .ZN(n6024) );
  INV_X1 U7602 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7603 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7604 ( .A1(n6036), .A2(n6021), .ZN(n7651) );
  OR2_X1 U7605 ( .A1(n5774), .A2(n7651), .ZN(n6023) );
  INV_X1 U7606 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9399) );
  OR2_X1 U7607 ( .A1(n8771), .A2(n9399), .ZN(n6022) );
  NAND4_X1 U7608 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .ZN(n9297)
         );
  NAND2_X1 U7609 ( .A1(n9297), .A2(n6168), .ZN(n6026) );
  NAND2_X1 U7610 ( .A1(n6027), .A2(n6026), .ZN(n6028) );
  XNOR2_X1 U7611 ( .A(n6028), .B(n6241), .ZN(n6047) );
  AND2_X1 U7612 ( .A1(n9297), .A2(n6219), .ZN(n6029) );
  AOI21_X1 U7613 ( .B1(n7650), .B2(n6168), .A(n6029), .ZN(n8499) );
  NAND2_X1 U7614 ( .A1(n6745), .A2(n5758), .ZN(n6034) );
  NAND2_X1 U7615 ( .A1(n6030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6032) );
  XNOR2_X1 U7616 ( .A(n6032), .B(n6031), .ZN(n7367) );
  INV_X1 U7617 ( .A(n7367), .ZN(n9880) );
  AOI22_X1 U7618 ( .A1(n5759), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5780), .B2(
        n9880), .ZN(n6033) );
  NAND2_X1 U7619 ( .A1(n9308), .A2(n6239), .ZN(n6043) );
  NAND2_X1 U7620 ( .A1(n5773), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6041) );
  INV_X1 U7621 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9874) );
  OR2_X1 U7622 ( .A1(n8771), .A2(n9874), .ZN(n6040) );
  INV_X1 U7623 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7624 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7625 ( .A1(n6056), .A2(n6037), .ZN(n9310) );
  OR2_X1 U7626 ( .A1(n5774), .A2(n9310), .ZN(n6039) );
  INV_X1 U7627 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9311) );
  OR2_X1 U7628 ( .A1(n5775), .A2(n9311), .ZN(n6038) );
  NAND4_X1 U7629 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9282)
         );
  NAND2_X1 U7630 ( .A1(n9282), .A2(n6168), .ZN(n6042) );
  NAND2_X1 U7631 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  XNOR2_X1 U7632 ( .A(n6044), .B(n6241), .ZN(n8571) );
  NAND2_X1 U7633 ( .A1(n9308), .A2(n6168), .ZN(n6046) );
  NAND2_X1 U7634 ( .A1(n9282), .A2(n6219), .ZN(n6045) );
  NAND2_X1 U7635 ( .A1(n6046), .A2(n6045), .ZN(n8634) );
  NOR2_X1 U7636 ( .A1(n8571), .A2(n8634), .ZN(n6065) );
  INV_X1 U7637 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7638 ( .A1(n6786), .A2(n5758), .ZN(n6054) );
  NAND2_X1 U7639 ( .A1(n6049), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6050) );
  MUX2_X1 U7640 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6050), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n6052) );
  NAND2_X1 U7641 ( .A1(n6052), .A2(n6051), .ZN(n7369) );
  INV_X1 U7642 ( .A(n7369), .ZN(n7392) );
  AOI22_X1 U7643 ( .A1(n5759), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4271), .B2(
        n7392), .ZN(n6053) );
  NAND2_X1 U7644 ( .A1(n5773), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6061) );
  INV_X1 U7645 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7362) );
  OR2_X1 U7646 ( .A1(n8771), .A2(n7362), .ZN(n6060) );
  NAND2_X1 U7647 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7648 ( .A1(n6074), .A2(n6057), .ZN(n9275) );
  OR2_X1 U7649 ( .A1(n5774), .A2(n9275), .ZN(n6059) );
  INV_X1 U7650 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9276) );
  OR2_X1 U7651 ( .A1(n5775), .A2(n9276), .ZN(n6058) );
  NOR2_X1 U7652 ( .A1(n9260), .A2(n8531), .ZN(n6062) );
  AOI21_X1 U7653 ( .B1(n9389), .B2(n6168), .A(n6062), .ZN(n6068) );
  INV_X1 U7654 ( .A(n9389), .ZN(n9274) );
  OAI22_X1 U7655 ( .A1(n9274), .A2(n5735), .B1(n9260), .B2(n8532), .ZN(n6063)
         );
  XNOR2_X1 U7656 ( .A(n6063), .B(n6241), .ZN(n6067) );
  XOR2_X1 U7657 ( .A(n6068), .B(n6067), .Z(n8575) );
  AOI21_X1 U7658 ( .B1(n8571), .B2(n8634), .A(n8575), .ZN(n6064) );
  INV_X1 U7659 ( .A(n6067), .ZN(n6069) );
  NAND2_X1 U7660 ( .A1(n6790), .A2(n5758), .ZN(n6072) );
  XNOR2_X1 U7661 ( .A(n6070), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7440) );
  AOI22_X1 U7662 ( .A1(n5759), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4271), .B2(
        n7440), .ZN(n6071) );
  NAND2_X1 U7663 ( .A1(n9384), .A2(n6239), .ZN(n6081) );
  NAND2_X1 U7664 ( .A1(n5773), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6079) );
  INV_X1 U7665 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7666 ( .A1(n8771), .A2(n6073), .ZN(n6078) );
  INV_X1 U7667 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U7668 ( .A1(n6074), .A2(n9989), .ZN(n6075) );
  NAND2_X1 U7669 ( .A1(n6092), .A2(n6075), .ZN(n9253) );
  OR2_X1 U7670 ( .A1(n5774), .A2(n9253), .ZN(n6077) );
  INV_X1 U7671 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9254) );
  OR2_X1 U7672 ( .A1(n5775), .A2(n9254), .ZN(n6076) );
  OR2_X1 U7673 ( .A1(n9240), .A2(n8532), .ZN(n6080) );
  NAND2_X1 U7674 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  XNOR2_X1 U7675 ( .A(n6082), .B(n6241), .ZN(n6084) );
  OAI22_X1 U7676 ( .A1(n6392), .A2(n8532), .B1(n9240), .B2(n8531), .ZN(n6083)
         );
  XNOR2_X1 U7677 ( .A(n6084), .B(n6083), .ZN(n8582) );
  OR2_X1 U7678 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  OAI21_X2 U7679 ( .B1(n8583), .B2(n8582), .A(n6085), .ZN(n8623) );
  NAND2_X1 U7680 ( .A1(n6810), .A2(n5758), .ZN(n6091) );
  OR2_X1 U7681 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  AND2_X1 U7682 ( .A1(n6089), .A2(n6088), .ZN(n7443) );
  AOI22_X1 U7683 ( .A1(n5759), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5780), .B2(
        n7443), .ZN(n6090) );
  NAND2_X1 U7684 ( .A1(n6092), .A2(n7431), .ZN(n6093) );
  NAND2_X1 U7685 ( .A1(n6105), .A2(n6093), .ZN(n9243) );
  NAND2_X1 U7686 ( .A1(n6094), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7687 ( .B1(n9243), .B2(n5774), .A(n6095), .ZN(n6099) );
  INV_X1 U7688 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7689 ( .A1(n5773), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7690 ( .B1(n8771), .B2(n6097), .A(n6096), .ZN(n6098) );
  AOI22_X1 U7691 ( .A1(n9379), .A2(n6239), .B1(n6168), .B2(n8940), .ZN(n6100)
         );
  XNOR2_X1 U7692 ( .A(n6100), .B(n6241), .ZN(n6101) );
  OAI22_X1 U7693 ( .A1(n9247), .A2(n8532), .B1(n9262), .B2(n8531), .ZN(n8620)
         );
  INV_X1 U7694 ( .A(n6101), .ZN(n8621) );
  NAND2_X1 U7695 ( .A1(n6971), .A2(n5758), .ZN(n6103) );
  AOI22_X1 U7696 ( .A1(n5759), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5780), .B2(
        n9045), .ZN(n6102) );
  NAND2_X1 U7697 ( .A1(n9233), .A2(n6239), .ZN(n6110) );
  INV_X1 U7698 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9375) );
  INV_X1 U7699 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7700 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  NAND2_X1 U7701 ( .A1(n6119), .A2(n6106), .ZN(n9226) );
  OR2_X1 U7702 ( .A1(n9226), .A2(n5774), .ZN(n6108) );
  AOI22_X1 U7703 ( .A1(n6094), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5773), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7704 ( .C1(n8771), .C2(n9375), .A(n6108), .B(n6107), .ZN(n8939)
         );
  NAND2_X1 U7705 ( .A1(n8939), .A2(n6168), .ZN(n6109) );
  NAND2_X1 U7706 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  XNOR2_X1 U7707 ( .A(n6111), .B(n8529), .ZN(n8521) );
  AND2_X1 U7708 ( .A1(n8939), .A2(n6219), .ZN(n6112) );
  AOI21_X1 U7709 ( .B1(n9233), .B2(n6168), .A(n6112), .ZN(n8520) );
  INV_X1 U7710 ( .A(n8521), .ZN(n6114) );
  INV_X1 U7711 ( .A(n8520), .ZN(n6113) );
  NAND2_X1 U7712 ( .A1(n7061), .A2(n5758), .ZN(n6117) );
  NAND2_X1 U7713 ( .A1(n5759), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7714 ( .A1(n9368), .A2(n6239), .ZN(n6126) );
  NAND2_X1 U7715 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  AND2_X1 U7716 ( .A1(n6121), .A2(n6120), .ZN(n9214) );
  INV_X1 U7717 ( .A(n5774), .ZN(n6232) );
  NAND2_X1 U7718 ( .A1(n9214), .A2(n6232), .ZN(n6124) );
  AOI22_X1 U7719 ( .A1(n6413), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5773), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7720 ( .A1(n6094), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6122) );
  OR2_X1 U7721 ( .A1(n9221), .A2(n8532), .ZN(n6125) );
  NAND2_X1 U7722 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  XNOR2_X1 U7723 ( .A(n6127), .B(n8529), .ZN(n6130) );
  INV_X1 U7724 ( .A(n6130), .ZN(n6132) );
  NOR2_X1 U7725 ( .A1(n9221), .A2(n8531), .ZN(n6128) );
  AOI21_X1 U7726 ( .B1(n9368), .B2(n6168), .A(n6128), .ZN(n6129) );
  INV_X1 U7727 ( .A(n6129), .ZN(n6131) );
  AND2_X1 U7728 ( .A1(n6130), .A2(n6129), .ZN(n6133) );
  AOI21_X1 U7729 ( .B1(n6132), .B2(n6131), .A(n6133), .ZN(n8601) );
  XOR2_X1 U7730 ( .A(n6136), .B(n6137), .Z(n8555) );
  AND2_X1 U7731 ( .A1(n8601), .A2(n8555), .ZN(n6135) );
  INV_X1 U7732 ( .A(n8555), .ZN(n6134) );
  INV_X1 U7733 ( .A(n6133), .ZN(n8552) );
  INV_X1 U7734 ( .A(n6152), .ZN(n6150) );
  NAND2_X1 U7735 ( .A1(n5759), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6138) );
  INV_X1 U7736 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U7737 ( .A1(n6140), .A2(n8614), .ZN(n6141) );
  NAND2_X1 U7738 ( .A1(n6157), .A2(n6141), .ZN(n9175) );
  OR2_X1 U7739 ( .A1(n9175), .A2(n5774), .ZN(n6147) );
  INV_X1 U7740 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7741 ( .A1(n5773), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7742 ( .A1(n6413), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6142) );
  OAI211_X1 U7743 ( .C1(n5775), .C2(n6144), .A(n6143), .B(n6142), .ZN(n6145)
         );
  INV_X1 U7744 ( .A(n6145), .ZN(n6146) );
  AOI22_X1 U7745 ( .A1(n9357), .A2(n6239), .B1(n6168), .B2(n9194), .ZN(n6148)
         );
  XNOR2_X1 U7746 ( .A(n6148), .B(n6241), .ZN(n6151) );
  INV_X1 U7747 ( .A(n6151), .ZN(n6149) );
  NAND2_X1 U7748 ( .A1(n6150), .A2(n6149), .ZN(n6153) );
  NAND2_X2 U7749 ( .A1(n6152), .A2(n6151), .ZN(n8513) );
  OAI22_X1 U7750 ( .A1(n9178), .A2(n8532), .B1(n9156), .B2(n8531), .ZN(n8613)
         );
  NAND2_X1 U7751 ( .A1(n7421), .A2(n5758), .ZN(n6156) );
  NAND2_X1 U7752 ( .A1(n5759), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7753 ( .A1(n9171), .A2(n6239), .ZN(n6165) );
  INV_X1 U7754 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U7755 ( .A1(n6157), .A2(n8515), .ZN(n6158) );
  NAND2_X1 U7756 ( .A1(n6177), .A2(n6158), .ZN(n9166) );
  OR2_X1 U7757 ( .A1(n9166), .A2(n5774), .ZN(n6163) );
  INV_X1 U7758 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U7759 ( .A1(n5773), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7760 ( .A1(n6413), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7761 ( .C1(n5775), .C2(n9165), .A(n6160), .B(n6159), .ZN(n6161)
         );
  INV_X1 U7762 ( .A(n6161), .ZN(n6162) );
  NAND2_X1 U7763 ( .A1(n8937), .A2(n6168), .ZN(n6164) );
  NAND2_X1 U7764 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  XNOR2_X1 U7765 ( .A(n6166), .B(n8529), .ZN(n6169) );
  AND2_X1 U7766 ( .A1(n8937), .A2(n6219), .ZN(n6167) );
  AOI21_X1 U7767 ( .B1(n9171), .B2(n6168), .A(n6167), .ZN(n6170) );
  NAND2_X1 U7768 ( .A1(n6169), .A2(n6170), .ZN(n6174) );
  INV_X1 U7769 ( .A(n6169), .ZN(n6172) );
  INV_X1 U7770 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7771 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7772 ( .A1(n6174), .A2(n6173), .ZN(n8512) );
  INV_X1 U7773 ( .A(n6174), .ZN(n8592) );
  NAND2_X1 U7774 ( .A1(n7510), .A2(n5758), .ZN(n6176) );
  NAND2_X1 U7775 ( .A1(n5759), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6175) );
  INV_X1 U7776 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U7777 ( .A1(n6177), .A2(n8595), .ZN(n6178) );
  AND2_X1 U7778 ( .A1(n6197), .A2(n6178), .ZN(n9149) );
  NAND2_X1 U7779 ( .A1(n9149), .A2(n6232), .ZN(n6184) );
  INV_X1 U7780 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7781 ( .A1(n5773), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7782 ( .A1(n6413), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6179) );
  OAI211_X1 U7783 ( .C1(n5775), .C2(n6181), .A(n6180), .B(n6179), .ZN(n6182)
         );
  INV_X1 U7784 ( .A(n6182), .ZN(n6183) );
  AND2_X2 U7785 ( .A1(n6184), .A2(n6183), .ZN(n9157) );
  OAI22_X1 U7786 ( .A1(n9152), .A2(n5735), .B1(n9157), .B2(n8532), .ZN(n6185)
         );
  XNOR2_X1 U7787 ( .A(n6185), .B(n8529), .ZN(n6188) );
  OR2_X1 U7788 ( .A1(n9152), .A2(n8532), .ZN(n6187) );
  INV_X1 U7789 ( .A(n9157), .ZN(n8936) );
  NAND2_X1 U7790 ( .A1(n8936), .A2(n6219), .ZN(n6186) );
  NAND2_X1 U7791 ( .A1(n6188), .A2(n6189), .ZN(n6193) );
  INV_X1 U7792 ( .A(n6188), .ZN(n6191) );
  INV_X1 U7793 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7794 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  NAND2_X1 U7795 ( .A1(n7589), .A2(n5758), .ZN(n6195) );
  NAND2_X1 U7796 ( .A1(n5759), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6194) );
  INV_X1 U7797 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U7798 ( .A1(n6197), .A2(n8565), .ZN(n6198) );
  NAND2_X1 U7799 ( .A1(n6211), .A2(n6198), .ZN(n9135) );
  INV_X1 U7800 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U7801 ( .A1(n6413), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7802 ( .A1(n5773), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6199) );
  OAI211_X1 U7803 ( .C1(n9126), .C2(n5775), .A(n6200), .B(n6199), .ZN(n6201)
         );
  INV_X1 U7804 ( .A(n6201), .ZN(n6202) );
  OAI22_X1 U7805 ( .A1(n9127), .A2(n8532), .B1(n9147), .B2(n8531), .ZN(n6224)
         );
  NAND2_X1 U7806 ( .A1(n9343), .A2(n6239), .ZN(n6205) );
  NAND2_X1 U7807 ( .A1(n9116), .A2(n6168), .ZN(n6204) );
  NAND2_X1 U7808 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  XNOR2_X1 U7809 ( .A(n6206), .B(n6241), .ZN(n6223) );
  XOR2_X1 U7810 ( .A(n6224), .B(n6223), .Z(n8563) );
  NAND2_X1 U7811 ( .A1(n7608), .A2(n5758), .ZN(n6208) );
  NAND2_X1 U7812 ( .A1(n5759), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7813 ( .A1(n9112), .A2(n8532), .ZN(n6221) );
  INV_X1 U7814 ( .A(n6211), .ZN(n6209) );
  INV_X1 U7815 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7816 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U7817 ( .A1(n6230), .A2(n6212), .ZN(n6304) );
  INV_X1 U7818 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7819 ( .A1(n6413), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7820 ( .A1(n5773), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6213) );
  OAI211_X1 U7821 ( .C1(n6215), .C2(n5775), .A(n6214), .B(n6213), .ZN(n6216)
         );
  INV_X1 U7822 ( .A(n6216), .ZN(n6217) );
  INV_X1 U7823 ( .A(n9134), .ZN(n8935) );
  NAND2_X1 U7824 ( .A1(n8935), .A2(n6219), .ZN(n6220) );
  NAND2_X1 U7825 ( .A1(n6221), .A2(n6220), .ZN(n6244) );
  OAI22_X1 U7826 ( .A1(n9112), .A2(n5735), .B1(n9134), .B2(n8532), .ZN(n6222)
         );
  XNOR2_X1 U7827 ( .A(n6222), .B(n6241), .ZN(n6245) );
  XOR2_X1 U7828 ( .A(n6244), .B(n6245), .Z(n6301) );
  INV_X1 U7829 ( .A(n6223), .ZN(n6226) );
  INV_X1 U7830 ( .A(n6224), .ZN(n6225) );
  NAND2_X1 U7831 ( .A1(n6226), .A2(n6225), .ZN(n6300) );
  NAND2_X1 U7832 ( .A1(n7640), .A2(n5758), .ZN(n6229) );
  NAND2_X1 U7833 ( .A1(n5759), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6228) );
  INV_X1 U7834 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U7835 ( .A1(n6230), .A2(n9906), .ZN(n6231) );
  NAND2_X1 U7836 ( .A1(n9102), .A2(n6232), .ZN(n6238) );
  INV_X1 U7837 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7838 ( .A1(n5773), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7839 ( .A1(n6413), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U7840 ( .C1(n6235), .C2(n5775), .A(n6234), .B(n6233), .ZN(n6236)
         );
  INV_X1 U7841 ( .A(n6236), .ZN(n6237) );
  AOI22_X1 U7842 ( .A1(n9101), .A2(n6239), .B1(n6168), .B2(n9117), .ZN(n6240)
         );
  XOR2_X1 U7843 ( .A(n6241), .B(n6240), .Z(n6243) );
  OAI22_X1 U7844 ( .A1(n6394), .A2(n8532), .B1(n8540), .B2(n8531), .ZN(n6242)
         );
  NOR2_X1 U7845 ( .A1(n6243), .A2(n6242), .ZN(n8546) );
  AOI21_X1 U7846 ( .B1(n6243), .B2(n6242), .A(n8546), .ZN(n6247) );
  NAND2_X1 U7847 ( .A1(n6245), .A2(n6244), .ZN(n6248) );
  INV_X1 U7848 ( .A(n8539), .ZN(n8536) );
  NOR2_X1 U7849 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n10009) );
  NOR4_X1 U7850 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6251) );
  NOR4_X1 U7851 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6250) );
  NOR4_X1 U7852 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6249) );
  NAND4_X1 U7853 ( .A1(n10009), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n6257)
         );
  NOR4_X1 U7854 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U7855 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U7856 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6253) );
  NOR4_X1 U7857 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6252) );
  NAND4_X1 U7858 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n6256)
         );
  NOR2_X1 U7859 ( .A1(n6257), .A2(n6256), .ZN(n6422) );
  NAND2_X1 U7860 ( .A1(n7591), .A2(P1_B_REG_SCAN_IN), .ZN(n6258) );
  MUX2_X1 U7861 ( .A(P1_B_REG_SCAN_IN), .B(n6258), .S(n7512), .Z(n6259) );
  INV_X1 U7862 ( .A(n6260), .ZN(n7612) );
  NAND2_X1 U7863 ( .A1(n7612), .A2(n7512), .ZN(n9443) );
  INV_X1 U7864 ( .A(n6814), .ZN(n6431) );
  NAND2_X1 U7865 ( .A1(n7612), .A2(n7591), .ZN(n9442) );
  OAI21_X1 U7866 ( .B1(n6421), .B2(P1_D_REG_1__SCAN_IN), .A(n9442), .ZN(n6426)
         );
  INV_X1 U7867 ( .A(n6426), .ZN(n6815) );
  OAI211_X1 U7868 ( .C1(n6422), .C2(n6421), .A(n6431), .B(n6815), .ZN(n6288)
         );
  NAND2_X1 U7869 ( .A1(n6261), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6263) );
  INV_X1 U7870 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6262) );
  INV_X1 U7871 ( .A(n6531), .ZN(n6295) );
  NOR2_X1 U7872 ( .A1(n6288), .A2(n6295), .ZN(n6293) );
  NOR2_X1 U7873 ( .A1(n9567), .A2(n8905), .ZN(n6267) );
  OAI21_X1 U7874 ( .B1(n8536), .B2(n6268), .A(n8603), .ZN(n6298) );
  INV_X1 U7875 ( .A(n6271), .ZN(n6269) );
  NAND2_X1 U7876 ( .A1(n6269), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9065) );
  INV_X1 U7877 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7878 ( .A1(n6271), .A2(n6270), .ZN(n6272) );
  NAND2_X1 U7879 ( .A1(n9065), .A2(n6272), .ZN(n8541) );
  OR2_X1 U7880 ( .A1(n8541), .A2(n5774), .ZN(n6277) );
  INV_X1 U7881 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U7882 ( .A1(n6413), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7883 ( .A1(n5773), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6273) );
  OAI211_X1 U7884 ( .C1(n9084), .C2(n5775), .A(n6274), .B(n6273), .ZN(n6275)
         );
  INV_X1 U7885 ( .A(n6275), .ZN(n6276) );
  INV_X1 U7886 ( .A(n6288), .ZN(n6283) );
  NOR2_X1 U7887 ( .A1(n6278), .A2(n6389), .ZN(n6279) );
  NAND2_X1 U7888 ( .A1(n6531), .A2(n6279), .ZN(n8911) );
  INV_X1 U7889 ( .A(n6280), .ZN(n8960) );
  NOR2_X1 U7890 ( .A1(n8911), .A2(n8960), .ZN(n6281) );
  NOR2_X1 U7891 ( .A1(n8911), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U7892 ( .A1(n6283), .A2(n6282), .ZN(n8624) );
  INV_X1 U7893 ( .A(n9567), .ZN(n9592) );
  NAND2_X1 U7894 ( .A1(n6288), .A2(n9592), .ZN(n6284) );
  NAND2_X1 U7895 ( .A1(n8905), .A2(n6266), .ZN(n6424) );
  NAND3_X1 U7896 ( .A1(n6284), .A2(n6441), .A3(n6424), .ZN(n6285) );
  NAND2_X1 U7897 ( .A1(n6285), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6290) );
  INV_X1 U7898 ( .A(n8893), .ZN(n8907) );
  NAND2_X1 U7899 ( .A1(n9557), .A2(n8907), .ZN(n6828) );
  NOR2_X1 U7900 ( .A1(n6828), .A2(P1_U3086), .ZN(n6287) );
  OR2_X1 U7901 ( .A1(n6532), .A2(P1_U3086), .ZN(n8924) );
  INV_X1 U7902 ( .A(n8924), .ZN(n8915) );
  AOI21_X1 U7903 ( .B1(n6288), .B2(n6287), .A(n8915), .ZN(n6289) );
  NAND2_X1 U7904 ( .A1(n6290), .A2(n6289), .ZN(n8607) );
  AOI22_X1 U7905 ( .A1(n9102), .A2(n8607), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6291) );
  OAI21_X1 U7906 ( .B1(n9134), .B2(n8624), .A(n6291), .ZN(n6292) );
  AOI21_X1 U7907 ( .B1(n8934), .B2(n8627), .A(n6292), .ZN(n6297) );
  INV_X1 U7908 ( .A(n6293), .ZN(n6294) );
  OR2_X1 U7909 ( .A1(n6294), .A2(n6828), .ZN(n6296) );
  NAND2_X1 U7910 ( .A1(n9229), .A2(n9045), .ZN(n6427) );
  NAND3_X1 U7911 ( .A1(n6298), .A2(n6297), .A3(n4846), .ZN(P1_U3214) );
  AND2_X1 U7912 ( .A1(n6299), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7913 ( .A1(n6303), .A2(n8603), .ZN(n6310) );
  INV_X1 U7914 ( .A(n6304), .ZN(n9110) );
  AOI22_X1 U7915 ( .A1(n9110), .A2(n8607), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n6305) );
  OAI21_X1 U7916 ( .B1(n9147), .B2(n8624), .A(n6305), .ZN(n6306) );
  AOI21_X1 U7917 ( .B1(n9117), .B2(n8627), .A(n6306), .ZN(n6307) );
  OAI21_X1 U7918 ( .B1(n6311), .B2(n6310), .A(n6309), .ZN(P1_U3240) );
  NAND2_X1 U7919 ( .A1(n7854), .A2(n6328), .ZN(n6312) );
  NAND2_X1 U7920 ( .A1(n6315), .A2(n6314), .ZN(n6325) );
  AND2_X1 U7921 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  INV_X1 U7922 ( .A(SI_28_), .ZN(n6320) );
  INV_X1 U7923 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6323) );
  INV_X1 U7924 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U7925 ( .A(n6323), .B(n6322), .S(n7731), .Z(n7708) );
  OR2_X1 U7926 ( .A1(n7737), .A2(n6323), .ZN(n6324) );
  NAND2_X1 U7927 ( .A1(n6345), .A2(n7009), .ZN(n7719) );
  NAND2_X1 U7928 ( .A1(n7856), .A2(n7719), .ZN(n7850) );
  XNOR2_X1 U7929 ( .A(n6325), .B(n7915), .ZN(n6341) );
  NAND2_X1 U7930 ( .A1(n8260), .A2(n6328), .ZN(n6326) );
  OR2_X1 U7931 ( .A1(n8260), .A2(n6328), .ZN(n6329) );
  NAND2_X1 U7932 ( .A1(n6330), .A2(n6329), .ZN(n7705) );
  INV_X1 U7933 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7934 ( .A1(n5164), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U7935 ( .A1(n5408), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6331) );
  OAI211_X1 U7936 ( .C1(n6334), .C2(n6333), .A(n6332), .B(n6331), .ZN(n6335)
         );
  INV_X1 U7937 ( .A(n6335), .ZN(n6336) );
  NAND2_X1 U7938 ( .A1(n7726), .A2(n6336), .ZN(n8129) );
  NAND2_X1 U7939 ( .A1(n6337), .A2(P2_B_REG_SCAN_IN), .ZN(n6338) );
  AND2_X1 U7940 ( .A1(n8362), .A2(n6338), .ZN(n8249) );
  AOI22_X1 U7941 ( .A1(n8130), .A2(n8360), .B1(n8129), .B2(n8249), .ZN(n6339)
         );
  OAI21_X1 U7942 ( .B1(n7995), .B2(n7031), .A(n6339), .ZN(n6340) );
  NAND2_X1 U7943 ( .A1(n7994), .A2(n6342), .ZN(n6349) );
  INV_X1 U7944 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7945 ( .A1(n9848), .A2(n6343), .ZN(n6344) );
  OAI21_X1 U7946 ( .B1(n6349), .B2(n9848), .A(n6344), .ZN(n6346) );
  INV_X1 U7947 ( .A(n6345), .ZN(n7999) );
  NAND2_X1 U7948 ( .A1(n6346), .A2(n4842), .ZN(P2_U3488) );
  NAND2_X1 U7949 ( .A1(n9831), .A2(n6347), .ZN(n6348) );
  OAI21_X1 U7950 ( .B1(n6349), .B2(n9831), .A(n6348), .ZN(n6350) );
  NAND2_X1 U7951 ( .A1(n6350), .A2(n4848), .ZN(P2_U3456) );
  NAND2_X1 U7952 ( .A1(n6351), .A2(n9556), .ZN(n6813) );
  NAND2_X1 U7953 ( .A1(n6397), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U7954 ( .A1(n6822), .A2(n6897), .ZN(n8671) );
  NAND2_X1 U7955 ( .A1(n5757), .A2(n9560), .ZN(n8821) );
  NAND2_X1 U7956 ( .A1(n6885), .A2(n8784), .ZN(n6884) );
  NAND2_X1 U7957 ( .A1(n6884), .A2(n6352), .ZN(n6850) );
  NAND2_X1 U7958 ( .A1(n6886), .A2(n6854), .ZN(n8823) );
  INV_X1 U7959 ( .A(n6886), .ZN(n8946) );
  NAND2_X1 U7960 ( .A1(n8946), .A2(n6941), .ZN(n8825) );
  NAND2_X1 U7961 ( .A1(n8823), .A2(n8825), .ZN(n6852) );
  NAND2_X1 U7962 ( .A1(n6850), .A2(n6852), .ZN(n6851) );
  NAND2_X1 U7963 ( .A1(n6851), .A2(n4856), .ZN(n6946) );
  NAND2_X1 U7964 ( .A1(n8663), .A2(n9566), .ZN(n7101) );
  NAND2_X1 U7965 ( .A1(n7101), .A2(n8826), .ZN(n8787) );
  NAND2_X1 U7966 ( .A1(n6946), .A2(n8787), .ZN(n6945) );
  NAND2_X1 U7967 ( .A1(n6945), .A2(n6353), .ZN(n7097) );
  NAND2_X1 U7968 ( .A1(n6959), .A2(n7107), .ZN(n8676) );
  NAND2_X1 U7969 ( .A1(n7073), .A2(n9543), .ZN(n8829) );
  NAND2_X1 U7970 ( .A1(n8676), .A2(n8829), .ZN(n8789) );
  NAND2_X1 U7971 ( .A1(n7050), .A2(n7074), .ZN(n8679) );
  NAND2_X1 U7972 ( .A1(n8944), .A2(n9575), .ZN(n7042) );
  NAND2_X1 U7973 ( .A1(n8679), .A2(n7042), .ZN(n8790) );
  NAND2_X1 U7974 ( .A1(n7085), .A2(n7051), .ZN(n8680) );
  INV_X1 U7975 ( .A(n7051), .ZN(n7198) );
  NAND2_X1 U7976 ( .A1(n7198), .A2(n5866), .ZN(n8687) );
  NAND2_X1 U7977 ( .A1(n8680), .A2(n8687), .ZN(n7041) );
  NAND2_X1 U7978 ( .A1(n7040), .A2(n7041), .ZN(n7039) );
  OAI21_X1 U7979 ( .B1(n5866), .B2(n7051), .A(n7039), .ZN(n7092) );
  OR2_X1 U7980 ( .A1(n7206), .A2(n7331), .ZN(n8692) );
  NAND2_X1 U7981 ( .A1(n7206), .A2(n7331), .ZN(n8683) );
  NAND2_X1 U7982 ( .A1(n8692), .A2(n8683), .ZN(n7091) );
  NAND2_X1 U7983 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  INV_X1 U7984 ( .A(n7331), .ZN(n6993) );
  NAND2_X1 U7985 ( .A1(n6391), .A2(n7331), .ZN(n6354) );
  NAND2_X1 U7986 ( .A1(n7090), .A2(n6354), .ZN(n7305) );
  NAND2_X1 U7987 ( .A1(n7307), .A2(n7401), .ZN(n8702) );
  NAND2_X1 U7988 ( .A1(n8701), .A2(n8702), .ZN(n7304) );
  NAND2_X1 U7989 ( .A1(n7305), .A2(n7304), .ZN(n7303) );
  NAND2_X1 U7990 ( .A1(n7303), .A2(n6355), .ZN(n7396) );
  OR2_X1 U7991 ( .A1(n7523), .A2(n7600), .ZN(n8835) );
  NAND2_X1 U7992 ( .A1(n7523), .A2(n7600), .ZN(n8705) );
  NAND2_X1 U7993 ( .A1(n8835), .A2(n8705), .ZN(n8783) );
  NAND2_X1 U7994 ( .A1(n7396), .A2(n8783), .ZN(n7395) );
  INV_X1 U7995 ( .A(n7600), .ZN(n8943) );
  NAND2_X1 U7996 ( .A1(n6356), .A2(n7600), .ZN(n6357) );
  NAND2_X1 U7997 ( .A1(n7395), .A2(n6357), .ZN(n7475) );
  NAND2_X1 U7998 ( .A1(n7605), .A2(n7632), .ZN(n8706) );
  NAND2_X1 U7999 ( .A1(n8709), .A2(n8706), .ZN(n8798) );
  INV_X1 U8000 ( .A(n7605), .ZN(n9593) );
  INV_X1 U8001 ( .A(n7632), .ZN(n6358) );
  AOI21_X2 U8002 ( .B1(n7475), .B2(n8798), .A(n6359), .ZN(n7533) );
  OR2_X1 U8003 ( .A1(n7637), .A2(n8942), .ZN(n6360) );
  NAND2_X1 U8004 ( .A1(n7533), .A2(n6360), .ZN(n6361) );
  INV_X1 U8005 ( .A(n7637), .ZN(n7577) );
  OR2_X1 U8006 ( .A1(n7674), .A2(n7529), .ZN(n8845) );
  NAND2_X1 U8007 ( .A1(n7674), .A2(n7529), .ZN(n8719) );
  NAND2_X1 U8008 ( .A1(n8845), .A2(n8719), .ZN(n8803) );
  INV_X1 U8009 ( .A(n7529), .ZN(n8941) );
  NOR2_X1 U8010 ( .A1(n7650), .A2(n9297), .ZN(n6362) );
  INV_X1 U8011 ( .A(n9297), .ZN(n7660) );
  INV_X1 U8012 ( .A(n9282), .ZN(n8505) );
  NAND2_X1 U8013 ( .A1(n9389), .A2(n9260), .ZN(n8855) );
  NAND2_X1 U8014 ( .A1(n8723), .A2(n8855), .ZN(n9271) );
  NAND2_X1 U8015 ( .A1(n9272), .A2(n9271), .ZN(n9270) );
  NAND2_X1 U8016 ( .A1(n9270), .A2(n4849), .ZN(n9252) );
  NAND2_X1 U8017 ( .A1(n9384), .A2(n9240), .ZN(n8733) );
  NAND2_X1 U8018 ( .A1(n8737), .A2(n8733), .ZN(n9251) );
  NAND2_X1 U8019 ( .A1(n9225), .A2(n6365), .ZN(n6366) );
  INV_X1 U8020 ( .A(n8939), .ZN(n9241) );
  NAND2_X1 U8021 ( .A1(n6366), .A2(n4850), .ZN(n9209) );
  NAND2_X1 U8022 ( .A1(n9368), .A2(n9221), .ZN(n9188) );
  NAND2_X1 U8023 ( .A1(n9189), .A2(n9188), .ZN(n9210) );
  NAND2_X1 U8024 ( .A1(n9209), .A2(n9210), .ZN(n6368) );
  INV_X1 U8025 ( .A(n9221), .ZN(n9193) );
  NAND2_X1 U8026 ( .A1(n9368), .A2(n9193), .ZN(n6367) );
  NAND2_X1 U8027 ( .A1(n6368), .A2(n6367), .ZN(n9197) );
  NOR2_X1 U8028 ( .A1(n9424), .A2(n9212), .ZN(n6369) );
  INV_X1 U8029 ( .A(n9212), .ZN(n8938) );
  NOR2_X1 U8030 ( .A1(n9357), .A2(n9194), .ZN(n9160) );
  OR2_X1 U8031 ( .A1(n9171), .A2(n8937), .ZN(n8653) );
  INV_X1 U8032 ( .A(n8653), .ZN(n6371) );
  OR2_X1 U8033 ( .A1(n9160), .A2(n6371), .ZN(n9139) );
  AND2_X1 U8034 ( .A1(n9152), .A2(n9157), .ZN(n6374) );
  OR2_X1 U8035 ( .A1(n9152), .A2(n9157), .ZN(n6372) );
  NAND2_X1 U8036 ( .A1(n9357), .A2(n9194), .ZN(n9161) );
  NAND2_X1 U8037 ( .A1(n9171), .A2(n8937), .ZN(n8652) );
  AND2_X1 U8038 ( .A1(n9161), .A2(n8652), .ZN(n6370) );
  AND2_X1 U8039 ( .A1(n6372), .A2(n9140), .ZN(n6373) );
  NOR2_X1 U8040 ( .A1(n9112), .A2(n9134), .ZN(n6375) );
  NAND2_X1 U8041 ( .A1(n9112), .A2(n9134), .ZN(n6376) );
  NAND2_X1 U8042 ( .A1(n9101), .A2(n8540), .ZN(n8757) );
  NAND2_X1 U8043 ( .A1(n8886), .A2(n8757), .ZN(n9089) );
  NOR2_X1 U8044 ( .A1(n9101), .A2(n9117), .ZN(n6378) );
  NAND2_X1 U8045 ( .A1(n7961), .A2(n5758), .ZN(n6380) );
  NAND2_X1 U8046 ( .A1(n5759), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8047 ( .A1(n7958), .A2(n5758), .ZN(n6382) );
  NAND2_X1 U8048 ( .A1(n5759), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6381) );
  OR2_X1 U8049 ( .A1(n9065), .A2(n5774), .ZN(n6387) );
  INV_X1 U8050 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U8051 ( .A1(n6094), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8052 ( .A1(n5773), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6383) );
  OAI211_X1 U8053 ( .C1(n9929), .C2(n8771), .A(n6384), .B(n6383), .ZN(n6385)
         );
  INV_X1 U8054 ( .A(n6385), .ZN(n6386) );
  NAND2_X1 U8055 ( .A1(n6396), .A2(n8543), .ZN(n8888) );
  INV_X1 U8056 ( .A(n6266), .ZN(n6388) );
  MUX2_X1 U8057 ( .A(n6389), .B(n6388), .S(n6278), .Z(n6390) );
  INV_X1 U8058 ( .A(n9557), .ZN(n6925) );
  NAND2_X1 U8059 ( .A1(n6390), .A2(n6925), .ZN(n6848) );
  NAND2_X1 U8060 ( .A1(n9064), .A2(n9595), .ZN(n6420) );
  NAND2_X1 U8061 ( .A1(n6894), .A2(n9560), .ZN(n6893) );
  NOR2_X1 U8062 ( .A1(n6952), .A2(n9566), .ZN(n7098) );
  AND2_X1 U8063 ( .A1(n7098), .A2(n9543), .ZN(n7099) );
  NAND2_X1 U8064 ( .A1(n7402), .A2(n6356), .ZN(n7477) );
  INV_X1 U8065 ( .A(n7674), .ZN(n7622) );
  NAND2_X1 U8066 ( .A1(n9127), .A2(n9148), .ZN(n9123) );
  INV_X1 U8067 ( .A(n9081), .ZN(n6395) );
  AOI211_X1 U8068 ( .C1(n6396), .C2(n6395), .A(n9306), .B(n4293), .ZN(n9070)
         );
  INV_X1 U8069 ( .A(n6397), .ZN(n6821) );
  INV_X1 U8070 ( .A(n5743), .ZN(n6887) );
  NAND2_X1 U8071 ( .A1(n6887), .A2(n7952), .ZN(n6398) );
  NAND2_X1 U8072 ( .A1(n6820), .A2(n6398), .ZN(n8670) );
  INV_X1 U8073 ( .A(n8671), .ZN(n6399) );
  AND2_X1 U8074 ( .A1(n8661), .A2(n8821), .ZN(n8828) );
  INV_X1 U8075 ( .A(n6852), .ZN(n8786) );
  NAND2_X1 U8076 ( .A1(n8828), .A2(n8786), .ZN(n6844) );
  NAND2_X1 U8077 ( .A1(n6844), .A2(n8823), .ZN(n6948) );
  INV_X1 U8078 ( .A(n8787), .ZN(n6949) );
  AND2_X1 U8079 ( .A1(n7101), .A2(n8676), .ZN(n8831) );
  NAND2_X1 U8080 ( .A1(n7102), .A2(n8831), .ZN(n7043) );
  NAND2_X1 U8081 ( .A1(n7043), .A2(n8829), .ZN(n6957) );
  AND2_X1 U8082 ( .A1(n8683), .A2(n8680), .ZN(n8690) );
  INV_X1 U8083 ( .A(n8679), .ZN(n8688) );
  NOR2_X1 U8084 ( .A1(n6400), .A2(n8688), .ZN(n8833) );
  INV_X1 U8085 ( .A(n6400), .ZN(n8797) );
  INV_X1 U8086 ( .A(n8687), .ZN(n8791) );
  INV_X1 U8087 ( .A(n7042), .ZN(n6401) );
  NAND2_X1 U8088 ( .A1(n7397), .A2(n8705), .ZN(n7471) );
  NAND2_X1 U8089 ( .A1(n7637), .A2(n7616), .ZN(n8841) );
  AND2_X1 U8090 ( .A1(n8841), .A2(n8706), .ZN(n8697) );
  NAND2_X1 U8091 ( .A1(n7526), .A2(n8697), .ZN(n6403) );
  OR2_X1 U8092 ( .A1(n7637), .A2(n7616), .ZN(n8710) );
  OR2_X1 U8093 ( .A1(n7650), .A2(n7660), .ZN(n8846) );
  NAND2_X1 U8094 ( .A1(n7650), .A2(n7660), .ZN(n8722) );
  NAND2_X1 U8095 ( .A1(n8846), .A2(n8722), .ZN(n7643) );
  INV_X1 U8096 ( .A(n8719), .ZN(n8843) );
  NOR2_X1 U8097 ( .A1(n7643), .A2(n8843), .ZN(n6404) );
  NAND2_X1 U8098 ( .A1(n6405), .A2(n8846), .ZN(n9292) );
  OR2_X1 U8099 ( .A1(n9308), .A2(n8505), .ZN(n8728) );
  NAND2_X1 U8100 ( .A1(n9308), .A2(n8505), .ZN(n9281) );
  NAND2_X1 U8101 ( .A1(n8728), .A2(n9281), .ZN(n9291) );
  OR2_X2 U8102 ( .A1(n9292), .A2(n9291), .ZN(n9294) );
  INV_X1 U8103 ( .A(n9281), .ZN(n8716) );
  NOR2_X1 U8104 ( .A1(n9271), .A2(n8716), .ZN(n6406) );
  INV_X1 U8105 ( .A(n9251), .ZN(n9257) );
  OR2_X1 U8106 ( .A1(n9379), .A2(n9262), .ZN(n8738) );
  NAND2_X1 U8107 ( .A1(n9379), .A2(n9262), .ZN(n8736) );
  NAND2_X1 U8108 ( .A1(n8738), .A2(n8736), .ZN(n9237) );
  OR2_X1 U8109 ( .A1(n9233), .A2(n9241), .ZN(n8660) );
  NAND2_X1 U8110 ( .A1(n9233), .A2(n9241), .ZN(n8872) );
  NAND2_X1 U8111 ( .A1(n9220), .A2(n9224), .ZN(n9219) );
  AND2_X1 U8112 ( .A1(n8782), .A2(n9189), .ZN(n8868) );
  NAND2_X1 U8113 ( .A1(n8897), .A2(n8868), .ZN(n6407) );
  NAND2_X1 U8114 ( .A1(n9201), .A2(n9212), .ZN(n8781) );
  NAND2_X1 U8115 ( .A1(n8781), .A2(n9188), .ZN(n8735) );
  NAND2_X1 U8116 ( .A1(n8735), .A2(n8782), .ZN(n8876) );
  NAND2_X1 U8117 ( .A1(n6407), .A2(n8876), .ZN(n9180) );
  OR2_X1 U8118 ( .A1(n9357), .A2(n9156), .ZN(n8863) );
  NAND2_X1 U8119 ( .A1(n9357), .A2(n9156), .ZN(n8875) );
  NAND2_X1 U8120 ( .A1(n8863), .A2(n8875), .ZN(n9179) );
  OR2_X1 U8121 ( .A1(n9171), .A2(n9181), .ZN(n8864) );
  NAND2_X1 U8122 ( .A1(n9171), .A2(n9181), .ZN(n8861) );
  NAND2_X1 U8123 ( .A1(n9348), .A2(n9157), .ZN(n8862) );
  OR2_X1 U8124 ( .A1(n9343), .A2(n9147), .ZN(n8780) );
  AND2_X1 U8125 ( .A1(n8780), .A2(n9129), .ZN(n8867) );
  NAND2_X1 U8126 ( .A1(n9343), .A2(n9147), .ZN(n8779) );
  NAND2_X1 U8127 ( .A1(n9337), .A2(n9134), .ZN(n8881) );
  NAND2_X1 U8128 ( .A1(n9092), .A2(n4546), .ZN(n9091) );
  NAND2_X1 U8129 ( .A1(n9091), .A2(n8757), .ZN(n9077) );
  NAND2_X1 U8130 ( .A1(n9327), .A2(n9094), .ZN(n8759) );
  NAND2_X1 U8131 ( .A1(n9077), .A2(n9078), .ZN(n9076) );
  NAND2_X1 U8132 ( .A1(n9076), .A2(n8759), .ZN(n6408) );
  XNOR2_X1 U8133 ( .A(n6408), .B(n8815), .ZN(n6410) );
  NAND2_X1 U8134 ( .A1(n8921), .A2(n9045), .ZN(n6409) );
  NAND2_X1 U8135 ( .A1(n6265), .A2(n8907), .ZN(n8923) );
  OR2_X1 U8136 ( .A1(n6410), .A2(n9553), .ZN(n6418) );
  INV_X1 U8137 ( .A(n8905), .ZN(n6411) );
  INV_X1 U8138 ( .A(n8959), .ZN(n6609) );
  NAND2_X1 U8139 ( .A1(n6609), .A2(P1_B_REG_SCAN_IN), .ZN(n6412) );
  AND2_X1 U8140 ( .A1(n9299), .A2(n6412), .ZN(n9054) );
  INV_X1 U8141 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8142 ( .A1(n6094), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8143 ( .A1(n6413), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6414) );
  OAI211_X1 U8144 ( .C1(n5751), .C2(n6416), .A(n6415), .B(n6414), .ZN(n8933)
         );
  AOI22_X1 U8145 ( .A1(n8934), .A2(n9298), .B1(n9054), .B2(n8933), .ZN(n6417)
         );
  NAND2_X1 U8146 ( .A1(n6418), .A2(n6417), .ZN(n9063) );
  NOR2_X1 U8147 ( .A1(n9070), .A2(n9063), .ZN(n6419) );
  NAND2_X1 U8148 ( .A1(n6420), .A2(n6419), .ZN(n6433) );
  NAND2_X1 U8149 ( .A1(n6531), .A2(n6422), .ZN(n6423) );
  NAND2_X1 U8150 ( .A1(n9550), .A2(n6423), .ZN(n6425) );
  NAND2_X1 U8151 ( .A1(n6425), .A2(n6424), .ZN(n6817) );
  NAND2_X1 U8152 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  OR2_X1 U8153 ( .A1(n6433), .A2(n9605), .ZN(n6429) );
  NAND2_X1 U8154 ( .A1(n6429), .A2(n4836), .ZN(n6430) );
  NAND2_X1 U8155 ( .A1(n6430), .A2(n4843), .ZN(P1_U3551) );
  OR2_X1 U8156 ( .A1(n6433), .A2(n9589), .ZN(n6434) );
  NAND2_X1 U8157 ( .A1(n6434), .A2(n4835), .ZN(n6435) );
  NAND2_X1 U8158 ( .A1(n6435), .A2(n4847), .ZN(P1_U3519) );
  INV_X1 U8159 ( .A(n6493), .ZN(n6436) );
  NOR2_X2 U8160 ( .A1(n6437), .A2(n6436), .ZN(P2_U3893) );
  INV_X1 U8161 ( .A(n6437), .ZN(n6438) );
  NAND2_X1 U8162 ( .A1(n6438), .A2(n7422), .ZN(n6446) );
  NAND2_X1 U8163 ( .A1(n7422), .A2(n7865), .ZN(n6439) );
  NAND2_X1 U8164 ( .A1(n6446), .A2(n6439), .ZN(n6455) );
  OAI21_X1 U8165 ( .B1(n6455), .B2(n6440), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  NOR2_X1 U8166 ( .A1(n6441), .A2(P1_U3086), .ZN(n6442) );
  AND2_X2 U8167 ( .A1(n6532), .A2(n6442), .ZN(P1_U3973) );
  XNOR2_X1 U8168 ( .A(n6517), .B(n6525), .ZN(n6445) );
  INV_X1 U8169 ( .A(n6510), .ZN(n6479) );
  XOR2_X1 U8170 ( .A(n6510), .B(n6443), .Z(n6505) );
  INV_X1 U8171 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9832) );
  INV_X1 U8172 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U8173 ( .A1(n9609), .A2(n9614), .ZN(n6504) );
  NOR2_X1 U8174 ( .A1(n6505), .A2(n6504), .ZN(n6503) );
  AOI21_X1 U8175 ( .B1(n6443), .B2(n6479), .A(n6503), .ZN(n6444) );
  NAND2_X1 U8176 ( .A1(P2_U3893), .A2(n7928), .ZN(n9622) );
  NOR2_X1 U8177 ( .A1(n6444), .A2(n6445), .ZN(n6516) );
  AOI211_X1 U8178 ( .C1(n6445), .C2(n6444), .A(n9622), .B(n6516), .ZN(n6471)
         );
  INV_X1 U8179 ( .A(n6446), .ZN(n6450) );
  INV_X1 U8180 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7130) );
  NOR2_X1 U8181 ( .A1(n9664), .A2(n7130), .ZN(n6470) );
  NAND2_X1 U8182 ( .A1(n7928), .A2(n6447), .ZN(n6448) );
  OR2_X1 U8183 ( .A1(n6455), .A2(n6448), .ZN(n6452) );
  NOR2_X1 U8184 ( .A1(n7928), .A2(P2_U3151), .ZN(n6454) );
  NAND2_X1 U8185 ( .A1(n6450), .A2(n6454), .ZN(n6451) );
  NAND2_X1 U8186 ( .A1(n6452), .A2(n6451), .ZN(n9696) );
  INV_X1 U8187 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6453) );
  OAI22_X1 U8188 ( .A1(n9766), .A2(n6525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6453), .ZN(n6469) );
  INV_X1 U8189 ( .A(n6454), .ZN(n7678) );
  OR2_X1 U8190 ( .A1(n6455), .A2(n7678), .ZN(n6465) );
  NOR2_X2 U8191 ( .A1(n6465), .A2(n4433), .ZN(n9762) );
  INV_X1 U8192 ( .A(n9762), .ZN(n7292) );
  NAND2_X1 U8193 ( .A1(n9614), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6457) );
  INV_X1 U8194 ( .A(n5085), .ZN(n6459) );
  OAI21_X1 U8195 ( .B1(n9832), .B2(n6459), .A(n6479), .ZN(n6456) );
  OAI21_X1 U8196 ( .B1(n5085), .B2(n6457), .A(n6456), .ZN(n6507) );
  AOI22_X1 U8197 ( .A1(n6507), .A2(P2_REG1_REG_1__SCAN_IN), .B1(n5085), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n6523) );
  XOR2_X1 U8198 ( .A(n6522), .B(n6523), .Z(n6467) );
  INV_X1 U8199 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8200 ( .A1(n9614), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6462) );
  INV_X1 U8201 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6460) );
  OAI21_X1 U8202 ( .B1(n6460), .B2(n6459), .A(n6479), .ZN(n6461) );
  OAI21_X1 U8203 ( .B1(n5085), .B2(n6462), .A(n6461), .ZN(n6506) );
  AOI22_X1 U8204 ( .A1(n6506), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n5085), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6463) );
  AOI21_X1 U8205 ( .B1(n6464), .B2(n6463), .A(n6524), .ZN(n6466) );
  INV_X1 U8206 ( .A(n6465), .ZN(n9611) );
  NAND2_X1 U8207 ( .A1(n9611), .A2(n4433), .ZN(n9755) );
  OAI22_X1 U8208 ( .A1(n7292), .A2(n6467), .B1(n6466), .B2(n9755), .ZN(n6468)
         );
  OR4_X1 U8209 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(P2_U3184)
         );
  NOR2_X1 U8210 ( .A1(n7731), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9446) );
  AOI22_X1 U8211 ( .A1(n8971), .A2(P1_STATE_REG_SCAN_IN), .B1(n9446), .B2(
        P2_DATAO_REG_2__SCAN_IN), .ZN(n6472) );
  OAI21_X1 U8212 ( .B1(n6476), .B2(n7960), .A(n6472), .ZN(P1_U3353) );
  AOI22_X1 U8213 ( .A1(n8984), .A2(P1_STATE_REG_SCAN_IN), .B1(n9446), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6473) );
  OAI21_X1 U8214 ( .B1(n6475), .B2(n7960), .A(n6473), .ZN(P1_U3352) );
  INV_X1 U8215 ( .A(n9446), .ZN(n7964) );
  OAI222_X1 U8216 ( .A1(P1_U3086), .A2(n6561), .B1(n7960), .B2(n4481), .C1(
        n4484), .C2(n7964), .ZN(P1_U3354) );
  AND2_X1 U8217 ( .A1(n7731), .A2(P2_U3151), .ZN(n8487) );
  AND2_X1 U8218 ( .A1(n4266), .A2(P2_U3151), .ZN(n7677) );
  INV_X2 U8219 ( .A(n7677), .ZN(n8492) );
  OAI222_X1 U8220 ( .A1(n8494), .A2(n9974), .B1(n8492), .B2(n6475), .C1(
        P2_U3151), .C2(n6597), .ZN(P2_U3292) );
  OAI222_X1 U8221 ( .A1(n8494), .A2(n6477), .B1(n8492), .B2(n6476), .C1(
        P2_U3151), .C2(n6525), .ZN(P2_U3293) );
  OAI222_X1 U8222 ( .A1(n6479), .A2(P2_U3151), .B1(n8492), .B2(n4481), .C1(
        n6478), .C2(n8494), .ZN(P2_U3294) );
  INV_X1 U8223 ( .A(n6566), .ZN(n8994) );
  OAI222_X1 U8224 ( .A1(n7964), .A2(n6480), .B1(n7960), .B2(n6481), .C1(
        P1_U3086), .C2(n8994), .ZN(P1_U3351) );
  OAI222_X1 U8225 ( .A1(n8494), .A2(n6482), .B1(n8492), .B2(n6481), .C1(
        P2_U3151), .C2(n7270), .ZN(P2_U3291) );
  AOI22_X1 U8226 ( .A1(n9011), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9446), .ZN(n6483) );
  OAI21_X1 U8227 ( .B1(n6484), .B2(n7960), .A(n6483), .ZN(P1_U3350) );
  OAI222_X1 U8228 ( .A1(n8494), .A2(n6618), .B1(n8492), .B2(n6484), .C1(
        P2_U3151), .C2(n7242), .ZN(P2_U3290) );
  OAI222_X1 U8229 ( .A1(n8494), .A2(n6485), .B1(n8492), .B2(n6486), .C1(
        P2_U3151), .C2(n7275), .ZN(P2_U3289) );
  OAI222_X1 U8230 ( .A1(n7964), .A2(n6487), .B1(n7960), .B2(n6486), .C1(
        P1_U3086), .C2(n6570), .ZN(P1_U3349) );
  INV_X1 U8231 ( .A(n5469), .ZN(n6488) );
  INV_X1 U8232 ( .A(n6490), .ZN(n6491) );
  AOI22_X1 U8233 ( .A1(n6498), .A2(n6492), .B1(n6493), .B2(n6491), .ZN(
        P2_U3377) );
  AOI22_X1 U8234 ( .A1(n6498), .A2(n6494), .B1(n4852), .B2(n6493), .ZN(
        P2_U3376) );
  AND2_X1 U8235 ( .A1(n6498), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8236 ( .A1(n6498), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8237 ( .A1(n6498), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8238 ( .A1(n6498), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8239 ( .A1(n6498), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8240 ( .A1(n6498), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8241 ( .A1(n6498), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8242 ( .A1(n6498), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8243 ( .A1(n6498), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8244 ( .A1(n6498), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8245 ( .A1(n6498), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8246 ( .A1(n6498), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8247 ( .A1(n6498), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8248 ( .A1(n6498), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8249 ( .A1(n6498), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8250 ( .A1(n6498), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8251 ( .A1(n6498), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8252 ( .A1(n6498), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8253 ( .A1(n6498), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8254 ( .A1(n6498), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8255 ( .A1(n6498), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8256 ( .A1(n6498), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8257 ( .A1(n6498), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8258 ( .A1(n6498), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8259 ( .A(n6574), .ZN(n9466) );
  OAI222_X1 U8260 ( .A1(n7964), .A2(n6495), .B1(n7960), .B2(n6496), .C1(
        P1_U3086), .C2(n9466), .ZN(P1_U3348) );
  OAI222_X1 U8261 ( .A1(n8494), .A2(n6497), .B1(n8492), .B2(n6496), .C1(
        P2_U3151), .C2(n7265), .ZN(P2_U3288) );
  INV_X1 U8262 ( .A(n6498), .ZN(n6499) );
  INV_X1 U8263 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9894) );
  NOR2_X1 U8264 ( .A1(n6499), .A2(n9894), .ZN(P2_U3242) );
  INV_X1 U8265 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U8266 ( .A1(n6499), .A2(n9944), .ZN(P2_U3252) );
  INV_X1 U8267 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U8268 ( .A1(n6499), .A2(n9912), .ZN(P2_U3256) );
  INV_X1 U8269 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U8270 ( .A1(n6499), .A2(n9953), .ZN(P2_U3255) );
  INV_X1 U8271 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U8272 ( .A1(n6499), .A2(n9896), .ZN(P2_U3257) );
  INV_X1 U8273 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9973) );
  NOR2_X1 U8274 ( .A1(n6499), .A2(n9973), .ZN(P2_U3248) );
  INV_X1 U8275 ( .A(n6500), .ZN(n6502) );
  OAI222_X1 U8276 ( .A1(n8494), .A2(n6620), .B1(n8492), .B2(n6502), .C1(
        P2_U3151), .C2(n7263), .ZN(P2_U3287) );
  INV_X1 U8277 ( .A(n9480), .ZN(n6501) );
  OAI222_X1 U8278 ( .A1(n7964), .A2(n9991), .B1(n7960), .B2(n6502), .C1(
        P1_U3086), .C2(n6501), .ZN(P1_U3347) );
  AOI211_X1 U8279 ( .C1(n6505), .C2(n6504), .A(n9622), .B(n6503), .ZN(n6515)
         );
  INV_X1 U8280 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6513) );
  INV_X1 U8281 ( .A(n9755), .ZN(n9737) );
  XNOR2_X1 U8282 ( .A(n6506), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n6509) );
  XNOR2_X1 U8283 ( .A(n6507), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6508) );
  AOI22_X1 U8284 ( .A1(n9737), .A2(n6509), .B1(n9762), .B2(n6508), .ZN(n6512)
         );
  AOI22_X1 U8285 ( .A1(n9696), .A2(n6510), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n6511) );
  OAI211_X1 U8286 ( .C1(n6513), .C2(n9664), .A(n6512), .B(n6511), .ZN(n6514)
         );
  OR2_X1 U8287 ( .A1(n6515), .A2(n6514), .ZN(P2_U3183) );
  INV_X1 U8288 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7126) );
  AOI21_X1 U8289 ( .B1(n6517), .B2(n6525), .A(n6516), .ZN(n6519) );
  XOR2_X1 U8290 ( .A(n6597), .B(n6588), .Z(n6518) );
  NAND2_X1 U8291 ( .A1(n6519), .A2(n6518), .ZN(n6587) );
  OAI21_X1 U8292 ( .B1(n6519), .B2(n6518), .A(n6587), .ZN(n6520) );
  NAND2_X1 U8293 ( .A1(n6520), .A2(n9750), .ZN(n6530) );
  NOR2_X1 U8294 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5091), .ZN(n6645) );
  INV_X1 U8295 ( .A(n6525), .ZN(n6521) );
  INV_X1 U8296 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9834) );
  XOR2_X1 U8297 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6592), .Z(n6527) );
  XNOR2_X1 U8298 ( .A(n6595), .B(n6597), .ZN(n6598) );
  INV_X1 U8299 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U8300 ( .A(n6598), .B(n6723), .ZN(n6526) );
  OAI22_X1 U8301 ( .A1(n7292), .A2(n6527), .B1(n6526), .B2(n9755), .ZN(n6528)
         );
  AOI211_X1 U8302 ( .C1(n4475), .C2(n9696), .A(n6645), .B(n6528), .ZN(n6529)
         );
  OAI211_X1 U8303 ( .C1(n7126), .C2(n9664), .A(n6530), .B(n6529), .ZN(P2_U3185) );
  OR2_X1 U8304 ( .A1(n8915), .A2(n6531), .ZN(n6543) );
  NAND2_X1 U8305 ( .A1(n6532), .A2(n8905), .ZN(n6533) );
  NAND2_X1 U8306 ( .A1(n5835), .A2(n6533), .ZN(n6541) );
  INV_X1 U8307 ( .A(n9892), .ZN(n8997) );
  NOR2_X1 U8308 ( .A1(n8997), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8309 ( .A(n6534), .ZN(n6536) );
  INV_X1 U8310 ( .A(n6673), .ZN(n6583) );
  OAI222_X1 U8311 ( .A1(n7964), .A2(n6535), .B1(n7960), .B2(n6536), .C1(n6583), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U8312 ( .A1(n8494), .A2(n6622), .B1(n8492), .B2(n6536), .C1(n9695), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8313 ( .A(n6537), .ZN(n6539) );
  INV_X1 U8314 ( .A(n9458), .ZN(n6665) );
  OAI222_X1 U8315 ( .A1(n7964), .A2(n6538), .B1(n7960), .B2(n6539), .C1(n6665), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8316 ( .A(n9697), .ZN(n7259) );
  OAI222_X1 U8317 ( .A1(n8494), .A2(n6540), .B1(n8492), .B2(n6539), .C1(n7259), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8318 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8319 ( .A1(n6611), .A2(n8959), .ZN(n9522) );
  INV_X1 U8320 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9603) );
  AOI22_X1 U8321 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6673), .B1(n6583), .B2(
        n9603), .ZN(n6559) );
  XNOR2_X1 U8322 ( .A(n8971), .B(n6544), .ZN(n8977) );
  XNOR2_X1 U8323 ( .A(n6561), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n8952) );
  AND2_X1 U8324 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8951) );
  NAND2_X1 U8325 ( .A1(n8952), .A2(n8951), .ZN(n8950) );
  NAND2_X1 U8326 ( .A1(n8949), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8327 ( .A1(n8950), .A2(n6545), .ZN(n8976) );
  NAND2_X1 U8328 ( .A1(n8977), .A2(n8976), .ZN(n8975) );
  NAND2_X1 U8329 ( .A1(n8971), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8330 ( .A1(n8975), .A2(n6546), .ZN(n8989) );
  XNOR2_X1 U8331 ( .A(n8984), .B(n6547), .ZN(n8990) );
  NAND2_X1 U8332 ( .A1(n8989), .A2(n8990), .ZN(n8988) );
  NAND2_X1 U8333 ( .A1(n8984), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U8334 ( .A1(n8988), .A2(n6548), .ZN(n8999) );
  MUX2_X1 U8335 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5793), .S(n6566), .Z(n9000)
         );
  NAND2_X1 U8336 ( .A1(n8999), .A2(n9000), .ZN(n8998) );
  NAND2_X1 U8337 ( .A1(n6566), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8338 ( .A1(n8998), .A2(n6549), .ZN(n9016) );
  XNOR2_X1 U8339 ( .A(n9011), .B(n10019), .ZN(n9017) );
  NAND2_X1 U8340 ( .A1(n9016), .A2(n9017), .ZN(n9015) );
  NAND2_X1 U8341 ( .A1(n9011), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8342 ( .A1(n9015), .A2(n6550), .ZN(n9029) );
  XNOR2_X1 U8343 ( .A(n6570), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U8344 ( .A1(n9029), .A2(n9030), .ZN(n9028) );
  INV_X1 U8345 ( .A(n6570), .ZN(n9024) );
  NAND2_X1 U8346 ( .A1(n9024), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6551) );
  AND2_X1 U8347 ( .A1(n9028), .A2(n6551), .ZN(n9463) );
  INV_X1 U8348 ( .A(n9463), .ZN(n6554) );
  OR2_X1 U8349 ( .A1(n6574), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8350 ( .A1(n6574), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U8351 ( .A1(n6552), .A2(n6555), .ZN(n9462) );
  INV_X1 U8352 ( .A(n9462), .ZN(n6553) );
  NAND2_X1 U8353 ( .A1(n6554), .A2(n6553), .ZN(n9470) );
  AND2_X1 U8354 ( .A1(n9470), .A2(n6555), .ZN(n9476) );
  OR2_X1 U8355 ( .A1(n9480), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U8356 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9480), .ZN(n6556) );
  NAND2_X1 U8357 ( .A1(n6557), .A2(n6556), .ZN(n9475) );
  NOR2_X1 U8358 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  AOI21_X1 U8359 ( .B1(n9480), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9477), .ZN(
        n6558) );
  NAND2_X1 U8360 ( .A1(n6559), .A2(n6558), .ZN(n6672) );
  OAI21_X1 U8361 ( .B1(n6559), .B2(n6558), .A(n6672), .ZN(n6585) );
  NAND2_X1 U8362 ( .A1(n6611), .A2(n6280), .ZN(n9502) );
  NOR2_X1 U8363 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6673), .ZN(n6560) );
  AOI21_X1 U8364 ( .B1(n6673), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6560), .ZN(
        n6577) );
  XNOR2_X1 U8365 ( .A(n8971), .B(n6892), .ZN(n8974) );
  XNOR2_X1 U8366 ( .A(n6561), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U8367 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n8962) );
  INV_X1 U8368 ( .A(n8962), .ZN(n8954) );
  NAND2_X1 U8369 ( .A1(n8955), .A2(n8954), .ZN(n8953) );
  NAND2_X1 U8370 ( .A1(n8949), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8371 ( .A1(n8953), .A2(n6562), .ZN(n8973) );
  NAND2_X1 U8372 ( .A1(n8974), .A2(n8973), .ZN(n8972) );
  NAND2_X1 U8373 ( .A1(n8971), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8374 ( .A1(n8972), .A2(n6563), .ZN(n8986) );
  XNOR2_X1 U8375 ( .A(n8984), .B(n6564), .ZN(n8987) );
  NAND2_X1 U8376 ( .A1(n8986), .A2(n8987), .ZN(n8985) );
  NAND2_X1 U8377 ( .A1(n8984), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8378 ( .A1(n8985), .A2(n6565), .ZN(n9002) );
  MUX2_X1 U8379 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6951), .S(n6566), .Z(n9003)
         );
  NAND2_X1 U8380 ( .A1(n9002), .A2(n9003), .ZN(n9001) );
  NAND2_X1 U8381 ( .A1(n6566), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8382 ( .A1(n9001), .A2(n6567), .ZN(n9013) );
  XNOR2_X1 U8383 ( .A(n9011), .B(n6568), .ZN(n9014) );
  NAND2_X1 U8384 ( .A1(n9013), .A2(n9014), .ZN(n9012) );
  NAND2_X1 U8385 ( .A1(n9011), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8386 ( .A1(n9012), .A2(n6569), .ZN(n9026) );
  XNOR2_X1 U8387 ( .A(n6570), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U8388 ( .A1(n9026), .A2(n9027), .ZN(n9025) );
  NAND2_X1 U8389 ( .A1(n9024), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8390 ( .A1(n9025), .A2(n6571), .ZN(n9464) );
  OR2_X1 U8391 ( .A1(n6574), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8392 ( .A1(n6574), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6572) );
  AND2_X1 U8393 ( .A1(n6573), .A2(n6572), .ZN(n9465) );
  AND2_X1 U8394 ( .A1(n9464), .A2(n9465), .ZN(n9467) );
  AOI21_X1 U8395 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6574), .A(n9467), .ZN(
        n9482) );
  NAND2_X1 U8396 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9480), .ZN(n6575) );
  OAI21_X1 U8397 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9480), .A(n6575), .ZN(
        n9483) );
  NOR2_X1 U8398 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  AOI21_X1 U8399 ( .B1(n9480), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9481), .ZN(
        n6576) );
  NAND2_X1 U8400 ( .A1(n6577), .A2(n6576), .ZN(n6666) );
  OAI21_X1 U8401 ( .B1(n6577), .B2(n6576), .A(n6666), .ZN(n6579) );
  NAND2_X1 U8402 ( .A1(n8960), .A2(n6609), .ZN(n8963) );
  INV_X1 U8403 ( .A(n8963), .ZN(n6578) );
  NAND2_X1 U8404 ( .A1(n6579), .A2(n9885), .ZN(n6582) );
  NOR2_X1 U8405 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6580), .ZN(n7329) );
  AOI21_X1 U8406 ( .B1(n8997), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7329), .ZN(
        n6581) );
  OAI211_X1 U8407 ( .C1(n9502), .C2(n6583), .A(n6582), .B(n6581), .ZN(n6584)
         );
  AOI21_X1 U8408 ( .B1(n9879), .B2(n6585), .A(n6584), .ZN(n6586) );
  INV_X1 U8409 ( .A(n6586), .ZN(P1_U3252) );
  INV_X1 U8410 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9959) );
  XNOR2_X1 U8411 ( .A(n7271), .B(n7270), .ZN(n6590) );
  OAI21_X1 U8412 ( .B1(n6588), .B2(n6597), .A(n6587), .ZN(n6589) );
  NOR2_X1 U8413 ( .A1(n6589), .A2(n6590), .ZN(n7269) );
  AOI211_X1 U8414 ( .C1(n6590), .C2(n6589), .A(n9622), .B(n7269), .ZN(n6591)
         );
  INV_X1 U8415 ( .A(n6591), .ZN(n6605) );
  INV_X1 U8416 ( .A(n7270), .ZN(n7241) );
  AND2_X1 U8417 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6689) );
  INV_X1 U8418 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9951) );
  MUX2_X1 U8419 ( .A(n9951), .B(P2_REG1_REG_4__SCAN_IN), .S(n7270), .Z(n6594)
         );
  NOR2_X1 U8420 ( .A1(n6593), .A2(n6594), .ZN(n7224) );
  AOI21_X1 U8421 ( .B1(n6594), .B2(n6593), .A(n7224), .ZN(n6602) );
  INV_X1 U8422 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7240) );
  MUX2_X1 U8423 ( .A(n7240), .B(P2_REG2_REG_4__SCAN_IN), .S(n7270), .Z(n6600)
         );
  INV_X1 U8424 ( .A(n6595), .ZN(n6596) );
  AOI22_X1 U8425 ( .A1(n6598), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n6597), .B2(
        n6596), .ZN(n6599) );
  AOI21_X1 U8426 ( .B1(n6600), .B2(n6599), .A(n7239), .ZN(n6601) );
  OAI22_X1 U8427 ( .A1(n7292), .A2(n6602), .B1(n6601), .B2(n9755), .ZN(n6603)
         );
  AOI211_X1 U8428 ( .C1(n7241), .C2(n9696), .A(n6689), .B(n6603), .ZN(n6604)
         );
  OAI211_X1 U8429 ( .C1(n9959), .C2(n9664), .A(n6605), .B(n6604), .ZN(P2_U3186) );
  INV_X1 U8430 ( .A(n6606), .ZN(n6607) );
  INV_X1 U8431 ( .A(n6675), .ZN(n9501) );
  OAI222_X1 U8432 ( .A1(n7964), .A2(n9945), .B1(n7960), .B2(n6607), .C1(
        P1_U3086), .C2(n9501), .ZN(P1_U3344) );
  OAI222_X1 U8433 ( .A1(n8494), .A2(n6624), .B1(n8492), .B2(n6607), .C1(
        P2_U3151), .C2(n9726), .ZN(P2_U3284) );
  NOR2_X1 U8434 ( .A1(n8959), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6608) );
  NOR2_X1 U8435 ( .A1(n6608), .A2(n6280), .ZN(n8967) );
  OAI21_X1 U8436 ( .B1(n6609), .B2(P1_REG1_REG_0__SCAN_IN), .A(n8967), .ZN(
        n6610) );
  MUX2_X1 U8437 ( .A(n6610), .B(n8967), .S(P1_IR_REG_0__SCAN_IN), .Z(n6617) );
  INV_X1 U8438 ( .A(n6611), .ZN(n6616) );
  NAND3_X1 U8439 ( .A1(n9879), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5723), .ZN(
        n6615) );
  INV_X1 U8440 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6612) );
  OAI22_X1 U8441 ( .A1(n9892), .A2(n6612), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6928), .ZN(n6613) );
  INV_X1 U8442 ( .A(n6613), .ZN(n6614) );
  OAI211_X1 U8443 ( .C1(n6617), .C2(n6616), .A(n6615), .B(n6614), .ZN(P1_U3243) );
  MUX2_X1 U8444 ( .A(n6618), .B(n6959), .S(P1_U3973), .Z(n6619) );
  INV_X1 U8445 ( .A(n6619), .ZN(P1_U3559) );
  MUX2_X1 U8446 ( .A(n6620), .B(n7331), .S(P1_U3973), .Z(n6621) );
  INV_X1 U8447 ( .A(n6621), .ZN(P1_U3562) );
  MUX2_X1 U8448 ( .A(n6622), .B(n7401), .S(P1_U3973), .Z(n6623) );
  INV_X1 U8449 ( .A(n6623), .ZN(P1_U3563) );
  MUX2_X1 U8450 ( .A(n6624), .B(n7632), .S(P1_U3973), .Z(n6625) );
  INV_X1 U8451 ( .A(n6625), .ZN(P1_U3565) );
  INV_X1 U8452 ( .A(n6626), .ZN(n6628) );
  INV_X1 U8453 ( .A(n7365), .ZN(n6679) );
  OAI222_X1 U8454 ( .A1(n7964), .A2(n6627), .B1(n7960), .B2(n6628), .C1(n6679), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8455 ( .A(n7548), .ZN(n7558) );
  OAI222_X1 U8456 ( .A1(n8494), .A2(n9963), .B1(n8492), .B2(n6628), .C1(n7558), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  NAND2_X1 U8457 ( .A1(n6629), .A2(n6632), .ZN(n6630) );
  OAI211_X1 U8458 ( .C1(n5534), .C2(n6632), .A(n6631), .B(n6630), .ZN(n6636)
         );
  INV_X1 U8459 ( .A(n6636), .ZN(n6633) );
  INV_X1 U8460 ( .A(n8276), .ZN(n8269) );
  NAND2_X1 U8461 ( .A1(n6633), .A2(n8269), .ZN(n8330) );
  NAND2_X1 U8462 ( .A1(n8149), .A2(n6640), .ZN(n7746) );
  NAND2_X1 U8463 ( .A1(n6634), .A2(n7746), .ZN(n7883) );
  INV_X1 U8464 ( .A(n7883), .ZN(n9767) );
  NOR3_X1 U8465 ( .A1(n9767), .A2(n9828), .A3(n6635), .ZN(n6637) );
  NOR2_X1 U8466 ( .A1(n7703), .A2(n8300), .ZN(n9770) );
  OAI21_X1 U8467 ( .B1(n6637), .B2(n9770), .A(n8366), .ZN(n6639) );
  INV_X2 U8468 ( .A(n7996), .ZN(n8368) );
  AOI22_X1 U8469 ( .A1(n8336), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n8368), .ZN(n6638) );
  OAI211_X1 U8470 ( .C1(n8330), .C2(n6640), .A(n6639), .B(n6638), .ZN(P2_U3233) );
  INV_X1 U8471 ( .A(n8124), .ZN(n8010) );
  OAI211_X1 U8472 ( .C1(n6643), .C2(n6642), .A(n6641), .B(n8117), .ZN(n6647)
         );
  INV_X1 U8473 ( .A(n8119), .ZN(n8109) );
  OAI22_X1 U8474 ( .A1(n8109), .A2(n6703), .B1(n6759), .B2(n8121), .ZN(n6644)
         );
  AOI211_X1 U8475 ( .C1(n6724), .C2(n8072), .A(n6645), .B(n6644), .ZN(n6646)
         );
  OAI211_X1 U8476 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8010), .A(n6647), .B(
        n6646), .ZN(P2_U3158) );
  INV_X1 U8477 ( .A(n8603), .ZN(n8643) );
  AOI22_X1 U8478 ( .A1(n8641), .A2(n9556), .B1(n8627), .B2(n5743), .ZN(n6651)
         );
  NAND2_X1 U8479 ( .A1(n8635), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7945) );
  NAND2_X1 U8480 ( .A1(n7945), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6650) );
  OAI211_X1 U8481 ( .C1(n8961), .C2(n8643), .A(n6651), .B(n6650), .ZN(P1_U3232) );
  INV_X1 U8482 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6653) );
  INV_X1 U8483 ( .A(n6652), .ZN(n6654) );
  OAI222_X1 U8484 ( .A1(n7964), .A2(n6653), .B1(n7960), .B2(n6654), .C1(
        P1_U3086), .C2(n7358), .ZN(P1_U3342) );
  INV_X1 U8485 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9981) );
  OAI222_X1 U8486 ( .A1(n8494), .A2(n9981), .B1(n8492), .B2(n6654), .C1(
        P2_U3151), .C2(n9741), .ZN(P2_U3282) );
  OAI21_X1 U8487 ( .B1(n7744), .B2(n4267), .A(n6655), .ZN(n8417) );
  INV_X1 U8488 ( .A(n8417), .ZN(n6663) );
  OR2_X1 U8489 ( .A1(n7743), .A2(n7174), .ZN(n6709) );
  NOR2_X1 U8490 ( .A1(n8336), .A2(n6709), .ZN(n8001) );
  INV_X1 U8491 ( .A(n8001), .ZN(n7038) );
  INV_X1 U8492 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6660) );
  INV_X1 U8493 ( .A(n7031), .ZN(n6975) );
  OAI22_X1 U8494 ( .A1(n6703), .A2(n8300), .B1(n4636), .B2(n8302), .ZN(n6659)
         );
  XNOR2_X1 U8495 ( .A(n7744), .B(n6656), .ZN(n6657) );
  NOR2_X1 U8496 ( .A1(n6657), .A2(n9768), .ZN(n6658) );
  AOI211_X1 U8497 ( .C1(n6975), .C2(n8417), .A(n6659), .B(n6658), .ZN(n8419)
         );
  MUX2_X1 U8498 ( .A(n6660), .B(n8419), .S(n8366), .Z(n6662) );
  AOI22_X1 U8499 ( .A1(n8369), .A2(n5536), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8368), .ZN(n6661) );
  OAI211_X1 U8500 ( .C1(n6663), .C2(n7038), .A(n6662), .B(n6661), .ZN(P2_U3232) );
  NOR2_X1 U8501 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7365), .ZN(n6664) );
  AOI21_X1 U8502 ( .B1(n7365), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6664), .ZN(
        n6669) );
  AOI22_X1 U8503 ( .A1(n9458), .A2(n5927), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6665), .ZN(n9454) );
  OAI21_X1 U8504 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6673), .A(n6666), .ZN(
        n9455) );
  NOR2_X1 U8505 ( .A1(n9454), .A2(n9455), .ZN(n9453) );
  AOI21_X1 U8506 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9458), .A(n9453), .ZN(
        n9494) );
  NAND2_X1 U8507 ( .A1(n6675), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U8508 ( .B1(n6675), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6667), .ZN(
        n9495) );
  NOR2_X1 U8509 ( .A1(n9494), .A2(n9495), .ZN(n9496) );
  AOI21_X1 U8510 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6675), .A(n9496), .ZN(
        n6668) );
  NAND2_X1 U8511 ( .A1(n6669), .A2(n6668), .ZN(n7364) );
  OAI21_X1 U8512 ( .B1(n6669), .B2(n6668), .A(n7364), .ZN(n6670) );
  NAND2_X1 U8513 ( .A1(n6670), .A2(n9885), .ZN(n6683) );
  INV_X1 U8514 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6671) );
  MUX2_X1 U8515 ( .A(n6671), .B(P1_REG1_REG_10__SCAN_IN), .S(n9458), .Z(n9451)
         );
  OAI21_X1 U8516 ( .B1(n6673), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6672), .ZN(
        n9452) );
  NOR2_X1 U8517 ( .A1(n9451), .A2(n9452), .ZN(n9450) );
  AOI21_X1 U8518 ( .B1(n9458), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9450), .ZN(
        n9491) );
  MUX2_X1 U8519 ( .A(n6674), .B(P1_REG1_REG_11__SCAN_IN), .S(n6675), .Z(n9492)
         );
  NOR2_X1 U8520 ( .A1(n9491), .A2(n9492), .ZN(n9490) );
  AOI21_X1 U8521 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6675), .A(n9490), .ZN(
        n6677) );
  AOI22_X1 U8522 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7365), .B1(n6679), .B2(
        n5967), .ZN(n6676) );
  NAND2_X1 U8523 ( .A1(n6677), .A2(n6676), .ZN(n7355) );
  OAI21_X1 U8524 ( .B1(n6677), .B2(n6676), .A(n7355), .ZN(n6681) );
  NAND2_X1 U8525 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U8526 ( .A1(n8997), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6678) );
  OAI211_X1 U8527 ( .C1(n9502), .C2(n6679), .A(n7631), .B(n6678), .ZN(n6680)
         );
  AOI21_X1 U8528 ( .B1(n6681), .B2(n9879), .A(n6680), .ZN(n6682) );
  NAND2_X1 U8529 ( .A1(n6683), .A2(n6682), .ZN(P1_U3255) );
  AOI21_X1 U8530 ( .B1(n6686), .B2(n6685), .A(n6684), .ZN(n6692) );
  OAI22_X1 U8531 ( .A1(n8109), .A2(n6732), .B1(n6687), .B2(n8121), .ZN(n6688)
         );
  AOI211_X1 U8532 ( .C1(n6715), .C2(n8072), .A(n6689), .B(n6688), .ZN(n6691)
         );
  NAND2_X1 U8533 ( .A1(n8124), .A2(n6714), .ZN(n6690) );
  OAI211_X1 U8534 ( .C1(n6692), .C2(n8052), .A(n6691), .B(n6690), .ZN(P2_U3170) );
  XOR2_X1 U8535 ( .A(n6694), .B(n6693), .Z(n6699) );
  NAND2_X1 U8536 ( .A1(n8010), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7700) );
  AOI22_X1 U8537 ( .A1(n8119), .A2(n8148), .B1(n6695), .B2(n8072), .ZN(n6696)
         );
  OAI21_X1 U8538 ( .B1(n6732), .B2(n8121), .A(n6696), .ZN(n6697) );
  AOI21_X1 U8539 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7700), .A(n6697), .ZN(
        n6698) );
  OAI21_X1 U8540 ( .B1(n6699), .B2(n8052), .A(n6698), .ZN(P2_U3177) );
  XOR2_X1 U8541 ( .A(n6701), .B(n6700), .Z(n6706) );
  AOI22_X1 U8542 ( .A1(n8119), .A2(n8149), .B1(n5536), .B2(n8072), .ZN(n6702)
         );
  OAI21_X1 U8543 ( .B1(n6703), .B2(n8121), .A(n6702), .ZN(n6704) );
  AOI21_X1 U8544 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7700), .A(n6704), .ZN(
        n6705) );
  OAI21_X1 U8545 ( .B1(n6706), .B2(n8052), .A(n6705), .ZN(P2_U3162) );
  INV_X1 U8546 ( .A(n6707), .ZN(n6727) );
  AOI22_X1 U8547 ( .A1(n9532), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9446), .ZN(n6708) );
  OAI21_X1 U8548 ( .B1(n6727), .B2(n7960), .A(n6708), .ZN(P1_U3341) );
  NAND2_X1 U8549 ( .A1(n7031), .A2(n6709), .ZN(n6710) );
  NAND2_X1 U8550 ( .A1(n7756), .A2(n7761), .ZN(n7882) );
  XNOR2_X1 U8551 ( .A(n6711), .B(n7882), .ZN(n9784) );
  XNOR2_X1 U8552 ( .A(n6712), .B(n7882), .ZN(n6713) );
  AOI222_X1 U8553 ( .A1(n8365), .A2(n6713), .B1(n8146), .B2(n8360), .C1(n8144), 
        .C2(n8362), .ZN(n9783) );
  MUX2_X1 U8554 ( .A(n7240), .B(n9783), .S(n8366), .Z(n6717) );
  AOI22_X1 U8555 ( .A1(n8369), .A2(n6715), .B1(n8368), .B2(n6714), .ZN(n6716)
         );
  OAI211_X1 U8556 ( .C1(n8372), .C2(n9784), .A(n6717), .B(n6716), .ZN(P2_U3229) );
  XNOR2_X1 U8557 ( .A(n6718), .B(n7880), .ZN(n9779) );
  NAND2_X1 U8558 ( .A1(n6720), .A2(n6719), .ZN(n6721) );
  XNOR2_X1 U8559 ( .A(n6721), .B(n7880), .ZN(n6722) );
  AOI222_X1 U8560 ( .A1(n8365), .A2(n6722), .B1(n8145), .B2(n8362), .C1(n8147), 
        .C2(n8360), .ZN(n9777) );
  MUX2_X1 U8561 ( .A(n6723), .B(n9777), .S(n8366), .Z(n6726) );
  AOI22_X1 U8562 ( .A1(n8369), .A2(n6724), .B1(n5091), .B2(n8368), .ZN(n6725)
         );
  OAI211_X1 U8563 ( .C1(n8372), .C2(n9779), .A(n6726), .B(n6725), .ZN(P2_U3230) );
  INV_X1 U8564 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6728) );
  INV_X1 U8565 ( .A(n9754), .ZN(n9765) );
  OAI222_X1 U8566 ( .A1(n8494), .A2(n6728), .B1(n8492), .B2(n6727), .C1(
        P2_U3151), .C2(n9765), .ZN(P2_U3281) );
  XNOR2_X1 U8567 ( .A(n6729), .B(n6731), .ZN(n9774) );
  NOR2_X1 U8568 ( .A1(n9773), .A2(n8276), .ZN(n6736) );
  XNOR2_X1 U8569 ( .A(n6730), .B(n6731), .ZN(n6734) );
  OAI22_X1 U8570 ( .A1(n7703), .A2(n8302), .B1(n6732), .B2(n8300), .ZN(n6733)
         );
  AOI21_X1 U8571 ( .B1(n6734), .B2(n8365), .A(n6733), .ZN(n6735) );
  OAI21_X1 U8572 ( .B1(n9774), .B2(n7031), .A(n6735), .ZN(n9776) );
  AOI211_X1 U8573 ( .C1(n8368), .C2(P2_REG3_REG_2__SCAN_IN), .A(n6736), .B(
        n9776), .ZN(n6737) );
  MUX2_X1 U8574 ( .A(n6458), .B(n6737), .S(n8366), .Z(n6738) );
  OAI21_X1 U8575 ( .B1(n9774), .B2(n7038), .A(n6738), .ZN(P2_U3231) );
  XOR2_X1 U8576 ( .A(n6739), .B(n6740), .Z(n6744) );
  INV_X1 U8577 ( .A(n8624), .ZN(n8636) );
  AOI22_X1 U8578 ( .A1(n8946), .A2(n8627), .B1(n8636), .B2(n5743), .ZN(n6741)
         );
  OAI21_X1 U8579 ( .B1(n9560), .B2(n8610), .A(n6741), .ZN(n6742) );
  AOI21_X1 U8580 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7945), .A(n6742), .ZN(
        n6743) );
  OAI21_X1 U8581 ( .B1(n6744), .B2(n8643), .A(n6743), .ZN(P1_U3237) );
  INV_X1 U8582 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6746) );
  INV_X1 U8583 ( .A(n6745), .ZN(n6747) );
  INV_X1 U8584 ( .A(n8151), .ZN(n8166) );
  OAI222_X1 U8585 ( .A1(n8494), .A2(n6746), .B1(n8492), .B2(n6747), .C1(
        P2_U3151), .C2(n8166), .ZN(P2_U3280) );
  INV_X1 U8586 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6748) );
  OAI222_X1 U8587 ( .A1(n7964), .A2(n6748), .B1(n7960), .B2(n6747), .C1(
        P1_U3086), .C2(n7367), .ZN(P1_U3340) );
  NAND2_X1 U8588 ( .A1(n6750), .A2(n6749), .ZN(n7884) );
  XOR2_X1 U8589 ( .A(n6751), .B(n7884), .Z(n9789) );
  INV_X1 U8590 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7268) );
  XNOR2_X1 U8591 ( .A(n6752), .B(n7884), .ZN(n6754) );
  OAI22_X1 U8592 ( .A1(n6759), .A2(n8302), .B1(n6874), .B2(n8300), .ZN(n6753)
         );
  AOI21_X1 U8593 ( .B1(n6754), .B2(n8365), .A(n6753), .ZN(n9790) );
  MUX2_X1 U8594 ( .A(n7268), .B(n9790), .S(n8366), .Z(n6756) );
  AOI22_X1 U8595 ( .A1(n8369), .A2(n6761), .B1(n8368), .B2(n6762), .ZN(n6755)
         );
  OAI211_X1 U8596 ( .C1(n9789), .C2(n8372), .A(n6756), .B(n6755), .ZN(P2_U3228) );
  XOR2_X1 U8597 ( .A(n6758), .B(n6757), .Z(n6765) );
  AND2_X1 U8598 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9626) );
  OAI22_X1 U8599 ( .A1(n8109), .A2(n6759), .B1(n6874), .B2(n8121), .ZN(n6760)
         );
  AOI211_X1 U8600 ( .C1(n6761), .C2(n8072), .A(n9626), .B(n6760), .ZN(n6764)
         );
  NAND2_X1 U8601 ( .A1(n8124), .A2(n6762), .ZN(n6763) );
  OAI211_X1 U8602 ( .C1(n6765), .C2(n8052), .A(n6764), .B(n6763), .ZN(P2_U3167) );
  INV_X1 U8603 ( .A(n6766), .ZN(n7766) );
  NAND2_X1 U8604 ( .A1(n7766), .A2(n7760), .ZN(n7888) );
  XOR2_X1 U8605 ( .A(n7888), .B(n6767), .Z(n9795) );
  INV_X1 U8606 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7238) );
  INV_X1 U8607 ( .A(n6768), .ZN(n6797) );
  OAI22_X1 U8608 ( .A1(n8366), .A2(n7238), .B1(n6797), .B2(n7996), .ZN(n6769)
         );
  AOI21_X1 U8609 ( .B1(n8369), .B2(n6770), .A(n6769), .ZN(n6777) );
  INV_X1 U8610 ( .A(n7888), .ZN(n6771) );
  XNOR2_X1 U8611 ( .A(n6772), .B(n6771), .ZN(n6773) );
  NAND2_X1 U8612 ( .A1(n6773), .A2(n8365), .ZN(n6775) );
  AOI22_X1 U8613 ( .A1(n8144), .A2(n8360), .B1(n8362), .B2(n8142), .ZN(n6774)
         );
  NAND2_X1 U8614 ( .A1(n6775), .A2(n6774), .ZN(n9796) );
  NAND2_X1 U8615 ( .A1(n9796), .A2(n8366), .ZN(n6776) );
  OAI211_X1 U8616 ( .C1(n9795), .C2(n8372), .A(n6777), .B(n6776), .ZN(P2_U3227) );
  XOR2_X1 U8617 ( .A(n6778), .B(n6779), .Z(n6785) );
  NOR2_X1 U8618 ( .A1(n8635), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6783) );
  INV_X1 U8619 ( .A(n8627), .ZN(n8638) );
  NAND2_X1 U8620 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8981) );
  INV_X1 U8621 ( .A(n8981), .ZN(n6780) );
  AOI21_X1 U8622 ( .B1(n5757), .B2(n8636), .A(n6780), .ZN(n6781) );
  OAI21_X1 U8623 ( .B1(n8663), .B2(n8638), .A(n6781), .ZN(n6782) );
  AOI211_X1 U8624 ( .C1(n6854), .C2(n8641), .A(n6783), .B(n6782), .ZN(n6784)
         );
  OAI21_X1 U8625 ( .B1(n6785), .B2(n8643), .A(n6784), .ZN(P1_U3218) );
  INV_X1 U8626 ( .A(n6786), .ZN(n6789) );
  OAI222_X1 U8627 ( .A1(n8494), .A2(n6787), .B1(n8492), .B2(n6789), .C1(n8178), 
        .C2(P2_U3151), .ZN(P2_U3279) );
  OAI222_X1 U8628 ( .A1(P1_U3086), .A2(n7369), .B1(n7960), .B2(n6789), .C1(
        n6788), .C2(n7964), .ZN(P1_U3339) );
  INV_X1 U8629 ( .A(n6790), .ZN(n6791) );
  INV_X1 U8630 ( .A(n7440), .ZN(n7374) );
  OAI222_X1 U8631 ( .A1(n7964), .A2(n9948), .B1(n7960), .B2(n6791), .C1(
        P1_U3086), .C2(n7374), .ZN(P1_U3338) );
  INV_X1 U8632 ( .A(n8210), .ZN(n8204) );
  OAI222_X1 U8633 ( .A1(n8494), .A2(n6792), .B1(n8492), .B2(n6791), .C1(
        P2_U3151), .C2(n8204), .ZN(P2_U3278) );
  AOI211_X1 U8634 ( .C1(n6795), .C2(n6794), .A(n8052), .B(n6793), .ZN(n6800)
         );
  NAND2_X1 U8635 ( .A1(n8119), .A2(n8144), .ZN(n6796) );
  NAND2_X1 U8636 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n9645) );
  OAI211_X1 U8637 ( .C1(n8121), .C2(n5548), .A(n6796), .B(n9645), .ZN(n6799)
         );
  OAI22_X1 U8638 ( .A1(n8010), .A2(n6797), .B1(n8128), .B2(n9794), .ZN(n6798)
         );
  OR3_X1 U8639 ( .A1(n6800), .A2(n6799), .A3(n6798), .ZN(P2_U3179) );
  AOI21_X1 U8640 ( .B1(n6801), .B2(n6802), .A(n8643), .ZN(n6804) );
  NAND2_X1 U8641 ( .A1(n6804), .A2(n6803), .ZN(n6809) );
  NOR2_X1 U8642 ( .A1(n6886), .A2(n8624), .ZN(n6807) );
  AND2_X1 U8643 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n8996) );
  INV_X1 U8644 ( .A(n8996), .ZN(n6805) );
  OAI21_X1 U8645 ( .B1(n6959), .B2(n8638), .A(n6805), .ZN(n6806) );
  AOI211_X1 U8646 ( .C1(n9566), .C2(n8641), .A(n6807), .B(n6806), .ZN(n6808)
         );
  OAI211_X1 U8647 ( .C1(n8635), .C2(n6953), .A(n6809), .B(n6808), .ZN(P1_U3230) );
  INV_X1 U8648 ( .A(n6810), .ZN(n6871) );
  AOI22_X1 U8649 ( .A1(n7443), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9446), .ZN(n6811) );
  OAI21_X1 U8650 ( .B1(n6871), .B2(n7960), .A(n6811), .ZN(P1_U3337) );
  OAI21_X1 U8651 ( .B1(n6397), .B2(n6813), .A(n6812), .ZN(n6864) );
  INV_X1 U8652 ( .A(n6864), .ZN(n6834) );
  NAND2_X1 U8653 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  INV_X1 U8654 ( .A(n6818), .ZN(n6819) );
  NAND2_X1 U8655 ( .A1(n9287), .A2(n6819), .ZN(n6900) );
  OAI21_X1 U8656 ( .B1(n6821), .B2(n6924), .A(n6820), .ZN(n6824) );
  INV_X1 U8657 ( .A(n6351), .ZN(n7950) );
  OAI22_X1 U8658 ( .A1(n7950), .A2(n9261), .B1(n6822), .B2(n9263), .ZN(n6823)
         );
  AOI21_X1 U8659 ( .B1(n6824), .B2(n9295), .A(n6823), .ZN(n6825) );
  OAI21_X1 U8660 ( .B1(n6834), .B2(n6848), .A(n6825), .ZN(n6862) );
  NAND2_X1 U8661 ( .A1(n6862), .A2(n9287), .ZN(n6833) );
  AOI211_X1 U8662 ( .C1(n9556), .C2(n7952), .A(n9306), .B(n6894), .ZN(n6863)
         );
  INV_X1 U8663 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6827) );
  OAI22_X1 U8664 ( .A1(n9287), .A2(n6827), .B1(n8947), .B2(n9309), .ZN(n6831)
         );
  INV_X1 U8665 ( .A(n6828), .ZN(n6829) );
  NAND2_X2 U8666 ( .A1(n9287), .A2(n6829), .ZN(n9542) );
  NOR2_X1 U8667 ( .A1(n9542), .A2(n5744), .ZN(n6830) );
  AOI211_X1 U8668 ( .C1(n6863), .C2(n4265), .A(n6831), .B(n6830), .ZN(n6832)
         );
  OAI211_X1 U8669 ( .C1(n6834), .C2(n6900), .A(n6833), .B(n6832), .ZN(P1_U3292) );
  OAI21_X1 U8670 ( .B1(n4354), .B2(n6836), .A(n6835), .ZN(n6842) );
  AND2_X1 U8671 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9659) );
  AOI21_X1 U8672 ( .B1(n8119), .B2(n8143), .A(n9659), .ZN(n6840) );
  NAND2_X1 U8673 ( .A1(n8072), .A2(n6881), .ZN(n6839) );
  NAND2_X1 U8674 ( .A1(n8124), .A2(n6877), .ZN(n6838) );
  OR2_X1 U8675 ( .A1(n8121), .A2(n6978), .ZN(n6837) );
  NAND4_X1 U8676 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n6841)
         );
  AOI21_X1 U8677 ( .B1(n6842), .B2(n8117), .A(n6841), .ZN(n6843) );
  INV_X1 U8678 ( .A(n6843), .ZN(P2_U3153) );
  INV_X1 U8679 ( .A(n8828), .ZN(n6846) );
  INV_X1 U8680 ( .A(n6844), .ZN(n6845) );
  AOI21_X1 U8681 ( .B1(n6852), .B2(n6846), .A(n6845), .ZN(n6847) );
  OAI222_X1 U8682 ( .A1(n9263), .A2(n8663), .B1(n9261), .B2(n6822), .C1(n9553), 
        .C2(n6847), .ZN(n6935) );
  INV_X1 U8683 ( .A(n6935), .ZN(n6860) );
  INV_X2 U8684 ( .A(n9287), .ZN(n9317) );
  INV_X1 U8685 ( .A(n6848), .ZN(n6889) );
  NAND2_X1 U8686 ( .A1(n9287), .A2(n6889), .ZN(n6849) );
  OAI21_X1 U8687 ( .B1(n6850), .B2(n6852), .A(n6851), .ZN(n6937) );
  INV_X1 U8688 ( .A(n6952), .ZN(n6853) );
  AOI211_X1 U8689 ( .C1(n6854), .C2(n6893), .A(n9306), .B(n6853), .ZN(n6936)
         );
  NAND2_X1 U8690 ( .A1(n6936), .A2(n4265), .ZN(n6857) );
  INV_X1 U8691 ( .A(n9309), .ZN(n9538) );
  INV_X1 U8692 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U8693 ( .A1(n9317), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9538), .B2(
        n6855), .ZN(n6856) );
  OAI211_X1 U8694 ( .C1(n6941), .C2(n9542), .A(n6857), .B(n6856), .ZN(n6858)
         );
  AOI21_X1 U8695 ( .B1(n9545), .B2(n6937), .A(n6858), .ZN(n6859) );
  OAI21_X1 U8696 ( .B1(n6860), .B2(n9317), .A(n6859), .ZN(P1_U3290) );
  INV_X1 U8697 ( .A(n6861), .ZN(n9564) );
  AOI211_X1 U8698 ( .C1(n9564), .C2(n6864), .A(n6863), .B(n6862), .ZN(n6869)
         );
  OAI22_X1 U8699 ( .A1(n9440), .A2(n5744), .B1(n9598), .B2(n5736), .ZN(n6865)
         );
  INV_X1 U8700 ( .A(n6865), .ZN(n6866) );
  OAI21_X1 U8701 ( .B1(n6869), .B2(n9589), .A(n6866), .ZN(P1_U3456) );
  OAI22_X1 U8702 ( .A1(n9401), .A2(n5744), .B1(n9608), .B2(n5739), .ZN(n6867)
         );
  INV_X1 U8703 ( .A(n6867), .ZN(n6868) );
  OAI21_X1 U8704 ( .B1(n6869), .B2(n9605), .A(n6868), .ZN(P1_U3523) );
  INV_X1 U8705 ( .A(n8220), .ZN(n8230) );
  OAI222_X1 U8706 ( .A1(P2_U3151), .A2(n8230), .B1(n8492), .B2(n6871), .C1(
        n6870), .C2(n8494), .ZN(P2_U3277) );
  INV_X1 U8707 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8708 ( .A1(n6872), .A2(n7768), .ZN(n6873) );
  AOI21_X1 U8709 ( .B1(n6905), .B2(n6873), .A(n9768), .ZN(n6876) );
  OAI22_X1 U8710 ( .A1(n6978), .A2(n8300), .B1(n6874), .B2(n8302), .ZN(n6875)
         );
  OR2_X1 U8711 ( .A1(n6876), .A2(n6875), .ZN(n9799) );
  AOI21_X1 U8712 ( .B1(n8368), .B2(n6877), .A(n9799), .ZN(n6878) );
  MUX2_X1 U8713 ( .A(n6879), .B(n6878), .S(n8366), .Z(n6883) );
  XNOR2_X1 U8714 ( .A(n6880), .B(n7768), .ZN(n9801) );
  AOI22_X1 U8715 ( .A1(n9801), .A2(n8333), .B1(n8369), .B2(n6881), .ZN(n6882)
         );
  NAND2_X1 U8716 ( .A1(n6883), .A2(n6882), .ZN(P2_U3226) );
  OAI21_X1 U8717 ( .B1(n6885), .B2(n8784), .A(n6884), .ZN(n9563) );
  INV_X1 U8718 ( .A(n9563), .ZN(n6901) );
  XNOR2_X1 U8719 ( .A(n8784), .B(n8670), .ZN(n6891) );
  OAI22_X1 U8720 ( .A1(n6887), .A2(n9261), .B1(n6886), .B2(n9263), .ZN(n6888)
         );
  AOI21_X1 U8721 ( .B1(n9563), .B2(n6889), .A(n6888), .ZN(n6890) );
  OAI21_X1 U8722 ( .B1(n9553), .B2(n6891), .A(n6890), .ZN(n9561) );
  NAND2_X1 U8723 ( .A1(n9561), .A2(n9287), .ZN(n6899) );
  INV_X1 U8724 ( .A(n9542), .ZN(n9268) );
  OAI22_X1 U8725 ( .A1(n9287), .A2(n6892), .B1(n8968), .B2(n9309), .ZN(n6896)
         );
  OAI211_X1 U8726 ( .C1(n6894), .C2(n9560), .A(n6893), .B(n9229), .ZN(n9559)
         );
  INV_X1 U8727 ( .A(n4265), .ZN(n9230) );
  NOR2_X1 U8728 ( .A1(n9559), .A2(n9230), .ZN(n6895) );
  AOI211_X1 U8729 ( .C1(n9268), .C2(n6897), .A(n6896), .B(n6895), .ZN(n6898)
         );
  OAI211_X1 U8730 ( .C1(n6901), .C2(n6900), .A(n6899), .B(n6898), .ZN(P1_U3291) );
  XOR2_X1 U8731 ( .A(n6902), .B(n7889), .Z(n9803) );
  INV_X1 U8732 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6910) );
  INV_X1 U8733 ( .A(n6903), .ZN(n6907) );
  AOI21_X1 U8734 ( .B1(n6905), .B2(n6904), .A(n7889), .ZN(n6906) );
  NOR3_X1 U8735 ( .A1(n6907), .A2(n6906), .A3(n9768), .ZN(n6909) );
  OAI22_X1 U8736 ( .A1(n5548), .A2(n8302), .B1(n7027), .B2(n8300), .ZN(n6908)
         );
  NOR2_X1 U8737 ( .A1(n6909), .A2(n6908), .ZN(n9804) );
  MUX2_X1 U8738 ( .A(n6910), .B(n9804), .S(n8366), .Z(n6913) );
  AOI22_X1 U8739 ( .A1(n8369), .A2(n6911), .B1(n8368), .B2(n6919), .ZN(n6912)
         );
  OAI211_X1 U8740 ( .C1(n9803), .C2(n8372), .A(n6913), .B(n6912), .ZN(P2_U3225) );
  XOR2_X1 U8741 ( .A(n6915), .B(n6914), .Z(n6921) );
  NOR2_X1 U8742 ( .A1(n8128), .A2(n9805), .ZN(n6918) );
  NAND2_X1 U8743 ( .A1(n8119), .A2(n8142), .ZN(n6916) );
  NAND2_X1 U8744 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n9679) );
  OAI211_X1 U8745 ( .C1(n8121), .C2(n7027), .A(n6916), .B(n9679), .ZN(n6917)
         );
  AOI211_X1 U8746 ( .C1(n6919), .C2(n8124), .A(n6918), .B(n6917), .ZN(n6920)
         );
  OAI21_X1 U8747 ( .B1(n6921), .B2(n8052), .A(n6920), .ZN(P2_U3161) );
  NAND2_X1 U8748 ( .A1(n6351), .A2(n6922), .ZN(n8820) );
  INV_X1 U8749 ( .A(n8820), .ZN(n6923) );
  NOR2_X1 U8750 ( .A1(n6924), .A2(n6923), .ZN(n9552) );
  INV_X1 U8751 ( .A(n9552), .ZN(n6926) );
  NAND3_X1 U8752 ( .A1(n6926), .A2(n6278), .A3(n6925), .ZN(n6927) );
  NAND2_X1 U8753 ( .A1(n5743), .A2(n9299), .ZN(n9551) );
  OAI211_X1 U8754 ( .C1(n9309), .C2(n6928), .A(n6927), .B(n9551), .ZN(n6931)
         );
  NOR3_X1 U8755 ( .A1(n9552), .A2(n6929), .A3(n9557), .ZN(n6930) );
  OAI21_X1 U8756 ( .B1(n6931), .B2(n6930), .A(n9287), .ZN(n6934) );
  OAI21_X1 U8757 ( .B1(n9230), .B2(n9306), .A(n9542), .ZN(n6932) );
  AOI22_X1 U8758 ( .A1(n6932), .A2(n9556), .B1(P1_REG2_REG_0__SCAN_IN), .B2(
        n9317), .ZN(n6933) );
  NAND2_X1 U8759 ( .A1(n6934), .A2(n6933), .ZN(P1_U3293) );
  AOI211_X1 U8760 ( .C1(n9595), .C2(n6937), .A(n6936), .B(n6935), .ZN(n6944)
         );
  INV_X1 U8761 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6938) );
  OAI22_X1 U8762 ( .A1(n9440), .A2(n6941), .B1(n9598), .B2(n6938), .ZN(n6939)
         );
  INV_X1 U8763 ( .A(n6939), .ZN(n6940) );
  OAI21_X1 U8764 ( .B1(n6944), .B2(n9589), .A(n6940), .ZN(P1_U3462) );
  OAI22_X1 U8765 ( .A1(n9401), .A2(n6941), .B1(n9608), .B2(n6547), .ZN(n6942)
         );
  INV_X1 U8766 ( .A(n6942), .ZN(n6943) );
  OAI21_X1 U8767 ( .B1(n6944), .B2(n9605), .A(n6943), .ZN(P1_U3525) );
  OAI21_X1 U8768 ( .B1(n6946), .B2(n8787), .A(n6945), .ZN(n6947) );
  INV_X1 U8769 ( .A(n6947), .ZN(n9570) );
  OAI21_X1 U8770 ( .B1(n6949), .B2(n6948), .A(n7102), .ZN(n6950) );
  AOI222_X1 U8771 ( .A1(n9295), .A2(n6950), .B1(n7073), .B2(n9299), .C1(n8946), 
        .C2(n9298), .ZN(n9569) );
  MUX2_X1 U8772 ( .A(n6951), .B(n9569), .S(n9287), .Z(n6956) );
  AOI211_X1 U8773 ( .C1(n9566), .C2(n6952), .A(n9306), .B(n7098), .ZN(n9565)
         );
  OAI22_X1 U8774 ( .A1(n9542), .A2(n8664), .B1(n9309), .B2(n6953), .ZN(n6954)
         );
  AOI21_X1 U8775 ( .B1(n9565), .B2(n4265), .A(n6954), .ZN(n6955) );
  OAI211_X1 U8776 ( .C1(n9290), .C2(n9570), .A(n6956), .B(n6955), .ZN(P1_U3289) );
  XNOR2_X1 U8777 ( .A(n6957), .B(n8790), .ZN(n6958) );
  NAND2_X1 U8778 ( .A1(n6958), .A2(n9295), .ZN(n6962) );
  OAI22_X1 U8779 ( .A1(n6959), .A2(n9261), .B1(n7085), .B2(n9263), .ZN(n6960)
         );
  INV_X1 U8780 ( .A(n6960), .ZN(n6961) );
  NAND2_X1 U8781 ( .A1(n6962), .A2(n6961), .ZN(n9576) );
  INV_X1 U8782 ( .A(n9576), .ZN(n6970) );
  OAI21_X1 U8783 ( .B1(n6964), .B2(n8790), .A(n6963), .ZN(n9578) );
  OAI211_X1 U8784 ( .C1(n7099), .C2(n9575), .A(n9229), .B(n7052), .ZN(n9574)
         );
  INV_X1 U8785 ( .A(n6965), .ZN(n7075) );
  AOI22_X1 U8786 ( .A1(n9317), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7075), .B2(
        n9538), .ZN(n6967) );
  NAND2_X1 U8787 ( .A1(n9268), .A2(n7074), .ZN(n6966) );
  OAI211_X1 U8788 ( .C1(n9574), .C2(n9230), .A(n6967), .B(n6966), .ZN(n6968)
         );
  AOI21_X1 U8789 ( .B1(n9578), .B2(n9545), .A(n6968), .ZN(n6969) );
  OAI21_X1 U8790 ( .B1(n9317), .B2(n6970), .A(n6969), .ZN(P1_U3287) );
  INV_X1 U8791 ( .A(n6971), .ZN(n7956) );
  OAI222_X1 U8792 ( .A1(n7964), .A2(n6972), .B1(n7960), .B2(n7956), .C1(n9264), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U8793 ( .A(n6973), .ZN(n7892) );
  XNOR2_X1 U8794 ( .A(n6974), .B(n7892), .ZN(n9813) );
  NAND2_X1 U8795 ( .A1(n9813), .A2(n6975), .ZN(n6982) );
  XNOR2_X1 U8796 ( .A(n6976), .B(n7892), .ZN(n6980) );
  NAND2_X1 U8797 ( .A1(n8139), .A2(n8362), .ZN(n6977) );
  OAI21_X1 U8798 ( .B1(n6978), .B2(n8302), .A(n6977), .ZN(n6979) );
  AOI21_X1 U8799 ( .B1(n6980), .B2(n8365), .A(n6979), .ZN(n6981) );
  AND2_X1 U8800 ( .A1(n6982), .A2(n6981), .ZN(n9815) );
  AOI22_X1 U8801 ( .A1(n8336), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8368), .B2(
        n8074), .ZN(n6983) );
  OAI21_X1 U8802 ( .B1(n9810), .B2(n8330), .A(n6983), .ZN(n6984) );
  AOI21_X1 U8803 ( .B1(n9813), .B2(n8001), .A(n6984), .ZN(n6985) );
  OAI21_X1 U8804 ( .B1(n9815), .B2(n8336), .A(n6985), .ZN(P2_U3224) );
  INV_X1 U8805 ( .A(n8543), .ZN(n9079) );
  NAND2_X1 U8806 ( .A1(n9079), .A2(P1_U3973), .ZN(n6986) );
  OAI21_X1 U8807 ( .B1(n6323), .B2(P1_U3973), .A(n6986), .ZN(P1_U3583) );
  INV_X1 U8808 ( .A(n6988), .ZN(n6989) );
  AOI21_X1 U8809 ( .B1(n6990), .B2(n6987), .A(n6989), .ZN(n6997) );
  NAND2_X1 U8810 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9472) );
  INV_X1 U8811 ( .A(n9472), .ZN(n6992) );
  NOR2_X1 U8812 ( .A1(n7050), .A2(n8624), .ZN(n6991) );
  AOI211_X1 U8813 ( .C1(n8627), .C2(n6993), .A(n6992), .B(n6991), .ZN(n6994)
         );
  OAI21_X1 U8814 ( .B1(n8635), .B2(n7054), .A(n6994), .ZN(n6995) );
  AOI21_X1 U8815 ( .B1(n7051), .B2(n8641), .A(n6995), .ZN(n6996) );
  OAI21_X1 U8816 ( .B1(n6997), .B2(n8643), .A(n6996), .ZN(P1_U3213) );
  XNOR2_X1 U8817 ( .A(n6998), .B(n6999), .ZN(n7000) );
  NAND2_X1 U8818 ( .A1(n7000), .A2(n7001), .ZN(n7066) );
  OAI21_X1 U8819 ( .B1(n7001), .B2(n7000), .A(n7066), .ZN(n7002) );
  NAND2_X1 U8820 ( .A1(n7002), .A2(n8603), .ZN(n7008) );
  INV_X1 U8821 ( .A(n7003), .ZN(n9539) );
  NAND2_X1 U8822 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9008) );
  INV_X1 U8823 ( .A(n9008), .ZN(n7004) );
  AOI21_X1 U8824 ( .B1(n8945), .B2(n8636), .A(n7004), .ZN(n7005) );
  OAI21_X1 U8825 ( .B1(n7050), .B2(n8638), .A(n7005), .ZN(n7006) );
  AOI21_X1 U8826 ( .B1(n9539), .B2(n8607), .A(n7006), .ZN(n7007) );
  OAI211_X1 U8827 ( .C1(n9543), .C2(n8610), .A(n7008), .B(n7007), .ZN(P1_U3227) );
  NAND2_X1 U8828 ( .A1(n4659), .A2(P2_U3893), .ZN(n7010) );
  OAI21_X1 U8829 ( .B1(n6322), .B2(P2_U3893), .A(n7010), .ZN(P2_U3520) );
  NAND2_X1 U8830 ( .A1(n7011), .A2(n7780), .ZN(n7013) );
  XNOR2_X1 U8831 ( .A(n7013), .B(n7012), .ZN(n9824) );
  INV_X1 U8832 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7015) );
  INV_X1 U8833 ( .A(n7318), .ZN(n7014) );
  OAI22_X1 U8834 ( .A1(n8366), .A2(n7015), .B1(n7014), .B2(n7996), .ZN(n7016)
         );
  AOI21_X1 U8835 ( .B1(n8369), .B2(n9827), .A(n7016), .ZN(n7022) );
  XNOR2_X1 U8836 ( .A(n7017), .B(n7894), .ZN(n7018) );
  NAND2_X1 U8837 ( .A1(n7018), .A2(n8365), .ZN(n7020) );
  AOI22_X1 U8838 ( .A1(n8360), .A2(n8139), .B1(n8137), .B2(n8362), .ZN(n7019)
         );
  NAND2_X1 U8839 ( .A1(n7020), .A2(n7019), .ZN(n9826) );
  NAND2_X1 U8840 ( .A1(n9826), .A2(n8366), .ZN(n7021) );
  OAI211_X1 U8841 ( .C1(n9824), .C2(n8372), .A(n7022), .B(n7021), .ZN(P2_U3222) );
  NAND2_X1 U8842 ( .A1(n7025), .A2(n7024), .ZN(n7893) );
  XNOR2_X1 U8843 ( .A(n7023), .B(n7893), .ZN(n9819) );
  XNOR2_X1 U8844 ( .A(n7026), .B(n7893), .ZN(n7029) );
  OAI22_X1 U8845 ( .A1(n7027), .A2(n8302), .B1(n7217), .B2(n8300), .ZN(n7028)
         );
  AOI21_X1 U8846 ( .B1(n7029), .B2(n8365), .A(n7028), .ZN(n7030) );
  OAI21_X1 U8847 ( .B1(n9819), .B2(n7031), .A(n7030), .ZN(n9821) );
  NAND2_X1 U8848 ( .A1(n9821), .A2(n8366), .ZN(n7037) );
  INV_X1 U8849 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7033) );
  INV_X1 U8850 ( .A(n7220), .ZN(n7032) );
  OAI22_X1 U8851 ( .A1(n8366), .A2(n7033), .B1(n7032), .B2(n7996), .ZN(n7034)
         );
  AOI21_X1 U8852 ( .B1(n8369), .B2(n7035), .A(n7034), .ZN(n7036) );
  OAI211_X1 U8853 ( .C1(n9819), .C2(n7038), .A(n7037), .B(n7036), .ZN(P2_U3223) );
  OAI21_X1 U8854 ( .B1(n7040), .B2(n7041), .A(n7039), .ZN(n7194) );
  INV_X1 U8855 ( .A(n7194), .ZN(n7060) );
  INV_X1 U8856 ( .A(n7041), .ZN(n7044) );
  NOR2_X1 U8857 ( .A1(n7044), .A2(n8688), .ZN(n7048) );
  NAND2_X1 U8858 ( .A1(n8829), .A2(n7042), .ZN(n8685) );
  INV_X1 U8859 ( .A(n8685), .ZN(n8677) );
  NAND2_X1 U8860 ( .A1(n7043), .A2(n8677), .ZN(n7047) );
  NAND2_X1 U8861 ( .A1(n7047), .A2(n8679), .ZN(n7045) );
  NAND2_X1 U8862 ( .A1(n7045), .A2(n7044), .ZN(n7296) );
  INV_X1 U8863 ( .A(n7296), .ZN(n7046) );
  AOI21_X1 U8864 ( .B1(n7048), .B2(n7047), .A(n7046), .ZN(n7049) );
  OAI222_X1 U8865 ( .A1(n9263), .A2(n7331), .B1(n9261), .B2(n7050), .C1(n9553), 
        .C2(n7049), .ZN(n7192) );
  NAND2_X1 U8866 ( .A1(n7192), .A2(n9287), .ZN(n7059) );
  AOI21_X1 U8867 ( .B1(n7052), .B2(n7051), .A(n9306), .ZN(n7053) );
  AND2_X1 U8868 ( .A1(n7053), .A2(n4352), .ZN(n7193) );
  NOR2_X1 U8869 ( .A1(n9309), .A2(n7054), .ZN(n7055) );
  AOI21_X1 U8870 ( .B1(n9317), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7055), .ZN(
        n7056) );
  OAI21_X1 U8871 ( .B1(n9542), .B2(n7198), .A(n7056), .ZN(n7057) );
  AOI21_X1 U8872 ( .B1(n7193), .B2(n4265), .A(n7057), .ZN(n7058) );
  OAI211_X1 U8873 ( .C1(n9290), .C2(n7060), .A(n7059), .B(n7058), .ZN(P1_U3286) );
  INV_X1 U8874 ( .A(n7061), .ZN(n7065) );
  OAI222_X1 U8875 ( .A1(n8494), .A2(n7063), .B1(n8492), .B2(n7065), .C1(n7062), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7064) );
  OAI222_X1 U8877 ( .A1(n8893), .A2(P1_U3086), .B1(n7960), .B2(n7065), .C1(
        n7064), .C2(n7964), .ZN(P1_U3335) );
  OAI21_X1 U8878 ( .B1(n7067), .B2(n6998), .A(n7066), .ZN(n7071) );
  XNOR2_X1 U8879 ( .A(n7069), .B(n7068), .ZN(n7070) );
  XNOR2_X1 U8880 ( .A(n7071), .B(n7070), .ZN(n7081) );
  NAND2_X1 U8881 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9021) );
  INV_X1 U8882 ( .A(n9021), .ZN(n7072) );
  AOI21_X1 U8883 ( .B1(n7073), .B2(n8636), .A(n7072), .ZN(n7079) );
  NAND2_X1 U8884 ( .A1(n8641), .A2(n7074), .ZN(n7078) );
  NAND2_X1 U8885 ( .A1(n8607), .A2(n7075), .ZN(n7077) );
  OR2_X1 U8886 ( .A1(n7085), .A2(n8638), .ZN(n7076) );
  NAND4_X1 U8887 ( .A1(n7079), .A2(n7078), .A3(n7077), .A4(n7076), .ZN(n7080)
         );
  AOI21_X1 U8888 ( .B1(n7081), .B2(n8603), .A(n7080), .ZN(n7082) );
  INV_X1 U8889 ( .A(n7082), .ZN(P1_U3239) );
  NAND2_X1 U8890 ( .A1(n7296), .A2(n8680), .ZN(n7083) );
  XNOR2_X1 U8891 ( .A(n7083), .B(n7091), .ZN(n7084) );
  OAI222_X1 U8892 ( .A1(n9263), .A2(n7401), .B1(n9261), .B2(n7085), .C1(n7084), 
        .C2(n9553), .ZN(n7183) );
  INV_X1 U8893 ( .A(n7183), .ZN(n7095) );
  AOI21_X1 U8894 ( .B1(n4352), .B2(n7206), .A(n9306), .ZN(n7086) );
  AND2_X1 U8895 ( .A1(n7293), .A2(n7086), .ZN(n7184) );
  NOR2_X1 U8896 ( .A1(n9309), .A2(n7207), .ZN(n7087) );
  AOI21_X1 U8897 ( .B1(n9317), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7087), .ZN(
        n7088) );
  OAI21_X1 U8898 ( .B1(n9542), .B2(n6391), .A(n7088), .ZN(n7089) );
  AOI21_X1 U8899 ( .B1(n7184), .B2(n4265), .A(n7089), .ZN(n7094) );
  OAI21_X1 U8900 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7185) );
  NAND2_X1 U8901 ( .A1(n7185), .A2(n9545), .ZN(n7093) );
  OAI211_X1 U8902 ( .C1(n7095), .C2(n9317), .A(n7094), .B(n7093), .ZN(P1_U3285) );
  OAI21_X1 U8903 ( .B1(n7097), .B2(n8789), .A(n7096), .ZN(n9546) );
  INV_X1 U8904 ( .A(n7098), .ZN(n7100) );
  AOI211_X1 U8905 ( .C1(n7107), .C2(n7100), .A(n9306), .B(n7099), .ZN(n9537)
         );
  NAND2_X1 U8906 ( .A1(n7102), .A2(n7101), .ZN(n7103) );
  XOR2_X1 U8907 ( .A(n8789), .B(n7103), .Z(n7104) );
  AOI222_X1 U8908 ( .A1(n9295), .A2(n7104), .B1(n8944), .B2(n9299), .C1(n8945), 
        .C2(n9298), .ZN(n9548) );
  INV_X1 U8909 ( .A(n9548), .ZN(n7105) );
  AOI211_X1 U8910 ( .C1(n9595), .C2(n9546), .A(n9537), .B(n7105), .ZN(n7109)
         );
  INV_X1 U8911 ( .A(n9401), .ZN(n7673) );
  AOI22_X1 U8912 ( .A1(n7673), .A2(n7107), .B1(n9605), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7106) );
  OAI21_X1 U8913 ( .B1(n7109), .B2(n9605), .A(n7106), .ZN(P1_U3527) );
  INV_X1 U8914 ( .A(n9440), .ZN(n7671) );
  AOI22_X1 U8915 ( .A1(n7671), .A2(n7107), .B1(n9589), .B2(
        P1_REG0_REG_5__SCAN_IN), .ZN(n7108) );
  OAI21_X1 U8916 ( .B1(n7109), .B2(n9589), .A(n7108), .ZN(P1_U3468) );
  XNOR2_X1 U8917 ( .A(n7110), .B(n8137), .ZN(n7111) );
  XNOR2_X1 U8918 ( .A(n4360), .B(n7111), .ZN(n7117) );
  NOR2_X1 U8919 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7112), .ZN(n7256) );
  AOI21_X1 U8920 ( .B1(n8107), .B2(n8136), .A(n7256), .ZN(n7114) );
  NAND2_X1 U8921 ( .A1(n8124), .A2(n7179), .ZN(n7113) );
  OAI211_X1 U8922 ( .C1(n7217), .C2(n8109), .A(n7114), .B(n7113), .ZN(n7115)
         );
  AOI21_X1 U8923 ( .B1(n7790), .B2(n8072), .A(n7115), .ZN(n7116) );
  OAI21_X1 U8924 ( .B1(n7117), .B2(n8052), .A(n7116), .ZN(P2_U3164) );
  INV_X1 U8925 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7120) );
  XNOR2_X1 U8926 ( .A(n7118), .B(n7796), .ZN(n7119) );
  AOI222_X1 U8927 ( .A1(n8365), .A2(n7119), .B1(n8136), .B2(n8362), .C1(n8138), 
        .C2(n8360), .ZN(n7178) );
  MUX2_X1 U8928 ( .A(n7120), .B(n7178), .S(n9829), .Z(n7123) );
  INV_X1 U8929 ( .A(n7796), .ZN(n7897) );
  XNOR2_X1 U8930 ( .A(n7121), .B(n7897), .ZN(n7177) );
  INV_X1 U8931 ( .A(n8481), .ZN(n8459) );
  AOI22_X1 U8932 ( .A1(n7177), .A2(n8459), .B1(n8477), .B2(n7790), .ZN(n7122)
         );
  NAND2_X1 U8933 ( .A1(n7123), .A2(n7122), .ZN(P2_U3426) );
  INV_X1 U8934 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7547) );
  MUX2_X1 U8935 ( .A(n7547), .B(n7178), .S(n9851), .Z(n7125) );
  INV_X1 U8936 ( .A(n8416), .ZN(n8403) );
  AOI22_X1 U8937 ( .A1(n7177), .A2(n8403), .B1(n8413), .B2(n7790), .ZN(n7124)
         );
  NAND2_X1 U8938 ( .A1(n7125), .A2(n7124), .ZN(P2_U3471) );
  NOR2_X1 U8939 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7167) );
  NOR2_X1 U8940 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7164) );
  NOR2_X1 U8941 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7161) );
  NOR2_X1 U8942 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7158) );
  NOR2_X1 U8943 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7156) );
  NOR2_X1 U8944 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7154) );
  NOR2_X1 U8945 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7152) );
  NOR2_X1 U8946 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7150) );
  NOR2_X1 U8947 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7148) );
  NOR2_X1 U8948 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7146) );
  NOR2_X1 U8949 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7143) );
  NOR2_X1 U8950 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7141) );
  NOR2_X1 U8951 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7139) );
  NOR2_X1 U8952 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7137) );
  NAND2_X1 U8953 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7134) );
  XNOR2_X1 U8954 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n7126), .ZN(n10052) );
  NAND2_X1 U8955 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7132) );
  AOI21_X1 U8956 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9852) );
  INV_X1 U8957 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U8958 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7127) );
  NOR2_X1 U8959 ( .A1(n7128), .A2(n7127), .ZN(n9853) );
  NOR2_X1 U8960 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9853), .ZN(n7129) );
  NOR2_X1 U8961 ( .A1(n9852), .A2(n7129), .ZN(n10050) );
  XNOR2_X1 U8962 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n7130), .ZN(n10049) );
  NAND2_X1 U8963 ( .A1(n10050), .A2(n10049), .ZN(n7131) );
  NAND2_X1 U8964 ( .A1(n7132), .A2(n7131), .ZN(n10051) );
  NAND2_X1 U8965 ( .A1(n10052), .A2(n10051), .ZN(n7133) );
  NAND2_X1 U8966 ( .A1(n7134), .A2(n7133), .ZN(n10054) );
  INV_X1 U8967 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7135) );
  AOI22_X1 U8968 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n7135), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n9959), .ZN(n10053) );
  NOR2_X1 U8969 ( .A1(n10054), .A2(n10053), .ZN(n7136) );
  NOR2_X1 U8970 ( .A1(n7137), .A2(n7136), .ZN(n10042) );
  INV_X1 U8971 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9630) );
  XOR2_X1 U8972 ( .A(n9630), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10041) );
  NOR2_X1 U8973 ( .A1(n10042), .A2(n10041), .ZN(n7138) );
  NOR2_X1 U8974 ( .A1(n7139), .A2(n7138), .ZN(n10040) );
  INV_X1 U8975 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9022) );
  XOR2_X1 U8976 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n9022), .Z(n10039) );
  NOR2_X1 U8977 ( .A1(n10040), .A2(n10039), .ZN(n7140) );
  NOR2_X1 U8978 ( .A1(n7141), .A2(n7140), .ZN(n10046) );
  INV_X1 U8979 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9474) );
  INV_X1 U8980 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9663) );
  AOI22_X1 U8981 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9474), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n9663), .ZN(n10045) );
  NOR2_X1 U8982 ( .A1(n10046), .A2(n10045), .ZN(n7142) );
  NOR2_X1 U8983 ( .A1(n7143), .A2(n7142), .ZN(n10048) );
  INV_X1 U8984 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9905) );
  INV_X1 U8985 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7144) );
  AOI22_X1 U8986 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9905), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n7144), .ZN(n10047) );
  NOR2_X1 U8987 ( .A1(n10048), .A2(n10047), .ZN(n7145) );
  NOR2_X1 U8988 ( .A1(n7146), .A2(n7145), .ZN(n10044) );
  XNOR2_X1 U8989 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10043) );
  NOR2_X1 U8990 ( .A1(n10044), .A2(n10043), .ZN(n7147) );
  NOR2_X1 U8991 ( .A1(n7148), .A2(n7147), .ZN(n9873) );
  INV_X1 U8992 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9461) );
  XOR2_X1 U8993 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n9461), .Z(n9872) );
  NOR2_X1 U8994 ( .A1(n9873), .A2(n9872), .ZN(n7149) );
  NOR2_X1 U8995 ( .A1(n7150), .A2(n7149), .ZN(n9871) );
  XNOR2_X1 U8996 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9870) );
  NOR2_X1 U8997 ( .A1(n9871), .A2(n9870), .ZN(n7151) );
  NOR2_X1 U8998 ( .A1(n7152), .A2(n7151), .ZN(n9869) );
  XNOR2_X1 U8999 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9868) );
  NOR2_X1 U9000 ( .A1(n9869), .A2(n9868), .ZN(n7153) );
  NOR2_X1 U9001 ( .A1(n7154), .A2(n7153), .ZN(n9867) );
  INV_X1 U9002 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9519) );
  XOR2_X1 U9003 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9519), .Z(n9866) );
  NOR2_X1 U9004 ( .A1(n9867), .A2(n9866), .ZN(n7155) );
  NOR2_X1 U9005 ( .A1(n7156), .A2(n7155), .ZN(n9865) );
  INV_X1 U9006 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9535) );
  XOR2_X1 U9007 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9535), .Z(n9864) );
  NOR2_X1 U9008 ( .A1(n9865), .A2(n9864), .ZN(n7157) );
  NOR2_X1 U9009 ( .A1(n7158), .A2(n7157), .ZN(n9863) );
  INV_X1 U9010 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9891) );
  INV_X1 U9011 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7159) );
  AOI22_X1 U9012 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9891), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n7159), .ZN(n9862) );
  NOR2_X1 U9013 ( .A1(n9863), .A2(n9862), .ZN(n7160) );
  NOR2_X1 U9014 ( .A1(n7161), .A2(n7160), .ZN(n9861) );
  INV_X1 U9015 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7162) );
  INV_X1 U9016 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8162) );
  AOI22_X1 U9017 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7162), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8162), .ZN(n9860) );
  NOR2_X1 U9018 ( .A1(n9861), .A2(n9860), .ZN(n7163) );
  NOR2_X1 U9019 ( .A1(n7164), .A2(n7163), .ZN(n9859) );
  INV_X1 U9020 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7165) );
  INV_X1 U9021 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8191) );
  AOI22_X1 U9022 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7165), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8191), .ZN(n9858) );
  NOR2_X1 U9023 ( .A1(n9859), .A2(n9858), .ZN(n7166) );
  NOR2_X1 U9024 ( .A1(n7167), .A2(n7166), .ZN(n7168) );
  NOR2_X1 U9025 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7168), .ZN(n9855) );
  AND2_X1 U9026 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7168), .ZN(n9856) );
  NOR2_X1 U9027 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9856), .ZN(n7169) );
  NOR2_X1 U9028 ( .A1(n9855), .A2(n7169), .ZN(n7171) );
  XNOR2_X1 U9029 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n7170) );
  XNOR2_X1 U9030 ( .A(n7171), .B(n7170), .ZN(ADD_1068_U4) );
  INV_X1 U9031 ( .A(n7172), .ZN(n7175) );
  OAI222_X1 U9032 ( .A1(n8819), .A2(P1_U3086), .B1(n7960), .B2(n7175), .C1(
        n7173), .C2(n7964), .ZN(P1_U3334) );
  OAI222_X1 U9033 ( .A1(n8494), .A2(n7176), .B1(n8492), .B2(n7175), .C1(n7174), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U9034 ( .A(n7177), .ZN(n7182) );
  INV_X1 U9035 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7236) );
  MUX2_X1 U9036 ( .A(n7236), .B(n7178), .S(n8366), .Z(n7181) );
  AOI22_X1 U9037 ( .A1(n7790), .A2(n8369), .B1(n8368), .B2(n7179), .ZN(n7180)
         );
  OAI211_X1 U9038 ( .C1(n7182), .C2(n8372), .A(n7181), .B(n7180), .ZN(P2_U3221) );
  AOI211_X1 U9039 ( .C1(n9595), .C2(n7185), .A(n7184), .B(n7183), .ZN(n7191)
         );
  NOR2_X1 U9040 ( .A1(n9608), .A2(n5883), .ZN(n7186) );
  AOI21_X1 U9041 ( .B1(n7673), .B2(n7206), .A(n7186), .ZN(n7187) );
  OAI21_X1 U9042 ( .B1(n7191), .B2(n9605), .A(n7187), .ZN(P1_U3530) );
  INV_X1 U9043 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7188) );
  NOR2_X1 U9044 ( .A1(n9598), .A2(n7188), .ZN(n7189) );
  AOI21_X1 U9045 ( .B1(n7671), .B2(n7206), .A(n7189), .ZN(n7190) );
  OAI21_X1 U9046 ( .B1(n7191), .B2(n9589), .A(n7190), .ZN(P1_U3477) );
  AOI211_X1 U9047 ( .C1(n9595), .C2(n7194), .A(n7193), .B(n7192), .ZN(n7201)
         );
  OAI22_X1 U9048 ( .A1(n9401), .A2(n7198), .B1(n9608), .B2(n5861), .ZN(n7195)
         );
  INV_X1 U9049 ( .A(n7195), .ZN(n7196) );
  OAI21_X1 U9050 ( .B1(n7201), .B2(n9605), .A(n7196), .ZN(P1_U3529) );
  INV_X1 U9051 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7197) );
  OAI22_X1 U9052 ( .A1(n9440), .A2(n7198), .B1(n9598), .B2(n7197), .ZN(n7199)
         );
  INV_X1 U9053 ( .A(n7199), .ZN(n7200) );
  OAI21_X1 U9054 ( .B1(n7201), .B2(n9589), .A(n7200), .ZN(P1_U3474) );
  OAI21_X1 U9055 ( .B1(n7204), .B2(n7202), .A(n7203), .ZN(n7214) );
  NAND2_X1 U9056 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9488) );
  INV_X1 U9057 ( .A(n9488), .ZN(n7205) );
  AOI21_X1 U9058 ( .B1(n5866), .B2(n8636), .A(n7205), .ZN(n7212) );
  NAND2_X1 U9059 ( .A1(n8641), .A2(n7206), .ZN(n7211) );
  INV_X1 U9060 ( .A(n7207), .ZN(n7208) );
  NAND2_X1 U9061 ( .A1(n8607), .A2(n7208), .ZN(n7210) );
  OR2_X1 U9062 ( .A1(n7401), .A2(n8638), .ZN(n7209) );
  NAND4_X1 U9063 ( .A1(n7212), .A2(n7211), .A3(n7210), .A4(n7209), .ZN(n7213)
         );
  AOI21_X1 U9064 ( .B1(n7214), .B2(n8603), .A(n7213), .ZN(n7215) );
  INV_X1 U9065 ( .A(n7215), .ZN(P1_U3221) );
  XNOR2_X1 U9066 ( .A(n7312), .B(n8139), .ZN(n7314) );
  XNOR2_X1 U9067 ( .A(n7314), .B(n7311), .ZN(n7222) );
  NOR2_X1 U9068 ( .A1(n9817), .A2(n8128), .ZN(n7219) );
  NAND2_X1 U9069 ( .A1(n8119), .A2(n8140), .ZN(n7216) );
  NAND2_X1 U9070 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n9710) );
  OAI211_X1 U9071 ( .C1(n8121), .C2(n7217), .A(n7216), .B(n9710), .ZN(n7218)
         );
  AOI211_X1 U9072 ( .C1(n7220), .C2(n8124), .A(n7219), .B(n7218), .ZN(n7221)
         );
  OAI21_X1 U9073 ( .B1(n7222), .B2(n8052), .A(n7221), .ZN(P2_U3157) );
  NAND2_X1 U9074 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7259), .ZN(n7233) );
  INV_X1 U9075 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7223) );
  MUX2_X1 U9076 ( .A(n7223), .B(P2_REG1_REG_10__SCAN_IN), .S(n9697), .Z(n9702)
         );
  NAND2_X1 U9077 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7263), .ZN(n7230) );
  INV_X1 U9078 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U9079 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7263), .B1(n9668), .B2(
        n9844), .ZN(n9675) );
  NAND2_X1 U9080 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n7275), .ZN(n7227) );
  INV_X1 U9081 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U9082 ( .A1(n9643), .A2(n9840), .B1(P2_REG1_REG_6__SCAN_IN), .B2(
        n7275), .ZN(n9636) );
  AOI21_X1 U9083 ( .B1(n7270), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7224), .ZN(
        n7225) );
  OR2_X1 U9084 ( .A1(n7225), .A2(n9627), .ZN(n7226) );
  XNOR2_X1 U9085 ( .A(n7225), .B(n7242), .ZN(n9618) );
  NAND2_X1 U9086 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(n9618), .ZN(n9617) );
  NAND2_X1 U9087 ( .A1(n7265), .A2(n7228), .ZN(n7229) );
  NAND2_X1 U9088 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n9651), .ZN(n9650) );
  NAND2_X1 U9089 ( .A1(n7229), .A2(n9650), .ZN(n9676) );
  NAND2_X1 U9090 ( .A1(n9675), .A2(n9676), .ZN(n9674) );
  NAND2_X1 U9091 ( .A1(n7230), .A2(n9674), .ZN(n7231) );
  NAND2_X1 U9092 ( .A1(n9695), .A2(n7231), .ZN(n7232) );
  XNOR2_X1 U9093 ( .A(n7231), .B(n7261), .ZN(n9686) );
  NAND2_X1 U9094 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n9686), .ZN(n9685) );
  NAND2_X1 U9095 ( .A1(n7232), .A2(n9685), .ZN(n9703) );
  NAND2_X1 U9096 ( .A1(n9702), .A2(n9703), .ZN(n9701) );
  NAND2_X1 U9097 ( .A1(n7233), .A2(n9701), .ZN(n7234) );
  NAND2_X1 U9098 ( .A1(n9726), .A2(n7234), .ZN(n7235) );
  XNOR2_X1 U9099 ( .A(n7234), .B(n7257), .ZN(n9717) );
  NAND2_X1 U9100 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9717), .ZN(n9716) );
  XNOR2_X1 U9101 ( .A(n7548), .B(n7547), .ZN(n7549) );
  XNOR2_X1 U9102 ( .A(n7546), .B(n7549), .ZN(n7291) );
  NOR2_X1 U9103 ( .A1(n7548), .A2(n7236), .ZN(n7237) );
  AOI21_X1 U9104 ( .B1(n7548), .B2(n7236), .A(n7237), .ZN(n7255) );
  NAND2_X1 U9105 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7259), .ZN(n7251) );
  MUX2_X1 U9106 ( .A(n7033), .B(P2_REG2_REG_10__SCAN_IN), .S(n9697), .Z(n9699)
         );
  NAND2_X1 U9107 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7263), .ZN(n7248) );
  AOI22_X1 U9108 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7263), .B1(n9668), .B2(
        n6910), .ZN(n9667) );
  NAND2_X1 U9109 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n7275), .ZN(n7245) );
  AOI22_X1 U9110 ( .A1(n9643), .A2(n7238), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n7275), .ZN(n9633) );
  NAND2_X1 U9111 ( .A1(n7243), .A2(n7242), .ZN(n7244) );
  NAND2_X1 U9112 ( .A1(n7265), .A2(n7246), .ZN(n7247) );
  NAND2_X1 U9113 ( .A1(n9695), .A2(n7249), .ZN(n7250) );
  XNOR2_X1 U9114 ( .A(n7249), .B(n7261), .ZN(n9684) );
  NAND2_X1 U9115 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n9684), .ZN(n9683) );
  NAND2_X1 U9116 ( .A1(n7250), .A2(n9683), .ZN(n9700) );
  NAND2_X1 U9117 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  NAND2_X1 U9118 ( .A1(n7251), .A2(n9698), .ZN(n7252) );
  NAND2_X1 U9119 ( .A1(n9726), .A2(n7252), .ZN(n7253) );
  XNOR2_X1 U9120 ( .A(n7252), .B(n7257), .ZN(n9715) );
  NAND2_X1 U9121 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n9715), .ZN(n9714) );
  NAND2_X1 U9122 ( .A1(n7253), .A2(n9714), .ZN(n7254) );
  NAND2_X1 U9123 ( .A1(n7254), .A2(n7255), .ZN(n7541) );
  OAI21_X1 U9124 ( .B1(n7255), .B2(n7254), .A(n7541), .ZN(n7289) );
  INV_X1 U9125 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7287) );
  AOI21_X1 U9126 ( .B1(n9696), .B2(n7548), .A(n7256), .ZN(n7286) );
  XNOR2_X1 U9127 ( .A(n7559), .B(n7548), .ZN(n7283) );
  OR2_X1 U9128 ( .A1(n7258), .A2(n9726), .ZN(n7281) );
  XNOR2_X1 U9129 ( .A(n7258), .B(n7257), .ZN(n9720) );
  OR2_X1 U9130 ( .A1(n7260), .A2(n7259), .ZN(n7280) );
  XNOR2_X1 U9131 ( .A(n7260), .B(n9697), .ZN(n9706) );
  OR2_X1 U9132 ( .A1(n7262), .A2(n9695), .ZN(n7279) );
  XNOR2_X1 U9133 ( .A(n7262), .B(n7261), .ZN(n9689) );
  OR2_X1 U9134 ( .A1(n7264), .A2(n7263), .ZN(n7278) );
  XNOR2_X1 U9135 ( .A(n7264), .B(n9668), .ZN(n9672) );
  OR2_X1 U9136 ( .A1(n7266), .A2(n7265), .ZN(n7277) );
  XNOR2_X1 U9137 ( .A(n7266), .B(n9660), .ZN(n9655) );
  XNOR2_X1 U9138 ( .A(n7276), .B(n9643), .ZN(n9641) );
  INV_X1 U9139 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7267) );
  NOR2_X1 U9140 ( .A1(n7272), .A2(n9627), .ZN(n7274) );
  AOI21_X1 U9141 ( .B1(n7271), .B2(n7270), .A(n7269), .ZN(n9624) );
  AOI21_X1 U9142 ( .B1(n9627), .B2(n7272), .A(n7274), .ZN(n7273) );
  INV_X1 U9143 ( .A(n7273), .ZN(n9623) );
  NOR2_X1 U9144 ( .A1(n9624), .A2(n9623), .ZN(n9621) );
  NOR2_X1 U9145 ( .A1(n7274), .A2(n9621), .ZN(n9640) );
  NAND2_X1 U9146 ( .A1(n9641), .A2(n9640), .ZN(n9639) );
  OAI21_X1 U9147 ( .B1(n7276), .B2(n7275), .A(n9639), .ZN(n9656) );
  NAND2_X1 U9148 ( .A1(n9655), .A2(n9656), .ZN(n9654) );
  NAND2_X1 U9149 ( .A1(n7277), .A2(n9654), .ZN(n9671) );
  NAND2_X1 U9150 ( .A1(n9672), .A2(n9671), .ZN(n9670) );
  NAND2_X1 U9151 ( .A1(n7278), .A2(n9670), .ZN(n9688) );
  NAND2_X1 U9152 ( .A1(n9689), .A2(n9688), .ZN(n9687) );
  NAND2_X1 U9153 ( .A1(n7279), .A2(n9687), .ZN(n9705) );
  NAND2_X1 U9154 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  NAND2_X1 U9155 ( .A1(n7280), .A2(n9704), .ZN(n9719) );
  NAND2_X1 U9156 ( .A1(n9720), .A2(n9719), .ZN(n9718) );
  NAND2_X1 U9157 ( .A1(n7281), .A2(n9718), .ZN(n7282) );
  NAND2_X1 U9158 ( .A1(n7283), .A2(n7282), .ZN(n7560) );
  OAI21_X1 U9159 ( .B1(n7283), .B2(n7282), .A(n7560), .ZN(n7284) );
  NAND2_X1 U9160 ( .A1(n7284), .A2(n9750), .ZN(n7285) );
  OAI211_X1 U9161 ( .C1(n9664), .C2(n7287), .A(n7286), .B(n7285), .ZN(n7288)
         );
  AOI21_X1 U9162 ( .B1(n7289), .B2(n9737), .A(n7288), .ZN(n7290) );
  OAI21_X1 U9163 ( .B1(n7292), .B2(n7291), .A(n7290), .ZN(P2_U3194) );
  XNOR2_X1 U9164 ( .A(n7293), .B(n4515), .ZN(n7295) );
  NOR2_X1 U9165 ( .A1(n7600), .A2(n9263), .ZN(n7294) );
  AOI21_X1 U9166 ( .B1(n7295), .B2(n9229), .A(n7294), .ZN(n9580) );
  INV_X1 U9167 ( .A(n9580), .ZN(n7302) );
  NAND2_X1 U9168 ( .A1(n7296), .A2(n8690), .ZN(n7297) );
  NAND2_X1 U9169 ( .A1(n7297), .A2(n8692), .ZN(n7298) );
  XNOR2_X1 U9170 ( .A(n7298), .B(n7304), .ZN(n7299) );
  NAND2_X1 U9171 ( .A1(n7299), .A2(n9295), .ZN(n7301) );
  OR2_X1 U9172 ( .A1(n7331), .A2(n9261), .ZN(n7300) );
  NAND2_X1 U9173 ( .A1(n7301), .A2(n7300), .ZN(n9582) );
  AOI21_X1 U9174 ( .B1(n9264), .B2(n7302), .A(n9582), .ZN(n7310) );
  OAI21_X1 U9175 ( .B1(n7305), .B2(n7304), .A(n7303), .ZN(n9583) );
  NAND2_X1 U9176 ( .A1(n9583), .A2(n9545), .ZN(n7309) );
  OAI22_X1 U9177 ( .A1(n9287), .A2(n5906), .B1(n7328), .B2(n9309), .ZN(n7306)
         );
  AOI21_X1 U9178 ( .B1(n9268), .B2(n7307), .A(n7306), .ZN(n7308) );
  OAI211_X1 U9179 ( .C1(n9317), .C2(n7310), .A(n7309), .B(n7308), .ZN(P1_U3284) );
  INV_X1 U9180 ( .A(n7311), .ZN(n7313) );
  OAI22_X1 U9181 ( .A1(n7314), .A2(n7313), .B1(n8139), .B2(n7312), .ZN(n7316)
         );
  XNOR2_X1 U9182 ( .A(n7316), .B(n7315), .ZN(n7323) );
  NOR2_X1 U9183 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7317), .ZN(n9713) );
  AOI21_X1 U9184 ( .B1(n8119), .B2(n8139), .A(n9713), .ZN(n7320) );
  NAND2_X1 U9185 ( .A1(n8124), .A2(n7318), .ZN(n7319) );
  OAI211_X1 U9186 ( .C1(n7792), .C2(n8121), .A(n7320), .B(n7319), .ZN(n7321)
         );
  AOI21_X1 U9187 ( .B1(n9827), .B2(n8072), .A(n7321), .ZN(n7322) );
  OAI21_X1 U9188 ( .B1(n7323), .B2(n8052), .A(n7322), .ZN(P2_U3176) );
  AND2_X1 U9189 ( .A1(n7203), .A2(n7324), .ZN(n7327) );
  OAI211_X1 U9190 ( .C1(n7327), .C2(n7326), .A(n8603), .B(n7325), .ZN(n7335)
         );
  INV_X1 U9191 ( .A(n7328), .ZN(n7333) );
  AOI21_X1 U9192 ( .B1(n8943), .B2(n8627), .A(n7329), .ZN(n7330) );
  OAI21_X1 U9193 ( .B1(n7331), .B2(n8624), .A(n7330), .ZN(n7332) );
  AOI21_X1 U9194 ( .B1(n7333), .B2(n8607), .A(n7332), .ZN(n7334) );
  OAI211_X1 U9195 ( .C1(n4515), .C2(n8610), .A(n7335), .B(n7334), .ZN(P1_U3231) );
  INV_X1 U9196 ( .A(n7351), .ZN(n7449) );
  OAI21_X1 U9197 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7339) );
  NAND2_X1 U9198 ( .A1(n7339), .A2(n8117), .ZN(n7343) );
  AND2_X1 U9199 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9727) );
  AOI21_X1 U9200 ( .B1(n8107), .B2(n8135), .A(n9727), .ZN(n7340) );
  OAI21_X1 U9201 ( .B1(n7792), .B2(n8109), .A(n7340), .ZN(n7341) );
  AOI21_X1 U9202 ( .B1(n7453), .B2(n8124), .A(n7341), .ZN(n7342) );
  OAI211_X1 U9203 ( .C1(n7449), .C2(n8128), .A(n7343), .B(n7342), .ZN(P2_U3174) );
  INV_X1 U9204 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7346) );
  XNOR2_X1 U9205 ( .A(n7344), .B(n7898), .ZN(n7345) );
  AOI222_X1 U9206 ( .A1(n8365), .A2(n7345), .B1(n8135), .B2(n8362), .C1(n8137), 
        .C2(n8360), .ZN(n7450) );
  MUX2_X1 U9207 ( .A(n7346), .B(n7450), .S(n9829), .Z(n7349) );
  XNOR2_X1 U9208 ( .A(n7347), .B(n7898), .ZN(n7454) );
  AOI22_X1 U9209 ( .A1(n7454), .A2(n8459), .B1(n8477), .B2(n7351), .ZN(n7348)
         );
  NAND2_X1 U9210 ( .A1(n7349), .A2(n7348), .ZN(P2_U3429) );
  INV_X1 U9211 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7350) );
  MUX2_X1 U9212 ( .A(n7350), .B(n7450), .S(n9851), .Z(n7353) );
  AOI22_X1 U9213 ( .A1(n7454), .A2(n8403), .B1(n8413), .B2(n7351), .ZN(n7352)
         );
  NAND2_X1 U9214 ( .A1(n7353), .A2(n7352), .ZN(P2_U3472) );
  XNOR2_X1 U9215 ( .A(n7440), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7434) );
  XNOR2_X1 U9216 ( .A(n9532), .B(n9399), .ZN(n9521) );
  NOR2_X1 U9217 ( .A1(n7358), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7354) );
  AOI21_X1 U9218 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7358), .A(n7354), .ZN(
        n9509) );
  OAI21_X1 U9219 ( .B1(n7365), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7355), .ZN(
        n9510) );
  NOR2_X1 U9220 ( .A1(n9509), .A2(n9510), .ZN(n9508) );
  INV_X1 U9221 ( .A(n9508), .ZN(n7356) );
  OAI21_X1 U9222 ( .B1(n7358), .B2(n7357), .A(n7356), .ZN(n9520) );
  AND2_X1 U9223 ( .A1(n9532), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7359) );
  NOR2_X1 U9224 ( .A1(n9523), .A2(n7359), .ZN(n7360) );
  NOR2_X1 U9225 ( .A1(n7360), .A2(n7367), .ZN(n7361) );
  XNOR2_X1 U9226 ( .A(n7360), .B(n7367), .ZN(n9875) );
  NOR2_X1 U9227 ( .A1(n9874), .A2(n9875), .ZN(n9876) );
  NOR2_X1 U9228 ( .A1(n7361), .A2(n9876), .ZN(n7384) );
  XNOR2_X1 U9229 ( .A(n7369), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7385) );
  AOI22_X1 U9230 ( .A1(n7384), .A2(n7385), .B1(n7369), .B2(n7362), .ZN(n7435)
         );
  XOR2_X1 U9231 ( .A(n7434), .B(n7435), .Z(n7378) );
  XNOR2_X1 U9232 ( .A(n7440), .B(n9254), .ZN(n7372) );
  XNOR2_X1 U9233 ( .A(n9532), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U9234 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9516), .ZN(n7363) );
  OAI21_X1 U9235 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9516), .A(n7363), .ZN(
        n9512) );
  OAI21_X1 U9236 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7365), .A(n7364), .ZN(
        n9513) );
  NOR2_X1 U9237 ( .A1(n9512), .A2(n9513), .ZN(n9511) );
  AOI21_X1 U9238 ( .B1(n9516), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9511), .ZN(
        n9529) );
  NOR2_X1 U9239 ( .A1(n9528), .A2(n9529), .ZN(n9527) );
  AOI21_X1 U9240 ( .B1(n9532), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9527), .ZN(
        n7366) );
  NOR2_X1 U9241 ( .A1(n7366), .A2(n7367), .ZN(n7368) );
  XNOR2_X1 U9242 ( .A(n7367), .B(n7366), .ZN(n9883) );
  NOR2_X1 U9243 ( .A1(n9311), .A2(n9883), .ZN(n9882) );
  NOR2_X1 U9244 ( .A1(n7368), .A2(n9882), .ZN(n7389) );
  XNOR2_X1 U9245 ( .A(n7369), .B(n9276), .ZN(n7388) );
  NAND2_X1 U9246 ( .A1(n7392), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7370) );
  NAND2_X1 U9247 ( .A1(n7371), .A2(n7372), .ZN(n7442) );
  OAI21_X1 U9248 ( .B1(n7372), .B2(n7371), .A(n7442), .ZN(n7373) );
  NAND2_X1 U9249 ( .A1(n7373), .A2(n9885), .ZN(n7377) );
  NOR2_X1 U9250 ( .A1(n9989), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8585) );
  NOR2_X1 U9251 ( .A1(n9502), .A2(n7374), .ZN(n7375) );
  AOI211_X1 U9252 ( .C1(n8997), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n8585), .B(
        n7375), .ZN(n7376) );
  OAI211_X1 U9253 ( .C1(n9522), .C2(n7378), .A(n7377), .B(n7376), .ZN(P1_U3260) );
  INV_X1 U9254 ( .A(n7379), .ZN(n7382) );
  OAI222_X1 U9255 ( .A1(n7964), .A2(n7380), .B1(n7960), .B2(n7382), .C1(n8914), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U9256 ( .A1(n8494), .A2(n7383), .B1(n8492), .B2(n7382), .C1(n7381), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  XOR2_X1 U9257 ( .A(n7385), .B(n7384), .Z(n7394) );
  INV_X1 U9258 ( .A(n9502), .ZN(n9881) );
  NAND2_X1 U9259 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8576) );
  OAI21_X1 U9260 ( .B1(n9892), .B2(n7162), .A(n8576), .ZN(n7391) );
  INV_X1 U9261 ( .A(n9885), .ZN(n9526) );
  INV_X1 U9262 ( .A(n7386), .ZN(n7387) );
  AOI211_X1 U9263 ( .C1(n7389), .C2(n7388), .A(n9526), .B(n7387), .ZN(n7390)
         );
  AOI211_X1 U9264 ( .C1(n9881), .C2(n7392), .A(n7391), .B(n7390), .ZN(n7393)
         );
  OAI21_X1 U9265 ( .B1(n7394), .B2(n9522), .A(n7393), .ZN(P1_U3259) );
  OAI21_X1 U9266 ( .B1(n7396), .B2(n8783), .A(n7395), .ZN(n9588) );
  INV_X1 U9267 ( .A(n9588), .ZN(n7407) );
  INV_X1 U9268 ( .A(n7397), .ZN(n7398) );
  AOI21_X1 U9269 ( .B1(n8783), .B2(n7399), .A(n7398), .ZN(n7400) );
  OAI222_X1 U9270 ( .A1(n9263), .A2(n7632), .B1(n9261), .B2(n7401), .C1(n9553), 
        .C2(n7400), .ZN(n9587) );
  OAI211_X1 U9271 ( .C1(n7402), .C2(n6356), .A(n9229), .B(n7477), .ZN(n9585)
         );
  OAI22_X1 U9272 ( .A1(n9287), .A2(n5927), .B1(n7521), .B2(n9309), .ZN(n7403)
         );
  AOI21_X1 U9273 ( .B1(n7523), .B2(n9268), .A(n7403), .ZN(n7404) );
  OAI21_X1 U9274 ( .B1(n9585), .B2(n9230), .A(n7404), .ZN(n7405) );
  AOI21_X1 U9275 ( .B1(n9587), .B2(n9287), .A(n7405), .ZN(n7406) );
  OAI21_X1 U9276 ( .B1(n7407), .B2(n9290), .A(n7406), .ZN(P1_U3283) );
  INV_X1 U9277 ( .A(n7421), .ZN(n7409) );
  AOI21_X1 U9278 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9446), .A(n8915), .ZN(
        n7408) );
  OAI21_X1 U9279 ( .B1(n7409), .B2(n7960), .A(n7408), .ZN(P1_U3332) );
  INV_X1 U9280 ( .A(n7410), .ZN(n7469) );
  NOR2_X1 U9281 ( .A1(n7469), .A2(n8276), .ZN(n7416) );
  NAND2_X1 U9282 ( .A1(n7411), .A2(n7900), .ZN(n7412) );
  NAND3_X1 U9283 ( .A1(n7413), .A2(n8365), .A3(n7412), .ZN(n7415) );
  AOI22_X1 U9284 ( .A1(n8136), .A2(n8360), .B1(n8362), .B2(n8361), .ZN(n7414)
         );
  NAND2_X1 U9285 ( .A1(n7415), .A2(n7414), .ZN(n7427) );
  AOI211_X1 U9286 ( .C1(n8368), .C2(n7466), .A(n7416), .B(n7427), .ZN(n7420)
         );
  XNOR2_X1 U9287 ( .A(n7417), .B(n7900), .ZN(n7428) );
  INV_X1 U9288 ( .A(n7428), .ZN(n7418) );
  AOI22_X1 U9289 ( .A1(n7418), .A2(n8333), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8336), .ZN(n7419) );
  OAI21_X1 U9290 ( .B1(n7420), .B2(n8336), .A(n7419), .ZN(P2_U3219) );
  NAND2_X1 U9291 ( .A1(n7421), .A2(n7677), .ZN(n7423) );
  OR2_X1 U9292 ( .A1(n7422), .A2(P2_U3151), .ZN(n7933) );
  OAI211_X1 U9293 ( .C1(n7424), .C2(n8494), .A(n7423), .B(n7933), .ZN(P2_U3272) );
  MUX2_X1 U9294 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n7427), .S(n9851), .Z(n7426)
         );
  OAI22_X1 U9295 ( .A1(n7428), .A2(n8416), .B1(n7469), .B2(n8386), .ZN(n7425)
         );
  OR2_X1 U9296 ( .A1(n7426), .A2(n7425), .ZN(P2_U3473) );
  MUX2_X1 U9297 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n7427), .S(n9829), .Z(n7430)
         );
  OAI22_X1 U9298 ( .A1(n7428), .A2(n8481), .B1(n7469), .B2(n8428), .ZN(n7429)
         );
  OR2_X1 U9299 ( .A1(n7430), .A2(n7429), .ZN(P2_U3432) );
  INV_X1 U9300 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n7433) );
  NOR2_X1 U9301 ( .A1(n7431), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8626) );
  INV_X1 U9302 ( .A(n8626), .ZN(n7432) );
  OAI21_X1 U9303 ( .B1(n9892), .B2(n7433), .A(n7432), .ZN(n7439) );
  NAND2_X1 U9304 ( .A1(n7443), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9034) );
  OAI21_X1 U9305 ( .B1(n7443), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9034), .ZN(
        n7437) );
  OAI22_X1 U9306 ( .A1(n7435), .A2(n7434), .B1(n7440), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n7436) );
  NOR2_X1 U9307 ( .A1(n7436), .A2(n7437), .ZN(n9036) );
  AOI211_X1 U9308 ( .C1(n7437), .C2(n7436), .A(n9522), .B(n9036), .ZN(n7438)
         );
  AOI211_X1 U9309 ( .C1(n9881), .C2(n7443), .A(n7439), .B(n7438), .ZN(n7448)
         );
  OR2_X1 U9310 ( .A1(n7440), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9311 ( .A1(n7443), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9038) );
  OR2_X1 U9312 ( .A1(n7443), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7444) );
  AND2_X1 U9313 ( .A1(n9038), .A2(n7444), .ZN(n7445) );
  NAND2_X1 U9314 ( .A1(n7446), .A2(n7445), .ZN(n9039) );
  OAI211_X1 U9315 ( .C1(n7446), .C2(n7445), .A(n9039), .B(n9885), .ZN(n7447)
         );
  NAND2_X1 U9316 ( .A1(n7448), .A2(n7447), .ZN(P1_U3261) );
  NOR2_X1 U9317 ( .A1(n7449), .A2(n8276), .ZN(n7452) );
  INV_X1 U9318 ( .A(n7450), .ZN(n7451) );
  AOI211_X1 U9319 ( .C1(n8368), .C2(n7453), .A(n7452), .B(n7451), .ZN(n7456)
         );
  AOI22_X1 U9320 ( .A1(n7454), .A2(n8333), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8336), .ZN(n7455) );
  OAI21_X1 U9321 ( .B1(n7456), .B2(n8336), .A(n7455), .ZN(P2_U3220) );
  INV_X1 U9322 ( .A(n7336), .ZN(n7459) );
  NOR3_X1 U9323 ( .A1(n7459), .A2(n7458), .A3(n7457), .ZN(n7462) );
  INV_X1 U9324 ( .A(n7460), .ZN(n7461) );
  OAI21_X1 U9325 ( .B1(n7462), .B2(n7461), .A(n8117), .ZN(n7468) );
  AND2_X1 U9326 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9742) );
  AOI21_X1 U9327 ( .B1(n8107), .B2(n8361), .A(n9742), .ZN(n7463) );
  OAI21_X1 U9328 ( .B1(n7464), .B2(n8109), .A(n7463), .ZN(n7465) );
  AOI21_X1 U9329 ( .B1(n7466), .B2(n8124), .A(n7465), .ZN(n7467) );
  OAI211_X1 U9330 ( .C1(n7469), .C2(n8128), .A(n7468), .B(n7467), .ZN(P2_U3155) );
  INV_X1 U9331 ( .A(n8798), .ZN(n7470) );
  XNOR2_X1 U9332 ( .A(n7471), .B(n7470), .ZN(n7474) );
  NAND2_X1 U9333 ( .A1(n8942), .A2(n9299), .ZN(n7472) );
  OAI21_X1 U9334 ( .B1(n7600), .B2(n9261), .A(n7472), .ZN(n7473) );
  AOI21_X1 U9335 ( .B1(n7474), .B2(n9295), .A(n7473), .ZN(n9591) );
  XNOR2_X1 U9336 ( .A(n7475), .B(n8798), .ZN(n9596) );
  NAND2_X1 U9337 ( .A1(n9596), .A2(n9545), .ZN(n7482) );
  OAI22_X1 U9338 ( .A1(n9287), .A2(n7476), .B1(n7603), .B2(n9309), .ZN(n7480)
         );
  INV_X1 U9339 ( .A(n7477), .ZN(n7478) );
  OAI211_X1 U9340 ( .C1(n7478), .C2(n9593), .A(n9229), .B(n7534), .ZN(n9590)
         );
  NOR2_X1 U9341 ( .A1(n9590), .A2(n9230), .ZN(n7479) );
  AOI211_X1 U9342 ( .C1(n9268), .C2(n7605), .A(n7480), .B(n7479), .ZN(n7481)
         );
  OAI211_X1 U9343 ( .C1(n9317), .C2(n9591), .A(n7482), .B(n7481), .ZN(P1_U3282) );
  INV_X1 U9344 ( .A(n8356), .ZN(n7485) );
  XNOR2_X1 U9345 ( .A(n7483), .B(n7899), .ZN(n7497) );
  INV_X1 U9346 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7488) );
  XNOR2_X1 U9347 ( .A(n7486), .B(n7899), .ZN(n7487) );
  AOI222_X1 U9348 ( .A1(n8365), .A2(n7487), .B1(n8135), .B2(n8360), .C1(n8349), 
        .C2(n8362), .ZN(n7494) );
  MUX2_X1 U9349 ( .A(n7488), .B(n7494), .S(n9829), .Z(n7490) );
  NAND2_X1 U9350 ( .A1(n7498), .A2(n8477), .ZN(n7489) );
  OAI211_X1 U9351 ( .C1(n7497), .C2(n8481), .A(n7490), .B(n7489), .ZN(P2_U3435) );
  INV_X1 U9352 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7491) );
  MUX2_X1 U9353 ( .A(n7491), .B(n7494), .S(n9851), .Z(n7493) );
  NAND2_X1 U9354 ( .A1(n7498), .A2(n8413), .ZN(n7492) );
  OAI211_X1 U9355 ( .C1(n8416), .C2(n7497), .A(n7493), .B(n7492), .ZN(P2_U3474) );
  INV_X1 U9356 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7545) );
  MUX2_X1 U9357 ( .A(n7545), .B(n7494), .S(n8366), .Z(n7496) );
  AOI22_X1 U9358 ( .A1(n7498), .A2(n8369), .B1(n8368), .B2(n7506), .ZN(n7495)
         );
  OAI211_X1 U9359 ( .C1(n7497), .C2(n8372), .A(n7496), .B(n7495), .ZN(P2_U3218) );
  INV_X1 U9360 ( .A(n7498), .ZN(n7509) );
  AOI21_X1 U9361 ( .B1(n7500), .B2(n7499), .A(n8052), .ZN(n7502) );
  NAND2_X1 U9362 ( .A1(n7502), .A2(n7501), .ZN(n7508) );
  AND2_X1 U9363 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7554) );
  AOI21_X1 U9364 ( .B1(n8107), .B2(n8349), .A(n7554), .ZN(n7503) );
  OAI21_X1 U9365 ( .B1(n7504), .B2(n8109), .A(n7503), .ZN(n7505) );
  AOI21_X1 U9366 ( .B1(n7506), .B2(n8124), .A(n7505), .ZN(n7507) );
  OAI211_X1 U9367 ( .C1(n7509), .C2(n8128), .A(n7508), .B(n7507), .ZN(P2_U3181) );
  INV_X1 U9368 ( .A(n7510), .ZN(n7514) );
  OAI222_X1 U9369 ( .A1(n7512), .A2(P1_U3086), .B1(n7960), .B2(n7514), .C1(
        n7511), .C2(n7964), .ZN(P1_U3331) );
  OAI222_X1 U9370 ( .A1(n8494), .A2(n7515), .B1(n8492), .B2(n7514), .C1(n7513), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  AOI21_X1 U9371 ( .B1(n7517), .B2(n7516), .A(n4346), .ZN(n7525) );
  NAND2_X1 U9372 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9459) );
  INV_X1 U9373 ( .A(n9459), .ZN(n7519) );
  NOR2_X1 U9374 ( .A1(n7632), .A2(n8638), .ZN(n7518) );
  AOI211_X1 U9375 ( .C1(n8636), .C2(n4514), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI21_X1 U9376 ( .B1(n8635), .B2(n7521), .A(n7520), .ZN(n7522) );
  AOI21_X1 U9377 ( .B1(n7523), .B2(n8641), .A(n7522), .ZN(n7524) );
  OAI21_X1 U9378 ( .B1(n7525), .B2(n8643), .A(n7524), .ZN(P1_U3217) );
  NAND2_X1 U9379 ( .A1(n7526), .A2(n8706), .ZN(n7527) );
  XNOR2_X1 U9380 ( .A(n7527), .B(n8801), .ZN(n7528) );
  NAND2_X1 U9381 ( .A1(n7528), .A2(n9295), .ZN(n7532) );
  OAI22_X1 U9382 ( .A1(n7632), .A2(n9261), .B1(n7529), .B2(n9263), .ZN(n7530)
         );
  INV_X1 U9383 ( .A(n7530), .ZN(n7531) );
  NAND2_X1 U9384 ( .A1(n7532), .A2(n7531), .ZN(n7573) );
  INV_X1 U9385 ( .A(n7573), .ZN(n7540) );
  XNOR2_X1 U9386 ( .A(n7533), .B(n8801), .ZN(n7575) );
  NAND2_X1 U9387 ( .A1(n7575), .A2(n9545), .ZN(n7539) );
  AOI211_X1 U9388 ( .C1(n7637), .C2(n7534), .A(n9306), .B(n7619), .ZN(n7574)
         );
  NOR2_X1 U9389 ( .A1(n7577), .A2(n9542), .ZN(n7537) );
  OAI22_X1 U9390 ( .A1(n9287), .A2(n7535), .B1(n7635), .B2(n9309), .ZN(n7536)
         );
  AOI211_X1 U9391 ( .C1(n7574), .C2(n4265), .A(n7537), .B(n7536), .ZN(n7538)
         );
  OAI211_X1 U9392 ( .C1(n9317), .C2(n7540), .A(n7539), .B(n7538), .ZN(P1_U3281) );
  INV_X1 U9393 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9753) );
  NAND2_X1 U9394 ( .A1(n9754), .A2(n9753), .ZN(n9752) );
  OAI21_X1 U9395 ( .B1(n7548), .B2(n7236), .A(n7541), .ZN(n7542) );
  NAND2_X1 U9396 ( .A1(n9741), .A2(n7542), .ZN(n7543) );
  AOI21_X1 U9397 ( .B1(n7545), .B2(n7544), .A(n8152), .ZN(n7572) );
  XNOR2_X1 U9398 ( .A(n9754), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U9399 ( .A1(n9741), .A2(n7550), .ZN(n7551) );
  NAND2_X1 U9400 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9731), .ZN(n9730) );
  NAND2_X1 U9401 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7552), .ZN(n8158) );
  OAI21_X1 U9402 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n7552), .A(n8158), .ZN(
        n7570) );
  NOR2_X1 U9403 ( .A1(n9766), .A2(n8166), .ZN(n7553) );
  AOI211_X1 U9404 ( .C1(n9743), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7554), .B(
        n7553), .ZN(n7568) );
  XNOR2_X1 U9405 ( .A(n8167), .B(n8151), .ZN(n7565) );
  OR2_X1 U9406 ( .A1(n7555), .A2(n9765), .ZN(n7563) );
  XNOR2_X1 U9407 ( .A(n7555), .B(n9754), .ZN(n9749) );
  OR2_X1 U9408 ( .A1(n7557), .A2(n9741), .ZN(n7562) );
  XNOR2_X1 U9409 ( .A(n7557), .B(n7556), .ZN(n9734) );
  OR2_X1 U9410 ( .A1(n7559), .A2(n7558), .ZN(n7561) );
  NAND2_X1 U9411 ( .A1(n7561), .A2(n7560), .ZN(n9733) );
  NAND2_X1 U9412 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  NAND2_X1 U9413 ( .A1(n7562), .A2(n9732), .ZN(n9748) );
  NAND2_X1 U9414 ( .A1(n9749), .A2(n9748), .ZN(n9747) );
  NAND2_X1 U9415 ( .A1(n7563), .A2(n9747), .ZN(n7564) );
  NAND2_X1 U9416 ( .A1(n7565), .A2(n7564), .ZN(n8165) );
  OAI21_X1 U9417 ( .B1(n7565), .B2(n7564), .A(n8165), .ZN(n7566) );
  NAND2_X1 U9418 ( .A1(n7566), .A2(n9750), .ZN(n7567) );
  NAND2_X1 U9419 ( .A1(n7568), .A2(n7567), .ZN(n7569) );
  AOI21_X1 U9420 ( .B1(n7570), .B2(n9762), .A(n7569), .ZN(n7571) );
  OAI21_X1 U9421 ( .B1(n7572), .B2(n9755), .A(n7571), .ZN(P2_U3197) );
  AOI211_X1 U9422 ( .C1(n7575), .C2(n9595), .A(n7574), .B(n7573), .ZN(n7581)
         );
  INV_X1 U9423 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7576) );
  OAI22_X1 U9424 ( .A1(n7577), .A2(n9440), .B1(n9598), .B2(n7576), .ZN(n7578)
         );
  INV_X1 U9425 ( .A(n7578), .ZN(n7579) );
  OAI21_X1 U9426 ( .B1(n7581), .B2(n9589), .A(n7579), .ZN(P1_U3489) );
  AOI22_X1 U9427 ( .A1(n7637), .A2(n7673), .B1(n9605), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7580) );
  OAI21_X1 U9428 ( .B1(n7581), .B2(n9605), .A(n7580), .ZN(P1_U3534) );
  XNOR2_X1 U9429 ( .A(n7583), .B(n7582), .ZN(n7588) );
  NAND2_X1 U9430 ( .A1(n8119), .A2(n8361), .ZN(n7584) );
  NAND2_X1 U9431 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8170) );
  OAI211_X1 U9432 ( .C1(n8121), .C2(n8110), .A(n7584), .B(n8170), .ZN(n7585)
         );
  AOI21_X1 U9433 ( .B1(n8367), .B2(n8124), .A(n7585), .ZN(n7587) );
  NAND2_X1 U9434 ( .A1(n8478), .A2(n8072), .ZN(n7586) );
  OAI211_X1 U9435 ( .C1(n7588), .C2(n8052), .A(n7587), .B(n7586), .ZN(P2_U3166) );
  INV_X1 U9436 ( .A(n7589), .ZN(n7593) );
  OAI222_X1 U9437 ( .A1(n7591), .A2(P1_U3086), .B1(n7960), .B2(n7593), .C1(
        n7590), .C2(n7964), .ZN(P1_U3330) );
  OAI222_X1 U9438 ( .A1(n8494), .A2(n7594), .B1(n8492), .B2(n7593), .C1(n7592), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  NAND2_X1 U9439 ( .A1(n7595), .A2(n7596), .ZN(n7628) );
  INV_X1 U9440 ( .A(n7628), .ZN(n7598) );
  AOI21_X1 U9441 ( .B1(n7596), .B2(n7627), .A(n7595), .ZN(n7597) );
  AOI21_X1 U9442 ( .B1(n7598), .B2(n7627), .A(n7597), .ZN(n7607) );
  NOR2_X1 U9443 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7599), .ZN(n9504) );
  NOR2_X1 U9444 ( .A1(n7600), .A2(n8624), .ZN(n7601) );
  AOI211_X1 U9445 ( .C1(n8627), .C2(n8942), .A(n9504), .B(n7601), .ZN(n7602)
         );
  OAI21_X1 U9446 ( .B1(n8635), .B2(n7603), .A(n7602), .ZN(n7604) );
  AOI21_X1 U9447 ( .B1(n7605), .B2(n8641), .A(n7604), .ZN(n7606) );
  OAI21_X1 U9448 ( .B1(n7607), .B2(n8643), .A(n7606), .ZN(P1_U3236) );
  INV_X1 U9449 ( .A(n7608), .ZN(n7611) );
  OAI222_X1 U9450 ( .A1(n8494), .A2(n7610), .B1(n8492), .B2(n7611), .C1(n7609), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  OAI222_X1 U9451 ( .A1(n7612), .A2(P1_U3086), .B1(n7960), .B2(n7611), .C1(
        n9964), .C2(n7964), .ZN(P1_U3329) );
  INV_X1 U9452 ( .A(n7663), .ZN(n7617) );
  INV_X1 U9453 ( .A(n7642), .ZN(n7613) );
  AOI21_X1 U9454 ( .B1(n8803), .B2(n7614), .A(n7613), .ZN(n7615) );
  OAI222_X1 U9455 ( .A1(n9261), .A2(n7616), .B1(n9263), .B2(n7660), .C1(n9553), 
        .C2(n7615), .ZN(n7668) );
  AOI21_X1 U9456 ( .B1(n7617), .B2(n9538), .A(n7668), .ZN(n7626) );
  XOR2_X1 U9457 ( .A(n7618), .B(n8803), .Z(n7670) );
  NAND2_X1 U9458 ( .A1(n7670), .A2(n9545), .ZN(n7625) );
  INV_X1 U9459 ( .A(n7619), .ZN(n7620) );
  AOI211_X1 U9460 ( .C1(n7674), .C2(n7620), .A(n9306), .B(n7648), .ZN(n7669)
         );
  OAI22_X1 U9461 ( .A1(n7622), .A2(n9542), .B1(n7621), .B2(n9287), .ZN(n7623)
         );
  AOI21_X1 U9462 ( .B1(n7669), .B2(n4265), .A(n7623), .ZN(n7624) );
  OAI211_X1 U9463 ( .C1(n9317), .C2(n7626), .A(n7625), .B(n7624), .ZN(P1_U3280) );
  NAND2_X1 U9464 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  XOR2_X1 U9465 ( .A(n7630), .B(n7629), .Z(n7639) );
  OAI21_X1 U9466 ( .B1(n7632), .B2(n8624), .A(n7631), .ZN(n7633) );
  AOI21_X1 U9467 ( .B1(n8627), .B2(n8941), .A(n7633), .ZN(n7634) );
  OAI21_X1 U9468 ( .B1(n8635), .B2(n7635), .A(n7634), .ZN(n7636) );
  AOI21_X1 U9469 ( .B1(n7637), .B2(n8641), .A(n7636), .ZN(n7638) );
  OAI21_X1 U9470 ( .B1(n7639), .B2(n8643), .A(n7638), .ZN(P1_U3224) );
  INV_X1 U9471 ( .A(n7640), .ZN(n7667) );
  XNOR2_X1 U9472 ( .A(n7641), .B(n7643), .ZN(n9398) );
  INV_X1 U9473 ( .A(n9398), .ZN(n7656) );
  NAND2_X1 U9474 ( .A1(n7642), .A2(n8719), .ZN(n7644) );
  INV_X1 U9475 ( .A(n7643), .ZN(n8805) );
  XNOR2_X1 U9476 ( .A(n7644), .B(n8805), .ZN(n7645) );
  NAND2_X1 U9477 ( .A1(n7645), .A2(n9295), .ZN(n7647) );
  AOI22_X1 U9478 ( .A1(n8941), .A2(n9298), .B1(n9299), .B2(n9282), .ZN(n7646)
         );
  NAND2_X1 U9479 ( .A1(n7647), .A2(n7646), .ZN(n9396) );
  INV_X1 U9480 ( .A(n7648), .ZN(n7649) );
  AOI211_X1 U9481 ( .C1(n7650), .C2(n7649), .A(n9306), .B(n4487), .ZN(n9397)
         );
  NAND2_X1 U9482 ( .A1(n9397), .A2(n4265), .ZN(n7653) );
  INV_X1 U9483 ( .A(n7651), .ZN(n8507) );
  AOI22_X1 U9484 ( .A1(n9317), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8507), .B2(
        n9538), .ZN(n7652) );
  OAI211_X1 U9485 ( .C1(n9441), .C2(n9542), .A(n7653), .B(n7652), .ZN(n7654)
         );
  AOI21_X1 U9486 ( .B1(n9287), .B2(n9396), .A(n7654), .ZN(n7655) );
  OAI21_X1 U9487 ( .B1(n7656), .B2(n9290), .A(n7655), .ZN(P1_U3279) );
  XOR2_X1 U9488 ( .A(n7658), .B(n7657), .Z(n7666) );
  OAI22_X1 U9489 ( .A1(n7660), .A2(n8638), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7659), .ZN(n7661) );
  AOI21_X1 U9490 ( .B1(n8636), .B2(n8942), .A(n7661), .ZN(n7662) );
  OAI21_X1 U9491 ( .B1(n8635), .B2(n7663), .A(n7662), .ZN(n7664) );
  AOI21_X1 U9492 ( .B1(n7674), .B2(n8641), .A(n7664), .ZN(n7665) );
  OAI21_X1 U9493 ( .B1(n7666), .B2(n8643), .A(n7665), .ZN(P1_U3234) );
  AOI211_X1 U9494 ( .C1(n7670), .C2(n9595), .A(n7669), .B(n7668), .ZN(n7676)
         );
  AOI22_X1 U9495 ( .A1(n7674), .A2(n7671), .B1(n9589), .B2(
        P1_REG0_REG_13__SCAN_IN), .ZN(n7672) );
  OAI21_X1 U9496 ( .B1(n7676), .B2(n9589), .A(n7672), .ZN(P1_U3492) );
  AOI22_X1 U9497 ( .A1(n7674), .A2(n7673), .B1(n9605), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7675) );
  OAI21_X1 U9498 ( .B1(n7676), .B2(n9605), .A(n7675), .ZN(P1_U3535) );
  NAND2_X1 U9499 ( .A1(n7961), .A2(n7677), .ZN(n7679) );
  OAI211_X1 U9500 ( .C1(n8494), .C2(n7680), .A(n7679), .B(n7678), .ZN(P2_U3267) );
  NOR2_X1 U9501 ( .A1(n7681), .A2(n7903), .ZN(n7683) );
  AOI22_X1 U9502 ( .A1(n8313), .A2(n8362), .B1(n8360), .B2(n8350), .ZN(n7684)
         );
  NAND2_X1 U9503 ( .A1(n7685), .A2(n7684), .ZN(n8456) );
  MUX2_X1 U9504 ( .A(n8456), .B(P2_REG2_REG_19__SCAN_IN), .S(n8336), .Z(n7690)
         );
  INV_X1 U9505 ( .A(n7903), .ZN(n7686) );
  XNOR2_X1 U9506 ( .A(n8323), .B(n7686), .ZN(n8460) );
  NAND2_X1 U9507 ( .A1(n8460), .A2(n8333), .ZN(n7688) );
  AOI22_X1 U9508 ( .A1(n8458), .A2(n8369), .B1(n8368), .B2(n7941), .ZN(n7687)
         );
  NAND2_X1 U9509 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  OR2_X1 U9510 ( .A1(n7690), .A2(n7689), .ZN(P2_U3214) );
  INV_X1 U9511 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U9512 ( .A1(n7832), .A2(n8282), .ZN(n7907) );
  XOR2_X1 U9513 ( .A(n7691), .B(n7907), .Z(n8294) );
  XOR2_X1 U9514 ( .A(n7907), .B(n7692), .Z(n7693) );
  OAI222_X1 U9515 ( .A1(n8300), .A2(n8266), .B1(n8302), .B2(n7694), .C1(n9768), 
        .C2(n7693), .ZN(n8289) );
  AOI21_X1 U9516 ( .B1(n9808), .B2(n8294), .A(n8289), .ZN(n7697) );
  MUX2_X1 U9517 ( .A(n7695), .B(n7697), .S(n9851), .Z(n7696) );
  OAI21_X1 U9518 ( .B1(n8292), .B2(n8386), .A(n7696), .ZN(P2_U3482) );
  INV_X1 U9519 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n7698) );
  MUX2_X1 U9520 ( .A(n7698), .B(n7697), .S(n9829), .Z(n7699) );
  OAI21_X1 U9521 ( .B1(n8292), .B2(n8428), .A(n7699), .ZN(P2_U3450) );
  AOI22_X1 U9522 ( .A1(n8117), .A2(n7883), .B1(n9771), .B2(n8072), .ZN(n7702)
         );
  NAND2_X1 U9523 ( .A1(n7700), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7701) );
  OAI211_X1 U9524 ( .C1(n7703), .C2(n8121), .A(n7702), .B(n7701), .ZN(P2_U3172) );
  INV_X1 U9525 ( .A(n7856), .ZN(n7704) );
  INV_X1 U9526 ( .A(SI_29_), .ZN(n7706) );
  INV_X1 U9527 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8489) );
  INV_X1 U9528 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7712) );
  MUX2_X1 U9529 ( .A(n8489), .B(n7712), .S(n7731), .Z(n7714) );
  INV_X1 U9530 ( .A(SI_30_), .ZN(n7713) );
  NAND2_X1 U9531 ( .A1(n7714), .A2(n7713), .ZN(n7728) );
  INV_X1 U9532 ( .A(n7714), .ZN(n7715) );
  NAND2_X1 U9533 ( .A1(n7715), .A2(SI_30_), .ZN(n7716) );
  NAND2_X1 U9534 ( .A1(n7728), .A2(n7716), .ZN(n7729) );
  NAND2_X1 U9535 ( .A1(n8765), .A2(n7739), .ZN(n7718) );
  OR2_X1 U9536 ( .A1(n7737), .A2(n8489), .ZN(n7717) );
  INV_X1 U9537 ( .A(n8129), .ZN(n7858) );
  NAND2_X1 U9538 ( .A1(n8424), .A2(n7858), .ZN(n7912) );
  NAND2_X1 U9539 ( .A1(n7912), .A2(n7719), .ZN(n7864) );
  INV_X1 U9540 ( .A(n7864), .ZN(n7720) );
  NAND2_X1 U9541 ( .A1(n7721), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U9542 ( .A1(n5164), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U9543 ( .A1(n5408), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7722) );
  AND3_X1 U9544 ( .A1(n7724), .A2(n7723), .A3(n7722), .ZN(n7725) );
  NAND2_X1 U9545 ( .A1(n7726), .A2(n7725), .ZN(n8250) );
  OR2_X1 U9546 ( .A1(n8424), .A2(n8250), .ZN(n7727) );
  INV_X1 U9547 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7736) );
  INV_X1 U9548 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7732) );
  MUX2_X1 U9549 ( .A(n7736), .B(n7732), .S(n7731), .Z(n7733) );
  XNOR2_X1 U9550 ( .A(n7733), .B(SI_31_), .ZN(n7734) );
  NOR2_X1 U9551 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  OR2_X1 U9552 ( .A1(n8424), .A2(n7858), .ZN(n7913) );
  INV_X1 U9553 ( .A(n7873), .ZN(n7740) );
  INV_X1 U9554 ( .A(n8374), .ZN(n8420) );
  INV_X1 U9555 ( .A(n8250), .ZN(n7741) );
  NOR2_X1 U9556 ( .A1(n7919), .A2(n7742), .ZN(n7872) );
  INV_X1 U9557 ( .A(n7743), .ZN(n7871) );
  NAND2_X1 U9558 ( .A1(n7764), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U9559 ( .A1(n8147), .A2(n9773), .ZN(n7750) );
  NAND2_X1 U9560 ( .A1(n7758), .A2(n7750), .ZN(n7751) );
  MUX2_X1 U9561 ( .A(n7752), .B(n7751), .S(n7865), .Z(n7753) );
  INV_X1 U9562 ( .A(n7756), .ZN(n7757) );
  NAND2_X1 U9563 ( .A1(n7766), .A2(n7759), .ZN(n7762) );
  INV_X1 U9564 ( .A(n7761), .ZN(n7763) );
  INV_X1 U9565 ( .A(n7768), .ZN(n7890) );
  NAND2_X1 U9566 ( .A1(n7773), .A2(n7769), .ZN(n7771) );
  OAI21_X1 U9567 ( .B1(n9798), .B2(n8142), .A(n7772), .ZN(n7770) );
  MUX2_X1 U9568 ( .A(n7771), .B(n7770), .S(n7865), .Z(n7775) );
  MUX2_X1 U9569 ( .A(n7773), .B(n7772), .S(n7857), .Z(n7774) );
  INV_X1 U9570 ( .A(n7778), .ZN(n7779) );
  OR2_X1 U9571 ( .A1(n7785), .A2(n7779), .ZN(n7782) );
  OAI21_X1 U9572 ( .B1(n9810), .B2(n8140), .A(n7780), .ZN(n7781) );
  MUX2_X1 U9573 ( .A(n7782), .B(n7781), .S(n7865), .Z(n7783) );
  INV_X1 U9574 ( .A(n7784), .ZN(n7786) );
  NOR2_X1 U9575 ( .A1(n7790), .A2(n7857), .ZN(n7794) );
  NOR2_X1 U9576 ( .A1(n7791), .A2(n7865), .ZN(n7793) );
  MUX2_X1 U9577 ( .A(n7794), .B(n7793), .S(n7792), .Z(n7795) );
  MUX2_X1 U9578 ( .A(n7798), .B(n7797), .S(n7857), .Z(n7799) );
  MUX2_X1 U9579 ( .A(n7801), .B(n7800), .S(n7865), .Z(n7802) );
  NAND2_X1 U9580 ( .A1(n7812), .A2(n7803), .ZN(n7806) );
  NAND2_X1 U9581 ( .A1(n8359), .A2(n7804), .ZN(n7805) );
  MUX2_X1 U9582 ( .A(n7806), .B(n7805), .S(n7857), .Z(n7807) );
  INV_X1 U9583 ( .A(n7807), .ZN(n7808) );
  NAND2_X1 U9584 ( .A1(n7813), .A2(n7878), .ZN(n7815) );
  OAI21_X1 U9585 ( .B1(n7816), .B2(n7815), .A(n7814), .ZN(n7817) );
  NAND2_X1 U9586 ( .A1(n7823), .A2(n7818), .ZN(n7821) );
  NAND2_X1 U9587 ( .A1(n7822), .A2(n7819), .ZN(n7820) );
  MUX2_X1 U9588 ( .A(n7821), .B(n7820), .S(n7865), .Z(n7825) );
  MUX2_X1 U9589 ( .A(n7823), .B(n7822), .S(n7857), .Z(n7824) );
  AND2_X1 U9590 ( .A1(n8282), .A2(n7826), .ZN(n7827) );
  INV_X1 U9591 ( .A(n7877), .ZN(n7830) );
  AOI21_X1 U9592 ( .B1(n7834), .B2(n7831), .A(n7830), .ZN(n7836) );
  MUX2_X1 U9593 ( .A(n7838), .B(n7837), .S(n7865), .Z(n7839) );
  INV_X1 U9594 ( .A(n7844), .ZN(n7841) );
  INV_X1 U9595 ( .A(n7842), .ZN(n7843) );
  MUX2_X1 U9596 ( .A(n7844), .B(n7843), .S(n7865), .Z(n7845) );
  NAND2_X1 U9597 ( .A1(n7847), .A2(n7848), .ZN(n7967) );
  MUX2_X1 U9598 ( .A(n7848), .B(n7847), .S(n7857), .Z(n7849) );
  INV_X1 U9599 ( .A(n7849), .ZN(n7851) );
  MUX2_X1 U9600 ( .A(n8130), .B(n8260), .S(n7857), .Z(n7853) );
  OAI21_X1 U9601 ( .B1(n7858), .B2(n7857), .A(n8424), .ZN(n7859) );
  INV_X1 U9602 ( .A(n7859), .ZN(n7861) );
  NOR2_X1 U9603 ( .A1(n8129), .A2(n7865), .ZN(n7860) );
  NAND2_X1 U9604 ( .A1(n7863), .A2(n7862), .ZN(n7870) );
  OAI21_X1 U9605 ( .B1(n7868), .B2(n8130), .A(n7867), .ZN(n7869) );
  NOR2_X1 U9606 ( .A1(n8243), .A2(n7873), .ZN(n7874) );
  NAND2_X1 U9607 ( .A1(n7875), .A2(n7874), .ZN(n7925) );
  INV_X1 U9608 ( .A(n7967), .ZN(n7965) );
  NAND2_X1 U9609 ( .A1(n7877), .A2(n7876), .ZN(n8284) );
  INV_X1 U9610 ( .A(n8310), .ZN(n7905) );
  INV_X1 U9611 ( .A(n8320), .ZN(n8326) );
  NAND2_X1 U9612 ( .A1(n7879), .A2(n7878), .ZN(n8338) );
  NOR2_X1 U9613 ( .A1(n7881), .A2(n7880), .ZN(n7887) );
  NOR2_X1 U9614 ( .A1(n7883), .A2(n7882), .ZN(n7886) );
  NAND4_X1 U9615 ( .A1(n7887), .A2(n7886), .A3(n7885), .A4(n7884), .ZN(n7891)
         );
  NOR4_X1 U9616 ( .A1(n7891), .A2(n7890), .A3(n7889), .A4(n7888), .ZN(n7895)
         );
  NAND4_X1 U9617 ( .A1(n7895), .A2(n7894), .A3(n7893), .A4(n7892), .ZN(n7896)
         );
  NAND4_X1 U9618 ( .A1(n8359), .A2(n7900), .A3(n4857), .A4(n7899), .ZN(n7901)
         );
  OR3_X1 U9619 ( .A1(n8338), .A2(n8347), .A3(n7901), .ZN(n7902) );
  NOR2_X1 U9620 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NAND4_X1 U9621 ( .A1(n8304), .A2(n7905), .A3(n8326), .A4(n7904), .ZN(n7906)
         );
  OR3_X1 U9622 ( .A1(n8284), .A2(n7907), .A3(n7906), .ZN(n7908) );
  NOR2_X1 U9623 ( .A1(n8271), .A2(n7908), .ZN(n7909) );
  NAND3_X1 U9624 ( .A1(n7965), .A2(n7983), .A3(n7909), .ZN(n7910) );
  NOR2_X1 U9625 ( .A1(n7911), .A2(n7910), .ZN(n7914) );
  AND4_X1 U9626 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n7916)
         );
  NAND2_X1 U9627 ( .A1(n7916), .A2(n4344), .ZN(n7920) );
  NAND3_X1 U9628 ( .A1(n7920), .A2(n8243), .A3(n7917), .ZN(n7922) );
  OR4_X1 U9629 ( .A1(n7920), .A2(n7919), .A3(n8243), .A4(n7918), .ZN(n7921) );
  OAI211_X1 U9630 ( .C1(n7875), .C2(n5487), .A(n7922), .B(n7921), .ZN(n7923)
         );
  INV_X1 U9631 ( .A(n7923), .ZN(n7924) );
  OAI21_X1 U9632 ( .B1(n7926), .B2(n7925), .A(n7924), .ZN(n7927) );
  NOR3_X1 U9633 ( .A1(n7929), .A2(n8236), .A3(n7928), .ZN(n7932) );
  OAI21_X1 U9634 ( .B1(n7933), .B2(n7930), .A(P2_B_REG_SCAN_IN), .ZN(n7931) );
  INV_X1 U9635 ( .A(n8765), .ZN(n8490) );
  AOI22_X1 U9636 ( .A1(n7934), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9446), .ZN(n7935) );
  OAI21_X1 U9637 ( .B1(n8490), .B2(n7960), .A(n7935), .ZN(P1_U3325) );
  INV_X1 U9638 ( .A(n8458), .ZN(n7944) );
  AOI21_X1 U9639 ( .B1(n7936), .B2(n7937), .A(n8052), .ZN(n7938) );
  NAND2_X1 U9640 ( .A1(n7938), .A2(n8081), .ZN(n7943) );
  AND2_X1 U9641 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8242) );
  AOI21_X1 U9642 ( .B1(n8107), .B2(n8313), .A(n8242), .ZN(n7939) );
  OAI21_X1 U9643 ( .B1(n5577), .B2(n8109), .A(n7939), .ZN(n7940) );
  AOI21_X1 U9644 ( .B1(n7941), .B2(n8124), .A(n7940), .ZN(n7942) );
  OAI211_X1 U9645 ( .C1(n7944), .C2(n8128), .A(n7943), .B(n7942), .ZN(P2_U3159) );
  INV_X1 U9646 ( .A(n7945), .ZN(n7955) );
  OAI21_X1 U9647 ( .B1(n7946), .B2(n7948), .A(n7947), .ZN(n7949) );
  NAND2_X1 U9648 ( .A1(n7949), .A2(n8603), .ZN(n7954) );
  OAI22_X1 U9649 ( .A1(n7950), .A2(n8624), .B1(n6822), .B2(n8638), .ZN(n7951)
         );
  AOI21_X1 U9650 ( .B1(n7952), .B2(n8641), .A(n7951), .ZN(n7953) );
  OAI211_X1 U9651 ( .C1(n7955), .C2(n8947), .A(n7954), .B(n7953), .ZN(P1_U3222) );
  OAI222_X1 U9652 ( .A1(n8494), .A2(n7957), .B1(n8492), .B2(n7956), .C1(
        P2_U3151), .C2(n5487), .ZN(P2_U3276) );
  INV_X1 U9653 ( .A(n7958), .ZN(n8493) );
  OAI222_X1 U9654 ( .A1(n7960), .A2(n8493), .B1(n7964), .B2(n6322), .C1(n7959), 
        .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U9655 ( .A(n7961), .ZN(n7962) );
  OAI222_X1 U9656 ( .A1(n7964), .A2(n7963), .B1(P1_U3086), .B2(n6280), .C1(
        n7960), .C2(n7962), .ZN(P1_U3327) );
  XNOR2_X1 U9657 ( .A(n7966), .B(n7965), .ZN(n7981) );
  XNOR2_X1 U9658 ( .A(n7968), .B(n7967), .ZN(n7969) );
  AOI222_X1 U9659 ( .A1(n8365), .A2(n7969), .B1(n8132), .B2(n8360), .C1(n8130), 
        .C2(n8362), .ZN(n7976) );
  MUX2_X1 U9660 ( .A(n7970), .B(n7976), .S(n9829), .Z(n7972) );
  NAND2_X1 U9661 ( .A1(n7978), .A2(n8477), .ZN(n7971) );
  OAI211_X1 U9662 ( .C1(n7981), .C2(n8481), .A(n7972), .B(n7971), .ZN(P2_U3454) );
  INV_X1 U9663 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7973) );
  MUX2_X1 U9664 ( .A(n7973), .B(n7976), .S(n9851), .Z(n7975) );
  NAND2_X1 U9665 ( .A1(n7978), .A2(n8413), .ZN(n7974) );
  OAI211_X1 U9666 ( .C1(n7981), .C2(n8416), .A(n7975), .B(n7974), .ZN(P2_U3486) );
  INV_X1 U9667 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7977) );
  MUX2_X1 U9668 ( .A(n7977), .B(n7976), .S(n8366), .Z(n7980) );
  AOI22_X1 U9669 ( .A1(n7978), .A2(n8369), .B1(n8368), .B2(n8008), .ZN(n7979)
         );
  OAI211_X1 U9670 ( .C1(n7981), .C2(n8372), .A(n7980), .B(n7979), .ZN(P2_U3206) );
  XOR2_X1 U9671 ( .A(n7982), .B(n7983), .Z(n8380) );
  XOR2_X1 U9672 ( .A(n7984), .B(n7983), .Z(n7985) );
  OAI222_X1 U9673 ( .A1(n8300), .A2(n8122), .B1(n8302), .B2(n8279), .C1(n9768), 
        .C2(n7985), .ZN(n8378) );
  INV_X1 U9674 ( .A(n8378), .ZN(n7989) );
  MUX2_X1 U9675 ( .A(n7986), .B(n7989), .S(n9829), .Z(n7988) );
  NAND2_X1 U9676 ( .A1(n7991), .A2(n8477), .ZN(n7987) );
  OAI211_X1 U9677 ( .C1(n8380), .C2(n8481), .A(n7988), .B(n7987), .ZN(P2_U3453) );
  INV_X1 U9678 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7990) );
  MUX2_X1 U9679 ( .A(n7990), .B(n7989), .S(n8366), .Z(n7993) );
  AOI22_X1 U9680 ( .A1(n7991), .A2(n8369), .B1(n8368), .B2(n8125), .ZN(n7992)
         );
  OAI211_X1 U9681 ( .C1(n8380), .C2(n8372), .A(n7993), .B(n7992), .ZN(P2_U3207) );
  INV_X1 U9682 ( .A(n7995), .ZN(n8002) );
  NOR2_X1 U9683 ( .A1(n7997), .A2(n7996), .ZN(n8251) );
  AOI21_X1 U9684 ( .B1(n8336), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8251), .ZN(
        n7998) );
  OAI21_X1 U9685 ( .B1(n7999), .B2(n8330), .A(n7998), .ZN(n8000) );
  AOI21_X1 U9686 ( .B1(n8002), .B2(n8001), .A(n8000), .ZN(n8003) );
  OAI21_X1 U9687 ( .B1(n7994), .B2(n8336), .A(n8003), .ZN(P2_U3204) );
  AOI21_X1 U9688 ( .B1(n8005), .B2(n8004), .A(n8052), .ZN(n8007) );
  NAND2_X1 U9689 ( .A1(n8007), .A2(n8006), .ZN(n8014) );
  INV_X1 U9690 ( .A(n8008), .ZN(n8011) );
  AOI22_X1 U9691 ( .A1(n8132), .A2(n8119), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8009) );
  OAI21_X1 U9692 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8012) );
  AOI21_X1 U9693 ( .B1(n8107), .B2(n8130), .A(n8012), .ZN(n8013) );
  OAI211_X1 U9694 ( .C1(n8015), .C2(n8128), .A(n8014), .B(n8013), .ZN(P2_U3154) );
  INV_X1 U9695 ( .A(n8017), .ZN(n8057) );
  AOI21_X1 U9696 ( .B1(n8134), .B2(n8016), .A(n8057), .ZN(n8023) );
  AOI22_X1 U9697 ( .A1(n8312), .A2(n8119), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8019) );
  NAND2_X1 U9698 ( .A1(n8124), .A2(n8290), .ZN(n8018) );
  OAI211_X1 U9699 ( .C1(n8266), .C2(n8121), .A(n8019), .B(n8018), .ZN(n8020)
         );
  AOI21_X1 U9700 ( .B1(n8021), .B2(n8072), .A(n8020), .ZN(n8022) );
  OAI21_X1 U9701 ( .B1(n8023), .B2(n8052), .A(n8022), .ZN(P2_U3156) );
  INV_X1 U9702 ( .A(n8024), .ZN(n8083) );
  NOR3_X1 U9703 ( .A1(n8083), .A2(n8026), .A3(n8025), .ZN(n8027) );
  OAI21_X1 U9704 ( .B1(n8027), .B2(n4342), .A(n8117), .ZN(n8032) );
  AOI22_X1 U9705 ( .A1(n8107), .A2(n8312), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8028) );
  OAI21_X1 U9706 ( .B1(n8029), .B2(n8109), .A(n8028), .ZN(n8030) );
  AOI21_X1 U9707 ( .B1(n8316), .B2(n8124), .A(n8030), .ZN(n8031) );
  OAI211_X1 U9708 ( .C1(n8033), .C2(n8128), .A(n8032), .B(n8031), .ZN(P2_U3163) );
  INV_X1 U9709 ( .A(n8034), .ZN(n8058) );
  INV_X1 U9710 ( .A(n8035), .ZN(n8037) );
  NOR3_X1 U9711 ( .A1(n8058), .A2(n8037), .A3(n8036), .ZN(n8040) );
  INV_X1 U9712 ( .A(n8038), .ZN(n8039) );
  OAI21_X1 U9713 ( .B1(n8040), .B2(n8039), .A(n8117), .ZN(n8044) );
  AOI22_X1 U9714 ( .A1(n8132), .A2(n8107), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8041) );
  OAI21_X1 U9715 ( .B1(n8266), .B2(n8109), .A(n8041), .ZN(n8042) );
  AOI21_X1 U9716 ( .B1(n8270), .B2(n8124), .A(n8042), .ZN(n8043) );
  OAI211_X1 U9717 ( .C1(n8429), .C2(n8128), .A(n8044), .B(n8043), .ZN(P2_U3165) );
  OR2_X1 U9718 ( .A1(n8045), .A2(n8047), .ZN(n8046) );
  INV_X1 U9719 ( .A(n8046), .ZN(n8102) );
  AOI21_X1 U9720 ( .B1(n8047), .B2(n8045), .A(n8102), .ZN(n8053) );
  NAND2_X1 U9721 ( .A1(n8119), .A2(n8349), .ZN(n8048) );
  NAND2_X1 U9722 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8190) );
  OAI211_X1 U9723 ( .C1(n8121), .C2(n5577), .A(n8048), .B(n8190), .ZN(n8049)
         );
  AOI21_X1 U9724 ( .B1(n8352), .B2(n8124), .A(n8049), .ZN(n8051) );
  NAND2_X1 U9725 ( .A1(n8471), .A2(n8072), .ZN(n8050) );
  OAI211_X1 U9726 ( .C1(n8053), .C2(n8052), .A(n8051), .B(n8050), .ZN(P2_U3168) );
  INV_X1 U9727 ( .A(n8054), .ZN(n8056) );
  NOR3_X1 U9728 ( .A1(n8057), .A2(n8056), .A3(n8055), .ZN(n8059) );
  OAI21_X1 U9729 ( .B1(n8059), .B2(n8058), .A(n8117), .ZN(n8063) );
  AOI22_X1 U9730 ( .A1(n4749), .A2(n8107), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8060) );
  OAI21_X1 U9731 ( .B1(n8299), .B2(n8109), .A(n8060), .ZN(n8061) );
  AOI21_X1 U9732 ( .B1(n8281), .B2(n8124), .A(n8061), .ZN(n8062) );
  OAI211_X1 U9733 ( .C1(n8387), .C2(n8128), .A(n8063), .B(n8062), .ZN(P2_U3169) );
  OAI211_X1 U9734 ( .C1(n8066), .C2(n8065), .A(n8064), .B(n8117), .ZN(n8078)
         );
  NAND2_X1 U9735 ( .A1(n8119), .A2(n8141), .ZN(n8069) );
  NOR2_X1 U9736 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8067), .ZN(n9682) );
  INV_X1 U9737 ( .A(n9682), .ZN(n8068) );
  OAI211_X1 U9738 ( .C1(n8121), .C2(n8070), .A(n8069), .B(n8068), .ZN(n8071)
         );
  INV_X1 U9739 ( .A(n8071), .ZN(n8077) );
  NAND2_X1 U9740 ( .A1(n8073), .A2(n8072), .ZN(n8076) );
  NAND2_X1 U9741 ( .A1(n8124), .A2(n8074), .ZN(n8075) );
  NAND4_X1 U9742 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(
        P2_U3171) );
  INV_X1 U9743 ( .A(n8399), .ZN(n8331) );
  AOI21_X1 U9744 ( .B1(n8081), .B2(n8080), .A(n8079), .ZN(n8082) );
  OAI21_X1 U9745 ( .B1(n8083), .B2(n8082), .A(n8117), .ZN(n8088) );
  AOI22_X1 U9746 ( .A1(n8107), .A2(n5351), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8084) );
  OAI21_X1 U9747 ( .B1(n8085), .B2(n8109), .A(n8084), .ZN(n8086) );
  AOI21_X1 U9748 ( .B1(n8328), .B2(n8124), .A(n8086), .ZN(n8087) );
  OAI211_X1 U9749 ( .C1(n8331), .C2(n8128), .A(n8088), .B(n8087), .ZN(P2_U3173) );
  INV_X1 U9750 ( .A(n8442), .ZN(n8098) );
  NOR3_X1 U9751 ( .A1(n4342), .A2(n4777), .A3(n8090), .ZN(n8093) );
  INV_X1 U9752 ( .A(n8091), .ZN(n8092) );
  OAI21_X1 U9753 ( .B1(n8093), .B2(n8092), .A(n8117), .ZN(n8097) );
  AOI22_X1 U9754 ( .A1(n8119), .A2(n5351), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8094) );
  OAI21_X1 U9755 ( .B1(n8299), .B2(n8121), .A(n8094), .ZN(n8095) );
  AOI21_X1 U9756 ( .B1(n8303), .B2(n8124), .A(n8095), .ZN(n8096) );
  OAI211_X1 U9757 ( .C1(n8098), .C2(n8128), .A(n8097), .B(n8096), .ZN(P2_U3175) );
  INV_X1 U9758 ( .A(n8465), .ZN(n8114) );
  INV_X1 U9759 ( .A(n8099), .ZN(n8101) );
  NOR3_X1 U9760 ( .A1(n8102), .A2(n8101), .A3(n8100), .ZN(n8106) );
  OR2_X1 U9761 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  OAI21_X1 U9762 ( .B1(n8106), .B2(n8105), .A(n8117), .ZN(n8113) );
  AND2_X1 U9763 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8219) );
  AOI21_X1 U9764 ( .B1(n8107), .B2(n8340), .A(n8219), .ZN(n8108) );
  OAI21_X1 U9765 ( .B1(n8110), .B2(n8109), .A(n8108), .ZN(n8111) );
  AOI21_X1 U9766 ( .B1(n8343), .B2(n8124), .A(n8111), .ZN(n8112) );
  OAI211_X1 U9767 ( .C1(n8114), .C2(n8128), .A(n8113), .B(n8112), .ZN(P2_U3178) );
  OAI21_X1 U9768 ( .B1(n8267), .B2(n8116), .A(n8115), .ZN(n8118) );
  NAND2_X1 U9769 ( .A1(n8118), .A2(n8117), .ZN(n8127) );
  AOI22_X1 U9770 ( .A1(n4749), .A2(n8119), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8120) );
  OAI21_X1 U9771 ( .B1(n8122), .B2(n8121), .A(n8120), .ZN(n8123) );
  AOI21_X1 U9772 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8126) );
  OAI211_X1 U9773 ( .C1(n8379), .C2(n8128), .A(n8127), .B(n8126), .ZN(P2_U3180) );
  MUX2_X1 U9774 ( .A(n8250), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8215), .Z(
        P2_U3522) );
  MUX2_X1 U9775 ( .A(n8129), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8215), .Z(
        P2_U3521) );
  MUX2_X1 U9776 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8130), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9777 ( .A(n8131), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8215), .Z(
        P2_U3518) );
  MUX2_X1 U9778 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8132), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9779 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n4749), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9780 ( .A(n8133), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8215), .Z(
        P2_U3515) );
  MUX2_X1 U9781 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8134), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9782 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8312), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9783 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n5351), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9784 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8313), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9785 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8340), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9786 ( .A(n8350), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8215), .Z(
        P2_U3509) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8363), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8349), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9789 ( .A(n8361), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8215), .Z(
        P2_U3506) );
  MUX2_X1 U9790 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8135), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9791 ( .A(n8136), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8215), .Z(
        P2_U3504) );
  MUX2_X1 U9792 ( .A(n8137), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8215), .Z(
        P2_U3503) );
  MUX2_X1 U9793 ( .A(n8138), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8215), .Z(
        P2_U3502) );
  MUX2_X1 U9794 ( .A(n8139), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8215), .Z(
        P2_U3501) );
  MUX2_X1 U9795 ( .A(n8140), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8215), .Z(
        P2_U3500) );
  MUX2_X1 U9796 ( .A(n8141), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8215), .Z(
        P2_U3499) );
  MUX2_X1 U9797 ( .A(n8142), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8215), .Z(
        P2_U3498) );
  MUX2_X1 U9798 ( .A(n8143), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8215), .Z(
        P2_U3497) );
  MUX2_X1 U9799 ( .A(n8144), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8215), .Z(
        P2_U3496) );
  MUX2_X1 U9800 ( .A(n8145), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8215), .Z(
        P2_U3495) );
  MUX2_X1 U9801 ( .A(n8146), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8215), .Z(
        P2_U3494) );
  MUX2_X1 U9802 ( .A(n8147), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8215), .Z(
        P2_U3493) );
  MUX2_X1 U9803 ( .A(n8148), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8215), .Z(
        P2_U3492) );
  MUX2_X1 U9804 ( .A(n8149), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8215), .Z(
        P2_U3491) );
  NOR2_X1 U9805 ( .A1(n8151), .A2(n8150), .ZN(n8153) );
  INV_X1 U9806 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8154) );
  AOI22_X1 U9807 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8181), .B1(n8178), .B2(
        n8154), .ZN(n8155) );
  AOI21_X1 U9808 ( .B1(n8156), .B2(n8155), .A(n8177), .ZN(n8176) );
  INV_X1 U9809 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8412) );
  AOI22_X1 U9810 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8178), .B1(n8181), .B2(
        n8412), .ZN(n8161) );
  NAND2_X1 U9811 ( .A1(n8166), .A2(n8157), .ZN(n8159) );
  OAI21_X1 U9812 ( .B1(n8161), .B2(n8160), .A(n8180), .ZN(n8174) );
  NOR2_X1 U9813 ( .A1(n9664), .A2(n8162), .ZN(n8173) );
  NOR2_X1 U9814 ( .A1(n8163), .A2(n8178), .ZN(n8183) );
  INV_X1 U9815 ( .A(n8183), .ZN(n8164) );
  NAND2_X1 U9816 ( .A1(n8163), .A2(n8178), .ZN(n8184) );
  NAND2_X1 U9817 ( .A1(n8164), .A2(n8184), .ZN(n8169) );
  OAI21_X1 U9818 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8185) );
  NAND2_X1 U9819 ( .A1(n8185), .A2(n8169), .ZN(n8168) );
  OAI211_X1 U9820 ( .C1(n8169), .C2(n8185), .A(n9750), .B(n8168), .ZN(n8171)
         );
  OAI211_X1 U9821 ( .C1(n9766), .C2(n8178), .A(n8171), .B(n8170), .ZN(n8172)
         );
  AOI211_X1 U9822 ( .C1(n8174), .C2(n9762), .A(n8173), .B(n8172), .ZN(n8175)
         );
  OAI21_X1 U9823 ( .B1(n8176), .B2(n9755), .A(n8175), .ZN(P2_U3198) );
  INV_X1 U9824 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9908) );
  XNOR2_X1 U9825 ( .A(n8198), .B(n8210), .ZN(n8179) );
  NOR2_X1 U9826 ( .A1(n9908), .A2(n8179), .ZN(n8199) );
  AOI21_X1 U9827 ( .B1(n9908), .B2(n8179), .A(n8199), .ZN(n8196) );
  NAND2_X1 U9828 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8182), .ZN(n8205) );
  OAI21_X1 U9829 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8182), .A(n8205), .ZN(
        n8194) );
  XNOR2_X1 U9830 ( .A(n8207), .B(n8204), .ZN(n8187) );
  AOI21_X1 U9831 ( .B1(n8185), .B2(n8184), .A(n8183), .ZN(n8186) );
  NOR2_X1 U9832 ( .A1(n8186), .A2(n8187), .ZN(n8208) );
  AOI21_X1 U9833 ( .B1(n8187), .B2(n8186), .A(n8208), .ZN(n8188) );
  NOR2_X1 U9834 ( .A1(n8188), .A2(n9622), .ZN(n8193) );
  NAND2_X1 U9835 ( .A1(n9696), .A2(n8210), .ZN(n8189) );
  OAI211_X1 U9836 ( .C1(n9664), .C2(n8191), .A(n8190), .B(n8189), .ZN(n8192)
         );
  AOI211_X1 U9837 ( .C1(n8194), .C2(n9762), .A(n8193), .B(n8192), .ZN(n8195)
         );
  OAI21_X1 U9838 ( .B1(n8196), .B2(n9755), .A(n8195), .ZN(P2_U3199) );
  NOR2_X1 U9839 ( .A1(n8220), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8197) );
  AOI21_X1 U9840 ( .B1(n8220), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8197), .ZN(
        n8202) );
  NOR2_X1 U9841 ( .A1(n8210), .A2(n8198), .ZN(n8200) );
  AOI21_X1 U9842 ( .B1(n8202), .B2(n8201), .A(n4337), .ZN(n8228) );
  NAND2_X1 U9843 ( .A1(n8204), .A2(n8203), .ZN(n8206) );
  NAND2_X1 U9844 ( .A1(n8206), .A2(n8205), .ZN(n8232) );
  XNOR2_X1 U9845 ( .A(n8220), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8231) );
  XNOR2_X1 U9846 ( .A(n8232), .B(n8231), .ZN(n8226) );
  INV_X1 U9847 ( .A(n8207), .ZN(n8209) );
  AOI21_X1 U9848 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8211) );
  NAND2_X1 U9849 ( .A1(n8211), .A2(n8212), .ZN(n8216) );
  NAND2_X1 U9850 ( .A1(n8216), .A2(n8220), .ZN(n8235) );
  INV_X1 U9851 ( .A(n8211), .ZN(n8214) );
  INV_X1 U9852 ( .A(n8212), .ZN(n8213) );
  NAND2_X1 U9853 ( .A1(n8214), .A2(n8213), .ZN(n8234) );
  INV_X1 U9854 ( .A(n8234), .ZN(n8217) );
  NOR3_X1 U9855 ( .A1(n8235), .A2(n8217), .A3(n8215), .ZN(n8225) );
  INV_X1 U9856 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8223) );
  INV_X1 U9857 ( .A(n8216), .ZN(n8218) );
  OAI211_X1 U9858 ( .C1(n8218), .C2(n8217), .A(n9750), .B(n8230), .ZN(n8222)
         );
  AOI21_X1 U9859 ( .B1(n9696), .B2(n8220), .A(n8219), .ZN(n8221) );
  OAI211_X1 U9860 ( .C1(n8223), .C2(n9664), .A(n8222), .B(n8221), .ZN(n8224)
         );
  AOI211_X1 U9861 ( .C1(n8226), .C2(n9762), .A(n8225), .B(n8224), .ZN(n8227)
         );
  OAI21_X1 U9862 ( .B1(n8228), .B2(n9755), .A(n8227), .ZN(P2_U3200) );
  INV_X1 U9863 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8229) );
  MUX2_X1 U9864 ( .A(n8229), .B(P2_REG2_REG_19__SCAN_IN), .S(n5487), .Z(n8237)
         );
  AOI22_X1 U9865 ( .A1(n8232), .A2(n8231), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8230), .ZN(n8233) );
  XNOR2_X1 U9866 ( .A(n5487), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8238) );
  XNOR2_X1 U9867 ( .A(n8233), .B(n8238), .ZN(n8247) );
  NAND2_X1 U9868 ( .A1(n8235), .A2(n8234), .ZN(n8240) );
  MUX2_X1 U9869 ( .A(n8238), .B(n8237), .S(n4433), .Z(n8239) );
  XNOR2_X1 U9870 ( .A(n8240), .B(n8239), .ZN(n8241) );
  NOR2_X1 U9871 ( .A1(n8241), .A2(n9622), .ZN(n8246) );
  AOI21_X1 U9872 ( .B1(n9696), .B2(n8243), .A(n8242), .ZN(n8244) );
  OAI21_X1 U9873 ( .B1(n9664), .B2(n4523), .A(n8244), .ZN(n8245) );
  AOI211_X1 U9874 ( .C1(n8247), .C2(n9762), .A(n8246), .B(n8245), .ZN(n8248)
         );
  AOI21_X1 U9875 ( .B1(n8421), .B2(n8366), .A(n8251), .ZN(n8254) );
  NAND2_X1 U9876 ( .A1(n8336), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8252) );
  OAI211_X1 U9877 ( .C1(n8374), .C2(n8330), .A(n8254), .B(n8252), .ZN(P2_U3202) );
  INV_X1 U9878 ( .A(n8424), .ZN(n8377) );
  NAND2_X1 U9879 ( .A1(n8336), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8253) );
  OAI211_X1 U9880 ( .C1(n8377), .C2(n8330), .A(n8254), .B(n8253), .ZN(P2_U3203) );
  OR2_X1 U9881 ( .A1(n8255), .A2(n8336), .ZN(n8258) );
  INV_X1 U9882 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U9883 ( .A1(n8336), .A2(n8256), .ZN(n8257) );
  NAND2_X1 U9884 ( .A1(n8258), .A2(n8257), .ZN(n8262) );
  AOI22_X1 U9885 ( .A1(n8260), .A2(n8369), .B1(n8368), .B2(n8259), .ZN(n8261)
         );
  OAI211_X1 U9886 ( .C1(n8263), .C2(n8372), .A(n8262), .B(n8261), .ZN(P2_U3205) );
  XOR2_X1 U9887 ( .A(n8271), .B(n8264), .Z(n8265) );
  OAI222_X1 U9888 ( .A1(n8300), .A2(n8267), .B1(n8302), .B2(n8266), .C1(n9768), 
        .C2(n8265), .ZN(n8427) );
  AOI21_X1 U9889 ( .B1(n8269), .B2(n8268), .A(n8427), .ZN(n8275) );
  AOI22_X1 U9890 ( .A1(n8270), .A2(n8368), .B1(n8336), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8274) );
  XNOR2_X1 U9891 ( .A(n8272), .B(n8271), .ZN(n8383) );
  NAND2_X1 U9892 ( .A1(n8383), .A2(n8333), .ZN(n8273) );
  OAI211_X1 U9893 ( .C1(n8275), .C2(n8336), .A(n8274), .B(n8273), .ZN(P2_U3208) );
  NOR2_X1 U9894 ( .A1(n8387), .A2(n8276), .ZN(n8280) );
  XOR2_X1 U9895 ( .A(n8284), .B(n8277), .Z(n8278) );
  OAI222_X1 U9896 ( .A1(n8302), .A2(n8299), .B1(n8300), .B2(n8279), .C1(n8278), 
        .C2(n9768), .ZN(n8433) );
  AOI211_X1 U9897 ( .C1(n8368), .C2(n8281), .A(n8280), .B(n8433), .ZN(n8288)
         );
  NAND2_X1 U9898 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  XNOR2_X1 U9899 ( .A(n8285), .B(n8284), .ZN(n8439) );
  INV_X1 U9900 ( .A(n8439), .ZN(n8286) );
  AOI22_X1 U9901 ( .A1(n8286), .A2(n8333), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8336), .ZN(n8287) );
  OAI21_X1 U9902 ( .B1(n8288), .B2(n8336), .A(n8287), .ZN(P2_U3209) );
  INV_X1 U9903 ( .A(n8289), .ZN(n8296) );
  AOI22_X1 U9904 ( .A1(n8336), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8290), .B2(
        n8368), .ZN(n8291) );
  OAI21_X1 U9905 ( .B1(n8292), .B2(n8330), .A(n8291), .ZN(n8293) );
  AOI21_X1 U9906 ( .B1(n8294), .B2(n8333), .A(n8293), .ZN(n8295) );
  OAI21_X1 U9907 ( .B1(n8296), .B2(n8336), .A(n8295), .ZN(P2_U3210) );
  XOR2_X1 U9908 ( .A(n8297), .B(n8304), .Z(n8298) );
  OAI222_X1 U9909 ( .A1(n8302), .A2(n8301), .B1(n8300), .B2(n8299), .C1(n9768), 
        .C2(n8298), .ZN(n8390) );
  AOI21_X1 U9910 ( .B1(n8368), .B2(n8303), .A(n8390), .ZN(n8308) );
  AOI22_X1 U9911 ( .A1(n8442), .A2(n8369), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n8336), .ZN(n8307) );
  XNOR2_X1 U9912 ( .A(n8305), .B(n4712), .ZN(n8443) );
  NAND2_X1 U9913 ( .A1(n8443), .A2(n8333), .ZN(n8306) );
  OAI211_X1 U9914 ( .C1(n8308), .C2(n8336), .A(n8307), .B(n8306), .ZN(P2_U3211) );
  XNOR2_X1 U9915 ( .A(n8309), .B(n8310), .ZN(n8451) );
  INV_X1 U9916 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8315) );
  XNOR2_X1 U9917 ( .A(n8311), .B(n8310), .ZN(n8314) );
  AOI222_X1 U9918 ( .A1(n8365), .A2(n8314), .B1(n8313), .B2(n8360), .C1(n8312), 
        .C2(n8362), .ZN(n8446) );
  MUX2_X1 U9919 ( .A(n8315), .B(n8446), .S(n8366), .Z(n8318) );
  AOI22_X1 U9920 ( .A1(n8448), .A2(n8369), .B1(n8368), .B2(n8316), .ZN(n8317)
         );
  OAI211_X1 U9921 ( .C1(n8451), .C2(n8372), .A(n8318), .B(n8317), .ZN(P2_U3212) );
  OAI21_X1 U9922 ( .B1(n8321), .B2(n8320), .A(n8319), .ZN(n8322) );
  AOI222_X1 U9923 ( .A1(n8365), .A2(n8322), .B1(n5351), .B2(n8362), .C1(n8340), 
        .C2(n8360), .ZN(n8397) );
  OR2_X1 U9924 ( .A1(n8323), .A2(n4586), .ZN(n8325) );
  NAND2_X1 U9925 ( .A1(n8325), .A2(n8324), .ZN(n8327) );
  XNOR2_X1 U9926 ( .A(n8327), .B(n8326), .ZN(n8455) );
  INV_X1 U9927 ( .A(n8455), .ZN(n8334) );
  AOI22_X1 U9928 ( .A1(n8336), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8368), .B2(
        n8328), .ZN(n8329) );
  OAI21_X1 U9929 ( .B1(n8331), .B2(n8330), .A(n8329), .ZN(n8332) );
  AOI21_X1 U9930 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8335) );
  OAI21_X1 U9931 ( .B1(n8397), .B2(n8336), .A(n8335), .ZN(P2_U3213) );
  XNOR2_X1 U9932 ( .A(n8337), .B(n8338), .ZN(n8468) );
  INV_X1 U9933 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8342) );
  XNOR2_X1 U9934 ( .A(n8339), .B(n8338), .ZN(n8341) );
  AOI222_X1 U9935 ( .A1(n8365), .A2(n8341), .B1(n8340), .B2(n8362), .C1(n8363), 
        .C2(n8360), .ZN(n8463) );
  MUX2_X1 U9936 ( .A(n8342), .B(n8463), .S(n8366), .Z(n8345) );
  AOI22_X1 U9937 ( .A1(n8465), .A2(n8369), .B1(n8368), .B2(n8343), .ZN(n8344)
         );
  OAI211_X1 U9938 ( .C1(n8468), .C2(n8372), .A(n8345), .B(n8344), .ZN(P2_U3215) );
  XOR2_X1 U9939 ( .A(n8346), .B(n8347), .Z(n8474) );
  XOR2_X1 U9940 ( .A(n8348), .B(n8347), .Z(n8351) );
  AOI222_X1 U9941 ( .A1(n8365), .A2(n8351), .B1(n8350), .B2(n8362), .C1(n8349), 
        .C2(n8360), .ZN(n8469) );
  MUX2_X1 U9942 ( .A(n9908), .B(n8469), .S(n8366), .Z(n8354) );
  AOI22_X1 U9943 ( .A1(n8471), .A2(n8369), .B1(n8368), .B2(n8352), .ZN(n8353)
         );
  OAI211_X1 U9944 ( .C1(n8474), .C2(n8372), .A(n8354), .B(n8353), .ZN(P2_U3216) );
  XNOR2_X1 U9945 ( .A(n8355), .B(n8359), .ZN(n8482) );
  NAND2_X1 U9946 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  XOR2_X1 U9947 ( .A(n8359), .B(n8358), .Z(n8364) );
  AOI222_X1 U9948 ( .A1(n8365), .A2(n8364), .B1(n8363), .B2(n8362), .C1(n8361), 
        .C2(n8360), .ZN(n8475) );
  MUX2_X1 U9949 ( .A(n8154), .B(n8475), .S(n8366), .Z(n8371) );
  AOI22_X1 U9950 ( .A1(n8478), .A2(n8369), .B1(n8368), .B2(n8367), .ZN(n8370)
         );
  OAI211_X1 U9951 ( .C1(n8482), .C2(n8372), .A(n8371), .B(n8370), .ZN(P2_U3217) );
  NAND2_X1 U9952 ( .A1(n9848), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U9953 ( .A1(n8421), .A2(n9851), .ZN(n8376) );
  OAI211_X1 U9954 ( .C1(n8374), .C2(n8386), .A(n8373), .B(n8376), .ZN(P2_U3490) );
  NAND2_X1 U9955 ( .A1(n9848), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8375) );
  OAI211_X1 U9956 ( .C1(n8377), .C2(n8386), .A(n8376), .B(n8375), .ZN(P2_U3489) );
  MUX2_X1 U9957 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8378), .S(n9851), .Z(n8382)
         );
  OAI22_X1 U9958 ( .A1(n8380), .A2(n8416), .B1(n8379), .B2(n8386), .ZN(n8381)
         );
  OR2_X1 U9959 ( .A1(n8382), .A2(n8381), .ZN(P2_U3485) );
  MUX2_X1 U9960 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8427), .S(n9851), .Z(n8385)
         );
  INV_X1 U9961 ( .A(n8383), .ZN(n8430) );
  OAI22_X1 U9962 ( .A1(n8430), .A2(n8416), .B1(n8429), .B2(n8386), .ZN(n8384)
         );
  OR2_X1 U9963 ( .A1(n8385), .A2(n8384), .ZN(P2_U3484) );
  MUX2_X1 U9964 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8433), .S(n9851), .Z(n8389)
         );
  OAI22_X1 U9965 ( .A1(n8439), .A2(n8416), .B1(n8387), .B2(n8386), .ZN(n8388)
         );
  OR2_X1 U9966 ( .A1(n8389), .A2(n8388), .ZN(P2_U3483) );
  INV_X1 U9967 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8391) );
  INV_X1 U9968 ( .A(n8390), .ZN(n8440) );
  MUX2_X1 U9969 ( .A(n8391), .B(n8440), .S(n9851), .Z(n8393) );
  AOI22_X1 U9970 ( .A1(n8443), .A2(n8403), .B1(n8413), .B2(n8442), .ZN(n8392)
         );
  NAND2_X1 U9971 ( .A1(n8393), .A2(n8392), .ZN(P2_U3481) );
  INV_X1 U9972 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8394) );
  MUX2_X1 U9973 ( .A(n8394), .B(n8446), .S(n9851), .Z(n8396) );
  NAND2_X1 U9974 ( .A1(n8448), .A2(n8413), .ZN(n8395) );
  OAI211_X1 U9975 ( .C1(n8416), .C2(n8451), .A(n8396), .B(n8395), .ZN(P2_U3480) );
  INV_X1 U9976 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8400) );
  INV_X1 U9977 ( .A(n8397), .ZN(n8398) );
  AOI21_X1 U9978 ( .B1(n9828), .B2(n8399), .A(n8398), .ZN(n8452) );
  MUX2_X1 U9979 ( .A(n8400), .B(n8452), .S(n9851), .Z(n8401) );
  OAI21_X1 U9980 ( .B1(n8455), .B2(n8416), .A(n8401), .ZN(P2_U3479) );
  MUX2_X1 U9981 ( .A(n8456), .B(P2_REG1_REG_19__SCAN_IN), .S(n9848), .Z(n8402)
         );
  INV_X1 U9982 ( .A(n8402), .ZN(n8405) );
  AOI22_X1 U9983 ( .A1(n8460), .A2(n8403), .B1(n8413), .B2(n8458), .ZN(n8404)
         );
  NAND2_X1 U9984 ( .A1(n8405), .A2(n8404), .ZN(P2_U3478) );
  INV_X1 U9985 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8406) );
  MUX2_X1 U9986 ( .A(n8406), .B(n8463), .S(n9851), .Z(n8408) );
  NAND2_X1 U9987 ( .A1(n8465), .A2(n8413), .ZN(n8407) );
  OAI211_X1 U9988 ( .C1(n8416), .C2(n8468), .A(n8408), .B(n8407), .ZN(P2_U3477) );
  INV_X1 U9989 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8409) );
  MUX2_X1 U9990 ( .A(n8409), .B(n8469), .S(n9851), .Z(n8411) );
  NAND2_X1 U9991 ( .A1(n8471), .A2(n8413), .ZN(n8410) );
  OAI211_X1 U9992 ( .C1(n8474), .C2(n8416), .A(n8411), .B(n8410), .ZN(P2_U3476) );
  MUX2_X1 U9993 ( .A(n8412), .B(n8475), .S(n9851), .Z(n8415) );
  NAND2_X1 U9994 ( .A1(n8478), .A2(n8413), .ZN(n8414) );
  OAI211_X1 U9995 ( .C1(n8482), .C2(n8416), .A(n8415), .B(n8414), .ZN(P2_U3475) );
  INV_X1 U9996 ( .A(n9818), .ZN(n9812) );
  AOI22_X1 U9997 ( .A1(n8417), .A2(n9812), .B1(n5536), .B2(n9828), .ZN(n8418)
         );
  NAND2_X1 U9998 ( .A1(n8419), .A2(n8418), .ZN(n8483) );
  MUX2_X1 U9999 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8483), .S(n9851), .Z(
        P2_U3460) );
  INV_X1 U10000 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10001 ( .A1(n8420), .A2(n8477), .ZN(n8422) );
  NAND2_X1 U10002 ( .A1(n8421), .A2(n9829), .ZN(n8425) );
  OAI211_X1 U10003 ( .C1(n8423), .C2(n9829), .A(n8422), .B(n8425), .ZN(
        P2_U3458) );
  NAND2_X1 U10004 ( .A1(n8424), .A2(n8477), .ZN(n8426) );
  OAI211_X1 U10005 ( .C1(n6334), .C2(n9829), .A(n8426), .B(n8425), .ZN(
        P2_U3457) );
  MUX2_X1 U10006 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8427), .S(n9829), .Z(n8432) );
  OAI22_X1 U10007 ( .A1(n8430), .A2(n8481), .B1(n8429), .B2(n8428), .ZN(n8431)
         );
  OR2_X1 U10008 ( .A1(n8432), .A2(n8431), .ZN(P2_U3452) );
  INV_X1 U10009 ( .A(n8433), .ZN(n8434) );
  MUX2_X1 U10010 ( .A(n8435), .B(n8434), .S(n9829), .Z(n8438) );
  NAND2_X1 U10011 ( .A1(n8436), .A2(n8477), .ZN(n8437) );
  OAI211_X1 U10012 ( .C1(n8439), .C2(n8481), .A(n8438), .B(n8437), .ZN(
        P2_U3451) );
  INV_X1 U10013 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8441) );
  MUX2_X1 U10014 ( .A(n8441), .B(n8440), .S(n9829), .Z(n8445) );
  AOI22_X1 U10015 ( .A1(n8443), .A2(n8459), .B1(n8477), .B2(n8442), .ZN(n8444)
         );
  NAND2_X1 U10016 ( .A1(n8445), .A2(n8444), .ZN(P2_U3449) );
  INV_X1 U10017 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8447) );
  MUX2_X1 U10018 ( .A(n8447), .B(n8446), .S(n9829), .Z(n8450) );
  NAND2_X1 U10019 ( .A1(n8448), .A2(n8477), .ZN(n8449) );
  OAI211_X1 U10020 ( .C1(n8451), .C2(n8481), .A(n8450), .B(n8449), .ZN(
        P2_U3448) );
  INV_X1 U10021 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8453) );
  MUX2_X1 U10022 ( .A(n8453), .B(n8452), .S(n9829), .Z(n8454) );
  OAI21_X1 U10023 ( .B1(n8455), .B2(n8481), .A(n8454), .ZN(P2_U3447) );
  MUX2_X1 U10024 ( .A(n8456), .B(P2_REG0_REG_19__SCAN_IN), .S(n9831), .Z(n8457) );
  INV_X1 U10025 ( .A(n8457), .ZN(n8462) );
  AOI22_X1 U10026 ( .A1(n8460), .A2(n8459), .B1(n8477), .B2(n8458), .ZN(n8461)
         );
  NAND2_X1 U10027 ( .A1(n8462), .A2(n8461), .ZN(P2_U3446) );
  INV_X1 U10028 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8464) );
  MUX2_X1 U10029 ( .A(n8464), .B(n8463), .S(n9829), .Z(n8467) );
  NAND2_X1 U10030 ( .A1(n8465), .A2(n8477), .ZN(n8466) );
  OAI211_X1 U10031 ( .C1(n8468), .C2(n8481), .A(n8467), .B(n8466), .ZN(
        P2_U3444) );
  INV_X1 U10032 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8470) );
  MUX2_X1 U10033 ( .A(n8470), .B(n8469), .S(n9829), .Z(n8473) );
  NAND2_X1 U10034 ( .A1(n8471), .A2(n8477), .ZN(n8472) );
  OAI211_X1 U10035 ( .C1(n8474), .C2(n8481), .A(n8473), .B(n8472), .ZN(
        P2_U3441) );
  INV_X1 U10036 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8476) );
  MUX2_X1 U10037 ( .A(n8476), .B(n8475), .S(n9829), .Z(n8480) );
  NAND2_X1 U10038 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  OAI211_X1 U10039 ( .C1(n8482), .C2(n8481), .A(n8480), .B(n8479), .ZN(
        P2_U3438) );
  MUX2_X1 U10040 ( .A(P2_REG0_REG_1__SCAN_IN), .B(n8483), .S(n9829), .Z(
        P2_U3393) );
  INV_X1 U10041 ( .A(n8768), .ZN(n9448) );
  NOR4_X1 U10042 ( .A1(n8484), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8485), .A4(
        P2_U3151), .ZN(n8486) );
  AOI21_X1 U10043 ( .B1(n8487), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8486), .ZN(
        n8488) );
  OAI21_X1 U10044 ( .B1(n9448), .B2(n8492), .A(n8488), .ZN(P2_U3264) );
  OAI222_X1 U10045 ( .A1(P2_U3151), .A2(n8491), .B1(n8492), .B2(n8490), .C1(
        n8489), .C2(n8494), .ZN(P2_U3265) );
  OAI222_X1 U10046 ( .A1(P2_U3151), .A2(n8495), .B1(n8494), .B2(n6323), .C1(
        n8493), .C2(n8492), .ZN(P2_U3266) );
  MUX2_X1 U10047 ( .A(n8496), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10048 ( .A(n8572), .ZN(n8502) );
  OAI21_X1 U10049 ( .B1(n8500), .B2(n8498), .A(n8499), .ZN(n8501) );
  OAI211_X1 U10050 ( .C1(n8502), .C2(n8498), .A(n8603), .B(n8501), .ZN(n8509)
         );
  NAND2_X1 U10051 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9533) );
  INV_X1 U10052 ( .A(n9533), .ZN(n8503) );
  AOI21_X1 U10053 ( .B1(n8941), .B2(n8636), .A(n8503), .ZN(n8504) );
  OAI21_X1 U10054 ( .B1(n8505), .B2(n8638), .A(n8504), .ZN(n8506) );
  AOI21_X1 U10055 ( .B1(n8507), .B2(n8607), .A(n8506), .ZN(n8508) );
  OAI211_X1 U10056 ( .C1(n9441), .C2(n8610), .A(n8509), .B(n8508), .ZN(
        P1_U3215) );
  AND3_X1 U10057 ( .A1(n8513), .A2(n8511), .A3(n8512), .ZN(n8514) );
  OAI21_X1 U10058 ( .B1(n8510), .B2(n8514), .A(n8603), .ZN(n8519) );
  NOR2_X1 U10059 ( .A1(n9166), .A2(n8635), .ZN(n8517) );
  OAI22_X1 U10060 ( .A1(n9156), .A2(n8624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8515), .ZN(n8516) );
  AOI211_X1 U10061 ( .C1(n8936), .C2(n8627), .A(n8517), .B(n8516), .ZN(n8518)
         );
  OAI211_X1 U10062 ( .C1(n6393), .C2(n8610), .A(n8519), .B(n8518), .ZN(
        P1_U3216) );
  XNOR2_X1 U10063 ( .A(n8521), .B(n8520), .ZN(n8522) );
  XNOR2_X1 U10064 ( .A(n8523), .B(n8522), .ZN(n8528) );
  NOR2_X1 U10065 ( .A1(n8635), .A2(n9226), .ZN(n8526) );
  NAND2_X1 U10066 ( .A1(n9193), .A2(n8627), .ZN(n8524) );
  NAND2_X1 U10067 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9048) );
  OAI211_X1 U10068 ( .C1(n9262), .C2(n8624), .A(n8524), .B(n9048), .ZN(n8525)
         );
  AOI211_X1 U10069 ( .C1(n9233), .C2(n8641), .A(n8526), .B(n8525), .ZN(n8527)
         );
  OAI21_X1 U10070 ( .B1(n8528), .B2(n8643), .A(n8527), .ZN(P1_U3219) );
  OAI22_X1 U10071 ( .A1(n9085), .A2(n5735), .B1(n9094), .B2(n8532), .ZN(n8530)
         );
  XNOR2_X1 U10072 ( .A(n8530), .B(n8529), .ZN(n8534) );
  OAI22_X1 U10073 ( .A1(n9085), .A2(n8532), .B1(n9094), .B2(n8531), .ZN(n8533)
         );
  XNOR2_X1 U10074 ( .A(n8534), .B(n8533), .ZN(n8547) );
  INV_X1 U10075 ( .A(n8546), .ZN(n8538) );
  INV_X1 U10076 ( .A(n8547), .ZN(n8537) );
  NAND4_X1 U10077 ( .A1(n8539), .A2(n8538), .A3(n8537), .A4(n8603), .ZN(n8550)
         );
  NOR2_X1 U10078 ( .A1(n8540), .A2(n8624), .ZN(n8545) );
  INV_X1 U10079 ( .A(n8541), .ZN(n9082) );
  AOI22_X1 U10080 ( .A1(n9082), .A2(n8607), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8542) );
  OAI21_X1 U10081 ( .B1(n8543), .B2(n8638), .A(n8542), .ZN(n8544) );
  AOI211_X1 U10082 ( .C1(n9327), .C2(n8641), .A(n8545), .B(n8544), .ZN(n8549)
         );
  NAND3_X1 U10083 ( .A1(n8547), .A2(n8603), .A3(n8546), .ZN(n8548) );
  NAND4_X1 U10084 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), .ZN(
        P1_U3220) );
  NAND2_X1 U10085 ( .A1(n8602), .A2(n8601), .ZN(n8600) );
  NAND2_X1 U10086 ( .A1(n8600), .A2(n8552), .ZN(n8554) );
  OAI21_X1 U10087 ( .B1(n8555), .B2(n8554), .A(n8553), .ZN(n8556) );
  NAND2_X1 U10088 ( .A1(n8556), .A2(n8603), .ZN(n8561) );
  NOR2_X1 U10089 ( .A1(n9203), .A2(n8635), .ZN(n8559) );
  OAI22_X1 U10090 ( .A1(n9221), .A2(n8624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8557), .ZN(n8558) );
  AOI211_X1 U10091 ( .C1(n8627), .C2(n9194), .A(n8559), .B(n8558), .ZN(n8560)
         );
  OAI211_X1 U10092 ( .C1(n9424), .C2(n8610), .A(n8561), .B(n8560), .ZN(
        P1_U3223) );
  OAI21_X1 U10093 ( .B1(n8563), .B2(n8562), .A(n6299), .ZN(n8564) );
  NAND2_X1 U10094 ( .A1(n8564), .A2(n8603), .ZN(n8569) );
  NOR2_X1 U10095 ( .A1(n9135), .A2(n8635), .ZN(n8567) );
  OAI22_X1 U10096 ( .A1(n9157), .A2(n8624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8565), .ZN(n8566) );
  AOI211_X1 U10097 ( .C1(n8935), .C2(n8627), .A(n8567), .B(n8566), .ZN(n8568)
         );
  OAI211_X1 U10098 ( .C1(n9127), .C2(n8610), .A(n8569), .B(n8568), .ZN(
        P1_U3225) );
  NOR2_X1 U10099 ( .A1(n8572), .A2(n8498), .ZN(n8570) );
  XOR2_X1 U10100 ( .A(n8571), .B(n8570), .Z(n8633) );
  NOR2_X1 U10101 ( .A1(n8633), .A2(n8634), .ZN(n8632) );
  NOR3_X1 U10102 ( .A1(n8572), .A2(n8498), .A3(n8571), .ZN(n8573) );
  NOR2_X1 U10103 ( .A1(n8632), .A2(n8573), .ZN(n8574) );
  XOR2_X1 U10104 ( .A(n8575), .B(n8574), .Z(n8581) );
  OAI21_X1 U10105 ( .B1(n9240), .B2(n8638), .A(n8576), .ZN(n8577) );
  AOI21_X1 U10106 ( .B1(n8636), .B2(n9282), .A(n8577), .ZN(n8578) );
  OAI21_X1 U10107 ( .B1(n8635), .B2(n9275), .A(n8578), .ZN(n8579) );
  AOI21_X1 U10108 ( .B1(n9389), .B2(n8641), .A(n8579), .ZN(n8580) );
  OAI21_X1 U10109 ( .B1(n8581), .B2(n8643), .A(n8580), .ZN(P1_U3226) );
  XOR2_X1 U10110 ( .A(n8583), .B(n8582), .Z(n8589) );
  NOR2_X1 U10111 ( .A1(n9260), .A2(n8624), .ZN(n8584) );
  AOI211_X1 U10112 ( .C1(n8627), .C2(n8940), .A(n8585), .B(n8584), .ZN(n8586)
         );
  OAI21_X1 U10113 ( .B1(n8635), .B2(n9253), .A(n8586), .ZN(n8587) );
  AOI21_X1 U10114 ( .B1(n9384), .B2(n8641), .A(n8587), .ZN(n8588) );
  OAI21_X1 U10115 ( .B1(n8589), .B2(n8643), .A(n8588), .ZN(P1_U3228) );
  INV_X1 U10116 ( .A(n8590), .ZN(n8594) );
  NOR3_X1 U10117 ( .A1(n8510), .A2(n8592), .A3(n8591), .ZN(n8593) );
  OAI21_X1 U10118 ( .B1(n8594), .B2(n8593), .A(n8603), .ZN(n8599) );
  OAI22_X1 U10119 ( .A1(n9181), .A2(n8624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8595), .ZN(n8597) );
  NOR2_X1 U10120 ( .A1(n9147), .A2(n8638), .ZN(n8596) );
  AOI211_X1 U10121 ( .C1(n9149), .C2(n8607), .A(n8597), .B(n8596), .ZN(n8598)
         );
  OAI211_X1 U10122 ( .C1(n9152), .C2(n8610), .A(n8599), .B(n8598), .ZN(
        P1_U3229) );
  OAI21_X1 U10123 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8604) );
  NAND2_X1 U10124 ( .A1(n8604), .A2(n8603), .ZN(n8609) );
  AOI22_X1 U10125 ( .A1(n8938), .A2(n8627), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8605) );
  OAI21_X1 U10126 ( .B1(n9241), .B2(n8624), .A(n8605), .ZN(n8606) );
  AOI21_X1 U10127 ( .B1(n9214), .B2(n8607), .A(n8606), .ZN(n8608) );
  OAI211_X1 U10128 ( .C1(n4496), .C2(n8610), .A(n8609), .B(n8608), .ZN(
        P1_U3233) );
  INV_X1 U10129 ( .A(n8511), .ZN(n8611) );
  AOI21_X1 U10130 ( .B1(n8613), .B2(n8612), .A(n8611), .ZN(n8619) );
  OAI22_X1 U10131 ( .A1(n9212), .A2(n8624), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8614), .ZN(n8615) );
  AOI21_X1 U10132 ( .B1(n8627), .B2(n8937), .A(n8615), .ZN(n8616) );
  OAI21_X1 U10133 ( .B1(n8635), .B2(n9175), .A(n8616), .ZN(n8617) );
  AOI21_X1 U10134 ( .B1(n9357), .B2(n8641), .A(n8617), .ZN(n8618) );
  OAI21_X1 U10135 ( .B1(n8619), .B2(n8643), .A(n8618), .ZN(P1_U3235) );
  XNOR2_X1 U10136 ( .A(n8621), .B(n8620), .ZN(n8622) );
  XNOR2_X1 U10137 ( .A(n8623), .B(n8622), .ZN(n8631) );
  NOR2_X1 U10138 ( .A1(n9240), .A2(n8624), .ZN(n8625) );
  AOI211_X1 U10139 ( .C1(n8627), .C2(n8939), .A(n8626), .B(n8625), .ZN(n8628)
         );
  OAI21_X1 U10140 ( .B1(n8635), .B2(n9243), .A(n8628), .ZN(n8629) );
  AOI21_X1 U10141 ( .B1(n9379), .B2(n8641), .A(n8629), .ZN(n8630) );
  OAI21_X1 U10142 ( .B1(n8631), .B2(n8643), .A(n8630), .ZN(P1_U3238) );
  AOI21_X1 U10143 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8644) );
  NOR2_X1 U10144 ( .A1(n8635), .A2(n9310), .ZN(n8640) );
  AOI22_X1 U10145 ( .A1(n9297), .A2(n8636), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8637) );
  OAI21_X1 U10146 ( .B1(n9260), .B2(n8638), .A(n8637), .ZN(n8639) );
  AOI211_X1 U10147 ( .C1(n9308), .C2(n8641), .A(n8640), .B(n8639), .ZN(n8642)
         );
  OAI21_X1 U10148 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(P1_U3241) );
  NOR2_X1 U10149 ( .A1(n9194), .A2(n8760), .ZN(n8646) );
  INV_X1 U10150 ( .A(n8646), .ZN(n8645) );
  OAI22_X1 U10151 ( .A1(n9178), .A2(n8645), .B1(n8760), .B2(n8937), .ZN(n8651)
         );
  AOI21_X1 U10152 ( .B1(n9181), .B2(n8646), .A(n9178), .ZN(n8650) );
  AND2_X1 U10153 ( .A1(n9194), .A2(n8760), .ZN(n8647) );
  AOI21_X1 U10154 ( .B1(n8647), .B2(n8937), .A(n9357), .ZN(n8649) );
  AOI22_X1 U10155 ( .A1(n9178), .A2(n8647), .B1(n8760), .B2(n8937), .ZN(n8648)
         );
  MUX2_X1 U10156 ( .A(n9129), .B(n8862), .S(n8919), .Z(n8748) );
  AOI21_X1 U10157 ( .B1(n8653), .B2(n8652), .A(n9179), .ZN(n8747) );
  OR2_X1 U10158 ( .A1(n8876), .A2(n8919), .ZN(n8659) );
  INV_X1 U10159 ( .A(n8781), .ZN(n8654) );
  INV_X1 U10160 ( .A(n8872), .ZN(n8655) );
  OR3_X1 U10161 ( .A1(n8735), .A2(n8760), .A3(n8655), .ZN(n8657) );
  NAND4_X1 U10162 ( .A1(n8782), .A2(n8760), .A3(n9189), .A4(n8660), .ZN(n8656)
         );
  NAND4_X1 U10163 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n8746)
         );
  AND2_X1 U10164 ( .A1(n8660), .A2(n8738), .ZN(n8856) );
  NAND4_X1 U10165 ( .A1(n8661), .A2(n8665), .A3(n8821), .A4(n8825), .ZN(n8675)
         );
  OAI21_X1 U10166 ( .B1(n8663), .B2(n8760), .A(n8664), .ZN(n8662) );
  OAI21_X1 U10167 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8668) );
  OR2_X1 U10168 ( .A1(n8666), .A2(n8823), .ZN(n8667) );
  OAI211_X1 U10169 ( .C1(n8760), .C2(n8825), .A(n8668), .B(n8667), .ZN(n8669)
         );
  INV_X1 U10170 ( .A(n8669), .ZN(n8674) );
  NAND2_X1 U10171 ( .A1(n8670), .A2(n8821), .ZN(n8672) );
  NAND4_X1 U10172 ( .A1(n8672), .A2(n8919), .A3(n8671), .A4(n8823), .ZN(n8673)
         );
  NAND3_X1 U10173 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n8686) );
  INV_X1 U10174 ( .A(n8676), .ZN(n8678) );
  OAI21_X1 U10175 ( .B1(n8686), .B2(n8678), .A(n8677), .ZN(n8681) );
  NAND3_X1 U10176 ( .A1(n8681), .A2(n8680), .A3(n8679), .ZN(n8682) );
  NAND3_X1 U10177 ( .A1(n8682), .A2(n8692), .A3(n8687), .ZN(n8684) );
  NAND3_X1 U10178 ( .A1(n8684), .A2(n8702), .A3(n8683), .ZN(n8695) );
  AOI21_X1 U10179 ( .B1(n8686), .B2(n8831), .A(n8685), .ZN(n8689) );
  OAI21_X1 U10180 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8691) );
  NAND2_X1 U10181 ( .A1(n8691), .A2(n8690), .ZN(n8693) );
  NAND2_X1 U10182 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  MUX2_X1 U10183 ( .A(n8695), .B(n8694), .S(n8919), .Z(n8704) );
  INV_X1 U10184 ( .A(n8705), .ZN(n8696) );
  AOI21_X1 U10185 ( .B1(n8704), .B2(n8701), .A(n8696), .ZN(n8699) );
  NAND2_X1 U10186 ( .A1(n8709), .A2(n8835), .ZN(n8698) );
  OAI21_X1 U10187 ( .B1(n8699), .B2(n8698), .A(n8697), .ZN(n8700) );
  NAND2_X1 U10188 ( .A1(n8700), .A2(n8710), .ZN(n8713) );
  INV_X1 U10189 ( .A(n8701), .ZN(n8703) );
  OAI21_X1 U10190 ( .B1(n8704), .B2(n8703), .A(n8702), .ZN(n8708) );
  AND2_X1 U10191 ( .A1(n8706), .A2(n8705), .ZN(n8839) );
  INV_X1 U10192 ( .A(n8839), .ZN(n8707) );
  AOI21_X1 U10193 ( .B1(n8708), .B2(n8835), .A(n8707), .ZN(n8711) );
  NAND2_X1 U10194 ( .A1(n8710), .A2(n8709), .ZN(n8838) );
  OAI21_X1 U10195 ( .B1(n8711), .B2(n8838), .A(n8841), .ZN(n8712) );
  MUX2_X1 U10196 ( .A(n8713), .B(n8712), .S(n8919), .Z(n8720) );
  NAND2_X1 U10197 ( .A1(n8720), .A2(n8845), .ZN(n8714) );
  NAND3_X1 U10198 ( .A1(n8714), .A2(n8719), .A3(n8722), .ZN(n8715) );
  AND2_X1 U10199 ( .A1(n8723), .A2(n8728), .ZN(n8850) );
  NAND3_X1 U10200 ( .A1(n8715), .A2(n8850), .A3(n8846), .ZN(n8718) );
  NAND2_X1 U10201 ( .A1(n8723), .A2(n8716), .ZN(n8717) );
  NAND3_X1 U10202 ( .A1(n8718), .A2(n8855), .A3(n8717), .ZN(n8731) );
  NAND2_X1 U10203 ( .A1(n8720), .A2(n8719), .ZN(n8721) );
  NAND3_X1 U10204 ( .A1(n8721), .A2(n8805), .A3(n8845), .ZN(n8726) );
  NAND2_X1 U10205 ( .A1(n9281), .A2(n8722), .ZN(n8851) );
  INV_X1 U10206 ( .A(n8851), .ZN(n8725) );
  INV_X1 U10207 ( .A(n8723), .ZN(n8724) );
  AOI21_X1 U10208 ( .B1(n8726), .B2(n8725), .A(n8724), .ZN(n8729) );
  INV_X1 U10209 ( .A(n8855), .ZN(n8727) );
  AOI21_X1 U10210 ( .B1(n8729), .B2(n8728), .A(n8727), .ZN(n8730) );
  MUX2_X1 U10211 ( .A(n8731), .B(n8730), .S(n8760), .Z(n8732) );
  NAND2_X1 U10212 ( .A1(n8732), .A2(n9257), .ZN(n8740) );
  NAND2_X1 U10213 ( .A1(n8736), .A2(n8733), .ZN(n8857) );
  INV_X1 U10214 ( .A(n8857), .ZN(n8808) );
  NAND2_X1 U10215 ( .A1(n8740), .A2(n8808), .ZN(n8734) );
  NAND4_X1 U10216 ( .A1(n8868), .A2(n8856), .A3(n8734), .A4(n8919), .ZN(n8745)
         );
  INV_X1 U10217 ( .A(n8735), .ZN(n8743) );
  AND2_X1 U10218 ( .A1(n8736), .A2(n8760), .ZN(n8742) );
  NAND2_X1 U10219 ( .A1(n8738), .A2(n8737), .ZN(n8853) );
  INV_X1 U10220 ( .A(n8853), .ZN(n8739) );
  NAND2_X1 U10221 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  NAND4_X1 U10222 ( .A1(n8743), .A2(n8742), .A3(n8741), .A4(n8872), .ZN(n8744)
         );
  INV_X1 U10223 ( .A(n8780), .ZN(n8749) );
  OAI211_X1 U10224 ( .C1(n8751), .C2(n8749), .A(n8881), .B(n8779), .ZN(n8750)
         );
  NAND2_X1 U10225 ( .A1(n8750), .A2(n8880), .ZN(n8754) );
  NAND2_X1 U10226 ( .A1(n8752), .A2(n8881), .ZN(n8753) );
  MUX2_X1 U10227 ( .A(n8754), .B(n8753), .S(n8919), .Z(n8756) );
  INV_X1 U10228 ( .A(n8886), .ZN(n8870) );
  NAND2_X1 U10229 ( .A1(n8759), .A2(n8757), .ZN(n8884) );
  INV_X1 U10230 ( .A(n8884), .ZN(n8755) );
  OAI21_X1 U10231 ( .B1(n8756), .B2(n8870), .A(n8755), .ZN(n8758) );
  AOI21_X1 U10232 ( .B1(n8859), .B2(n8886), .A(n8760), .ZN(n8761) );
  OAI22_X1 U10233 ( .A1(n8762), .A2(n8761), .B1(n8760), .B2(n8759), .ZN(n8764)
         );
  MUX2_X1 U10234 ( .A(n8888), .B(n8860), .S(n8919), .Z(n8763) );
  NAND2_X1 U10235 ( .A1(n8765), .A2(n5758), .ZN(n8767) );
  NAND2_X1 U10236 ( .A1(n5759), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U10237 ( .A1(n8768), .A2(n5758), .ZN(n8770) );
  NAND2_X1 U10238 ( .A1(n5759), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8769) );
  INV_X1 U10239 ( .A(n8933), .ZN(n8816) );
  NAND2_X1 U10240 ( .A1(n6094), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8774) );
  INV_X1 U10241 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9320) );
  OR2_X1 U10242 ( .A1(n8771), .A2(n9320), .ZN(n8773) );
  INV_X1 U10243 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9403) );
  OR2_X1 U10244 ( .A1(n5751), .A2(n9403), .ZN(n8772) );
  AND3_X1 U10245 ( .A1(n8774), .A2(n8773), .A3(n8772), .ZN(n9056) );
  AOI21_X1 U10246 ( .B1(n9052), .B2(n8816), .A(n9056), .ZN(n8778) );
  MUX2_X1 U10247 ( .A(n8919), .B(n8775), .S(n9051), .Z(n8776) );
  NAND3_X1 U10248 ( .A1(n8776), .A2(n8933), .A3(n9052), .ZN(n8777) );
  NAND2_X1 U10249 ( .A1(n9052), .A2(n9056), .ZN(n8920) );
  AOI21_X1 U10250 ( .B1(n8922), .B2(n8921), .A(n8819), .ZN(n8931) );
  OR2_X1 U10251 ( .A1(n9052), .A2(n9056), .ZN(n8904) );
  NAND2_X1 U10252 ( .A1(n8780), .A2(n8779), .ZN(n9132) );
  NAND2_X1 U10253 ( .A1(n8782), .A2(n8781), .ZN(n9198) );
  INV_X1 U10254 ( .A(n9271), .ZN(n9280) );
  INV_X1 U10255 ( .A(n9291), .ZN(n9303) );
  INV_X1 U10256 ( .A(n8783), .ZN(n8796) );
  INV_X1 U10257 ( .A(n8784), .ZN(n8785) );
  NAND4_X1 U10258 ( .A1(n9552), .A2(n8786), .A3(n8785), .A4(n8819), .ZN(n8788)
         );
  OR3_X1 U10259 ( .A1(n8788), .A2(n6397), .A3(n8787), .ZN(n8792) );
  NOR4_X1 U10260 ( .A1(n8792), .A2(n8791), .A3(n8790), .A4(n8789), .ZN(n8795)
         );
  INV_X1 U10261 ( .A(n8793), .ZN(n8794) );
  NAND4_X1 U10262 ( .A1(n8797), .A2(n8796), .A3(n8795), .A4(n8794), .ZN(n8799)
         );
  NOR2_X1 U10263 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  NAND2_X1 U10264 ( .A1(n8801), .A2(n8800), .ZN(n8802) );
  NOR2_X1 U10265 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  NAND4_X1 U10266 ( .A1(n9280), .A2(n8805), .A3(n9303), .A4(n8804), .ZN(n8806)
         );
  NOR2_X1 U10267 ( .A1(n8853), .A2(n8806), .ZN(n8807) );
  NAND3_X1 U10268 ( .A1(n9224), .A2(n8808), .A3(n8807), .ZN(n8809) );
  OR3_X1 U10269 ( .A1(n9198), .A2(n9210), .A3(n8809), .ZN(n8810) );
  NOR2_X1 U10270 ( .A1(n9179), .A2(n8810), .ZN(n8811) );
  NAND3_X1 U10271 ( .A1(n9144), .A2(n9164), .A3(n8811), .ZN(n8812) );
  NOR2_X1 U10272 ( .A1(n9132), .A2(n8812), .ZN(n8813) );
  NAND4_X1 U10273 ( .A1(n9078), .A2(n4546), .A3(n9115), .A4(n8813), .ZN(n8814)
         );
  NOR2_X1 U10274 ( .A1(n8815), .A2(n8814), .ZN(n8818) );
  OR2_X1 U10275 ( .A1(n9051), .A2(n8816), .ZN(n8900) );
  NAND2_X1 U10276 ( .A1(n9051), .A2(n8816), .ZN(n8887) );
  AND2_X1 U10277 ( .A1(n8900), .A2(n8887), .ZN(n8817) );
  NAND4_X1 U10278 ( .A1(n8904), .A2(n8920), .A3(n8818), .A4(n8817), .ZN(n8909)
         );
  NAND4_X1 U10279 ( .A1(n8909), .A2(n8915), .A3(n9045), .A4(n8907), .ZN(n8930)
         );
  AOI21_X1 U10280 ( .B1(n5743), .B2(n5744), .A(n8819), .ZN(n8822) );
  NAND3_X1 U10281 ( .A1(n8822), .A2(n8821), .A3(n8820), .ZN(n8824) );
  NAND2_X1 U10282 ( .A1(n8824), .A2(n8823), .ZN(n8827) );
  OAI211_X1 U10283 ( .C1(n8828), .C2(n8827), .A(n8826), .B(n8825), .ZN(n8832)
         );
  INV_X1 U10284 ( .A(n8829), .ZN(n8830) );
  AOI21_X1 U10285 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8837) );
  INV_X1 U10286 ( .A(n8833), .ZN(n8836) );
  OAI211_X1 U10287 ( .C1(n8837), .C2(n8836), .A(n8835), .B(n8834), .ZN(n8840)
         );
  AOI21_X1 U10288 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8844) );
  INV_X1 U10289 ( .A(n8841), .ZN(n8842) );
  NOR3_X1 U10290 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n8849) );
  INV_X1 U10291 ( .A(n8845), .ZN(n8848) );
  INV_X1 U10292 ( .A(n8846), .ZN(n8847) );
  NOR3_X1 U10293 ( .A1(n8849), .A2(n8848), .A3(n8847), .ZN(n8852) );
  OAI21_X1 U10294 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8854) );
  AOI21_X1 U10295 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n8858) );
  OAI21_X1 U10296 ( .B1(n8858), .B2(n8857), .A(n8856), .ZN(n8871) );
  NAND2_X1 U10297 ( .A1(n8860), .A2(n8859), .ZN(n8890) );
  NAND2_X1 U10298 ( .A1(n8862), .A2(n8861), .ZN(n8874) );
  AND2_X1 U10299 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  OR2_X1 U10300 ( .A1(n8874), .A2(n8865), .ZN(n8866) );
  NAND2_X1 U10301 ( .A1(n8867), .A2(n8866), .ZN(n8873) );
  NAND2_X1 U10302 ( .A1(n8880), .A2(n8868), .ZN(n8869) );
  OR4_X1 U10303 ( .A1(n8890), .A2(n8870), .A3(n8873), .A4(n8869), .ZN(n8896)
         );
  AOI21_X1 U10304 ( .B1(n8872), .B2(n8871), .A(n8896), .ZN(n8891) );
  INV_X1 U10305 ( .A(n8873), .ZN(n8879) );
  INV_X1 U10306 ( .A(n8874), .ZN(n8877) );
  NAND3_X1 U10307 ( .A1(n8877), .A2(n8876), .A3(n8875), .ZN(n8878) );
  AOI21_X1 U10308 ( .B1(n8879), .B2(n8878), .A(n4513), .ZN(n8883) );
  INV_X1 U10309 ( .A(n8880), .ZN(n8882) );
  OAI21_X1 U10310 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8885) );
  AOI21_X1 U10311 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n8889) );
  OAI211_X1 U10312 ( .C1(n8890), .C2(n8889), .A(n8888), .B(n8887), .ZN(n8899)
         );
  OAI211_X1 U10313 ( .C1(n8891), .C2(n8899), .A(n8920), .B(n8900), .ZN(n8892)
         );
  NAND2_X1 U10314 ( .A1(n8892), .A2(n8904), .ZN(n8895) );
  AOI21_X1 U10315 ( .B1(n9045), .B2(n8893), .A(n8895), .ZN(n8894) );
  AOI211_X1 U10316 ( .C1(n6266), .C2(n8895), .A(n8924), .B(n8894), .ZN(n8918)
         );
  INV_X1 U10317 ( .A(n8896), .ZN(n8898) );
  AOI22_X1 U10318 ( .A1(n8898), .A2(n8897), .B1(n9405), .B2(n9051), .ZN(n8903)
         );
  INV_X1 U10319 ( .A(n8899), .ZN(n8902) );
  INV_X1 U10320 ( .A(n8900), .ZN(n8901) );
  INV_X1 U10321 ( .A(n9056), .ZN(n8932) );
  AOI22_X1 U10322 ( .A1(n8903), .A2(n8902), .B1(n8901), .B2(n8932), .ZN(n8906)
         );
  INV_X1 U10323 ( .A(n8904), .ZN(n8925) );
  OAI211_X1 U10324 ( .C1(n8906), .C2(n8925), .A(n8905), .B(n8920), .ZN(n8910)
         );
  NAND3_X1 U10325 ( .A1(n8915), .A2(n8907), .A3(n9264), .ZN(n8908) );
  AOI21_X1 U10326 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8917) );
  INV_X1 U10327 ( .A(P1_B_REG_SCAN_IN), .ZN(n8913) );
  NOR2_X1 U10328 ( .A1(n8911), .A2(n8963), .ZN(n8912) );
  AOI211_X1 U10329 ( .C1(n8915), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8916)
         );
  NOR3_X1 U10330 ( .A1(n8918), .A2(n8917), .A3(n8916), .ZN(n8929) );
  OAI22_X1 U10331 ( .A1(n8922), .A2(n8921), .B1(n8920), .B2(n8919), .ZN(n8927)
         );
  AOI211_X1 U10332 ( .C1(n8925), .C2(n9045), .A(n8924), .B(n8923), .ZN(n8926)
         );
  NAND2_X1 U10333 ( .A1(n8927), .A2(n8926), .ZN(n8928) );
  OAI211_X1 U10334 ( .C1(n8931), .C2(n8930), .A(n8929), .B(n8928), .ZN(
        P1_U3242) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n8932), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10336 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8933), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8934), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9117), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8935), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10340 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9116), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10341 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8936), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10342 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8937), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n8938), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9193), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n8939), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8940), .S(P1_U3973), .Z(
        P1_U3572) );
  INV_X1 U10348 ( .A(n9240), .ZN(n9283) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9283), .S(P1_U3973), .Z(
        P1_U3571) );
  INV_X1 U10350 ( .A(n9260), .ZN(n9300) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9300), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9282), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9297), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8941), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8942), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8943), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n5866), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8944), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8945), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8946), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5757), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5743), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6351), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI22_X1 U10364 ( .A1(n9892), .A2(n7128), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8947), .ZN(n8948) );
  AOI21_X1 U10365 ( .B1(n9881), .B2(n8949), .A(n8948), .ZN(n8958) );
  OAI211_X1 U10366 ( .C1(n8952), .C2(n8951), .A(n9879), .B(n8950), .ZN(n8957)
         );
  OAI211_X1 U10367 ( .C1(n8955), .C2(n8954), .A(n9885), .B(n8953), .ZN(n8956)
         );
  NAND3_X1 U10368 ( .A1(n8958), .A2(n8957), .A3(n8956), .ZN(P1_U3244) );
  NAND3_X1 U10369 ( .A1(n8961), .A2(n8960), .A3(n8959), .ZN(n8966) );
  OAI21_X1 U10370 ( .B1(n8963), .B2(n8962), .A(P1_U3973), .ZN(n8964) );
  INV_X1 U10371 ( .A(n8964), .ZN(n8965) );
  OAI211_X1 U10372 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n8967), .A(n8966), .B(
        n8965), .ZN(n9007) );
  INV_X1 U10373 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8969) );
  OAI22_X1 U10374 ( .A1(n9892), .A2(n8969), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8968), .ZN(n8970) );
  AOI21_X1 U10375 ( .B1(n9881), .B2(n8971), .A(n8970), .ZN(n8980) );
  OAI211_X1 U10376 ( .C1(n8974), .C2(n8973), .A(n9885), .B(n8972), .ZN(n8979)
         );
  OAI211_X1 U10377 ( .C1(n8977), .C2(n8976), .A(n9879), .B(n8975), .ZN(n8978)
         );
  NAND4_X1 U10378 ( .A1(n9007), .A2(n8980), .A3(n8979), .A4(n8978), .ZN(
        P1_U3245) );
  INV_X1 U10379 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8982) );
  OAI21_X1 U10380 ( .B1(n9892), .B2(n8982), .A(n8981), .ZN(n8983) );
  AOI21_X1 U10381 ( .B1(n9881), .B2(n8984), .A(n8983), .ZN(n8993) );
  OAI211_X1 U10382 ( .C1(n8987), .C2(n8986), .A(n9885), .B(n8985), .ZN(n8992)
         );
  OAI211_X1 U10383 ( .C1(n8990), .C2(n8989), .A(n9879), .B(n8988), .ZN(n8991)
         );
  NAND3_X1 U10384 ( .A1(n8993), .A2(n8992), .A3(n8991), .ZN(P1_U3246) );
  NOR2_X1 U10385 ( .A1(n9502), .A2(n8994), .ZN(n8995) );
  AOI211_X1 U10386 ( .C1(n8997), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n8996), .B(
        n8995), .ZN(n9006) );
  OAI211_X1 U10387 ( .C1(n9000), .C2(n8999), .A(n9879), .B(n8998), .ZN(n9005)
         );
  OAI211_X1 U10388 ( .C1(n9003), .C2(n9002), .A(n9885), .B(n9001), .ZN(n9004)
         );
  NAND4_X1 U10389 ( .A1(n9007), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(
        P1_U3247) );
  INV_X1 U10390 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9009) );
  OAI21_X1 U10391 ( .B1(n9892), .B2(n9009), .A(n9008), .ZN(n9010) );
  AOI21_X1 U10392 ( .B1(n9881), .B2(n9011), .A(n9010), .ZN(n9020) );
  OAI211_X1 U10393 ( .C1(n9014), .C2(n9013), .A(n9885), .B(n9012), .ZN(n9019)
         );
  OAI211_X1 U10394 ( .C1(n9017), .C2(n9016), .A(n9879), .B(n9015), .ZN(n9018)
         );
  NAND3_X1 U10395 ( .A1(n9020), .A2(n9019), .A3(n9018), .ZN(P1_U3248) );
  OAI21_X1 U10396 ( .B1(n9892), .B2(n9022), .A(n9021), .ZN(n9023) );
  AOI21_X1 U10397 ( .B1(n9881), .B2(n9024), .A(n9023), .ZN(n9033) );
  OAI211_X1 U10398 ( .C1(n9027), .C2(n9026), .A(n9885), .B(n9025), .ZN(n9032)
         );
  OAI211_X1 U10399 ( .C1(n9030), .C2(n9029), .A(n9879), .B(n9028), .ZN(n9031)
         );
  NAND3_X1 U10400 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(P1_U3249) );
  INV_X1 U10401 ( .A(n9034), .ZN(n9035) );
  NOR2_X1 U10402 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  XNOR2_X1 U10403 ( .A(n9037), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U10404 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  XNOR2_X1 U10405 ( .A(n9040), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9044) );
  INV_X1 U10406 ( .A(n9044), .ZN(n9041) );
  AOI22_X1 U10407 ( .A1(n9879), .A2(n9042), .B1(n9041), .B2(n9885), .ZN(n9047)
         );
  OAI21_X1 U10408 ( .B1(n9042), .B2(n9522), .A(n9502), .ZN(n9043) );
  AOI21_X1 U10409 ( .B1(n9044), .B2(n9885), .A(n9043), .ZN(n9046) );
  MUX2_X1 U10410 ( .A(n9047), .B(n9046), .S(n9045), .Z(n9049) );
  OAI211_X1 U10411 ( .C1(n9050), .C2(n9892), .A(n9049), .B(n9048), .ZN(
        P1_U3262) );
  XNOR2_X1 U10412 ( .A(n9059), .B(n9052), .ZN(n9053) );
  NAND2_X1 U10413 ( .A1(n9319), .A2(n4265), .ZN(n9058) );
  INV_X1 U10414 ( .A(n9054), .ZN(n9055) );
  NOR2_X1 U10415 ( .A1(n9056), .A2(n9055), .ZN(n9318) );
  INV_X1 U10416 ( .A(n9318), .ZN(n9322) );
  NOR2_X1 U10417 ( .A1(n9322), .A2(n9317), .ZN(n9061) );
  AOI21_X1 U10418 ( .B1(n9317), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9061), .ZN(
        n9057) );
  OAI211_X1 U10419 ( .C1(n9405), .C2(n9542), .A(n9058), .B(n9057), .ZN(
        P1_U3263) );
  OAI211_X1 U10420 ( .C1(n9408), .C2(n4293), .A(n9229), .B(n9059), .ZN(n9323)
         );
  NOR2_X1 U10421 ( .A1(n9408), .A2(n9542), .ZN(n9060) );
  AOI211_X1 U10422 ( .C1(n9317), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9061), .B(
        n9060), .ZN(n9062) );
  OAI21_X1 U10423 ( .B1(n9230), .B2(n9323), .A(n9062), .ZN(P1_U3264) );
  INV_X1 U10424 ( .A(n9063), .ZN(n9073) );
  NAND2_X1 U10425 ( .A1(n9064), .A2(n9545), .ZN(n9072) );
  INV_X1 U10426 ( .A(n9065), .ZN(n9066) );
  AOI22_X1 U10427 ( .A1(n9066), .A2(n9538), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9317), .ZN(n9067) );
  OAI21_X1 U10428 ( .B1(n9068), .B2(n9542), .A(n9067), .ZN(n9069) );
  AOI21_X1 U10429 ( .B1(n9070), .B2(n4265), .A(n9069), .ZN(n9071) );
  OAI211_X1 U10430 ( .C1(n9073), .C2(n9317), .A(n9072), .B(n9071), .ZN(
        P1_U3356) );
  INV_X1 U10431 ( .A(n9078), .ZN(n9074) );
  XNOR2_X1 U10432 ( .A(n9075), .B(n9074), .ZN(n9330) );
  OAI21_X1 U10433 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9080) );
  AOI222_X1 U10434 ( .A1(n9295), .A2(n9080), .B1(n9079), .B2(n9299), .C1(n9117), .C2(n9298), .ZN(n9329) );
  AOI211_X1 U10435 ( .C1(n9327), .C2(n9099), .A(n9306), .B(n9081), .ZN(n9326)
         );
  AOI22_X1 U10436 ( .A1(n9326), .A2(n9264), .B1(n9082), .B2(n9538), .ZN(n9083)
         );
  AOI21_X1 U10437 ( .B1(n9329), .B2(n9083), .A(n9317), .ZN(n9087) );
  OAI22_X1 U10438 ( .A1(n9085), .A2(n9542), .B1(n9287), .B2(n9084), .ZN(n9086)
         );
  NOR2_X1 U10439 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  OAI21_X1 U10440 ( .B1(n9330), .B2(n9290), .A(n9088), .ZN(P1_U3265) );
  XNOR2_X1 U10441 ( .A(n9090), .B(n9089), .ZN(n9333) );
  INV_X1 U10442 ( .A(n9333), .ZN(n9107) );
  OAI21_X1 U10443 ( .B1(n4546), .B2(n9092), .A(n9091), .ZN(n9093) );
  NAND2_X1 U10444 ( .A1(n9093), .A2(n9295), .ZN(n9097) );
  OAI22_X1 U10445 ( .A1(n9094), .A2(n9263), .B1(n9134), .B2(n9261), .ZN(n9095)
         );
  INV_X1 U10446 ( .A(n9095), .ZN(n9096) );
  NAND2_X1 U10447 ( .A1(n9097), .A2(n9096), .ZN(n9331) );
  INV_X1 U10448 ( .A(n9099), .ZN(n9100) );
  AOI211_X1 U10449 ( .C1(n9101), .C2(n9109), .A(n9306), .B(n9100), .ZN(n9332)
         );
  NAND2_X1 U10450 ( .A1(n9332), .A2(n4265), .ZN(n9104) );
  AOI22_X1 U10451 ( .A1(n9102), .A2(n9538), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9317), .ZN(n9103) );
  OAI211_X1 U10452 ( .C1(n6394), .C2(n9542), .A(n9104), .B(n9103), .ZN(n9105)
         );
  AOI21_X1 U10453 ( .B1(n9331), .B2(n9287), .A(n9105), .ZN(n9106) );
  OAI21_X1 U10454 ( .B1(n9107), .B2(n9290), .A(n9106), .ZN(P1_U3266) );
  XOR2_X1 U10455 ( .A(n9115), .B(n9108), .Z(n9340) );
  AOI211_X1 U10456 ( .C1(n9337), .C2(n9123), .A(n9306), .B(n9098), .ZN(n9336)
         );
  AOI22_X1 U10457 ( .A1(n9110), .A2(n9538), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9317), .ZN(n9111) );
  OAI21_X1 U10458 ( .B1(n9112), .B2(n9542), .A(n9111), .ZN(n9120) );
  OAI21_X1 U10459 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9118) );
  AOI222_X1 U10460 ( .A1(n9295), .A2(n9118), .B1(n9117), .B2(n9299), .C1(n9116), .C2(n9298), .ZN(n9339) );
  NOR2_X1 U10461 ( .A1(n9339), .A2(n9317), .ZN(n9119) );
  AOI211_X1 U10462 ( .C1(n9336), .C2(n4265), .A(n9120), .B(n9119), .ZN(n9121)
         );
  OAI21_X1 U10463 ( .B1(n9340), .B2(n9290), .A(n9121), .ZN(P1_U3267) );
  XOR2_X1 U10464 ( .A(n9132), .B(n9122), .Z(n9345) );
  INV_X1 U10465 ( .A(n9148), .ZN(n9125) );
  INV_X1 U10466 ( .A(n9123), .ZN(n9124) );
  AOI211_X1 U10467 ( .C1(n9343), .C2(n9125), .A(n9306), .B(n9124), .ZN(n9342)
         );
  OAI22_X1 U10468 ( .A1(n9127), .A2(n9542), .B1(n9126), .B2(n9287), .ZN(n9128)
         );
  AOI21_X1 U10469 ( .B1(n9342), .B2(n4265), .A(n9128), .ZN(n9138) );
  NAND2_X1 U10470 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  XOR2_X1 U10471 ( .A(n9132), .B(n9131), .Z(n9133) );
  OAI222_X1 U10472 ( .A1(n9263), .A2(n9134), .B1(n9261), .B2(n9157), .C1(n9553), .C2(n9133), .ZN(n9341) );
  NOR2_X1 U10473 ( .A1(n9135), .A2(n9309), .ZN(n9136) );
  OAI21_X1 U10474 ( .B1(n9341), .B2(n9136), .A(n9287), .ZN(n9137) );
  OAI211_X1 U10475 ( .C1(n9345), .C2(n9290), .A(n9138), .B(n9137), .ZN(
        P1_U3268) );
  OR2_X1 U10476 ( .A1(n9174), .A2(n9139), .ZN(n9141) );
  NAND2_X1 U10477 ( .A1(n9141), .A2(n9140), .ZN(n9143) );
  XNOR2_X1 U10478 ( .A(n9143), .B(n9142), .ZN(n9350) );
  XNOR2_X1 U10479 ( .A(n9145), .B(n9144), .ZN(n9146) );
  OAI222_X1 U10480 ( .A1(n9263), .A2(n9147), .B1(n9261), .B2(n9181), .C1(n9146), .C2(n9553), .ZN(n9346) );
  AOI211_X1 U10481 ( .C1(n9348), .C2(n9168), .A(n9306), .B(n9148), .ZN(n9347)
         );
  NAND2_X1 U10482 ( .A1(n9347), .A2(n4265), .ZN(n9151) );
  AOI22_X1 U10483 ( .A1(n9149), .A2(n9538), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9317), .ZN(n9150) );
  OAI211_X1 U10484 ( .C1(n9152), .C2(n9542), .A(n9151), .B(n9150), .ZN(n9153)
         );
  AOI21_X1 U10485 ( .B1(n9346), .B2(n9287), .A(n9153), .ZN(n9154) );
  OAI21_X1 U10486 ( .B1(n9350), .B2(n9290), .A(n9154), .ZN(P1_U3269) );
  OAI21_X1 U10487 ( .B1(n9164), .B2(n4340), .A(n9155), .ZN(n9159) );
  OAI22_X1 U10488 ( .A1(n9157), .A2(n9263), .B1(n9156), .B2(n9261), .ZN(n9158)
         );
  AOI21_X1 U10489 ( .B1(n9159), .B2(n9295), .A(n9158), .ZN(n9352) );
  OR2_X1 U10490 ( .A1(n9174), .A2(n9160), .ZN(n9162) );
  NAND2_X1 U10491 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  XOR2_X1 U10492 ( .A(n9164), .B(n9163), .Z(n9353) );
  OR2_X1 U10493 ( .A1(n9353), .A2(n9290), .ZN(n9173) );
  OAI22_X1 U10494 ( .A1(n9166), .A2(n9309), .B1(n9165), .B2(n9287), .ZN(n9170)
         );
  OAI211_X1 U10495 ( .C1(n6393), .C2(n9167), .A(n9229), .B(n9168), .ZN(n9351)
         );
  NOR2_X1 U10496 ( .A1(n9351), .A2(n9230), .ZN(n9169) );
  AOI211_X1 U10497 ( .C1(n9268), .C2(n9171), .A(n9170), .B(n9169), .ZN(n9172)
         );
  OAI211_X1 U10498 ( .C1(n9317), .C2(n9352), .A(n9173), .B(n9172), .ZN(
        P1_U3270) );
  XOR2_X1 U10499 ( .A(n9179), .B(n9174), .Z(n9360) );
  AOI211_X1 U10500 ( .C1(n9357), .C2(n9199), .A(n9306), .B(n9167), .ZN(n9356)
         );
  INV_X1 U10501 ( .A(n9175), .ZN(n9176) );
  AOI22_X1 U10502 ( .A1(n9176), .A2(n9538), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9317), .ZN(n9177) );
  OAI21_X1 U10503 ( .B1(n9178), .B2(n9542), .A(n9177), .ZN(n9186) );
  AOI21_X1 U10504 ( .B1(n9180), .B2(n9179), .A(n9553), .ZN(n9184) );
  OAI22_X1 U10505 ( .A1(n9181), .A2(n9263), .B1(n9212), .B2(n9261), .ZN(n9182)
         );
  AOI21_X1 U10506 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9359) );
  NOR2_X1 U10507 ( .A1(n9359), .A2(n9317), .ZN(n9185) );
  AOI211_X1 U10508 ( .C1(n9356), .C2(n4265), .A(n9186), .B(n9185), .ZN(n9187)
         );
  OAI21_X1 U10509 ( .B1(n9360), .B2(n9290), .A(n9187), .ZN(P1_U3271) );
  INV_X1 U10510 ( .A(n9188), .ZN(n9190) );
  OAI21_X1 U10511 ( .B1(n8897), .B2(n9190), .A(n9189), .ZN(n9191) );
  XNOR2_X1 U10512 ( .A(n9191), .B(n9198), .ZN(n9192) );
  NAND2_X1 U10513 ( .A1(n9192), .A2(n9295), .ZN(n9196) );
  AOI22_X1 U10514 ( .A1(n9194), .A2(n9299), .B1(n9193), .B2(n9298), .ZN(n9195)
         );
  NAND2_X1 U10515 ( .A1(n9196), .A2(n9195), .ZN(n9361) );
  INV_X1 U10516 ( .A(n9361), .ZN(n9208) );
  XOR2_X1 U10517 ( .A(n9198), .B(n9197), .Z(n9363) );
  NAND2_X1 U10518 ( .A1(n9363), .A2(n9545), .ZN(n9207) );
  INV_X1 U10519 ( .A(n9199), .ZN(n9200) );
  AOI211_X1 U10520 ( .C1(n9201), .C2(n4498), .A(n9306), .B(n9200), .ZN(n9362)
         );
  NOR2_X1 U10521 ( .A1(n9424), .A2(n9542), .ZN(n9205) );
  OAI22_X1 U10522 ( .A1(n9203), .A2(n9309), .B1(n9287), .B2(n9202), .ZN(n9204)
         );
  AOI211_X1 U10523 ( .C1(n9362), .C2(n4265), .A(n9205), .B(n9204), .ZN(n9206)
         );
  OAI211_X1 U10524 ( .C1(n9317), .C2(n9208), .A(n9207), .B(n9206), .ZN(
        P1_U3272) );
  XNOR2_X1 U10525 ( .A(n9209), .B(n9210), .ZN(n9370) );
  XNOR2_X1 U10526 ( .A(n8897), .B(n9210), .ZN(n9211) );
  OAI222_X1 U10527 ( .A1(n9263), .A2(n9212), .B1(n9261), .B2(n9241), .C1(n9211), .C2(n9553), .ZN(n9366) );
  AOI211_X1 U10528 ( .C1(n9368), .C2(n9228), .A(n9306), .B(n9213), .ZN(n9367)
         );
  NAND2_X1 U10529 ( .A1(n9367), .A2(n4265), .ZN(n9216) );
  AOI22_X1 U10530 ( .A1(n9214), .A2(n9538), .B1(n9317), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9215) );
  OAI211_X1 U10531 ( .C1(n4496), .C2(n9542), .A(n9216), .B(n9215), .ZN(n9217)
         );
  AOI21_X1 U10532 ( .B1(n9366), .B2(n9287), .A(n9217), .ZN(n9218) );
  OAI21_X1 U10533 ( .B1(n9370), .B2(n9290), .A(n9218), .ZN(P1_U3273) );
  OAI21_X1 U10534 ( .B1(n9224), .B2(n9220), .A(n9219), .ZN(n9223) );
  OAI22_X1 U10535 ( .A1(n9221), .A2(n9263), .B1(n9262), .B2(n9261), .ZN(n9222)
         );
  AOI21_X1 U10536 ( .B1(n9223), .B2(n9295), .A(n9222), .ZN(n9372) );
  XOR2_X1 U10537 ( .A(n9225), .B(n9224), .Z(n9373) );
  OR2_X1 U10538 ( .A1(n9373), .A2(n9290), .ZN(n9235) );
  INV_X1 U10539 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9227) );
  OAI22_X1 U10540 ( .A1(n9287), .A2(n9227), .B1(n9226), .B2(n9309), .ZN(n9232)
         );
  OAI211_X1 U10541 ( .C1(n4343), .C2(n9429), .A(n9229), .B(n9228), .ZN(n9371)
         );
  NOR2_X1 U10542 ( .A1(n9371), .A2(n9230), .ZN(n9231) );
  AOI211_X1 U10543 ( .C1(n9268), .C2(n9233), .A(n9232), .B(n9231), .ZN(n9234)
         );
  OAI211_X1 U10544 ( .C1(n9317), .C2(n9372), .A(n9235), .B(n9234), .ZN(
        P1_U3274) );
  XNOR2_X1 U10545 ( .A(n9236), .B(n9237), .ZN(n9381) );
  AOI21_X1 U10546 ( .B1(n9238), .B2(n9237), .A(n4345), .ZN(n9239) );
  OAI222_X1 U10547 ( .A1(n9263), .A2(n9241), .B1(n9261), .B2(n9240), .C1(n9553), .C2(n9239), .ZN(n9377) );
  INV_X1 U10548 ( .A(n9255), .ZN(n9242) );
  AOI211_X1 U10549 ( .C1(n9379), .C2(n9242), .A(n9306), .B(n4343), .ZN(n9378)
         );
  NAND2_X1 U10550 ( .A1(n9378), .A2(n4265), .ZN(n9246) );
  INV_X1 U10551 ( .A(n9243), .ZN(n9244) );
  AOI22_X1 U10552 ( .A1(n9317), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9244), .B2(
        n9538), .ZN(n9245) );
  OAI211_X1 U10553 ( .C1(n9247), .C2(n9542), .A(n9246), .B(n9245), .ZN(n9248)
         );
  AOI21_X1 U10554 ( .B1(n9377), .B2(n9287), .A(n9248), .ZN(n9249) );
  OAI21_X1 U10555 ( .B1(n9381), .B2(n9290), .A(n9249), .ZN(P1_U3275) );
  OAI21_X1 U10556 ( .B1(n9252), .B2(n9251), .A(n9250), .ZN(n9386) );
  OAI22_X1 U10557 ( .A1(n9287), .A2(n9254), .B1(n9253), .B2(n9309), .ZN(n9267)
         );
  INV_X1 U10558 ( .A(n9273), .ZN(n9256) );
  AOI211_X1 U10559 ( .C1(n9384), .C2(n9256), .A(n9306), .B(n9255), .ZN(n9383)
         );
  XNOR2_X1 U10560 ( .A(n9258), .B(n9257), .ZN(n9259) );
  OAI222_X1 U10561 ( .A1(n9263), .A2(n9262), .B1(n9261), .B2(n9260), .C1(n9553), .C2(n9259), .ZN(n9382) );
  AOI21_X1 U10562 ( .B1(n9383), .B2(n9264), .A(n9382), .ZN(n9265) );
  NOR2_X1 U10563 ( .A1(n9265), .A2(n9317), .ZN(n9266) );
  AOI211_X1 U10564 ( .C1(n9268), .C2(n9384), .A(n9267), .B(n9266), .ZN(n9269)
         );
  OAI21_X1 U10565 ( .B1(n9386), .B2(n9290), .A(n9269), .ZN(P1_U3276) );
  OAI21_X1 U10566 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(n9391) );
  AOI211_X1 U10567 ( .C1(n9389), .C2(n9305), .A(n9306), .B(n9273), .ZN(n9388)
         );
  NOR2_X1 U10568 ( .A1(n9274), .A2(n9542), .ZN(n9278) );
  OAI22_X1 U10569 ( .A1(n9287), .A2(n9276), .B1(n9275), .B2(n9309), .ZN(n9277)
         );
  AOI211_X1 U10570 ( .C1(n9388), .C2(n4265), .A(n9278), .B(n9277), .ZN(n9289)
         );
  NAND2_X1 U10571 ( .A1(n9279), .A2(n9295), .ZN(n9286) );
  AOI21_X1 U10572 ( .B1(n9294), .B2(n9281), .A(n9280), .ZN(n9285) );
  AOI22_X1 U10573 ( .A1(n9283), .A2(n9299), .B1(n9298), .B2(n9282), .ZN(n9284)
         );
  OAI21_X1 U10574 ( .B1(n9286), .B2(n9285), .A(n9284), .ZN(n9387) );
  NAND2_X1 U10575 ( .A1(n9387), .A2(n9287), .ZN(n9288) );
  OAI211_X1 U10576 ( .C1(n9391), .C2(n9290), .A(n9289), .B(n9288), .ZN(
        P1_U3277) );
  NAND2_X1 U10577 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  NAND2_X1 U10578 ( .A1(n9294), .A2(n9293), .ZN(n9296) );
  NAND2_X1 U10579 ( .A1(n9296), .A2(n9295), .ZN(n9302) );
  AOI22_X1 U10580 ( .A1(n9300), .A2(n9299), .B1(n9298), .B2(n9297), .ZN(n9301)
         );
  NAND2_X1 U10581 ( .A1(n9302), .A2(n9301), .ZN(n9392) );
  INV_X1 U10582 ( .A(n9392), .ZN(n9316) );
  XNOR2_X1 U10583 ( .A(n9304), .B(n9303), .ZN(n9394) );
  NAND2_X1 U10584 ( .A1(n9394), .A2(n9545), .ZN(n9315) );
  AOI211_X1 U10585 ( .C1(n9308), .C2(n9307), .A(n9306), .B(n4486), .ZN(n9393)
         );
  NOR2_X1 U10586 ( .A1(n9436), .A2(n9542), .ZN(n9313) );
  OAI22_X1 U10587 ( .A1(n9287), .A2(n9311), .B1(n9310), .B2(n9309), .ZN(n9312)
         );
  AOI211_X1 U10588 ( .C1(n9393), .C2(n4265), .A(n9313), .B(n9312), .ZN(n9314)
         );
  OAI211_X1 U10589 ( .C1(n9317), .C2(n9316), .A(n9315), .B(n9314), .ZN(
        P1_U3278) );
  NOR2_X1 U10590 ( .A1(n9319), .A2(n9318), .ZN(n9402) );
  MUX2_X1 U10591 ( .A(n9320), .B(n9402), .S(n9608), .Z(n9321) );
  OAI21_X1 U10592 ( .B1(n9405), .B2(n9401), .A(n9321), .ZN(P1_U3553) );
  INV_X1 U10593 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9324) );
  AND2_X1 U10594 ( .A1(n9323), .A2(n9322), .ZN(n9406) );
  MUX2_X1 U10595 ( .A(n9324), .B(n9406), .S(n9608), .Z(n9325) );
  OAI21_X1 U10596 ( .B1(n9408), .B2(n9401), .A(n9325), .ZN(P1_U3552) );
  AOI21_X1 U10597 ( .B1(n9567), .B2(n9327), .A(n9326), .ZN(n9328) );
  OAI211_X1 U10598 ( .C1(n9330), .C2(n9571), .A(n9329), .B(n9328), .ZN(n9409)
         );
  MUX2_X1 U10599 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9409), .S(n9608), .Z(
        P1_U3550) );
  INV_X1 U10600 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9334) );
  AOI211_X1 U10601 ( .C1(n9333), .C2(n9595), .A(n9332), .B(n9331), .ZN(n9410)
         );
  MUX2_X1 U10602 ( .A(n9334), .B(n9410), .S(n9608), .Z(n9335) );
  OAI21_X1 U10603 ( .B1(n6394), .B2(n9401), .A(n9335), .ZN(P1_U3549) );
  AOI21_X1 U10604 ( .B1(n9567), .B2(n9337), .A(n9336), .ZN(n9338) );
  OAI211_X1 U10605 ( .C1(n9340), .C2(n9571), .A(n9339), .B(n9338), .ZN(n9413)
         );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9413), .S(n9608), .Z(
        P1_U3548) );
  AOI211_X1 U10607 ( .C1(n9567), .C2(n9343), .A(n9342), .B(n9341), .ZN(n9344)
         );
  OAI21_X1 U10608 ( .B1(n9345), .B2(n9571), .A(n9344), .ZN(n9414) );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9414), .S(n9608), .Z(
        P1_U3547) );
  AOI211_X1 U10610 ( .C1(n9567), .C2(n9348), .A(n9347), .B(n9346), .ZN(n9349)
         );
  OAI21_X1 U10611 ( .B1(n9350), .B2(n9571), .A(n9349), .ZN(n9415) );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9415), .S(n9608), .Z(
        P1_U3546) );
  OAI211_X1 U10613 ( .C1(n9353), .C2(n9571), .A(n9352), .B(n9351), .ZN(n9416)
         );
  MUX2_X1 U10614 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9416), .S(n9608), .Z(n9354) );
  INV_X1 U10615 ( .A(n9354), .ZN(n9355) );
  OAI21_X1 U10616 ( .B1(n6393), .B2(n9401), .A(n9355), .ZN(P1_U3545) );
  AOI21_X1 U10617 ( .B1(n9567), .B2(n9357), .A(n9356), .ZN(n9358) );
  OAI211_X1 U10618 ( .C1(n9360), .C2(n9571), .A(n9359), .B(n9358), .ZN(n9420)
         );
  MUX2_X1 U10619 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9420), .S(n9608), .Z(
        P1_U3544) );
  INV_X1 U10620 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9364) );
  AOI211_X1 U10621 ( .C1(n9363), .C2(n9595), .A(n9362), .B(n9361), .ZN(n9421)
         );
  MUX2_X1 U10622 ( .A(n9364), .B(n9421), .S(n9608), .Z(n9365) );
  OAI21_X1 U10623 ( .B1(n9424), .B2(n9401), .A(n9365), .ZN(P1_U3543) );
  AOI211_X1 U10624 ( .C1(n9567), .C2(n9368), .A(n9367), .B(n9366), .ZN(n9369)
         );
  OAI21_X1 U10625 ( .B1(n9370), .B2(n9571), .A(n9369), .ZN(n9425) );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9425), .S(n9608), .Z(
        P1_U3542) );
  OAI211_X1 U10627 ( .C1(n9373), .C2(n9571), .A(n9372), .B(n9371), .ZN(n9426)
         );
  INV_X1 U10628 ( .A(n9426), .ZN(n9374) );
  MUX2_X1 U10629 ( .A(n9375), .B(n9374), .S(n9608), .Z(n9376) );
  OAI21_X1 U10630 ( .B1(n9429), .B2(n9401), .A(n9376), .ZN(P1_U3541) );
  AOI211_X1 U10631 ( .C1(n9567), .C2(n9379), .A(n9378), .B(n9377), .ZN(n9380)
         );
  OAI21_X1 U10632 ( .B1(n9381), .B2(n9571), .A(n9380), .ZN(n9430) );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9430), .S(n9608), .Z(
        P1_U3540) );
  AOI211_X1 U10634 ( .C1(n9567), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9385)
         );
  OAI21_X1 U10635 ( .B1(n9386), .B2(n9571), .A(n9385), .ZN(n9431) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9431), .S(n9608), .Z(
        P1_U3539) );
  AOI211_X1 U10637 ( .C1(n9567), .C2(n9389), .A(n9388), .B(n9387), .ZN(n9390)
         );
  OAI21_X1 U10638 ( .B1(n9391), .B2(n9571), .A(n9390), .ZN(n9432) );
  MUX2_X1 U10639 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9432), .S(n9608), .Z(
        P1_U3538) );
  AOI211_X1 U10640 ( .C1(n9394), .C2(n9595), .A(n9393), .B(n9392), .ZN(n9433)
         );
  MUX2_X1 U10641 ( .A(n9874), .B(n9433), .S(n9608), .Z(n9395) );
  OAI21_X1 U10642 ( .B1(n9436), .B2(n9401), .A(n9395), .ZN(P1_U3537) );
  AOI211_X1 U10643 ( .C1(n9398), .C2(n9595), .A(n9397), .B(n9396), .ZN(n9437)
         );
  MUX2_X1 U10644 ( .A(n9399), .B(n9437), .S(n9608), .Z(n9400) );
  OAI21_X1 U10645 ( .B1(n9441), .B2(n9401), .A(n9400), .ZN(P1_U3536) );
  MUX2_X1 U10646 ( .A(n9403), .B(n9402), .S(n9598), .Z(n9404) );
  OAI21_X1 U10647 ( .B1(n9405), .B2(n9440), .A(n9404), .ZN(P1_U3521) );
  MUX2_X1 U10648 ( .A(n6416), .B(n9406), .S(n9598), .Z(n9407) );
  OAI21_X1 U10649 ( .B1(n9408), .B2(n9440), .A(n9407), .ZN(P1_U3520) );
  MUX2_X1 U10650 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9409), .S(n9598), .Z(
        P1_U3518) );
  INV_X1 U10651 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U10652 ( .A(n9411), .B(n9410), .S(n9598), .Z(n9412) );
  OAI21_X1 U10653 ( .B1(n6394), .B2(n9440), .A(n9412), .ZN(P1_U3517) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9413), .S(n9598), .Z(
        P1_U3516) );
  MUX2_X1 U10655 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9414), .S(n9598), .Z(
        P1_U3515) );
  MUX2_X1 U10656 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9415), .S(n9598), .Z(
        P1_U3514) );
  INV_X1 U10657 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9418) );
  INV_X1 U10658 ( .A(n9416), .ZN(n9417) );
  MUX2_X1 U10659 ( .A(n9418), .B(n9417), .S(n9598), .Z(n9419) );
  OAI21_X1 U10660 ( .B1(n6393), .B2(n9440), .A(n9419), .ZN(P1_U3513) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9420), .S(n9598), .Z(
        P1_U3512) );
  INV_X1 U10662 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9422) );
  MUX2_X1 U10663 ( .A(n9422), .B(n9421), .S(n9598), .Z(n9423) );
  OAI21_X1 U10664 ( .B1(n9424), .B2(n9440), .A(n9423), .ZN(P1_U3511) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9425), .S(n9598), .Z(
        P1_U3510) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9426), .S(n9598), .Z(n9427) );
  INV_X1 U10667 ( .A(n9427), .ZN(n9428) );
  OAI21_X1 U10668 ( .B1(n9429), .B2(n9440), .A(n9428), .ZN(P1_U3509) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9430), .S(n9598), .Z(
        P1_U3507) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9431), .S(n9598), .Z(
        P1_U3504) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9432), .S(n9598), .Z(
        P1_U3501) );
  INV_X1 U10672 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9434) );
  MUX2_X1 U10673 ( .A(n9434), .B(n9433), .S(n9598), .Z(n9435) );
  OAI21_X1 U10674 ( .B1(n9436), .B2(n9440), .A(n9435), .ZN(P1_U3498) );
  INV_X1 U10675 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U10676 ( .A(n9438), .B(n9437), .S(n9598), .Z(n9439) );
  OAI21_X1 U10677 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(P1_U3495) );
  MUX2_X1 U10678 ( .A(n9442), .B(P1_D_REG_1__SCAN_IN), .S(n9550), .Z(P1_U3440)
         );
  MUX2_X1 U10679 ( .A(n9443), .B(P1_D_REG_0__SCAN_IN), .S(n9550), .Z(P1_U3439)
         );
  NOR4_X1 U10680 ( .A1(n9444), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5992), .A4(
        P1_U3086), .ZN(n9445) );
  AOI21_X1 U10681 ( .B1(n9446), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9445), .ZN(
        n9447) );
  OAI21_X1 U10682 ( .B1(n9448), .B2(n7960), .A(n9447), .ZN(P1_U3324) );
  MUX2_X1 U10683 ( .A(n9449), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10684 ( .C1(n9452), .C2(n9451), .A(n9450), .B(n9522), .ZN(n9457)
         );
  AOI211_X1 U10685 ( .C1(n9455), .C2(n9454), .A(n9453), .B(n9526), .ZN(n9456)
         );
  AOI211_X1 U10686 ( .C1(n9881), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9460)
         );
  OAI211_X1 U10687 ( .C1(n9892), .C2(n9461), .A(n9460), .B(n9459), .ZN(
        P1_U3253) );
  AOI21_X1 U10688 ( .B1(n9463), .B2(n9462), .A(n9522), .ZN(n9471) );
  OAI21_X1 U10689 ( .B1(n9465), .B2(n9464), .A(n9885), .ZN(n9468) );
  OAI22_X1 U10690 ( .A1(n9468), .A2(n9467), .B1(n9466), .B2(n9502), .ZN(n9469)
         );
  AOI21_X1 U10691 ( .B1(n9471), .B2(n9470), .A(n9469), .ZN(n9473) );
  OAI211_X1 U10692 ( .C1(n9892), .C2(n9474), .A(n9473), .B(n9472), .ZN(
        P1_U3250) );
  NAND2_X1 U10693 ( .A1(n9476), .A2(n9475), .ZN(n9479) );
  INV_X1 U10694 ( .A(n9477), .ZN(n9478) );
  NAND3_X1 U10695 ( .A1(n9879), .A2(n9479), .A3(n9478), .ZN(n9487) );
  NAND2_X1 U10696 ( .A1(n9881), .A2(n9480), .ZN(n9486) );
  AOI21_X1 U10697 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9484) );
  NAND2_X1 U10698 ( .A1(n9885), .A2(n9484), .ZN(n9485) );
  AND3_X1 U10699 ( .A1(n9487), .A2(n9486), .A3(n9485), .ZN(n9489) );
  OAI211_X1 U10700 ( .C1(n9892), .C2(n9905), .A(n9489), .B(n9488), .ZN(
        P1_U3251) );
  INV_X1 U10701 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9950) );
  XOR2_X1 U10702 ( .A(n9950), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10703 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10704 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9507) );
  AOI21_X1 U10705 ( .B1(n9492), .B2(n9491), .A(n9490), .ZN(n9493) );
  NAND2_X1 U10706 ( .A1(n9879), .A2(n9493), .ZN(n9500) );
  NAND2_X1 U10707 ( .A1(n9495), .A2(n9494), .ZN(n9498) );
  INV_X1 U10708 ( .A(n9496), .ZN(n9497) );
  NAND3_X1 U10709 ( .A1(n9885), .A2(n9498), .A3(n9497), .ZN(n9499) );
  OAI211_X1 U10710 ( .C1(n9502), .C2(n9501), .A(n9500), .B(n9499), .ZN(n9503)
         );
  INV_X1 U10711 ( .A(n9503), .ZN(n9506) );
  INV_X1 U10712 ( .A(n9504), .ZN(n9505) );
  OAI211_X1 U10713 ( .C1(n9892), .C2(n9507), .A(n9506), .B(n9505), .ZN(
        P1_U3254) );
  AOI211_X1 U10714 ( .C1(n9510), .C2(n9509), .A(n9508), .B(n9522), .ZN(n9515)
         );
  AOI211_X1 U10715 ( .C1(n9513), .C2(n9512), .A(n9511), .B(n9526), .ZN(n9514)
         );
  AOI211_X1 U10716 ( .C1(n9881), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9518)
         );
  NAND2_X1 U10717 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9517) );
  OAI211_X1 U10718 ( .C1(n9892), .C2(n9519), .A(n9518), .B(n9517), .ZN(
        P1_U3256) );
  INV_X1 U10719 ( .A(n9520), .ZN(n9525) );
  INV_X1 U10720 ( .A(n9521), .ZN(n9524) );
  AOI211_X1 U10721 ( .C1(n9525), .C2(n9524), .A(n9523), .B(n9522), .ZN(n9531)
         );
  AOI211_X1 U10722 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9530)
         );
  AOI211_X1 U10723 ( .C1(n9881), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9534)
         );
  OAI211_X1 U10724 ( .C1(n9892), .C2(n9535), .A(n9534), .B(n9533), .ZN(
        P1_U3257) );
  NAND2_X1 U10725 ( .A1(n9537), .A2(n4265), .ZN(n9541) );
  AOI22_X1 U10726 ( .A1(n9317), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9539), .B2(
        n9538), .ZN(n9540) );
  OAI211_X1 U10727 ( .C1(n9543), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9544)
         );
  AOI21_X1 U10728 ( .B1(n9546), .B2(n9545), .A(n9544), .ZN(n9547) );
  OAI21_X1 U10729 ( .B1(n9317), .B2(n9548), .A(n9547), .ZN(P1_U3288) );
  INV_X1 U10730 ( .A(n9550), .ZN(n9549) );
  INV_X1 U10731 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9961) );
  NOR2_X1 U10732 ( .A1(n9549), .A2(n9961), .ZN(P1_U3294) );
  AND2_X1 U10733 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9550), .ZN(P1_U3295) );
  AND2_X1 U10734 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9550), .ZN(P1_U3296) );
  INV_X1 U10735 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10017) );
  NOR2_X1 U10736 ( .A1(n9549), .A2(n10017), .ZN(P1_U3297) );
  AND2_X1 U10737 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9550), .ZN(P1_U3298) );
  AND2_X1 U10738 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9550), .ZN(P1_U3299) );
  AND2_X1 U10739 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9550), .ZN(P1_U3300) );
  AND2_X1 U10740 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9550), .ZN(P1_U3301) );
  AND2_X1 U10741 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9550), .ZN(P1_U3302) );
  AND2_X1 U10742 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9550), .ZN(P1_U3303) );
  AND2_X1 U10743 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9550), .ZN(P1_U3304) );
  INV_X1 U10744 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U10745 ( .A1(n9549), .A2(n10018), .ZN(P1_U3305) );
  AND2_X1 U10746 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9550), .ZN(P1_U3306) );
  AND2_X1 U10747 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9550), .ZN(P1_U3307) );
  AND2_X1 U10748 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9550), .ZN(P1_U3308) );
  AND2_X1 U10749 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9550), .ZN(P1_U3309) );
  AND2_X1 U10750 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9550), .ZN(P1_U3310) );
  AND2_X1 U10751 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9550), .ZN(P1_U3311) );
  AND2_X1 U10752 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9550), .ZN(P1_U3312) );
  AND2_X1 U10753 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9550), .ZN(P1_U3313) );
  INV_X1 U10754 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U10755 ( .A1(n9549), .A2(n9982), .ZN(P1_U3314) );
  AND2_X1 U10756 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9550), .ZN(P1_U3315) );
  AND2_X1 U10757 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9550), .ZN(P1_U3316) );
  AND2_X1 U10758 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9550), .ZN(P1_U3317) );
  AND2_X1 U10759 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9550), .ZN(P1_U3318) );
  AND2_X1 U10760 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9550), .ZN(P1_U3319) );
  AND2_X1 U10761 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9550), .ZN(P1_U3320) );
  AND2_X1 U10762 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9550), .ZN(P1_U3321) );
  AND2_X1 U10763 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9550), .ZN(P1_U3322) );
  AND2_X1 U10764 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9550), .ZN(P1_U3323) );
  INV_X1 U10765 ( .A(n9551), .ZN(n9555) );
  AOI21_X1 U10766 ( .B1(n9571), .B2(n9553), .A(n9552), .ZN(n9554) );
  AOI211_X1 U10767 ( .C1(n9557), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9599)
         );
  INV_X1 U10768 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9558) );
  AOI22_X1 U10769 ( .A1(n9598), .A2(n9599), .B1(n9558), .B2(n9589), .ZN(
        P1_U3453) );
  OAI21_X1 U10770 ( .B1(n9560), .B2(n9592), .A(n9559), .ZN(n9562) );
  AOI211_X1 U10771 ( .C1(n9564), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9600)
         );
  AOI22_X1 U10772 ( .A1(n9598), .A2(n9600), .B1(n5752), .B2(n9589), .ZN(
        P1_U3459) );
  AOI21_X1 U10773 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(n9568) );
  OAI211_X1 U10774 ( .C1(n9571), .C2(n9570), .A(n9569), .B(n9568), .ZN(n9572)
         );
  INV_X1 U10775 ( .A(n9572), .ZN(n9601) );
  INV_X1 U10776 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9573) );
  AOI22_X1 U10777 ( .A1(n9598), .A2(n9601), .B1(n9573), .B2(n9589), .ZN(
        P1_U3465) );
  OAI21_X1 U10778 ( .B1(n9575), .B2(n9592), .A(n9574), .ZN(n9577) );
  AOI211_X1 U10779 ( .C1(n9595), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9602)
         );
  INV_X1 U10780 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9579) );
  AOI22_X1 U10781 ( .A1(n9598), .A2(n9602), .B1(n9579), .B2(n9589), .ZN(
        P1_U3471) );
  OAI21_X1 U10782 ( .B1(n4515), .B2(n9592), .A(n9580), .ZN(n9581) );
  AOI211_X1 U10783 ( .C1(n9583), .C2(n9595), .A(n9582), .B(n9581), .ZN(n9604)
         );
  INV_X1 U10784 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9584) );
  AOI22_X1 U10785 ( .A1(n9598), .A2(n9604), .B1(n9584), .B2(n9589), .ZN(
        P1_U3480) );
  OAI21_X1 U10786 ( .B1(n6356), .B2(n9592), .A(n9585), .ZN(n9586) );
  AOI211_X1 U10787 ( .C1(n9588), .C2(n9595), .A(n9587), .B(n9586), .ZN(n9606)
         );
  AOI22_X1 U10788 ( .A1(n9598), .A2(n9606), .B1(n5926), .B2(n9589), .ZN(
        P1_U3483) );
  OAI211_X1 U10789 ( .C1(n9593), .C2(n9592), .A(n9591), .B(n9590), .ZN(n9594)
         );
  AOI21_X1 U10790 ( .B1(n9596), .B2(n9595), .A(n9594), .ZN(n9607) );
  INV_X1 U10791 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9597) );
  AOI22_X1 U10792 ( .A1(n9598), .A2(n9607), .B1(n9597), .B2(n9589), .ZN(
        P1_U3486) );
  AOI22_X1 U10793 ( .A1(n9608), .A2(n9599), .B1(n5723), .B2(n9605), .ZN(
        P1_U3522) );
  AOI22_X1 U10794 ( .A1(n9608), .A2(n9600), .B1(n6544), .B2(n9605), .ZN(
        P1_U3524) );
  AOI22_X1 U10795 ( .A1(n9608), .A2(n9601), .B1(n5793), .B2(n9605), .ZN(
        P1_U3526) );
  AOI22_X1 U10796 ( .A1(n9608), .A2(n9602), .B1(n5830), .B2(n9605), .ZN(
        P1_U3528) );
  AOI22_X1 U10797 ( .A1(n9608), .A2(n9604), .B1(n9603), .B2(n9605), .ZN(
        P1_U3531) );
  AOI22_X1 U10798 ( .A1(n9608), .A2(n9606), .B1(n6671), .B2(n9605), .ZN(
        P1_U3532) );
  AOI22_X1 U10799 ( .A1(n9608), .A2(n9607), .B1(n6674), .B2(n9605), .ZN(
        P1_U3533) );
  AOI22_X1 U10800 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n9743), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9613) );
  XNOR2_X1 U10801 ( .A(n9609), .B(n9614), .ZN(n9610) );
  OAI21_X1 U10802 ( .B1(n9611), .B2(n9750), .A(n9610), .ZN(n9612) );
  OAI211_X1 U10803 ( .C1(n9766), .C2(n9614), .A(n9613), .B(n9612), .ZN(
        P2_U3182) );
  OAI21_X1 U10804 ( .B1(n9616), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9615), .ZN(
        n9620) );
  OAI21_X1 U10805 ( .B1(n9618), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9617), .ZN(
        n9619) );
  AOI22_X1 U10806 ( .A1(n9737), .A2(n9620), .B1(n9619), .B2(n9762), .ZN(n9629)
         );
  AOI211_X1 U10807 ( .C1(n9624), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9625)
         );
  AOI211_X1 U10808 ( .C1(n9627), .C2(n9696), .A(n9626), .B(n9625), .ZN(n9628)
         );
  OAI211_X1 U10809 ( .C1(n9664), .C2(n9630), .A(n9629), .B(n9628), .ZN(
        P2_U3187) );
  OAI21_X1 U10810 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9638) );
  OAI21_X1 U10811 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9637) );
  AOI22_X1 U10812 ( .A1(n9737), .A2(n9638), .B1(n9762), .B2(n9637), .ZN(n9647)
         );
  OAI21_X1 U10813 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9642) );
  AOI22_X1 U10814 ( .A1(n9743), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(n9750), .B2(
        n9642), .ZN(n9646) );
  NAND2_X1 U10815 ( .A1(n9643), .A2(n9696), .ZN(n9644) );
  NAND4_X1 U10816 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(
        P2_U3188) );
  OAI21_X1 U10817 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n9649), .A(n9648), .ZN(
        n9653) );
  OAI21_X1 U10818 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n9651), .A(n9650), .ZN(
        n9652) );
  AOI22_X1 U10819 ( .A1(n9653), .A2(n9737), .B1(n9652), .B2(n9762), .ZN(n9662)
         );
  OAI21_X1 U10820 ( .B1(n9656), .B2(n9655), .A(n9654), .ZN(n9657) );
  AND2_X1 U10821 ( .A1(n9657), .A2(n9750), .ZN(n9658) );
  AOI211_X1 U10822 ( .C1(n9660), .C2(n9696), .A(n9659), .B(n9658), .ZN(n9661)
         );
  OAI211_X1 U10823 ( .C1(n9664), .C2(n9663), .A(n9662), .B(n9661), .ZN(
        P2_U3189) );
  OAI21_X1 U10824 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9669) );
  AOI22_X1 U10825 ( .A1(n9669), .A2(n9737), .B1(n9668), .B2(n9696), .ZN(n9681)
         );
  OAI21_X1 U10826 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9673) );
  AOI22_X1 U10827 ( .A1(n9743), .A2(P2_ADDR_REG_8__SCAN_IN), .B1(n9750), .B2(
        n9673), .ZN(n9680) );
  OAI21_X1 U10828 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(n9677) );
  NAND2_X1 U10829 ( .A1(n9677), .A2(n9762), .ZN(n9678) );
  NAND4_X1 U10830 ( .A1(n9681), .A2(n9680), .A3(n9679), .A4(n9678), .ZN(
        P2_U3190) );
  AOI21_X1 U10831 ( .B1(n9743), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9682), .ZN(
        n9694) );
  OAI21_X1 U10832 ( .B1(n9684), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9683), .ZN(
        n9692) );
  OAI21_X1 U10833 ( .B1(n9686), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9685), .ZN(
        n9691) );
  OAI21_X1 U10834 ( .B1(n9689), .B2(n9688), .A(n9687), .ZN(n9690) );
  AOI222_X1 U10835 ( .A1(n9692), .A2(n9737), .B1(n9691), .B2(n9762), .C1(n9690), .C2(n9750), .ZN(n9693) );
  OAI211_X1 U10836 ( .C1(n9766), .C2(n9695), .A(n9694), .B(n9693), .ZN(
        P2_U3191) );
  AOI22_X1 U10837 ( .A1(n9697), .A2(n9696), .B1(n9743), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n9712) );
  OAI21_X1 U10838 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9709) );
  OAI21_X1 U10839 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9708) );
  OAI21_X1 U10840 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  AOI222_X1 U10841 ( .A1(n9709), .A2(n9737), .B1(n9708), .B2(n9762), .C1(n9707), .C2(n9750), .ZN(n9711) );
  NAND3_X1 U10842 ( .A1(n9712), .A2(n9711), .A3(n9710), .ZN(P2_U3192) );
  AOI21_X1 U10843 ( .B1(n9743), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9713), .ZN(
        n9725) );
  OAI21_X1 U10844 ( .B1(n9715), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9714), .ZN(
        n9723) );
  OAI21_X1 U10845 ( .B1(n9717), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9716), .ZN(
        n9722) );
  OAI21_X1 U10846 ( .B1(n9720), .B2(n9719), .A(n9718), .ZN(n9721) );
  AOI222_X1 U10847 ( .A1(n9723), .A2(n9737), .B1(n9722), .B2(n9762), .C1(n9721), .C2(n9750), .ZN(n9724) );
  OAI211_X1 U10848 ( .C1(n9766), .C2(n9726), .A(n9725), .B(n9724), .ZN(
        P2_U3193) );
  AOI21_X1 U10849 ( .B1(n9743), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n9727), .ZN(
        n9740) );
  OAI21_X1 U10850 ( .B1(n9729), .B2(P2_REG2_REG_13__SCAN_IN), .A(n9728), .ZN(
        n9738) );
  OAI21_X1 U10851 ( .B1(n9731), .B2(P2_REG1_REG_13__SCAN_IN), .A(n9730), .ZN(
        n9736) );
  OAI21_X1 U10852 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  AOI222_X1 U10853 ( .A1(n9738), .A2(n9737), .B1(n9736), .B2(n9762), .C1(n9735), .C2(n9750), .ZN(n9739) );
  OAI211_X1 U10854 ( .C1(n9766), .C2(n9741), .A(n9740), .B(n9739), .ZN(
        P2_U3195) );
  AOI21_X1 U10855 ( .B1(n9743), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n9742), .ZN(
        n9764) );
  OAI21_X1 U10856 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9761) );
  OAI21_X1 U10857 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9751) );
  AND2_X1 U10858 ( .A1(n9751), .A2(n9750), .ZN(n9760) );
  OAI21_X1 U10859 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9757) );
  NOR2_X1 U10860 ( .A1(n9758), .A2(n9757), .ZN(n9756) );
  AOI211_X1 U10861 ( .C1(n9758), .C2(n9757), .A(n9756), .B(n9755), .ZN(n9759)
         );
  AOI211_X1 U10862 ( .C1(n9762), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9763)
         );
  OAI211_X1 U10863 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(
        P2_U3196) );
  INV_X1 U10864 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9772) );
  INV_X1 U10865 ( .A(n9808), .ZN(n9823) );
  AOI21_X1 U10866 ( .B1(n9768), .B2(n9823), .A(n9767), .ZN(n9769) );
  AOI211_X1 U10867 ( .C1(n9828), .C2(n9771), .A(n9770), .B(n9769), .ZN(n9833)
         );
  AOI22_X1 U10868 ( .A1(n9831), .A2(n9772), .B1(n9833), .B2(n9829), .ZN(
        P2_U3390) );
  INV_X1 U10869 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9947) );
  OAI22_X1 U10870 ( .A1(n9774), .A2(n9818), .B1(n9773), .B2(n9816), .ZN(n9775)
         );
  NOR2_X1 U10871 ( .A1(n9776), .A2(n9775), .ZN(n9835) );
  AOI22_X1 U10872 ( .A1(n9831), .A2(n9947), .B1(n9835), .B2(n9829), .ZN(
        P2_U3396) );
  INV_X1 U10873 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9782) );
  INV_X1 U10874 ( .A(n9777), .ZN(n9781) );
  OAI22_X1 U10875 ( .A1(n9779), .A2(n9823), .B1(n9778), .B2(n9816), .ZN(n9780)
         );
  NOR2_X1 U10876 ( .A1(n9781), .A2(n9780), .ZN(n9837) );
  AOI22_X1 U10877 ( .A1(n9831), .A2(n9782), .B1(n9837), .B2(n9829), .ZN(
        P2_U3399) );
  INV_X1 U10878 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9787) );
  INV_X1 U10879 ( .A(n9783), .ZN(n9786) );
  OAI22_X1 U10880 ( .A1(n9784), .A2(n9823), .B1(n4735), .B2(n9816), .ZN(n9785)
         );
  NOR2_X1 U10881 ( .A1(n9786), .A2(n9785), .ZN(n9838) );
  AOI22_X1 U10882 ( .A1(n9831), .A2(n9787), .B1(n9838), .B2(n9829), .ZN(
        P2_U3402) );
  INV_X1 U10883 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9793) );
  OAI22_X1 U10884 ( .A1(n9789), .A2(n9823), .B1(n9788), .B2(n9816), .ZN(n9792)
         );
  INV_X1 U10885 ( .A(n9790), .ZN(n9791) );
  NOR2_X1 U10886 ( .A1(n9792), .A2(n9791), .ZN(n9839) );
  AOI22_X1 U10887 ( .A1(n9831), .A2(n9793), .B1(n9839), .B2(n9829), .ZN(
        P2_U3405) );
  INV_X1 U10888 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9931) );
  OAI22_X1 U10889 ( .A1(n9795), .A2(n9823), .B1(n9794), .B2(n9816), .ZN(n9797)
         );
  NOR2_X1 U10890 ( .A1(n9797), .A2(n9796), .ZN(n9841) );
  AOI22_X1 U10891 ( .A1(n9831), .A2(n9931), .B1(n9841), .B2(n9829), .ZN(
        P2_U3408) );
  INV_X1 U10892 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U10893 ( .A1(n9798), .A2(n9816), .ZN(n9800) );
  AOI211_X1 U10894 ( .C1(n9808), .C2(n9801), .A(n9800), .B(n9799), .ZN(n9843)
         );
  AOI22_X1 U10895 ( .A1(n9831), .A2(n9802), .B1(n9843), .B2(n9829), .ZN(
        P2_U3411) );
  INV_X1 U10896 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9809) );
  INV_X1 U10897 ( .A(n9803), .ZN(n9807) );
  OAI21_X1 U10898 ( .B1(n9805), .B2(n9816), .A(n9804), .ZN(n9806) );
  AOI21_X1 U10899 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9845) );
  AOI22_X1 U10900 ( .A1(n9831), .A2(n9809), .B1(n9845), .B2(n9829), .ZN(
        P2_U3414) );
  INV_X1 U10901 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9987) );
  NOR2_X1 U10902 ( .A1(n9810), .A2(n9816), .ZN(n9811) );
  AOI21_X1 U10903 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  AND2_X1 U10904 ( .A1(n9815), .A2(n9814), .ZN(n9846) );
  AOI22_X1 U10905 ( .A1(n9831), .A2(n9987), .B1(n9846), .B2(n9829), .ZN(
        P2_U3417) );
  INV_X1 U10906 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9822) );
  OAI22_X1 U10907 ( .A1(n9819), .A2(n9818), .B1(n9817), .B2(n9816), .ZN(n9820)
         );
  NOR2_X1 U10908 ( .A1(n9821), .A2(n9820), .ZN(n9847) );
  AOI22_X1 U10909 ( .A1(n9831), .A2(n9822), .B1(n9847), .B2(n9829), .ZN(
        P2_U3420) );
  INV_X1 U10910 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U10911 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  AOI211_X1 U10912 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9850)
         );
  AOI22_X1 U10913 ( .A1(n9831), .A2(n9830), .B1(n9850), .B2(n9829), .ZN(
        P2_U3423) );
  AOI22_X1 U10914 ( .A1(n9851), .A2(n9833), .B1(n9832), .B2(n9848), .ZN(
        P2_U3459) );
  AOI22_X1 U10915 ( .A1(n9851), .A2(n9835), .B1(n9834), .B2(n9848), .ZN(
        P2_U3461) );
  INV_X1 U10916 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10917 ( .A1(n9851), .A2(n9837), .B1(n9836), .B2(n9848), .ZN(
        P2_U3462) );
  AOI22_X1 U10918 ( .A1(n9851), .A2(n9838), .B1(n9951), .B2(n9848), .ZN(
        P2_U3463) );
  AOI22_X1 U10919 ( .A1(n9851), .A2(n9839), .B1(n7267), .B2(n9848), .ZN(
        P2_U3464) );
  AOI22_X1 U10920 ( .A1(n9851), .A2(n9841), .B1(n9840), .B2(n9848), .ZN(
        P2_U3465) );
  INV_X1 U10921 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10922 ( .A1(n9851), .A2(n9843), .B1(n9842), .B2(n9848), .ZN(
        P2_U3466) );
  AOI22_X1 U10923 ( .A1(n9851), .A2(n9845), .B1(n9844), .B2(n9848), .ZN(
        P2_U3467) );
  INV_X1 U10924 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U10925 ( .A1(n9851), .A2(n9846), .B1(n9917), .B2(n9848), .ZN(
        P2_U3468) );
  AOI22_X1 U10926 ( .A1(n9851), .A2(n9847), .B1(n7223), .B2(n9848), .ZN(
        P2_U3469) );
  INV_X1 U10927 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9849) );
  AOI22_X1 U10928 ( .A1(n9851), .A2(n9850), .B1(n9849), .B2(n9848), .ZN(
        P2_U3470) );
  NOR2_X1 U10929 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  XOR2_X1 U10930 ( .A(n9854), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  XOR2_X1 U10931 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10932 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  XOR2_X1 U10933 ( .A(n9857), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55) );
  XNOR2_X1 U10934 ( .A(n9859), .B(n9858), .ZN(ADD_1068_U56) );
  XNOR2_X1 U10935 ( .A(n9861), .B(n9860), .ZN(ADD_1068_U57) );
  XNOR2_X1 U10936 ( .A(n9863), .B(n9862), .ZN(ADD_1068_U58) );
  XNOR2_X1 U10937 ( .A(n9865), .B(n9864), .ZN(ADD_1068_U59) );
  XNOR2_X1 U10938 ( .A(n9867), .B(n9866), .ZN(ADD_1068_U60) );
  XNOR2_X1 U10939 ( .A(n9869), .B(n9868), .ZN(ADD_1068_U61) );
  XNOR2_X1 U10940 ( .A(n9871), .B(n9870), .ZN(ADD_1068_U62) );
  XNOR2_X1 U10941 ( .A(n9873), .B(n9872), .ZN(ADD_1068_U63) );
  NAND2_X1 U10942 ( .A1(n9875), .A2(n9874), .ZN(n9878) );
  INV_X1 U10943 ( .A(n9876), .ZN(n9877) );
  NAND3_X1 U10944 ( .A1(n9879), .A2(n9878), .A3(n9877), .ZN(n9888) );
  NAND2_X1 U10945 ( .A1(n9881), .A2(n9880), .ZN(n9887) );
  AOI21_X1 U10946 ( .B1(n9883), .B2(n9311), .A(n9882), .ZN(n9884) );
  NAND2_X1 U10947 ( .A1(n9885), .A2(n9884), .ZN(n9886) );
  AND3_X1 U10948 ( .A1(n9888), .A2(n9887), .A3(n9886), .ZN(n9890) );
  NAND2_X1 U10949 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9889) );
  OAI211_X1 U10950 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9889), .ZN(n10038)
         );
  AOI22_X1 U10951 ( .A1(n10012), .A2(keyinput46), .B1(keyinput55), .B2(n9894), 
        .ZN(n9893) );
  OAI221_X1 U10952 ( .B1(n10012), .B2(keyinput46), .C1(n9894), .C2(keyinput55), 
        .A(n9893), .ZN(n9903) );
  INV_X1 U10953 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10019) );
  AOI22_X1 U10954 ( .A1(n10019), .A2(keyinput33), .B1(keyinput21), .B2(n9896), 
        .ZN(n9895) );
  OAI221_X1 U10955 ( .B1(n10019), .B2(keyinput33), .C1(n9896), .C2(keyinput21), 
        .A(n9895), .ZN(n9902) );
  AOI22_X1 U10956 ( .A1(n10010), .A2(keyinput0), .B1(n5926), .B2(keyinput36), 
        .ZN(n9897) );
  OAI221_X1 U10957 ( .B1(n10010), .B2(keyinput0), .C1(n5926), .C2(keyinput36), 
        .A(n9897), .ZN(n9901) );
  XNOR2_X1 U10958 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput7), .ZN(n9899) );
  XNOR2_X1 U10959 ( .A(keyinput63), .B(P1_REG0_REG_13__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U10960 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  NOR4_X1 U10961 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9942)
         );
  AOI22_X1 U10962 ( .A1(n9906), .A2(keyinput4), .B1(keyinput19), .B2(n9905), 
        .ZN(n9904) );
  OAI221_X1 U10963 ( .B1(n9906), .B2(keyinput4), .C1(n9905), .C2(keyinput19), 
        .A(n9904), .ZN(n9916) );
  AOI22_X1 U10964 ( .A1(n9908), .A2(keyinput44), .B1(n8342), .B2(keyinput1), 
        .ZN(n9907) );
  OAI221_X1 U10965 ( .B1(n9908), .B2(keyinput44), .C1(n8342), .C2(keyinput1), 
        .A(n9907), .ZN(n9915) );
  XNOR2_X1 U10966 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput37), .ZN(n9911) );
  XNOR2_X1 U10967 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput27), .ZN(n9910) );
  XNOR2_X1 U10968 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput41), .ZN(n9909)
         );
  NAND3_X1 U10969 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(n9914) );
  XNOR2_X1 U10970 ( .A(n9912), .B(keyinput34), .ZN(n9913) );
  NOR4_X1 U10971 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n9941)
         );
  XOR2_X1 U10972 ( .A(n9917), .B(keyinput40), .Z(n9921) );
  XNOR2_X1 U10973 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput3), .ZN(n9920) );
  XNOR2_X1 U10974 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput15), .ZN(n9919) );
  XNOR2_X1 U10975 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput43), .ZN(n9918) );
  NAND4_X1 U10976 ( .A1(n9921), .A2(n9920), .A3(n9919), .A4(n9918), .ZN(n9927)
         );
  XNOR2_X1 U10977 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput48), .ZN(n9925) );
  XNOR2_X1 U10978 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput26), .ZN(n9924)
         );
  XNOR2_X1 U10979 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput22), .ZN(n9923) );
  XNOR2_X1 U10980 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput29), .ZN(n9922) );
  NAND4_X1 U10981 ( .A1(n9925), .A2(n9924), .A3(n9923), .A4(n9922), .ZN(n9926)
         );
  NOR2_X1 U10982 ( .A1(n9927), .A2(n9926), .ZN(n9940) );
  AOI22_X1 U10983 ( .A1(n9929), .A2(keyinput2), .B1(n9165), .B2(keyinput57), 
        .ZN(n9928) );
  OAI221_X1 U10984 ( .B1(n9929), .B2(keyinput2), .C1(n9165), .C2(keyinput57), 
        .A(n9928), .ZN(n9938) );
  AOI22_X1 U10985 ( .A1(n9931), .A2(keyinput17), .B1(n6181), .B2(keyinput39), 
        .ZN(n9930) );
  OAI221_X1 U10986 ( .B1(n9931), .B2(keyinput17), .C1(n6181), .C2(keyinput39), 
        .A(n9930), .ZN(n9937) );
  XNOR2_X1 U10987 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput10), .ZN(n9935) );
  XNOR2_X1 U10988 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput62), .ZN(n9934) );
  XNOR2_X1 U10989 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput49), .ZN(n9933) );
  XNOR2_X1 U10990 ( .A(P2_B_REG_SCAN_IN), .B(keyinput60), .ZN(n9932) );
  NAND4_X1 U10991 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(n9936)
         );
  NOR3_X1 U10992 ( .A1(n9938), .A2(n9937), .A3(n9936), .ZN(n9939) );
  NAND4_X1 U10993 ( .A1(n9942), .A2(n9941), .A3(n9940), .A4(n9939), .ZN(n10003) );
  AOI22_X1 U10994 ( .A1(n9945), .A2(keyinput28), .B1(keyinput54), .B2(n9944), 
        .ZN(n9943) );
  OAI221_X1 U10995 ( .B1(n9945), .B2(keyinput28), .C1(n9944), .C2(keyinput54), 
        .A(n9943), .ZN(n9957) );
  AOI22_X1 U10996 ( .A1(n9948), .A2(keyinput8), .B1(keyinput45), .B2(n9947), 
        .ZN(n9946) );
  OAI221_X1 U10997 ( .B1(n9948), .B2(keyinput8), .C1(n9947), .C2(keyinput45), 
        .A(n9946), .ZN(n9956) );
  AOI22_X1 U10998 ( .A1(n9951), .A2(keyinput23), .B1(keyinput24), .B2(n9950), 
        .ZN(n9949) );
  OAI221_X1 U10999 ( .B1(n9951), .B2(keyinput23), .C1(n9950), .C2(keyinput24), 
        .A(n9949), .ZN(n9955) );
  AOI22_X1 U11000 ( .A1(n9953), .A2(keyinput53), .B1(n9126), .B2(keyinput31), 
        .ZN(n9952) );
  OAI221_X1 U11001 ( .B1(n9953), .B2(keyinput53), .C1(n9126), .C2(keyinput31), 
        .A(n9952), .ZN(n9954) );
  NOR4_X1 U11002 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n9954), .ZN(n10001)
         );
  AOI22_X1 U11003 ( .A1(n5809), .A2(keyinput9), .B1(keyinput20), .B2(n9959), 
        .ZN(n9958) );
  OAI221_X1 U11004 ( .B1(n5809), .B2(keyinput9), .C1(n9959), .C2(keyinput20), 
        .A(n9958), .ZN(n9970) );
  AOI22_X1 U11005 ( .A1(n9961), .A2(keyinput30), .B1(keyinput58), .B2(n6416), 
        .ZN(n9960) );
  OAI221_X1 U11006 ( .B1(n9961), .B2(keyinput30), .C1(n6416), .C2(keyinput58), 
        .A(n9960), .ZN(n9969) );
  AOI22_X1 U11007 ( .A1(n9964), .A2(keyinput56), .B1(keyinput59), .B2(n9963), 
        .ZN(n9962) );
  OAI221_X1 U11008 ( .B1(n9964), .B2(keyinput56), .C1(n9963), .C2(keyinput59), 
        .A(n9962), .ZN(n9968) );
  XOR2_X1 U11009 ( .A(n6323), .B(keyinput61), .Z(n9966) );
  XNOR2_X1 U11010 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput47), .ZN(n9965) );
  NAND2_X1 U11011 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  NOR4_X1 U11012 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n9967), .ZN(n10000)
         );
  AOI22_X1 U11013 ( .A1(n7621), .A2(keyinput5), .B1(n9972), .B2(keyinput38), 
        .ZN(n9971) );
  OAI221_X1 U11014 ( .B1(n7621), .B2(keyinput5), .C1(n9972), .C2(keyinput38), 
        .A(n9971), .ZN(n9977) );
  XNOR2_X1 U11015 ( .A(n9973), .B(keyinput35), .ZN(n9976) );
  XNOR2_X1 U11016 ( .A(n9974), .B(keyinput14), .ZN(n9975) );
  OR3_X1 U11017 ( .A1(n9977), .A2(n9976), .A3(n9975), .ZN(n9985) );
  INV_X1 U11018 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11019 ( .A1(n7535), .A2(keyinput16), .B1(keyinput25), .B2(n9979), 
        .ZN(n9978) );
  OAI221_X1 U11020 ( .B1(n7535), .B2(keyinput16), .C1(n9979), .C2(keyinput25), 
        .A(n9978), .ZN(n9984) );
  AOI22_X1 U11021 ( .A1(n9982), .A2(keyinput12), .B1(keyinput51), .B2(n9981), 
        .ZN(n9980) );
  OAI221_X1 U11022 ( .B1(n9982), .B2(keyinput12), .C1(n9981), .C2(keyinput51), 
        .A(n9980), .ZN(n9983) );
  NOR3_X1 U11023 ( .A1(n9985), .A2(n9984), .A3(n9983), .ZN(n9999) );
  AOI22_X1 U11024 ( .A1(n9987), .A2(keyinput13), .B1(n10018), .B2(keyinput50), 
        .ZN(n9986) );
  OAI221_X1 U11025 ( .B1(n9987), .B2(keyinput13), .C1(n10018), .C2(keyinput50), 
        .A(n9986), .ZN(n9997) );
  AOI22_X1 U11026 ( .A1(n9989), .A2(keyinput6), .B1(n6118), .B2(keyinput52), 
        .ZN(n9988) );
  OAI221_X1 U11027 ( .B1(n9989), .B2(keyinput6), .C1(n6118), .C2(keyinput52), 
        .A(n9988), .ZN(n9996) );
  AOI22_X1 U11028 ( .A1(n10017), .A2(keyinput18), .B1(keyinput32), .B2(n9991), 
        .ZN(n9990) );
  OAI221_X1 U11029 ( .B1(n10017), .B2(keyinput18), .C1(n9991), .C2(keyinput32), 
        .A(n9990), .ZN(n9995) );
  XNOR2_X1 U11030 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput11), .ZN(n9993) );
  XNOR2_X1 U11031 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput42), .ZN(n9992) );
  NAND2_X1 U11032 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  NOR4_X1 U11033 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n9998)
         );
  NAND4_X1 U11034 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        n10002) );
  NOR2_X1 U11035 ( .A1(n10003), .A2(n10002), .ZN(n10036) );
  NOR3_X1 U11036 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(P1_IR_REG_21__SCAN_IN), .ZN(n10004) );
  NAND4_X1 U11037 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .A3(P1_IR_REG_18__SCAN_IN), .A4(n10004), .ZN(n10007) );
  INV_X1 U11038 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10006) );
  OR3_X1 U11039 ( .A1(n10007), .A2(n10006), .A3(n10005), .ZN(n10034) );
  NAND4_X1 U11040 ( .A1(n10009), .A2(n10008), .A3(P2_ADDR_REG_4__SCAN_IN), 
        .A4(P1_ADDR_REG_8__SCAN_IN), .ZN(n10033) );
  NOR4_X1 U11041 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P1_REG1_REG_29__SCAN_IN), 
        .A3(P2_REG1_REG_4__SCAN_IN), .A4(P1_REG0_REG_30__SCAN_IN), .ZN(n10016)
         );
  NOR4_X1 U11042 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(P2_IR_REG_30__SCAN_IN), .ZN(n10015)
         );
  NOR4_X1 U11043 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P2_REG2_REG_17__SCAN_IN), .A4(P2_REG2_REG_13__SCAN_IN), .ZN(n10014) );
  INV_X1 U11044 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10011) );
  NOR4_X1 U11045 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n8342), .ZN(
        n10013) );
  NAND4_X1 U11046 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10032) );
  NOR4_X1 U11047 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P2_DATAO_REG_5__SCAN_IN), .A4(P1_DATAO_REG_29__SCAN_IN), .ZN(
        n10030) );
  NOR4_X1 U11048 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(P2_REG0_REG_12__SCAN_IN), 
        .A3(P2_REG1_REG_9__SCAN_IN), .A4(P2_REG0_REG_6__SCAN_IN), .ZN(n10029)
         );
  NAND2_X1 U11049 ( .A1(n10018), .A2(n10017), .ZN(n10022) );
  NAND4_X1 U11050 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(P1_REG2_REG_12__SCAN_IN), 
        .A3(n10020), .A4(n10019), .ZN(n10021) );
  NOR4_X1 U11051 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(P2_WR_REG_SCAN_IN), .A3(
        n10022), .A4(n10021), .ZN(n10028) );
  NAND4_X1 U11052 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(P1_REG0_REG_23__SCAN_IN), 
        .A3(P1_REG3_REG_1__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n10026) );
  NAND4_X1 U11053 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(P1_REG0_REG_5__SCAN_IN), 
        .A3(P2_IR_REG_12__SCAN_IN), .A4(P2_IR_REG_27__SCAN_IN), .ZN(n10025) );
  NAND4_X1 U11054 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(P1_REG2_REG_25__SCAN_IN), .A3(P2_D_REG_10__SCAN_IN), .A4(P2_REG0_REG_2__SCAN_IN), .ZN(n10024) );
  NAND4_X1 U11055 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_13__SCAN_IN), .A3(P1_DATAO_REG_3__SCAN_IN), .A4(
        P2_REG0_REG_9__SCAN_IN), .ZN(n10023) );
  NOR4_X1 U11056 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10027) );
  NAND4_X1 U11057 ( .A1(n10030), .A2(n10029), .A3(n10028), .A4(n10027), .ZN(
        n10031) );
  NOR4_X1 U11058 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10035) );
  XNOR2_X1 U11059 ( .A(n10036), .B(n10035), .ZN(n10037) );
  XNOR2_X1 U11060 ( .A(n10038), .B(n10037), .ZN(P1_U3258) );
  XNOR2_X1 U11061 ( .A(n10040), .B(n10039), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11062 ( .A(n10042), .B(n10041), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11063 ( .A(n10044), .B(n10043), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11064 ( .A(n10046), .B(n10045), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11065 ( .A(n10048), .B(n10047), .ZN(ADD_1068_U48) );
  XOR2_X1 U11066 ( .A(n10050), .B(n10049), .Z(ADD_1068_U54) );
  XOR2_X1 U11067 ( .A(n10052), .B(n10051), .Z(ADD_1068_U53) );
  XNOR2_X1 U11068 ( .A(n10054), .B(n10053), .ZN(ADD_1068_U52) );
  NAND2_X1 U6508 ( .A1(n4266), .A2(n5048), .ZN(n5160) );
  NAND3_X2 U5832 ( .A1(n5742), .A2(n5741), .A3(n5740), .ZN(n5743) );
  NAND2_X1 U4796 ( .A1(n7764), .A2(n7758), .ZN(n7880) );
  CLKBUF_X1 U5768 ( .A(n5687), .Z(n9264) );
endmodule

