

module b22_C_SARLock_k_128_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6564, n6565, n6566, n6568, n6569, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554;

  AND2_X1 U7313 ( .A1(n13499), .A2(n13498), .ZN(n13705) );
  NAND2_X1 U7314 ( .A1(n11018), .A2(n11017), .ZN(n11052) );
  OR2_X1 U7315 ( .A1(n10618), .A2(n14660), .ZN(n14308) );
  CLKBUF_X2 U7316 ( .A(n7717), .Z(n6770) );
  NAND2_X1 U7317 ( .A1(n11983), .A2(n11982), .ZN(n10708) );
  INV_X1 U7318 ( .A(n10644), .ZN(n12749) );
  INV_X1 U7319 ( .A(n12076), .ZN(n12087) );
  AND2_X1 U7320 ( .A1(n8531), .A2(n8530), .ZN(n15084) );
  AND4_X1 U7322 ( .A1(n7710), .A2(n7709), .A3(n7708), .A4(n7707), .ZN(n10657)
         );
  NAND2_X1 U7323 ( .A1(n8574), .A2(n8575), .ZN(n10121) );
  INV_X1 U7324 ( .A(n8490), .ZN(n8449) );
  CLKBUF_X2 U7325 ( .A(n12322), .Z(n6569) );
  AND2_X1 U7326 ( .A1(n7948), .A2(n7645), .ZN(n7968) );
  CLKBUF_X2 U7328 ( .A(n11494), .Z(n6573) );
  INV_X1 U7329 ( .A(n11642), .ZN(n8436) );
  INV_X1 U7330 ( .A(n8438), .ZN(n8512) );
  INV_X1 U7331 ( .A(n11413), .ZN(n11338) );
  INV_X1 U7332 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U7333 ( .A1(n7038), .A2(n7520), .ZN(n7632) );
  OAI21_X1 U7335 ( .B1(n8420), .B2(n8421), .A(n8290), .ZN(n8461) );
  INV_X1 U7336 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14578) );
  CLKBUF_X1 U7337 ( .A(n13953), .Z(n6564) );
  OAI21_X1 U7338 ( .B1(n9373), .B2(n9363), .A(n14783), .ZN(n13953) );
  XNOR2_X1 U7339 ( .A(n6902), .B(n14519), .ZN(n14550) );
  OR2_X1 U7340 ( .A1(n14328), .A2(n7217), .ZN(n6565) );
  NAND2_X1 U7341 ( .A1(n6565), .A2(n7215), .ZN(P1_U3525) );
  XOR2_X1 U7342 ( .A(n6566), .B(P1_IR_REG_29__SCAN_IN), .Z(n9236) );
  NOR2_X1 U7343 ( .A1(n9233), .A2(n8966), .ZN(n6566) );
  NAND4_X4 U7344 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n12144)
         );
  NAND2_X2 U7345 ( .A1(n6991), .A2(n6990), .ZN(n12779) );
  NAND2_X2 U7346 ( .A1(n9571), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9615) );
  INV_X2 U7347 ( .A(n13225), .ZN(n7602) );
  INV_X2 U7348 ( .A(n11431), .ZN(n6799) );
  INV_X1 U7349 ( .A(n11351), .ZN(n11504) );
  OAI21_X1 U7350 ( .B1(n12882), .B2(n11943), .A(n10195), .ZN(n7649) );
  AOI21_X1 U7351 ( .B1(n12865), .B2(n12864), .A(n12863), .ZN(n12889) );
  INV_X1 U7352 ( .A(n7717), .ZN(n7752) );
  INV_X2 U7353 ( .A(n6770), .ZN(n9635) );
  NAND2_X1 U7354 ( .A1(n12070), .A2(n12069), .ZN(n12920) );
  INV_X1 U7355 ( .A(n11746), .ZN(n11787) );
  NAND2_X1 U7356 ( .A1(n10306), .A2(n11675), .ZN(n11190) );
  OAI21_X1 U7357 ( .B1(n7989), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7648) );
  OAI21_X1 U7359 ( .B1(n12249), .B2(n12251), .A(n11052), .ZN(n11079) );
  AND2_X1 U7360 ( .A1(n8559), .A2(n8558), .ZN(n15098) );
  INV_X1 U7361 ( .A(n11227), .ZN(n14868) );
  XNOR2_X1 U7362 ( .A(n8709), .B(SI_14_), .ZN(n8712) );
  AND3_X1 U7363 ( .A1(n7777), .A2(n7776), .A3(n7775), .ZN(n15209) );
  AND2_X1 U7364 ( .A1(n7767), .A2(n7766), .ZN(n10645) );
  NAND2_X1 U7365 ( .A1(n7992), .A2(n7991), .ZN(n13136) );
  MUX2_X1 U7366 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7624), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7628) );
  INV_X1 U7367 ( .A(n6586), .ZN(n13778) );
  INV_X2 U7368 ( .A(n8705), .ZN(n6577) );
  AND2_X1 U7369 ( .A1(n13486), .A2(n12396), .ZN(n13584) );
  NAND2_X1 U7370 ( .A1(n10118), .A2(n10117), .ZN(n11238) );
  NAND2_X2 U7371 ( .A1(n10124), .A2(n10123), .ZN(n14891) );
  NAND2_X1 U7372 ( .A1(n11464), .A2(n11463), .ZN(n14137) );
  NAND2_X1 U7373 ( .A1(n10578), .A2(n10577), .ZN(n14660) );
  NAND3_X1 U7374 ( .A1(n9313), .A2(n9314), .A3(n6627), .ZN(n11211) );
  XNOR2_X1 U7375 ( .A(n8838), .B(n8837), .ZN(n11428) );
  INV_X1 U7376 ( .A(n10645), .ZN(n12748) );
  INV_X1 U7377 ( .A(n10657), .ZN(n12750) );
  NAND2_X1 U7380 ( .A1(n13299), .A2(n12508), .ZN(n13230) );
  AOI21_X1 U7381 ( .B1(n13497), .B2(n13683), .A(n13496), .ZN(n13708) );
  INV_X1 U7382 ( .A(n8400), .ZN(n13805) );
  NAND2_X1 U7383 ( .A1(n8382), .A2(n8381), .ZN(n8879) );
  INV_X1 U7384 ( .A(n14402), .ZN(n6967) );
  BUF_X1 U7385 ( .A(n9298), .Z(n13986) );
  XNOR2_X1 U7386 ( .A(n8477), .B(n8476), .ZN(n9330) );
  NAND2_X1 U7387 ( .A1(n6588), .A2(n6576), .ZN(n8825) );
  CLKBUF_X1 U7388 ( .A(n8463), .Z(n6582) );
  AND2_X1 U7389 ( .A1(n12524), .A2(n13225), .ZN(n7758) );
  NAND4_X2 U7392 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n13985)
         );
  NAND4_X2 U7393 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n9282), .ZN(n9298)
         );
  AOI21_X2 U7394 ( .B1(n9653), .B2(n6582), .A(n7464), .ZN(n9826) );
  OAI22_X2 U7395 ( .A1(n13656), .A2(n13657), .B1(n13666), .B2(n13747), .ZN(
        n13635) );
  NAND2_X2 U7396 ( .A1(n12559), .A2(n12986), .ZN(n12558) );
  NOR2_X2 U7397 ( .A1(n8090), .A2(n8085), .ZN(n12559) );
  INV_X1 U7398 ( .A(n8399), .ZN(n11172) );
  AOI21_X2 U7399 ( .B1(n10797), .B2(n10796), .A(n6756), .ZN(n10857) );
  NAND2_X4 U7401 ( .A1(n6766), .A2(n7668), .ZN(n12752) );
  AND3_X2 U7402 ( .A1(n7670), .A2(n7667), .A3(n7669), .ZN(n6766) );
  CLKBUF_X3 U7403 ( .A(n8490), .Z(n8765) );
  NAND4_X2 U7404 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n13320)
         );
  XNOR2_X1 U7405 ( .A(n7858), .B(n7856), .ZN(n12690) );
  NAND2_X1 U7406 ( .A1(n12567), .A2(n7840), .ZN(n7858) );
  INV_X1 U7407 ( .A(n11746), .ZN(n6571) );
  INV_X1 U7408 ( .A(n11746), .ZN(n6572) );
  AND2_X1 U7409 ( .A1(n11195), .A2(n9251), .ZN(n11771) );
  BUF_X4 U7410 ( .A(n9660), .Z(n11387) );
  INV_X1 U7411 ( .A(n11181), .ZN(n11494) );
  NOR3_X2 U7412 ( .A1(n10733), .A2(n10732), .A3(n10731), .ZN(n10892) );
  NOR2_X2 U7413 ( .A1(n10544), .A2(n10543), .ZN(n10733) );
  CLKBUF_X1 U7415 ( .A(n9289), .Z(n6574) );
  XNOR2_X1 U7416 ( .A(n8908), .B(n8907), .ZN(n9289) );
  NOR2_X4 U7417 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7660) );
  NOR2_X2 U7418 ( .A1(n10546), .A2(n7301), .ZN(n10226) );
  AND2_X2 U7419 ( .A1(n7302), .A2(n10233), .ZN(n10546) );
  NAND2_X1 U7421 ( .A1(n7470), .A2(n7469), .ZN(n6575) );
  NAND2_X1 U7422 ( .A1(n7470), .A2(n7469), .ZN(n6576) );
  AOI21_X2 U7423 ( .B1(n12757), .B2(n12755), .A(n12756), .ZN(n12759) );
  NAND2_X2 U7424 ( .A1(n10226), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n12757) );
  NOR3_X2 U7425 ( .A1(n10892), .A2(n10891), .A3(n10890), .ZN(n10998) );
  OAI21_X1 U7426 ( .B1(n14119), .B2(n7342), .A(n7341), .ZN(n7340) );
  NAND2_X1 U7427 ( .A1(n14159), .A2(n6781), .ZN(n14131) );
  NAND2_X1 U7428 ( .A1(n13630), .A2(n13482), .ZN(n13614) );
  NOR2_X1 U7429 ( .A1(n14324), .A2(n14323), .ZN(n14327) );
  NAND2_X1 U7430 ( .A1(n13662), .A2(n13479), .ZN(n13647) );
  NAND2_X1 U7431 ( .A1(n12587), .A2(n8018), .ZN(n12683) );
  NAND2_X1 U7432 ( .A1(n14345), .A2(n14140), .ZN(n7341) );
  INV_X2 U7433 ( .A(n12470), .ZN(n12474) );
  OR2_X1 U7434 ( .A1(n13073), .A2(n7021), .ZN(n7018) );
  OR2_X1 U7435 ( .A1(n7314), .A2(n7313), .ZN(n7312) );
  NAND2_X1 U7436 ( .A1(n6967), .A2(n13976), .ZN(n11806) );
  AND2_X1 U7437 ( .A1(n10915), .A2(n10914), .ZN(n10956) );
  INV_X1 U7439 ( .A(n13571), .ZN(n13490) );
  AND2_X1 U7440 ( .A1(n7654), .A2(n7652), .ZN(n9637) );
  INV_X1 U7441 ( .A(n12600), .ZN(n10916) );
  INV_X2 U7442 ( .A(n14748), .ZN(n10149) );
  INV_X2 U7443 ( .A(n14860), .ZN(n10082) );
  INV_X1 U7444 ( .A(n14852), .ZN(n9708) );
  NAND2_X1 U7445 ( .A1(n9633), .A2(n15168), .ZN(n11949) );
  OAI211_X1 U7446 ( .C1(n11567), .C2(n9657), .A(n9656), .B(n9655), .ZN(n14860)
         );
  NOR2_X1 U7447 ( .A1(n12754), .A2(n10496), .ZN(n9632) );
  INV_X2 U7448 ( .A(n12225), .ZN(n12180) );
  INV_X1 U7449 ( .A(n9826), .ZN(n15075) );
  NAND2_X1 U7450 ( .A1(n8520), .A2(n8303), .ZN(n8539) );
  CLKBUF_X2 U7451 ( .A(n11390), .Z(n11491) );
  INV_X4 U7452 ( .A(n11692), .ZN(n11789) );
  XNOR2_X1 U7453 ( .A(n7648), .B(n7647), .ZN(n12882) );
  INV_X2 U7454 ( .A(n11381), .ZN(n11565) );
  INV_X2 U7455 ( .A(n11745), .ZN(n11788) );
  CLKBUF_X2 U7456 ( .A(n9324), .Z(n11390) );
  BUF_X2 U7457 ( .A(n9311), .Z(n11567) );
  BUF_X2 U7458 ( .A(n7690), .Z(n6590) );
  NAND2_X1 U7459 ( .A1(n6580), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8428) );
  INV_X1 U7460 ( .A(n15035), .ZN(n9128) );
  NAND2_X2 U7461 ( .A1(n9552), .A2(n6927), .ZN(n7843) );
  NAND2_X1 U7462 ( .A1(n8879), .A2(n12436), .ZN(n12351) );
  NAND2_X2 U7463 ( .A1(n8978), .A2(n8977), .ZN(n11413) );
  NOR2_X1 U7464 ( .A1(n7644), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7922) );
  CLKBUF_X2 U7465 ( .A(n7870), .Z(n6817) );
  INV_X2 U7466 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7467 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7299) );
  AOI21_X1 U7468 ( .B1(n12537), .B2(n11911), .A(n6675), .ZN(n12099) );
  OAI21_X1 U7469 ( .B1(n14326), .B2(n14908), .A(n7219), .ZN(n7214) );
  AND2_X1 U7470 ( .A1(n14327), .A2(n14326), .ZN(n6779) );
  AND2_X1 U7471 ( .A1(n7571), .A2(n12121), .ZN(n14342) );
  OR2_X1 U7472 ( .A1(n14339), .A2(n14556), .ZN(n7571) );
  OAI22_X1 U7473 ( .A1(n13170), .A2(n13212), .B1(n15225), .B2(n6823), .ZN(
        n6822) );
  NAND2_X1 U7474 ( .A1(n13541), .A2(n7390), .ZN(n13542) );
  AOI21_X1 U7475 ( .B1(n6833), .B2(n13683), .A(n6830), .ZN(n13724) );
  OAI21_X1 U7476 ( .B1(n13560), .B2(n7382), .A(n7381), .ZN(n13521) );
  NAND2_X1 U7477 ( .A1(n7203), .A2(n7201), .ZN(n14159) );
  NAND2_X1 U7478 ( .A1(n8063), .A2(n8062), .ZN(n8072) );
  OR2_X1 U7479 ( .A1(n8835), .A2(n6628), .ZN(n8836) );
  NAND2_X1 U7480 ( .A1(n12482), .A2(n12481), .ZN(n12984) );
  AND2_X1 U7481 ( .A1(n12480), .A2(n12479), .ZN(n12482) );
  NAND2_X1 U7482 ( .A1(n13597), .A2(n6655), .ZN(n13575) );
  NOR2_X1 U7483 ( .A1(n7385), .A2(n13526), .ZN(n7384) );
  AOI21_X1 U7484 ( .B1(n7474), .B2(n7477), .A(n6667), .ZN(n7471) );
  AOI21_X1 U7485 ( .B1(n13647), .B2(n13481), .A(n6672), .ZN(n13631) );
  NAND2_X1 U7486 ( .A1(n7563), .A2(n12287), .ZN(n12364) );
  NAND2_X1 U7487 ( .A1(n11833), .A2(n11832), .ZN(n14383) );
  AND2_X1 U7488 ( .A1(n13135), .A2(n12035), .ZN(n13033) );
  AND2_X1 U7489 ( .A1(n14125), .A2(n12118), .ZN(n7342) );
  NAND2_X1 U7490 ( .A1(n7284), .A2(n6630), .ZN(n13681) );
  NAND2_X1 U7491 ( .A1(n7296), .A2(n6738), .ZN(n12826) );
  NAND2_X1 U7492 ( .A1(n12282), .A2(n12281), .ZN(n13722) );
  NAND2_X1 U7493 ( .A1(n14296), .A2(n11804), .ZN(n14277) );
  NAND2_X1 U7494 ( .A1(n11483), .A2(n11482), .ZN(n14125) );
  NAND2_X1 U7495 ( .A1(n11503), .A2(n11502), .ZN(n14337) );
  NAND2_X1 U7496 ( .A1(n12318), .A2(n12317), .ZN(n13717) );
  AND2_X1 U7497 ( .A1(n13482), .A2(n12398), .ZN(n13636) );
  NAND2_X1 U7498 ( .A1(n11630), .A2(n11629), .ZN(n13727) );
  NOR2_X1 U7499 ( .A1(n13732), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U7500 ( .A1(n8369), .A2(n8368), .ZN(n13732) );
  INV_X1 U7501 ( .A(n13624), .ZN(n7056) );
  AND2_X1 U7502 ( .A1(n8827), .A2(n8826), .ZN(n13741) );
  INV_X1 U7503 ( .A(n7416), .ZN(n10860) );
  INV_X1 U7504 ( .A(n13655), .ZN(n13747) );
  XOR2_X1 U7505 ( .A(n12814), .B(n12806), .Z(n12784) );
  AND2_X1 U7506 ( .A1(n11700), .A2(n11688), .ZN(n7502) );
  NAND2_X1 U7507 ( .A1(n11413), .A2(n14437), .ZN(n14198) );
  NAND2_X1 U7508 ( .A1(n12783), .A2(n12782), .ZN(n12806) );
  AND2_X1 U7509 ( .A1(n8808), .A2(n8807), .ZN(n13655) );
  OAI21_X1 U7510 ( .B1(n10794), .B2(n7418), .A(n7417), .ZN(n7416) );
  INV_X1 U7511 ( .A(n7073), .ZN(n7072) );
  NAND2_X1 U7512 ( .A1(n11411), .A2(n8820), .ZN(n8824) );
  OAI21_X1 U7513 ( .B1(n10245), .B2(n10246), .A(n8631), .ZN(n10387) );
  NOR2_X1 U7514 ( .A1(n12841), .A2(n12842), .ZN(n12863) );
  NAND2_X1 U7515 ( .A1(n7312), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U7516 ( .A1(n10369), .A2(n10368), .ZN(n10374) );
  OAI21_X1 U7517 ( .B1(n10888), .B2(n14623), .A(n10884), .ZN(n10984) );
  AND2_X1 U7518 ( .A1(n8801), .A2(n8351), .ZN(n8352) );
  NAND2_X1 U7519 ( .A1(n8780), .A2(n8779), .ZN(n13757) );
  AND2_X1 U7520 ( .A1(n8419), .A2(n8418), .ZN(n13478) );
  NAND2_X1 U7521 ( .A1(n11304), .A2(n11303), .ZN(n11350) );
  NAND2_X2 U7522 ( .A1(n11283), .A2(n11282), .ZN(n11297) );
  AOI21_X1 U7523 ( .B1(n10504), .B2(n15332), .A(n10497), .ZN(n10498) );
  NAND2_X1 U7524 ( .A1(n7128), .A2(n14520), .ZN(n14552) );
  NAND2_X1 U7525 ( .A1(n12627), .A2(n12628), .ZN(n12626) );
  XNOR2_X1 U7526 ( .A(n8715), .B(n8714), .ZN(n11285) );
  AND2_X1 U7527 ( .A1(n8679), .A2(n8678), .ZN(n14634) );
  NAND2_X1 U7528 ( .A1(n11314), .A2(n11313), .ZN(n14397) );
  AOI21_X1 U7529 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8715) );
  OR2_X1 U7530 ( .A1(n10467), .A2(n11258), .ZN(n10458) );
  NAND2_X1 U7531 ( .A1(n10571), .A2(n10570), .ZN(n13877) );
  XNOR2_X1 U7532 ( .A(n8672), .B(n8671), .ZN(n10573) );
  NAND2_X1 U7533 ( .A1(n8635), .A2(n8634), .ZN(n10776) );
  NAND2_X1 U7534 ( .A1(n10411), .A2(n10410), .ZN(n11258) );
  OR2_X1 U7535 ( .A1(n10224), .A2(n6728), .ZN(n7302) );
  NAND2_X1 U7536 ( .A1(n8622), .A2(n8621), .ZN(n15119) );
  AOI21_X1 U7537 ( .B1(n10049), .B2(n10031), .A(n10032), .ZN(n10224) );
  NAND2_X1 U7538 ( .A1(n10050), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U7539 ( .A1(n7066), .A2(n8324), .ZN(n8652) );
  AOI21_X1 U7540 ( .B1(n14673), .B2(n9409), .A(n9404), .ZN(n9406) );
  INV_X2 U7541 ( .A(n15198), .ZN(n14582) );
  NOR2_X1 U7542 ( .A1(n10030), .A2(n6988), .ZN(n10050) );
  NOR2_X1 U7543 ( .A1(n14596), .A2(n15183), .ZN(n14583) );
  AOI21_X1 U7544 ( .B1(n6947), .B2(n6948), .A(n6647), .ZN(n6946) );
  OR2_X1 U7545 ( .A1(n7888), .A2(n10574), .ZN(n6807) );
  NOR2_X1 U7546 ( .A1(n6989), .A2(n10052), .ZN(n6988) );
  AND2_X1 U7547 ( .A1(n6989), .A2(n10052), .ZN(n10030) );
  NAND3_X1 U7548 ( .A1(n8320), .A2(n8321), .A3(SI_10_), .ZN(n8619) );
  NAND2_X1 U7549 ( .A1(n9687), .A2(n7339), .ZN(n14779) );
  OR2_X1 U7550 ( .A1(n10027), .A2(n6633), .ZN(n6989) );
  NAND2_X1 U7551 ( .A1(n8317), .A2(n8316), .ZN(n8320) );
  NAND2_X1 U7552 ( .A1(n8319), .A2(n8318), .ZN(n8321) );
  INV_X2 U7553 ( .A(n15045), .ZN(n6578) );
  AOI21_X1 U7554 ( .B1(n9998), .B2(n9996), .A(n9997), .ZN(n10027) );
  AND2_X1 U7555 ( .A1(n11956), .A2(n11957), .ZN(n11945) );
  NAND2_X1 U7556 ( .A1(n8596), .A2(n8315), .ZN(n8319) );
  XNOR2_X2 U7557 ( .A(n10082), .B(n13984), .ZN(n11590) );
  NAND2_X1 U7558 ( .A1(n7098), .A2(n7682), .ZN(n12751) );
  NAND2_X1 U7559 ( .A1(n15192), .A2(n10199), .ZN(n11955) );
  OAI22_X1 U7560 ( .A1(n9607), .A2(n9608), .B1(n9584), .B2(n9598), .ZN(n9588)
         );
  NAND4_X1 U7561 ( .A1(n9368), .A2(n9367), .A3(n9366), .A4(n9365), .ZN(n13984)
         );
  AND2_X1 U7562 ( .A1(n7304), .A2(n9585), .ZN(n9995) );
  AND4_X1 U7563 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n10644)
         );
  NOR2_X1 U7564 ( .A1(n6623), .A2(n7094), .ZN(n7098) );
  AND2_X2 U7565 ( .A1(n7192), .A2(n9333), .ZN(n14852) );
  BUF_X1 U7566 ( .A(n9634), .Z(n15168) );
  INV_X1 U7567 ( .A(n15062), .ZN(n9906) );
  NOR2_X1 U7568 ( .A1(n9904), .A2(n15062), .ZN(n9903) );
  AND2_X1 U7569 ( .A1(n6653), .A2(n8493), .ZN(n9528) );
  INV_X4 U7570 ( .A(n12180), .ZN(n12331) );
  OR2_X1 U7571 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  NAND2_X1 U7572 ( .A1(n6994), .A2(n6993), .ZN(n7306) );
  AND3_X1 U7573 ( .A1(n7679), .A2(n7678), .A3(n7677), .ZN(n12581) );
  OAI211_X1 U7574 ( .C1(n11413), .C2(n6574), .A(n9288), .B(n9287), .ZN(n14834)
         );
  AND3_X1 U7575 ( .A1(n7665), .A2(n7664), .A3(n7666), .ZN(n10199) );
  CLKBUF_X1 U7576 ( .A(n11181), .Z(n11538) );
  INV_X2 U7577 ( .A(n11567), .ZN(n11519) );
  OR2_X1 U7578 ( .A1(n11381), .A2(n9330), .ZN(n9333) );
  NOR2_X1 U7579 ( .A1(n9008), .A2(P2_U3088), .ZN(P2_U3947) );
  CLKBUF_X1 U7580 ( .A(n8463), .Z(n6581) );
  CLKBUF_X1 U7581 ( .A(n8451), .Z(n12357) );
  NAND2_X1 U7582 ( .A1(n12353), .A2(n8879), .ZN(n12140) );
  AND2_X1 U7583 ( .A1(n9238), .A2(n11162), .ZN(n11181) );
  OR2_X1 U7584 ( .A1(n8490), .A2(n9045), .ZN(n8441) );
  BUF_X1 U7585 ( .A(n9235), .Z(n12132) );
  INV_X1 U7586 ( .A(n7758), .ZN(n6579) );
  INV_X1 U7587 ( .A(n11574), .ZN(n11195) );
  INV_X1 U7588 ( .A(n8881), .ZN(n12353) );
  INV_X1 U7589 ( .A(n12348), .ZN(n8778) );
  NAND2_X1 U7590 ( .A1(n7574), .A2(n6928), .ZN(n6929) );
  AND2_X1 U7591 ( .A1(n7294), .A2(n9613), .ZN(n9571) );
  OR2_X1 U7592 ( .A1(n12348), .A2(n8917), .ZN(n8464) );
  INV_X2 U7593 ( .A(n8466), .ZN(n8484) );
  NAND2_X1 U7594 ( .A1(n8378), .A2(n8377), .ZN(n8881) );
  BUF_X2 U7595 ( .A(n11576), .Z(n6790) );
  INV_X2 U7596 ( .A(n12884), .ZN(n12862) );
  INV_X1 U7597 ( .A(n7536), .ZN(n7535) );
  INV_X1 U7598 ( .A(n8490), .ZN(n6580) );
  XNOR2_X1 U7599 ( .A(n9232), .B(n9231), .ZN(n9235) );
  XNOR2_X1 U7600 ( .A(n8967), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U7601 ( .A1(n14421), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U7602 ( .A1(n8381), .A2(n8374), .ZN(n8378) );
  CLKBUF_X1 U7603 ( .A(n8978), .Z(n12134) );
  XNOR2_X1 U7604 ( .A(n8390), .B(P2_IR_REG_19__SCAN_IN), .ZN(n12436) );
  MUX2_X1 U7605 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8380), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8382) );
  NOR2_X1 U7606 ( .A1(n7849), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U7607 ( .A1(n8387), .A2(n8386), .ZN(n12352) );
  XNOR2_X1 U7608 ( .A(n8243), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9339) );
  OR2_X1 U7609 ( .A1(n7115), .A2(n7662), .ZN(n7596) );
  NAND2_X1 U7610 ( .A1(n8242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8243) );
  AND2_X1 U7611 ( .A1(n8249), .A2(n6696), .ZN(n9233) );
  NOR2_X1 U7612 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U7613 ( .A1(n8394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8367) );
  NOR2_X1 U7614 ( .A1(n8394), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7615 ( .A1(n8240), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n8242) );
  NOR2_X1 U7616 ( .A1(n8416), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n8388) );
  NAND2_X2 U7617 ( .A1(n7300), .A2(n7297), .ZN(n9981) );
  NOR2_X1 U7618 ( .A1(n7528), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7527) );
  AND2_X1 U7619 ( .A1(n8234), .A2(n8232), .ZN(n7060) );
  INV_X1 U7620 ( .A(n7573), .ZN(n7039) );
  NAND2_X1 U7621 ( .A1(n8233), .A2(n8921), .ZN(n7235) );
  AND2_X1 U7622 ( .A1(n7645), .A2(n7646), .ZN(n7121) );
  NAND2_X1 U7623 ( .A1(n8248), .A2(n7529), .ZN(n7528) );
  AND3_X1 U7624 ( .A1(n8238), .A2(n8237), .A3(n8236), .ZN(n8245) );
  AND4_X1 U7625 ( .A1(n8257), .A2(n8256), .A3(n8480), .A4(n8525), .ZN(n8258)
         );
  NAND3_X1 U7626 ( .A1(n7257), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U7627 ( .A1(n7130), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7655) );
  AND2_X1 U7628 ( .A1(n6900), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14492) );
  AND4_X1 U7629 ( .A1(n7589), .A2(n7588), .A3(n7779), .A4(n7740), .ZN(n7590)
         );
  AND2_X1 U7630 ( .A1(n7523), .A2(n7591), .ZN(n7522) );
  INV_X1 U7631 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7529) );
  INV_X1 U7632 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8370) );
  INV_X1 U7633 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8929) );
  INV_X1 U7634 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8371) );
  INV_X1 U7635 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8384) );
  INV_X1 U7636 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9231) );
  INV_X4 U7637 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7638 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8268) );
  NOR2_X1 U7639 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8375) );
  INV_X1 U7640 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U7641 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8902) );
  NOR2_X1 U7642 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7003) );
  INV_X1 U7643 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8597) );
  INV_X1 U7644 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7779) );
  INV_X1 U7645 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8480) );
  INV_X1 U7646 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U7647 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14491) );
  INV_X1 U7648 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8653) );
  NOR2_X1 U7649 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7588) );
  NOR2_X1 U7650 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7589) );
  NOR2_X1 U7651 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8227) );
  NOR2_X1 U7652 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8228) );
  NOR2_X1 U7653 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8226) );
  INV_X1 U7654 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8525) );
  INV_X1 U7655 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8234) );
  NOR2_X1 U7656 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8257) );
  NOR2_X1 U7657 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7593) );
  NOR2_X1 U7658 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7592) );
  NOR2_X1 U7659 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8259) );
  NOR2_X1 U7660 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n8260) );
  INV_X1 U7661 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7645) );
  INV_X1 U7662 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7646) );
  OR2_X1 U7663 ( .A1(n10116), .A2(n11381), .ZN(n10118) );
  OAI21_X1 U7664 ( .B1(n8553), .B2(n8554), .A(n8555), .ZN(n10116) );
  OR2_X1 U7665 ( .A1(n8416), .A2(n8271), .ZN(n8383) );
  OR2_X1 U7666 ( .A1(n8451), .A2(n8427), .ZN(n8430) );
  OAI21_X1 U7667 ( .B1(n7959), .B2(n7962), .A(n7960), .ZN(n6769) );
  NAND2_X2 U7668 ( .A1(n13278), .A2(n8836), .ZN(n8852) );
  NOR2_X4 U7669 ( .A1(n11861), .A2(n11860), .ZN(n14335) );
  OAI21_X2 U7670 ( .B1(n13971), .B2(n14337), .A(n12112), .ZN(n11861) );
  OAI21_X2 U7671 ( .B1(n7363), .B2(n7361), .A(n7358), .ZN(n14235) );
  NAND2_X2 U7672 ( .A1(n12114), .A2(n12113), .ZN(n12112) );
  NOR2_X2 U7673 ( .A1(n13921), .A2(n13920), .ZN(n13919) );
  AOI21_X2 U7674 ( .B1(n7504), .B2(n7507), .A(n7503), .ZN(n13921) );
  INV_X4 U7675 ( .A(n11431), .ZN(n11351) );
  INV_X1 U7676 ( .A(n8825), .ZN(n8463) );
  XNOR2_X2 U7677 ( .A(n10149), .B(n14875), .ZN(n11591) );
  NOR2_X4 U7678 ( .A1(n6817), .A2(n7040), .ZN(n7621) );
  NAND2_X2 U7679 ( .A1(n8399), .A2(n8400), .ZN(n6583) );
  NAND2_X2 U7680 ( .A1(n8399), .A2(n8400), .ZN(n8438) );
  NOR2_X2 U7681 ( .A1(n12902), .A2(n12080), .ZN(n12491) );
  NOR2_X2 U7682 ( .A1(n13252), .A2(n7572), .ZN(n8834) );
  NAND2_X1 U7683 ( .A1(n9503), .A2(n10201), .ZN(n11950) );
  NOR2_X2 U7684 ( .A1(n7017), .A2(n7016), .ZN(n10201) );
  AND2_X1 U7685 ( .A1(n12524), .A2(n13225), .ZN(n6584) );
  OAI21_X1 U7686 ( .B1(n9842), .B2(n12100), .A(n7649), .ZN(n6585) );
  XNOR2_X2 U7687 ( .A(n12147), .B(n6929), .ZN(n9525) );
  XNOR2_X2 U7688 ( .A(n8904), .B(n8903), .ZN(n13998) );
  OR2_X4 U7689 ( .A1(n15033), .A2(n8407), .ZN(n8705) );
  BUF_X8 U7690 ( .A(n7761), .Z(n6587) );
  NAND2_X1 U7691 ( .A1(n9010), .A2(n9012), .ZN(n6588) );
  AND2_X2 U7692 ( .A1(n13672), .A2(n13655), .ZN(n13650) );
  NOR2_X2 U7693 ( .A1(n13752), .A2(n13693), .ZN(n13672) );
  AOI21_X2 U7694 ( .B1(n6812), .B2(n6606), .A(n6658), .ZN(n13476) );
  NOR2_X4 U7695 ( .A1(n14308), .A2(n11297), .ZN(n14282) );
  NAND2_X1 U7696 ( .A1(n8400), .A2(n11172), .ZN(n8490) );
  XNOR2_X2 U7697 ( .A(n8396), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8399) );
  NOR2_X2 U7698 ( .A1(n13548), .A2(n13712), .ZN(n7042) );
  AOI211_X1 U7699 ( .C1(n15103), .C2(n14943), .A(n9949), .B(n9948), .ZN(n9950)
         );
  CLKBUF_X3 U7700 ( .A(n9666), .Z(n11540) );
  NOR2_X1 U7701 ( .A1(n7538), .A2(n7082), .ZN(n7081) );
  NAND2_X1 U7702 ( .A1(n8332), .A2(n6591), .ZN(n7538) );
  NOR2_X1 U7703 ( .A1(n11874), .A2(n7092), .ZN(n7091) );
  INV_X1 U7704 ( .A(n11873), .ZN(n7092) );
  NAND2_X1 U7705 ( .A1(n13624), .A2(n13596), .ZN(n7431) );
  INV_X1 U7706 ( .A(n7290), .ZN(n11012) );
  INV_X1 U7707 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8269) );
  NOR3_X1 U7708 ( .A1(n12089), .A2(n11933), .A3(n12091), .ZN(n12101) );
  NAND2_X1 U7709 ( .A1(n6697), .A2(n12178), .ZN(n7336) );
  NAND2_X1 U7710 ( .A1(n6966), .A2(n6965), .ZN(n11300) );
  NAND2_X1 U7711 ( .A1(n11585), .A2(n11351), .ZN(n6965) );
  OAI21_X1 U7712 ( .B1(n7319), .B2(n7317), .A(n7315), .ZN(n12257) );
  NAND2_X1 U7713 ( .A1(n12252), .A2(n7316), .ZN(n7315) );
  AND2_X1 U7714 ( .A1(n12253), .A2(n7318), .ZN(n7317) );
  AND2_X1 U7715 ( .A1(n12248), .A2(n12247), .ZN(n7319) );
  NAND2_X1 U7716 ( .A1(n7331), .A2(n7332), .ZN(n7329) );
  MUX2_X1 U7717 ( .A(n14167), .B(n14359), .S(n11504), .Z(n11449) );
  NAND2_X1 U7718 ( .A1(n7320), .A2(n7321), .ZN(n12272) );
  NAND2_X1 U7719 ( .A1(n12271), .A2(n7322), .ZN(n7321) );
  NOR2_X1 U7720 ( .A1(n6665), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U7721 ( .A1(n12212), .A2(n13314), .ZN(n7264) );
  INV_X1 U7722 ( .A(n6968), .ZN(n6897) );
  AND2_X1 U7723 ( .A1(n8321), .A2(n7068), .ZN(n7067) );
  INV_X1 U7724 ( .A(n12984), .ZN(n7034) );
  INV_X1 U7725 ( .A(n7035), .ZN(n7031) );
  INV_X1 U7726 ( .A(n8059), .ZN(n7148) );
  INV_X1 U7727 ( .A(n7463), .ZN(n6941) );
  NOR2_X1 U7728 ( .A1(n12140), .A2(n12460), .ZN(n12388) );
  NOR2_X1 U7729 ( .A1(n12379), .A2(n7555), .ZN(n12342) );
  AND2_X1 U7730 ( .A1(n12343), .A2(n12344), .ZN(n7555) );
  AND2_X1 U7731 ( .A1(n7054), .A2(n7055), .ZN(n7053) );
  INV_X1 U7732 ( .A(n13636), .ZN(n7429) );
  NOR2_X1 U7733 ( .A1(n7412), .A2(n6617), .ZN(n7411) );
  NAND2_X1 U7734 ( .A1(n12235), .A2(n13311), .ZN(n7406) );
  OAI21_X1 U7735 ( .B1(n9760), .B2(n9533), .A(n9534), .ZN(n9743) );
  NAND2_X1 U7736 ( .A1(n9528), .A2(n15070), .ZN(n9815) );
  NOR2_X1 U7737 ( .A1(n8383), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8281) );
  OAI21_X1 U7738 ( .B1(n6888), .B2(n11842), .A(n7567), .ZN(n6886) );
  OR2_X1 U7739 ( .A1(n14353), .A2(n13972), .ZN(n7567) );
  AND2_X1 U7740 ( .A1(n14257), .A2(n6600), .ZN(n6878) );
  OR2_X1 U7741 ( .A1(n11290), .A2(n15522), .ZN(n11324) );
  NAND2_X1 U7742 ( .A1(n14402), .A2(n11299), .ZN(n11805) );
  NAND2_X1 U7743 ( .A1(n9708), .A2(n7338), .ZN(n11213) );
  AND2_X1 U7744 ( .A1(n11213), .A2(n11214), .ZN(n11588) );
  NOR2_X1 U7745 ( .A1(n8246), .A2(n7375), .ZN(n7374) );
  NAND2_X1 U7746 ( .A1(n7526), .A2(n8234), .ZN(n7375) );
  INV_X1 U7747 ( .A(n7528), .ZN(n7526) );
  XNOR2_X1 U7748 ( .A(n8349), .B(SI_20_), .ZN(n8788) );
  INV_X1 U7749 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U7750 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  AOI21_X1 U7751 ( .B1(n7078), .B2(n7080), .A(n7077), .ZN(n7076) );
  NOR2_X2 U7752 ( .A1(n7235), .A2(n7233), .ZN(n9896) );
  AND2_X1 U7753 ( .A1(n7234), .A2(n8234), .ZN(n7231) );
  INV_X1 U7754 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7234) );
  AND2_X1 U7755 ( .A1(n7535), .A2(n6876), .ZN(n6875) );
  NAND2_X1 U7756 ( .A1(n8305), .A2(n8306), .ZN(n6876) );
  AND4_X1 U7757 ( .A1(n7606), .A2(n7605), .A3(n7604), .A4(n7603), .ZN(n9634)
         );
  NAND2_X1 U7758 ( .A1(n12495), .A2(n6748), .ZN(n6747) );
  INV_X1 U7759 ( .A(n12909), .ZN(n6748) );
  NAND2_X1 U7760 ( .A1(n12077), .A2(n11878), .ZN(n12492) );
  NAND2_X1 U7761 ( .A1(n12485), .A2(n12492), .ZN(n12525) );
  AOI21_X1 U7762 ( .B1(n7091), .B2(n12942), .A(n7089), .ZN(n7088) );
  INV_X1 U7763 ( .A(n12070), .ZN(n7089) );
  INV_X1 U7764 ( .A(n7091), .ZN(n7090) );
  AND2_X1 U7765 ( .A1(n11876), .A2(n11875), .ZN(n12907) );
  AOI21_X1 U7766 ( .B1(n7110), .B2(n7108), .A(n7107), .ZN(n7106) );
  INV_X1 U7767 ( .A(n7113), .ZN(n7108) );
  NAND2_X1 U7768 ( .A1(n10206), .A2(n12102), .ZN(n15149) );
  NAND2_X1 U7769 ( .A1(n9552), .A2(n11550), .ZN(n7690) );
  NAND2_X1 U7770 ( .A1(n10348), .A2(n10347), .ZN(n10354) );
  INV_X1 U7771 ( .A(n7843), .ZN(n11897) );
  NAND2_X1 U7772 ( .A1(n8038), .A2(n8037), .ZN(n8040) );
  AOI21_X1 U7773 ( .B1(n13231), .B2(n7442), .A(n7441), .ZN(n7440) );
  NOR2_X1 U7774 ( .A1(n12515), .A2(n12511), .ZN(n7441) );
  XNOR2_X1 U7775 ( .A(n9906), .B(n8426), .ZN(n8470) );
  AND2_X1 U7776 ( .A1(n12387), .A2(n12386), .ZN(n12446) );
  INV_X1 U7777 ( .A(n8451), .ZN(n12319) );
  NAND2_X1 U7778 ( .A1(n12350), .A2(n12349), .ZN(n13469) );
  NAND2_X1 U7779 ( .A1(n13717), .A2(n13571), .ZN(n7393) );
  NAND2_X1 U7780 ( .A1(n6746), .A2(n6651), .ZN(n7380) );
  INV_X1 U7781 ( .A(n13575), .ZN(n6746) );
  NAND2_X1 U7782 ( .A1(n13613), .A2(n7428), .ZN(n7427) );
  INV_X1 U7783 ( .A(n7432), .ZN(n7428) );
  NAND2_X1 U7784 ( .A1(n7288), .A2(n7400), .ZN(n7290) );
  AND2_X1 U7785 ( .A1(n14944), .A2(n10795), .ZN(n6756) );
  NAND2_X1 U7786 ( .A1(n6787), .A2(n15062), .ZN(n9779) );
  AND2_X1 U7787 ( .A1(n8361), .A2(n8363), .ZN(n8364) );
  AND2_X1 U7788 ( .A1(n11738), .A2(n11739), .ZN(n6818) );
  NAND2_X1 U7789 ( .A1(n11177), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11435) );
  INV_X1 U7790 ( .A(n11390), .ZN(n11510) );
  NAND2_X1 U7791 ( .A1(n12132), .A2(n9236), .ZN(n9666) );
  INV_X1 U7792 ( .A(n14140), .ZN(n12118) );
  NAND2_X1 U7793 ( .A1(n14134), .A2(n6889), .ZN(n6888) );
  INV_X1 U7794 ( .A(n6890), .ZN(n6889) );
  NOR2_X1 U7795 ( .A1(n11842), .A2(n11859), .ZN(n7201) );
  AOI21_X1 U7796 ( .B1(n7367), .B2(n11841), .A(n6686), .ZN(n7365) );
  BUF_X1 U7797 ( .A(n9329), .Z(n11381) );
  NOR2_X2 U7798 ( .A1(n10108), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9293) );
  INV_X1 U7799 ( .A(n11550), .ZN(n6927) );
  AOI21_X1 U7800 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14466), .A(n14465), .ZN(
        n14479) );
  NOR2_X1 U7801 ( .A1(n14524), .A2(n14523), .ZN(n14465) );
  OR2_X1 U7802 ( .A1(n14534), .A2(n6641), .ZN(n6911) );
  OR2_X1 U7803 ( .A1(n14535), .A2(n6913), .ZN(n6912) );
  NAND2_X1 U7804 ( .A1(n14099), .A2(n14096), .ZN(n7347) );
  OAI21_X1 U7805 ( .B1(n14099), .B2(n6678), .A(n7346), .ZN(n7345) );
  NAND2_X1 U7806 ( .A1(n11206), .A2(n11207), .ZN(n7230) );
  INV_X1 U7807 ( .A(n11228), .ZN(n7224) );
  INV_X1 U7808 ( .A(n11230), .ZN(n6795) );
  OR2_X1 U7809 ( .A1(n11230), .A2(n7224), .ZN(n7223) );
  NAND2_X1 U7810 ( .A1(n12147), .A2(n12225), .ZN(n7394) );
  OR2_X1 U7811 ( .A1(n7256), .A2(n11240), .ZN(n6793) );
  INV_X1 U7812 ( .A(n11239), .ZN(n7256) );
  OR2_X1 U7813 ( .A1(n12190), .A2(n12191), .ZN(n6852) );
  OR2_X1 U7814 ( .A1(n12178), .A2(n6697), .ZN(n7335) );
  NOR2_X1 U7815 ( .A1(n7309), .A2(n12194), .ZN(n6853) );
  AND2_X1 U7816 ( .A1(n11300), .A2(n7238), .ZN(n6740) );
  NAND2_X1 U7817 ( .A1(n11300), .A2(n6671), .ZN(n7236) );
  NAND2_X1 U7818 ( .A1(n11368), .A2(n11367), .ZN(n11401) );
  NAND2_X1 U7819 ( .A1(n12224), .A2(n12223), .ZN(n6867) );
  NAND2_X1 U7820 ( .A1(n6864), .A2(n12226), .ZN(n6863) );
  INV_X1 U7821 ( .A(n6867), .ZN(n6864) );
  NOR2_X1 U7822 ( .A1(n6865), .A2(n6861), .ZN(n6860) );
  NOR2_X1 U7823 ( .A1(n6868), .A2(n6866), .ZN(n6865) );
  INV_X1 U7824 ( .A(n6863), .ZN(n6861) );
  AOI21_X1 U7825 ( .B1(n7246), .B2(n7244), .A(n7242), .ZN(n7241) );
  INV_X1 U7826 ( .A(n11449), .ZN(n7242) );
  OAI21_X1 U7827 ( .B1(n12257), .B2(n12256), .A(n12255), .ZN(n6849) );
  NAND2_X1 U7828 ( .A1(n12262), .A2(n12261), .ZN(n7328) );
  NAND2_X1 U7829 ( .A1(n7330), .A2(n7329), .ZN(n7327) );
  NOR2_X1 U7830 ( .A1(n7331), .A2(n7332), .ZN(n7330) );
  INV_X1 U7831 ( .A(n7329), .ZN(n7326) );
  MUX2_X1 U7832 ( .A(n14102), .B(n14330), .S(n11504), .Z(n11524) );
  INV_X1 U7833 ( .A(n6982), .ZN(n6981) );
  NOR2_X1 U7834 ( .A1(n7253), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U7835 ( .A1(n6753), .A2(n6752), .ZN(n12475) );
  INV_X1 U7836 ( .A(n13193), .ZN(n6753) );
  INV_X1 U7837 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7623) );
  INV_X1 U7838 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7591) );
  INV_X1 U7839 ( .A(n9674), .ZN(n7191) );
  NAND2_X1 U7840 ( .A1(n6734), .A2(n6614), .ZN(n7551) );
  NAND2_X1 U7841 ( .A1(n7072), .A2(n8837), .ZN(n7070) );
  NAND2_X1 U7842 ( .A1(n8824), .A2(n7072), .ZN(n7071) );
  AND2_X1 U7843 ( .A1(n7547), .A2(n11152), .ZN(n7546) );
  INV_X1 U7844 ( .A(n7551), .ZN(n7547) );
  NOR2_X1 U7845 ( .A1(n11461), .A2(n7553), .ZN(n7552) );
  INV_X1 U7846 ( .A(n11154), .ZN(n7553) );
  INV_X1 U7847 ( .A(n7559), .ZN(n7558) );
  OAI21_X1 U7848 ( .B1(n7561), .B2(n7562), .A(n7560), .ZN(n7559) );
  INV_X1 U7849 ( .A(n8777), .ZN(n7560) );
  NOR2_X1 U7850 ( .A1(n7082), .A2(n6899), .ZN(n6898) );
  INV_X1 U7851 ( .A(n8651), .ZN(n6899) );
  NAND2_X1 U7852 ( .A1(n14444), .A2(n14445), .ZN(n14446) );
  INV_X1 U7853 ( .A(n8072), .ZN(n6782) );
  AND2_X1 U7854 ( .A1(n10557), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6767) );
  OAI22_X1 U7855 ( .A1(n12832), .A2(n12831), .B1(n12830), .B2(n12829), .ZN(
        n12855) );
  OR2_X1 U7856 ( .A1(n12931), .A2(n12910), .ZN(n12070) );
  NAND2_X1 U7857 ( .A1(n7037), .A2(n7036), .ZN(n7035) );
  NAND2_X1 U7858 ( .A1(n7034), .A2(n7033), .ZN(n7032) );
  INV_X1 U7859 ( .A(n12047), .ZN(n7102) );
  INV_X1 U7860 ( .A(n7022), .ZN(n7021) );
  NAND2_X1 U7861 ( .A1(n7022), .A2(n7020), .ZN(n7019) );
  INV_X1 U7862 ( .A(n12465), .ZN(n7020) );
  NOR2_X1 U7863 ( .A1(n12010), .A2(n7111), .ZN(n7110) );
  NAND2_X1 U7864 ( .A1(n12751), .A2(n10216), .ZN(n11957) );
  INV_X1 U7865 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7119) );
  INV_X1 U7866 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7610) );
  NAND2_X1 U7867 ( .A1(n6773), .A2(n7160), .ZN(n6778) );
  NOR2_X1 U7868 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8091), .ZN(n7159) );
  AND2_X1 U7869 ( .A1(n7622), .A2(n7623), .ZN(n7531) );
  INV_X1 U7870 ( .A(n7520), .ZN(n7040) );
  NAND2_X1 U7871 ( .A1(n6690), .A2(n7821), .ZN(n7170) );
  NOR2_X1 U7872 ( .A1(n7170), .A2(n7166), .ZN(n7165) );
  INV_X1 U7873 ( .A(n7801), .ZN(n7166) );
  NOR2_X1 U7874 ( .A1(n9458), .A2(n6949), .ZN(n6948) );
  OR2_X1 U7875 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  OAI21_X1 U7876 ( .B1(n6661), .B2(n6842), .A(n6841), .ZN(n12278) );
  INV_X1 U7877 ( .A(n12274), .ZN(n6842) );
  OR2_X1 U7878 ( .A1(n12272), .A2(n12273), .ZN(n6841) );
  AOI21_X1 U7879 ( .B1(n7570), .B2(n13555), .A(n7273), .ZN(n7272) );
  INV_X1 U7880 ( .A(n13491), .ZN(n7273) );
  INV_X1 U7881 ( .A(n13741), .ZN(n13515) );
  NOR2_X1 U7882 ( .A1(n13757), .A2(n13668), .ZN(n13508) );
  NOR2_X1 U7883 ( .A1(n11022), .A2(n13773), .ZN(n7046) );
  AND2_X1 U7884 ( .A1(n7050), .A2(n12196), .ZN(n7049) );
  NAND2_X1 U7885 ( .A1(n9532), .A2(n9531), .ZN(n9760) );
  NOR2_X1 U7886 ( .A1(n9286), .A2(n7614), .ZN(n6926) );
  NOR2_X1 U7887 ( .A1(n7389), .A2(n7386), .ZN(n7385) );
  INV_X1 U7888 ( .A(n7391), .ZN(n7386) );
  AND2_X1 U7889 ( .A1(n12140), .A2(n12460), .ZN(n8391) );
  NAND2_X1 U7890 ( .A1(n9803), .A2(n9802), .ZN(n10066) );
  INV_X1 U7891 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8263) );
  INV_X1 U7892 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8262) );
  INV_X1 U7893 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8273) );
  INV_X1 U7894 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8256) );
  AOI21_X1 U7895 ( .B1(n7370), .B2(n11840), .A(n14166), .ZN(n7367) );
  INV_X1 U7896 ( .A(n14290), .ZN(n11824) );
  AND2_X1 U7897 ( .A1(n11597), .A2(n7180), .ZN(n7176) );
  INV_X1 U7898 ( .A(n10437), .ZN(n7180) );
  NAND2_X1 U7899 ( .A1(n10444), .A2(n10437), .ZN(n7179) );
  NOR2_X1 U7900 ( .A1(n11624), .A2(n9642), .ZN(n10315) );
  OAI21_X1 U7901 ( .B1(n11501), .B2(n11158), .A(n11157), .ZN(n11518) );
  NAND2_X1 U7902 ( .A1(n7554), .A2(n7552), .ZN(n7548) );
  INV_X1 U7903 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8248) );
  AND2_X1 U7904 ( .A1(n7083), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U7905 ( .A1(n6692), .A2(n6591), .ZN(n7083) );
  NAND2_X1 U7906 ( .A1(n7081), .A2(n6969), .ZN(n7079) );
  INV_X1 U7907 ( .A(n7081), .ZN(n7080) );
  INV_X1 U7908 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8231) );
  INV_X1 U7909 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8230) );
  OR2_X1 U7910 ( .A1(n6897), .A2(n6898), .ZN(n6896) );
  NOR2_X1 U7911 ( .A1(n6897), .A2(n6894), .ZN(n6893) );
  INV_X1 U7912 ( .A(n8324), .ZN(n6894) );
  NOR2_X1 U7913 ( .A1(n9100), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9102) );
  OAI211_X1 U7914 ( .C1(n7470), .C2(n8916), .A(n7468), .B(n7467), .ZN(n8288)
         );
  NAND2_X1 U7915 ( .A1(n6906), .A2(n6904), .ZN(n14443) );
  NAND2_X1 U7916 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6905), .ZN(n6904) );
  NAND2_X1 U7917 ( .A1(n14490), .A2(n14489), .ZN(n6906) );
  XNOR2_X1 U7918 ( .A(n14446), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14486) );
  OAI21_X1 U7919 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14464), .A(n14463), .ZN(
        n14523) );
  INV_X1 U7920 ( .A(n7885), .ZN(n7486) );
  AOI21_X1 U7921 ( .B1(n7514), .B2(n7984), .A(n6682), .ZN(n7513) );
  NAND2_X1 U7922 ( .A1(n12721), .A2(n8142), .ZN(n12552) );
  OR2_X1 U7923 ( .A1(n8065), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8086) );
  OR2_X1 U7924 ( .A1(n6813), .A2(n7984), .ZN(n7517) );
  OR2_X1 U7925 ( .A1(n7993), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8011) );
  NOR2_X1 U7926 ( .A1(n9854), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9558) );
  OAI21_X1 U7927 ( .B1(n9981), .B2(n9557), .A(n6810), .ZN(n9970) );
  NAND2_X1 U7928 ( .A1(n9981), .A2(n9557), .ZN(n6810) );
  NAND2_X1 U7929 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  AOI21_X1 U7930 ( .B1(n9723), .B2(n9547), .A(n9714), .ZN(n9977) );
  NAND2_X1 U7931 ( .A1(n10985), .A2(n10986), .ZN(n10988) );
  INV_X1 U7932 ( .A(n10996), .ZN(n6990) );
  NAND2_X1 U7933 ( .A1(n12826), .A2(n12825), .ZN(n6992) );
  NOR2_X1 U7934 ( .A1(n12866), .A2(n12867), .ZN(n12887) );
  NOR2_X1 U7935 ( .A1(n11916), .A2(n12086), .ZN(n12538) );
  AND2_X1 U7936 ( .A1(n7088), .A2(n12907), .ZN(n7086) );
  INV_X1 U7937 ( .A(n12939), .ZN(n12910) );
  NAND2_X1 U7938 ( .A1(n12918), .A2(n12931), .ZN(n7004) );
  OR2_X1 U7939 ( .A1(n12931), .A2(n12939), .ZN(n7006) );
  NAND2_X1 U7940 ( .A1(n12953), .A2(n6622), .ZN(n12937) );
  NAND2_X1 U7941 ( .A1(n8095), .A2(n12650), .ZN(n8115) );
  INV_X1 U7942 ( .A(n8096), .ZN(n8095) );
  AND2_X1 U7943 ( .A1(n8122), .A2(n8121), .ZN(n12951) );
  NAND2_X1 U7944 ( .A1(n11871), .A2(n12060), .ZN(n12955) );
  OR2_X1 U7945 ( .A1(n13111), .A2(n12738), .ZN(n6772) );
  INV_X1 U7946 ( .A(n13016), .ZN(n12987) );
  OR2_X1 U7947 ( .A1(n8025), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U7948 ( .A1(n11869), .A2(n12470), .ZN(n13021) );
  OR2_X1 U7949 ( .A1(n7953), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7976) );
  AND2_X1 U7950 ( .A1(n12016), .A2(n12024), .ZN(n13077) );
  INV_X1 U7951 ( .A(n7110), .ZN(n7109) );
  NOR2_X1 U7952 ( .A1(n12008), .A2(n7114), .ZN(n7113) );
  AOI21_X1 U7953 ( .B1(n7014), .B2(n15147), .A(n6668), .ZN(n7013) );
  AND2_X1 U7954 ( .A1(n12006), .A2(n12003), .ZN(n14594) );
  OR2_X1 U7955 ( .A1(n7830), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U7956 ( .A1(n11097), .A2(n11096), .ZN(n15152) );
  AND2_X1 U7957 ( .A1(n7762), .A2(n15525), .ZN(n7814) );
  NAND2_X1 U7958 ( .A1(n10653), .A2(n10641), .ZN(n10642) );
  NAND2_X1 U7959 ( .A1(n7011), .A2(n10208), .ZN(n10328) );
  OAI21_X1 U7960 ( .B1(n10644), .B2(n15193), .A(n7096), .ZN(n10330) );
  OAI21_X1 U7961 ( .B1(n10208), .B2(n7010), .A(n11918), .ZN(n7008) );
  NAND2_X1 U7962 ( .A1(n10202), .A2(n7001), .ZN(n15164) );
  NAND2_X1 U7963 ( .A1(n15181), .A2(n15188), .ZN(n7001) );
  INV_X1 U7964 ( .A(n15149), .ZN(n15191) );
  NAND2_X1 U7965 ( .A1(n8113), .A2(n8112), .ZN(n13103) );
  NAND2_X1 U7966 ( .A1(n8042), .A2(n8041), .ZN(n12611) );
  NAND2_X1 U7967 ( .A1(n11888), .A2(n11887), .ZN(n11896) );
  NAND2_X1 U7968 ( .A1(n7142), .A2(n7141), .ZN(n11888) );
  AND2_X1 U7969 ( .A1(n7143), .A2(n6739), .ZN(n7141) );
  NAND2_X1 U7970 ( .A1(n7132), .A2(n8130), .ZN(n8145) );
  INV_X1 U7971 ( .A(n7147), .ZN(n7146) );
  NOR2_X1 U7972 ( .A1(n8057), .A2(n7150), .ZN(n7149) );
  INV_X1 U7973 ( .A(n8039), .ZN(n7150) );
  NOR2_X1 U7974 ( .A1(n8019), .A2(n7163), .ZN(n7162) );
  NAND2_X1 U7975 ( .A1(n7968), .A2(n7646), .ZN(n7989) );
  AND2_X1 U7976 ( .A1(n7922), .A2(n7923), .ZN(n7948) );
  AND2_X1 U7977 ( .A1(n9158), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7862) );
  NOR2_X1 U7978 ( .A1(n7822), .A2(n7172), .ZN(n7171) );
  AND2_X1 U7979 ( .A1(n8990), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7822) );
  INV_X1 U7980 ( .A(n7803), .ZN(n7172) );
  NAND2_X1 U7981 ( .A1(n7771), .A2(n7748), .ZN(n7802) );
  CLKBUF_X1 U7982 ( .A(n7727), .Z(n7728) );
  NAND2_X1 U7983 ( .A1(n7155), .A2(n7693), .ZN(n7154) );
  INV_X1 U7984 ( .A(n7695), .ZN(n7155) );
  NAND2_X1 U7985 ( .A1(n7156), .A2(n7693), .ZN(n7696) );
  NAND2_X1 U7986 ( .A1(n7692), .A2(n7577), .ZN(n7156) );
  INV_X1 U7987 ( .A(n7663), .ZN(n7298) );
  AND2_X1 U7988 ( .A1(n10814), .A2(n8694), .ZN(n6942) );
  INV_X1 U7989 ( .A(n15070), .ZN(n9536) );
  XNOR2_X1 U7990 ( .A(n8426), .B(n9536), .ZN(n8495) );
  XNOR2_X1 U7991 ( .A(n8426), .B(n12148), .ZN(n8434) );
  NOR2_X1 U7992 ( .A1(n6957), .A2(n13254), .ZN(n6956) );
  INV_X1 U7993 ( .A(n6958), .ZN(n6957) );
  INV_X1 U7994 ( .A(n13269), .ZN(n7454) );
  INV_X1 U7995 ( .A(n8878), .ZN(n7447) );
  INV_X1 U7996 ( .A(n11042), .ZN(n7449) );
  NAND2_X1 U7997 ( .A1(n13236), .A2(n13237), .ZN(n7448) );
  NAND2_X1 U7998 ( .A1(n7448), .A2(n6595), .ZN(n11632) );
  XNOR2_X1 U7999 ( .A(n9826), .B(n8426), .ZN(n8507) );
  NAND2_X1 U8000 ( .A1(n6931), .A2(n6663), .ZN(n9266) );
  INV_X1 U8001 ( .A(n9268), .ZN(n6934) );
  INV_X1 U8002 ( .A(n7456), .ZN(n7455) );
  OAI21_X1 U8003 ( .B1(n7457), .B2(n7459), .A(n13243), .ZN(n7456) );
  AND2_X1 U8004 ( .A1(n8693), .A2(n8670), .ZN(n7463) );
  NAND2_X1 U8005 ( .A1(n6688), .A2(n6608), .ZN(n12379) );
  AND2_X1 U8006 ( .A1(n8817), .A2(n8816), .ZN(n13480) );
  AND4_X1 U8007 ( .A1(n8730), .A2(n8729), .A3(n8728), .A4(n8727), .ZN(n12239)
         );
  AND4_X1 U8008 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12195)
         );
  AND4_X1 U8009 ( .A1(n8550), .A2(n8549), .A3(n8548), .A4(n8547), .ZN(n12187)
         );
  NAND2_X1 U8010 ( .A1(n8436), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8442) );
  NOR2_X1 U8011 ( .A1(n13469), .A2(n13498), .ZN(n13470) );
  NAND2_X1 U8012 ( .A1(n7042), .A2(n7041), .ZN(n13498) );
  AOI21_X1 U8013 ( .B1(n7278), .B2(n7280), .A(n7276), .ZN(n7275) );
  INV_X1 U8014 ( .A(n13486), .ZN(n7276) );
  NAND2_X1 U8015 ( .A1(n13571), .A2(n13665), .ZN(n6832) );
  NOR2_X1 U8016 ( .A1(n13722), .A2(n7052), .ZN(n7051) );
  INV_X1 U8017 ( .A(n7053), .ZN(n7052) );
  NAND2_X1 U8018 ( .A1(n7380), .A2(n7377), .ZN(n13560) );
  INV_X1 U8019 ( .A(n7279), .ZN(n7278) );
  OAI21_X1 U8020 ( .B1(n13593), .B2(n7280), .A(n13584), .ZN(n7279) );
  INV_X1 U8021 ( .A(n13485), .ZN(n7280) );
  NAND2_X1 U8022 ( .A1(n7421), .A2(n7423), .ZN(n13597) );
  INV_X1 U8023 ( .A(n7424), .ZN(n7423) );
  OAI21_X1 U8024 ( .B1(n6625), .B2(n7425), .A(n13598), .ZN(n7424) );
  NAND2_X1 U8025 ( .A1(n13592), .A2(n13593), .ZN(n13591) );
  AND2_X1 U8026 ( .A1(n13741), .A2(n13650), .ZN(n13638) );
  AND2_X1 U8027 ( .A1(n13757), .A2(n13507), .ZN(n7283) );
  NAND2_X1 U8028 ( .A1(n13506), .A2(n13668), .ZN(n7282) );
  AOI21_X1 U8029 ( .B1(n7414), .B2(n12422), .A(n6685), .ZN(n7412) );
  INV_X1 U8030 ( .A(n7414), .ZN(n7413) );
  AND2_X1 U8031 ( .A1(n12426), .A2(n6636), .ZN(n7414) );
  INV_X1 U8032 ( .A(n7292), .ZN(n7291) );
  INV_X1 U8033 ( .A(n12424), .ZN(n7402) );
  NAND2_X1 U8034 ( .A1(n12227), .A2(n7408), .ZN(n7407) );
  OAI21_X1 U8035 ( .B1(n12227), .B2(n7408), .A(n10860), .ZN(n10861) );
  NOR2_X1 U8036 ( .A1(n14944), .A2(n10693), .ZN(n10801) );
  AOI21_X1 U8037 ( .B1(n10524), .B2(n7260), .A(n7259), .ZN(n7258) );
  INV_X1 U8038 ( .A(n10687), .ZN(n7259) );
  INV_X1 U8039 ( .A(n7261), .ZN(n7260) );
  OR2_X1 U8040 ( .A1(n13320), .A2(n9826), .ZN(n9766) );
  INV_X1 U8041 ( .A(n13352), .ZN(n7466) );
  OR2_X1 U8042 ( .A1(n9528), .A2(n15070), .ZN(n9512) );
  AND2_X1 U8043 ( .A1(n9006), .A2(n8885), .ZN(n13667) );
  NAND2_X1 U8044 ( .A1(n7387), .A2(n6624), .ZN(n13556) );
  NAND2_X1 U8045 ( .A1(n7380), .A2(n7378), .ZN(n7387) );
  NOR2_X1 U8046 ( .A1(n13518), .A2(n7379), .ZN(n7378) );
  AND2_X1 U8047 ( .A1(n8856), .A2(n8855), .ZN(n15048) );
  NAND2_X1 U8048 ( .A1(n8284), .A2(n8283), .ZN(n11007) );
  NOR2_X1 U8049 ( .A1(n8675), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8717) );
  INV_X1 U8050 ( .A(n10590), .ZN(n10587) );
  NAND2_X1 U8051 ( .A1(n10374), .A2(n6620), .ZN(n10403) );
  NAND2_X1 U8052 ( .A1(n10827), .A2(n6609), .ZN(n13871) );
  AOI21_X1 U8053 ( .B1(n7479), .B2(n6592), .A(n6677), .ZN(n7478) );
  OR2_X1 U8054 ( .A1(n10128), .A2(n10127), .ZN(n10141) );
  INV_X1 U8055 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10140) );
  INV_X1 U8056 ( .A(n13936), .ZN(n7506) );
  INV_X1 U8057 ( .A(n11731), .ZN(n7508) );
  OR2_X1 U8058 ( .A1(n11370), .A2(n11369), .ZN(n11385) );
  OR2_X1 U8059 ( .A1(n10450), .A2(n10449), .ZN(n10590) );
  NAND2_X1 U8060 ( .A1(n13926), .A2(n13927), .ZN(n13925) );
  INV_X1 U8061 ( .A(n6790), .ZN(n11570) );
  AND2_X1 U8062 ( .A1(n9251), .A2(n9055), .ZN(n9371) );
  NAND2_X1 U8063 ( .A1(n11707), .A2(n13958), .ZN(n7519) );
  AND2_X1 U8064 ( .A1(n11410), .A2(n11409), .ZN(n13861) );
  INV_X1 U8065 ( .A(n11541), .ZN(n9660) );
  NAND2_X1 U8066 ( .A1(n12132), .A2(n11162), .ZN(n9322) );
  NAND2_X1 U8067 ( .A1(n14790), .A2(n11573), .ZN(n10314) );
  AOI21_X1 U8068 ( .B1(n14134), .B2(n7211), .A(n14120), .ZN(n7210) );
  NOR2_X1 U8069 ( .A1(n14359), .A2(n6891), .ZN(n6890) );
  INV_X1 U8070 ( .A(n14167), .ZN(n6891) );
  OR2_X1 U8071 ( .A1(n14359), .A2(n14167), .ZN(n6781) );
  NOR2_X1 U8072 ( .A1(n14131), .A2(n14134), .ZN(n14130) );
  NOR2_X1 U8073 ( .A1(n14149), .A2(n14160), .ZN(n14148) );
  NAND2_X1 U8074 ( .A1(n14209), .A2(n7369), .ZN(n7368) );
  NAND2_X1 U8075 ( .A1(n7373), .A2(n13973), .ZN(n7372) );
  OR2_X1 U8076 ( .A1(n11572), .A2(n9369), .ZN(n14189) );
  INV_X1 U8077 ( .A(n14747), .ZN(n14191) );
  INV_X1 U8078 ( .A(n7368), .ZN(n14184) );
  AOI21_X1 U8079 ( .B1(n7196), .B2(n7198), .A(n6666), .ZN(n7193) );
  NOR2_X1 U8080 ( .A1(n11830), .A2(n7200), .ZN(n7199) );
  INV_X1 U8081 ( .A(n11828), .ZN(n7200) );
  INV_X1 U8082 ( .A(n11805), .ZN(n6880) );
  NAND2_X1 U8083 ( .A1(n7363), .A2(n6619), .ZN(n7362) );
  NAND2_X1 U8084 ( .A1(n14277), .A2(n14291), .ZN(n14276) );
  OR2_X1 U8085 ( .A1(n13877), .A2(n10844), .ZN(n10572) );
  NAND2_X1 U8086 ( .A1(n7357), .A2(n11593), .ZN(n7356) );
  INV_X1 U8087 ( .A(n11675), .ZN(n11573) );
  NAND2_X1 U8088 ( .A1(n14779), .A2(n11588), .ZN(n9688) );
  OAI21_X1 U8089 ( .B1(n9727), .B2(n9728), .A(n11204), .ZN(n9952) );
  INV_X1 U8090 ( .A(n14091), .ZN(n14319) );
  INV_X1 U8091 ( .A(n14837), .ZN(n14790) );
  NAND2_X1 U8092 ( .A1(n11382), .A2(n11565), .ZN(n11384) );
  OR2_X1 U8093 ( .A1(n9338), .A2(n9359), .ZN(n14899) );
  INV_X1 U8094 ( .A(n14902), .ZN(n14863) );
  AND2_X1 U8095 ( .A1(n9053), .A2(n9054), .ZN(n9354) );
  NAND2_X1 U8096 ( .A1(n7566), .A2(n7565), .ZN(n7564) );
  XNOR2_X1 U8097 ( .A(n11171), .B(n11170), .ZN(n12347) );
  XNOR2_X1 U8098 ( .A(n11167), .B(n11166), .ZN(n12291) );
  XNOR2_X1 U8099 ( .A(n7174), .B(n9230), .ZN(n8978) );
  NAND2_X1 U8100 ( .A1(n7061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8101 ( .A1(n8971), .A2(n7061), .ZN(n8977) );
  MUX2_X1 U8102 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8970), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8971) );
  NAND2_X1 U8103 ( .A1(n6789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U8104 ( .A(n9246), .B(n9245), .ZN(n11576) );
  NAND2_X1 U8105 ( .A1(n9292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9246) );
  XNOR2_X1 U8106 ( .A(n8652), .B(n8651), .ZN(n10568) );
  AOI21_X1 U8107 ( .B1(n7535), .B2(n7537), .A(n7534), .ZN(n7533) );
  NAND2_X1 U8108 ( .A1(n6875), .A2(n6877), .ZN(n6874) );
  INV_X1 U8109 ( .A(n6914), .ZN(n14505) );
  NAND2_X1 U8110 ( .A1(n7126), .A2(n14513), .ZN(n14514) );
  NAND2_X1 U8111 ( .A1(n15546), .A2(n15547), .ZN(n7126) );
  AOI21_X1 U8112 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14460), .A(n14459), .ZN(
        n14482) );
  NOR2_X1 U8113 ( .A1(n14517), .A2(n14516), .ZN(n14459) );
  OAI22_X1 U8114 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14477), .B1(n14479), 
        .B2(n14467), .ZN(n14528) );
  OAI211_X1 U8115 ( .C1(n14685), .C2(n6918), .A(n7122), .B(n6917), .ZN(n7125)
         );
  OR2_X1 U8116 ( .A1(n14687), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7122) );
  OR2_X1 U8117 ( .A1(n7123), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8118 ( .A1(n14527), .A2(n6915), .ZN(n6917) );
  AOI21_X1 U8119 ( .B1(n14540), .B2(n14539), .A(n14567), .ZN(n14573) );
  AND3_X1 U8120 ( .A1(n7829), .A2(n7828), .A3(n7827), .ZN(n15159) );
  NOR2_X1 U8121 ( .A1(n7496), .A2(n12699), .ZN(n7494) );
  NOR2_X1 U8122 ( .A1(n7497), .A2(n7499), .ZN(n7496) );
  INV_X1 U8123 ( .A(n7500), .ZN(n7497) );
  NAND2_X1 U8124 ( .A1(n7500), .A2(n7501), .ZN(n7498) );
  NAND2_X1 U8125 ( .A1(n12552), .A2(n12553), .ZN(n12551) );
  AND4_X1 U8126 ( .A1(n7998), .A2(n7997), .A3(n7996), .A4(n7995), .ZN(n13053)
         );
  AND3_X1 U8128 ( .A1(n7812), .A2(n7811), .A3(n7810), .ZN(n12675) );
  OR2_X1 U8129 ( .A1(n7843), .A2(n8936), .ZN(n7665) );
  AOI21_X1 U8130 ( .B1(n12488), .B2(n6587), .A(n8172), .ZN(n12909) );
  AND2_X1 U8131 ( .A1(n7311), .A2(n6999), .ZN(n10729) );
  INV_X1 U8132 ( .A(n12779), .ZN(n12778) );
  XNOR2_X1 U8133 ( .A(n6992), .B(n12864), .ZN(n12827) );
  AOI21_X1 U8134 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n12875), .A(n12874), .ZN(
        n12876) );
  NAND2_X1 U8135 ( .A1(n12877), .A2(n6809), .ZN(n12879) );
  OR2_X1 U8136 ( .A1(n12888), .A2(n13141), .ZN(n6809) );
  OAI21_X1 U8137 ( .B1(n12892), .B2(n12891), .A(n6763), .ZN(n6762) );
  INV_X1 U8138 ( .A(n12893), .ZN(n6763) );
  XNOR2_X1 U8139 ( .A(n6824), .B(n12890), .ZN(n12892) );
  AND2_X1 U8140 ( .A1(n12487), .A2(n12486), .ZN(n13091) );
  OR2_X1 U8141 ( .A1(n6590), .A2(n12499), .ZN(n8147) );
  AND2_X1 U8142 ( .A1(n8178), .A2(n8177), .ZN(n13214) );
  NOR2_X1 U8143 ( .A1(n6604), .A2(n14939), .ZN(n7436) );
  INV_X1 U8144 ( .A(n7442), .ZN(n7438) );
  NAND2_X1 U8145 ( .A1(n7444), .A2(n7440), .ZN(n7439) );
  OR2_X1 U8146 ( .A1(n13231), .A2(n12515), .ZN(n7444) );
  NAND2_X1 U8147 ( .A1(n8463), .A2(n8462), .ZN(n8465) );
  AND2_X1 U8148 ( .A1(n8471), .A2(n8472), .ZN(n9112) );
  NAND2_X1 U8149 ( .A1(n8883), .A2(n15037), .ZN(n14943) );
  INV_X1 U8150 ( .A(n12455), .ZN(n6750) );
  NAND2_X1 U8151 ( .A1(n12453), .A2(n12454), .ZN(n7543) );
  AND2_X1 U8152 ( .A1(n7542), .A2(n12456), .ZN(n7540) );
  INV_X1 U8153 ( .A(n12352), .ZN(n12460) );
  INV_X1 U8154 ( .A(n13469), .ZN(n13704) );
  XNOR2_X1 U8155 ( .A(n6786), .B(n13489), .ZN(n13710) );
  NAND2_X1 U8156 ( .A1(n7383), .A2(n7388), .ZN(n6786) );
  NAND2_X1 U8157 ( .A1(n8882), .A2(n15056), .ZN(n15037) );
  NAND2_X1 U8158 ( .A1(n11377), .A2(n11376), .ZN(n14381) );
  NAND2_X1 U8159 ( .A1(n6744), .A2(n6650), .ZN(n6743) );
  AND2_X1 U8160 ( .A1(n11580), .A2(n11581), .ZN(n6745) );
  NAND2_X1 U8161 ( .A1(n11497), .A2(n11496), .ZN(n13971) );
  NAND2_X1 U8162 ( .A1(n11477), .A2(n11476), .ZN(n14140) );
  NAND2_X1 U8163 ( .A1(n11460), .A2(n11459), .ZN(n13972) );
  NAND2_X1 U8164 ( .A1(n11427), .A2(n11426), .ZN(n14183) );
  OR2_X1 U8165 ( .A1(n10314), .A2(n9378), .ZN(n14783) );
  NAND2_X1 U8166 ( .A1(n6872), .A2(n11333), .ZN(n14271) );
  NAND2_X1 U8167 ( .A1(n11331), .A2(n11565), .ZN(n6872) );
  OAI211_X1 U8168 ( .C1(n14335), .C2(n6689), .A(n7218), .B(n7212), .ZN(n14328)
         );
  NAND2_X1 U8169 ( .A1(n7221), .A2(n14094), .ZN(n7218) );
  OR2_X1 U8170 ( .A1(n14909), .A2(n7220), .ZN(n7219) );
  INV_X1 U8171 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U8172 ( .A1(n7248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U8173 ( .A1(n14550), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7128) );
  OR2_X1 U8174 ( .A1(n14685), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6916) );
  AND2_X1 U8175 ( .A1(n6912), .A2(n6910), .ZN(n6909) );
  INV_X1 U8176 ( .A(n14697), .ZN(n6910) );
  XNOR2_X1 U8177 ( .A(n14573), .B(n14572), .ZN(n14571) );
  NAND2_X1 U8178 ( .A1(n6799), .A2(n11203), .ZN(n6798) );
  AND2_X1 U8179 ( .A1(n11212), .A2(n11211), .ZN(n7228) );
  OAI21_X1 U8180 ( .B1(n7230), .B2(n11212), .A(n11210), .ZN(n7229) );
  INV_X1 U8181 ( .A(n7222), .ZN(n11235) );
  NAND2_X1 U8182 ( .A1(n7225), .A2(n11233), .ZN(n11232) );
  NAND2_X1 U8183 ( .A1(n11249), .A2(n11248), .ZN(n11253) );
  NAND2_X1 U8184 ( .A1(n15075), .A2(n12275), .ZN(n6854) );
  NAND2_X1 U8185 ( .A1(n12331), .A2(n13320), .ZN(n6855) );
  NAND2_X1 U8186 ( .A1(n11268), .A2(n11270), .ZN(n6791) );
  NAND2_X1 U8187 ( .A1(n6851), .A2(n6850), .ZN(n12201) );
  NAND2_X1 U8188 ( .A1(n11279), .A2(n11284), .ZN(n7238) );
  INV_X1 U8189 ( .A(n12213), .ZN(n7308) );
  MUX2_X1 U8190 ( .A(n13974), .B(n14381), .S(n11351), .Z(n11379) );
  AND2_X1 U8191 ( .A1(n11336), .A2(n7581), .ZN(n11365) );
  OR2_X1 U8192 ( .A1(n11334), .A2(n11335), .ZN(n7581) );
  NAND2_X1 U8193 ( .A1(n6859), .A2(n6858), .ZN(n6862) );
  NAND2_X1 U8194 ( .A1(n12221), .A2(n12220), .ZN(n6858) );
  AOI21_X1 U8195 ( .B1(n12219), .B2(n6648), .A(n6860), .ZN(n6857) );
  NAND2_X1 U8196 ( .A1(n12221), .A2(n6639), .ZN(n6856) );
  AND2_X1 U8197 ( .A1(n12236), .A2(n12237), .ZN(n6840) );
  NAND2_X1 U8198 ( .A1(n6839), .A2(n6838), .ZN(n6837) );
  INV_X1 U8199 ( .A(n12237), .ZN(n6838) );
  INV_X1 U8200 ( .A(n12236), .ZN(n6839) );
  AOI21_X1 U8201 ( .B1(n12238), .B2(n6837), .A(n6835), .ZN(n6834) );
  NAND2_X1 U8202 ( .A1(n6836), .A2(n12244), .ZN(n6835) );
  NAND2_X1 U8203 ( .A1(n6840), .A2(n6837), .ZN(n6836) );
  MUX2_X1 U8204 ( .A(n14168), .B(n14370), .S(n11504), .Z(n11418) );
  MUX2_X1 U8205 ( .A(n14183), .B(n14364), .S(n11431), .Z(n11432) );
  INV_X1 U8206 ( .A(n12253), .ZN(n7316) );
  NAND2_X1 U8207 ( .A1(n7245), .A2(n11432), .ZN(n7244) );
  INV_X1 U8208 ( .A(n12259), .ZN(n7331) );
  NAND2_X1 U8209 ( .A1(n11468), .A2(n11465), .ZN(n6986) );
  NAND2_X1 U8210 ( .A1(n11484), .A2(n11487), .ZN(n7252) );
  INV_X1 U8211 ( .A(n6986), .ZN(n6985) );
  NAND2_X1 U8212 ( .A1(n6848), .A2(n7325), .ZN(n12265) );
  AOI21_X1 U8213 ( .B1(n6593), .B2(n7326), .A(n6676), .ZN(n7325) );
  NOR2_X1 U8214 ( .A1(n6847), .A2(n12269), .ZN(n6846) );
  AND2_X1 U8215 ( .A1(n11298), .A2(n11805), .ZN(n11585) );
  NOR2_X1 U8216 ( .A1(n11525), .A2(n11522), .ZN(n7255) );
  INV_X1 U8217 ( .A(n11522), .ZN(n7254) );
  INV_X1 U8218 ( .A(SI_16_), .ZN(n8337) );
  NAND2_X1 U8219 ( .A1(n7306), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U8220 ( .A1(n9598), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7305) );
  NOR2_X1 U8221 ( .A1(n12469), .A2(n7023), .ZN(n7022) );
  INV_X1 U8222 ( .A(n12467), .ZN(n7023) );
  INV_X1 U8223 ( .A(n11527), .ZN(n6978) );
  INV_X1 U8224 ( .A(n8754), .ZN(n7077) );
  NAND2_X1 U8225 ( .A1(n8332), .A2(n6611), .ZN(n7539) );
  AOI21_X1 U8226 ( .B1(n8671), .B2(n6969), .A(n6611), .ZN(n6968) );
  OAI21_X1 U8227 ( .B1(n7614), .B2(n8925), .A(n7293), .ZN(n8297) );
  NAND2_X1 U8228 ( .A1(n6927), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7293) );
  INV_X1 U8229 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7257) );
  NOR2_X1 U8230 ( .A1(n9995), .A2(n7303), .ZN(n9599) );
  NOR2_X1 U8231 ( .A1(n7304), .A2(n9585), .ZN(n7303) );
  NAND2_X1 U8232 ( .A1(n9599), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U8233 ( .A1(n12770), .A2(n6723), .ZN(n10736) );
  OR2_X1 U8234 ( .A1(n12495), .A2(n12909), .ZN(n12077) );
  OR2_X1 U8235 ( .A1(n13054), .A2(n12477), .ZN(n12996) );
  OR2_X1 U8236 ( .A1(n12473), .A2(n12472), .ZN(n13010) );
  OR2_X1 U8237 ( .A1(n13136), .A2(n13053), .ZN(n12035) );
  INV_X1 U8238 ( .A(n13077), .ZN(n7105) );
  NOR2_X1 U8239 ( .A1(n6659), .A2(n6602), .ZN(n7014) );
  INV_X1 U8240 ( .A(n11096), .ZN(n7015) );
  OAI21_X1 U8241 ( .B1(n7149), .B2(n7148), .A(n8074), .ZN(n7147) );
  INV_X1 U8242 ( .A(n8003), .ZN(n7163) );
  NAND2_X1 U8243 ( .A1(n7888), .A2(n10574), .ZN(n7905) );
  NAND2_X1 U8244 ( .A1(n6768), .A2(n7522), .ZN(n7644) );
  INV_X1 U8245 ( .A(n6817), .ZN(n6768) );
  INV_X1 U8246 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7587) );
  CLKBUF_X1 U8247 ( .A(n7698), .Z(n7699) );
  NAND2_X1 U8248 ( .A1(n7492), .A2(n7660), .ZN(n7675) );
  AND2_X1 U8249 ( .A1(n7586), .A2(n7299), .ZN(n7492) );
  INV_X1 U8250 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7586) );
  INV_X1 U8251 ( .A(n7460), .ZN(n7459) );
  AND2_X1 U8252 ( .A1(n12304), .A2(n12433), .ZN(n7582) );
  OR2_X1 U8253 ( .A1(n13487), .A2(n12431), .ZN(n12432) );
  INV_X1 U8254 ( .A(n7570), .ZN(n7274) );
  NAND2_X1 U8255 ( .A1(n7392), .A2(n13555), .ZN(n7391) );
  INV_X1 U8256 ( .A(n13518), .ZN(n7392) );
  NAND2_X1 U8257 ( .A1(n7074), .A2(n6603), .ZN(n13491) );
  OR2_X1 U8258 ( .A1(n13515), .A2(n13250), .ZN(n13482) );
  INV_X1 U8259 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U8260 ( .A1(n6691), .A2(n7264), .ZN(n7261) );
  NAND2_X1 U8261 ( .A1(n10254), .A2(n6649), .ZN(n7262) );
  OR2_X1 U8262 ( .A1(n8623), .A2(n15436), .ZN(n8637) );
  INV_X1 U8263 ( .A(n11074), .ZN(n7044) );
  NAND2_X1 U8264 ( .A1(n7043), .A2(n13506), .ZN(n13693) );
  INV_X1 U8265 ( .A(n7046), .ZN(n11055) );
  AOI21_X1 U8266 ( .B1(n7396), .B2(n12414), .A(n6656), .ZN(n7395) );
  INV_X1 U8267 ( .A(n10065), .ZN(n7396) );
  INV_X1 U8268 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8265) );
  OR2_X1 U8269 ( .A1(n8599), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U8270 ( .A1(n14096), .A2(n7351), .ZN(n7350) );
  INV_X1 U8271 ( .A(n11843), .ZN(n7351) );
  INV_X1 U8272 ( .A(n7372), .ZN(n7371) );
  INV_X1 U8273 ( .A(n11829), .ZN(n7198) );
  INV_X1 U8274 ( .A(n7197), .ZN(n7196) );
  OAI21_X1 U8275 ( .B1(n7199), .B2(n7198), .A(n11831), .ZN(n7197) );
  NOR2_X1 U8276 ( .A1(n14402), .A2(n14271), .ZN(n7063) );
  INV_X1 U8277 ( .A(n11238), .ZN(n7065) );
  NAND2_X1 U8278 ( .A1(n9659), .A2(n7188), .ZN(n7187) );
  INV_X1 U8279 ( .A(n9658), .ZN(n7189) );
  AND2_X2 U8280 ( .A1(n9247), .A2(n11576), .ZN(n11574) );
  CLKBUF_X1 U8281 ( .A(n11574), .Z(n6785) );
  OR2_X1 U8282 ( .A1(n14660), .A2(n11801), .ZN(n11802) );
  OR2_X1 U8283 ( .A1(n9338), .A2(n11570), .ZN(n9358) );
  INV_X1 U8284 ( .A(n11557), .ZN(n7566) );
  NOR2_X1 U8285 ( .A1(n11559), .A2(n11552), .ZN(n7565) );
  NAND2_X1 U8286 ( .A1(n11167), .A2(n11166), .ZN(n11557) );
  INV_X1 U8287 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9230) );
  INV_X1 U8288 ( .A(n7550), .ZN(n7549) );
  OAI21_X1 U8289 ( .B1(n7552), .B2(n7551), .A(n11156), .ZN(n7550) );
  OAI21_X1 U8290 ( .B1(n8824), .B2(n8837), .A(n7072), .ZN(n11153) );
  AOI21_X1 U8291 ( .B1(n7558), .B2(n7561), .A(n6727), .ZN(n7556) );
  OR2_X1 U8292 ( .A1(n8346), .A2(n9479), .ZN(n7562) );
  AND2_X1 U8293 ( .A1(n8346), .A2(n9479), .ZN(n7561) );
  NAND2_X1 U8294 ( .A1(n6895), .A2(n6968), .ZN(n8709) );
  NAND2_X1 U8295 ( .A1(n8652), .A2(n6898), .ZN(n6895) );
  INV_X1 U8296 ( .A(n8306), .ZN(n6877) );
  INV_X1 U8297 ( .A(n8312), .ZN(n7534) );
  OR2_X1 U8298 ( .A1(n8958), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8987) );
  OR2_X1 U8299 ( .A1(n8945), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U8300 ( .A1(n8297), .A2(SI_4_), .ZN(n8299) );
  NAND2_X1 U8301 ( .A1(n8294), .A2(SI_3_), .ZN(n8295) );
  NAND2_X1 U8302 ( .A1(n8288), .A2(SI_1_), .ZN(n8290) );
  NAND3_X1 U8303 ( .A1(n11679), .A2(n6870), .A3(n6869), .ZN(n7532) );
  INV_X1 U8304 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6870) );
  INV_X1 U8305 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6869) );
  OAI21_X1 U8306 ( .B1(n14486), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14447), .ZN(
        n14448) );
  XOR2_X1 U8307 ( .A(n14448), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n14502) );
  AOI22_X1 U8308 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14506), .B1(n14507), .B2(
        n14452), .ZN(n14454) );
  OR2_X1 U8309 ( .A1(n14506), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14452) );
  OAI21_X1 U8310 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14458), .A(n14457), .ZN(
        n14516) );
  INV_X1 U8311 ( .A(n7123), .ZN(n6915) );
  AND2_X1 U8312 ( .A1(n14687), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7123) );
  INV_X1 U8313 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6913) );
  NOR2_X1 U8314 ( .A1(n7787), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7762) );
  INV_X1 U8315 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15525) );
  AND2_X1 U8316 ( .A1(n8054), .A2(n8033), .ZN(n7524) );
  AND2_X1 U8317 ( .A1(n7873), .A2(n7872), .ZN(n11121) );
  AND2_X1 U8318 ( .A1(n8126), .A2(n8125), .ZN(n12618) );
  INV_X1 U8319 ( .A(n12659), .ZN(n7714) );
  NAND2_X1 U8320 ( .A1(n8044), .A2(n8043), .ZN(n8065) );
  INV_X1 U8321 ( .A(n8045), .ZN(n8044) );
  AND3_X1 U8322 ( .A1(n7848), .A2(n7847), .A3(n7846), .ZN(n14610) );
  AND4_X1 U8323 ( .A1(n7855), .A2(n7854), .A3(n7853), .A4(n7852), .ZN(n12691)
         );
  NAND2_X1 U8324 ( .A1(n7683), .A2(n7684), .ZN(n7094) );
  OAI21_X1 U8325 ( .B1(n9555), .B2(n15200), .A(n6827), .ZN(n9546) );
  NAND2_X1 U8326 ( .A1(n9555), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6827) );
  INV_X1 U8327 ( .A(n9570), .ZN(n7295) );
  AOI21_X1 U8328 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9598), .A(n9612), .ZN(
        n9990) );
  NOR2_X1 U8329 ( .A1(n7302), .A2(n10233), .ZN(n7301) );
  AOI21_X1 U8330 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10225), .A(n10223), .ZN(
        n10553) );
  OAI21_X1 U8331 ( .B1(n10238), .B2(n10237), .A(n10236), .ZN(n12766) );
  NAND2_X1 U8332 ( .A1(n12771), .A2(n12772), .ZN(n12770) );
  NAND2_X1 U8333 ( .A1(n6998), .A2(n6997), .ZN(n10978) );
  NAND2_X1 U8334 ( .A1(n10728), .A2(n7324), .ZN(n6997) );
  NOR2_X1 U8335 ( .A1(n12793), .A2(n12792), .ZN(n12800) );
  OAI21_X1 U8336 ( .B1(n12840), .B2(n12839), .A(n12838), .ZN(n12841) );
  NAND2_X1 U8337 ( .A1(n12858), .A2(n12859), .ZN(n12877) );
  NAND2_X1 U8338 ( .A1(n6826), .A2(n6825), .ZN(n6824) );
  OAI21_X1 U8339 ( .B1(n7028), .B2(n7030), .A(n12955), .ZN(n7027) );
  NAND2_X1 U8340 ( .A1(n12984), .A2(n7030), .ZN(n7025) );
  NAND2_X1 U8341 ( .A1(n7032), .A2(n7035), .ZN(n12969) );
  NAND2_X1 U8342 ( .A1(n7032), .A2(n7030), .ZN(n12971) );
  NAND2_X1 U8343 ( .A1(n7100), .A2(n7102), .ZN(n7099) );
  AND2_X1 U8344 ( .A1(n12055), .A2(n12054), .ZN(n12989) );
  INV_X1 U8345 ( .A(n8011), .ZN(n8010) );
  AND2_X1 U8346 ( .A1(n13008), .A2(n13007), .ZN(n13040) );
  NAND2_X1 U8347 ( .A1(n7018), .A2(n6598), .ZN(n12995) );
  AND2_X1 U8348 ( .A1(n12036), .A2(n12033), .ZN(n13054) );
  INV_X1 U8349 ( .A(n7929), .ZN(n7928) );
  INV_X1 U8350 ( .A(n11129), .ZN(n12005) );
  AND2_X1 U8351 ( .A1(n11939), .A2(n12001), .ZN(n14608) );
  INV_X1 U8352 ( .A(n12745), .ZN(n14603) );
  NAND2_X1 U8353 ( .A1(n15152), .A2(n15151), .ZN(n15150) );
  NAND2_X1 U8354 ( .A1(n10920), .A2(n10919), .ZN(n11097) );
  AND4_X1 U8355 ( .A1(n7835), .A2(n7834), .A3(n7833), .A4(n7832), .ZN(n14602)
         );
  NAND2_X1 U8356 ( .A1(n7814), .A2(n7813), .ZN(n7830) );
  AND4_X1 U8357 ( .A1(n7757), .A2(n7756), .A3(n7755), .A4(n7754), .ZN(n10921)
         );
  AND4_X1 U8358 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), .ZN(n10703)
         );
  NAND2_X1 U8359 ( .A1(n7000), .A2(n10643), .ZN(n10701) );
  AND2_X1 U8360 ( .A1(n11981), .A2(n11975), .ZN(n11919) );
  OR2_X1 U8361 ( .A1(n7785), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7787) );
  AND2_X1 U8362 ( .A1(n11971), .A2(n11974), .ZN(n11966) );
  INV_X1 U8363 ( .A(n10199), .ZN(n15173) );
  AND2_X1 U8364 ( .A1(n9846), .A2(n9845), .ZN(n10348) );
  AND2_X1 U8365 ( .A1(n11906), .A2(n10275), .ZN(n12899) );
  NAND2_X1 U8366 ( .A1(n8094), .A2(n8093), .ZN(n13107) );
  INV_X1 U8367 ( .A(n6590), .ZN(n8006) );
  AND2_X1 U8368 ( .A1(n12922), .A2(n13098), .ZN(n13112) );
  AND2_X1 U8369 ( .A1(n8286), .A2(n13215), .ZN(n9843) );
  NAND2_X1 U8370 ( .A1(n9849), .A2(n10350), .ZN(n15183) );
  INV_X1 U8371 ( .A(n15183), .ZN(n15210) );
  XNOR2_X1 U8372 ( .A(P3_IR_REG_0__SCAN_IN), .B(keyinput87), .ZN(n15424) );
  NAND2_X1 U8373 ( .A1(n7117), .A2(n7595), .ZN(n7116) );
  INV_X1 U8374 ( .A(n7118), .ZN(n7117) );
  AOI21_X1 U8375 ( .B1(n11880), .B2(n7144), .A(n6737), .ZN(n7143) );
  INV_X1 U8376 ( .A(n8163), .ZN(n7144) );
  NAND2_X1 U8377 ( .A1(n7131), .A2(n8146), .ZN(n8162) );
  AOI21_X1 U8378 ( .B1(n6736), .B2(n8080), .A(n7159), .ZN(n7158) );
  AND2_X1 U8379 ( .A1(n7531), .A2(n8192), .ZN(n7530) );
  NAND2_X1 U8380 ( .A1(n6774), .A2(n6773), .ZN(n8092) );
  XNOR2_X1 U8381 ( .A(n8193), .B(n8192), .ZN(n9550) );
  NAND2_X1 U8382 ( .A1(n7621), .A2(n7531), .ZN(n8191) );
  AND2_X1 U8383 ( .A1(n7640), .A2(n6631), .ZN(n11943) );
  INV_X1 U8384 ( .A(n7621), .ZN(n7642) );
  INV_X1 U8385 ( .A(n8001), .ZN(n6801) );
  AND2_X1 U8386 ( .A1(n7965), .A2(n7944), .ZN(n7945) );
  INV_X1 U8387 ( .A(n7169), .ZN(n7168) );
  OAI22_X1 U8388 ( .A1(n7171), .A2(n7170), .B1(n9106), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7169) );
  OR2_X1 U8389 ( .A1(n7772), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7742) );
  OR2_X1 U8390 ( .A1(n7742), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7806) );
  OAI22_X1 U8391 ( .A1(n7782), .A2(n7746), .B1(P1_DATAO_REG_6__SCAN_IN), .B2(
        n8947), .ZN(n7769) );
  XNOR2_X1 U8392 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7781) );
  NAND2_X1 U8393 ( .A1(n7154), .A2(n7718), .ZN(n7151) );
  INV_X1 U8394 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7130) );
  INV_X1 U8395 ( .A(n13260), .ZN(n6947) );
  INV_X1 U8396 ( .A(n6948), .ZN(n6944) );
  NOR2_X1 U8397 ( .A1(n8699), .A2(n10818), .ZN(n8725) );
  AND2_X1 U8398 ( .A1(n8781), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8791) );
  NOR2_X1 U8399 ( .A1(n7443), .A2(n7446), .ZN(n7442) );
  INV_X1 U8400 ( .A(n12511), .ZN(n7443) );
  NOR2_X1 U8401 ( .A1(n6594), .A2(n6959), .ZN(n6958) );
  INV_X1 U8402 ( .A(n8771), .ZN(n6959) );
  NAND2_X1 U8403 ( .A1(n8791), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8810) );
  AND2_X1 U8404 ( .A1(n8725), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U8405 ( .A1(n6937), .A2(n6936), .ZN(n6935) );
  INV_X1 U8406 ( .A(n8494), .ZN(n6936) );
  INV_X1 U8407 ( .A(n8495), .ZN(n6937) );
  NAND2_X1 U8408 ( .A1(n9110), .A2(n6932), .ZN(n6931) );
  INV_X1 U8409 ( .A(n8472), .ZN(n6933) );
  INV_X1 U8410 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8603) );
  OR2_X1 U8411 ( .A1(n8604), .A2(n8603), .ZN(n8623) );
  NAND2_X1 U8412 ( .A1(n7458), .A2(n6732), .ZN(n7457) );
  NAND2_X1 U8413 ( .A1(n7459), .A2(n13290), .ZN(n7458) );
  NOR2_X1 U8414 ( .A1(n8828), .A2(n13282), .ZN(n8841) );
  NOR2_X1 U8415 ( .A1(n13289), .A2(n13290), .ZN(n13288) );
  NAND2_X1 U8416 ( .A1(n11083), .A2(n8771), .ZN(n13289) );
  NAND2_X1 U8417 ( .A1(n13258), .A2(n13260), .ZN(n13259) );
  AND2_X1 U8418 ( .A1(n12353), .A2(n12460), .ZN(n9006) );
  AOI21_X1 U8419 ( .B1(n6942), .B2(n6941), .A(n6646), .ZN(n6940) );
  INV_X1 U8420 ( .A(n12278), .ZN(n12280) );
  AND3_X1 U8421 ( .A1(n12342), .A2(n12341), .A3(n12340), .ZN(n12382) );
  OR2_X1 U8422 ( .A1(n8451), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U8423 ( .A1(n13799), .A2(n6581), .ZN(n7563) );
  NOR2_X1 U8424 ( .A1(n13492), .A2(n7271), .ZN(n7270) );
  INV_X1 U8425 ( .A(n7272), .ZN(n7271) );
  INV_X1 U8426 ( .A(n7267), .ZN(n7265) );
  AOI21_X1 U8427 ( .B1(n7272), .B2(n7269), .A(n7268), .ZN(n7267) );
  NAND2_X1 U8428 ( .A1(n7274), .A2(n13520), .ZN(n7269) );
  NOR2_X1 U8429 ( .A1(n7272), .A2(n13492), .ZN(n7268) );
  NOR2_X1 U8430 ( .A1(n7391), .A2(n7379), .ZN(n7376) );
  INV_X1 U8431 ( .A(n12296), .ZN(n12321) );
  NAND2_X1 U8432 ( .A1(n13638), .A2(n7055), .ZN(n13603) );
  AND2_X1 U8433 ( .A1(n13515), .A2(n13514), .ZN(n7432) );
  NAND2_X1 U8434 ( .A1(n13638), .A2(n13624), .ZN(n13618) );
  NOR2_X1 U8435 ( .A1(n7411), .A2(n13508), .ZN(n7410) );
  NAND2_X1 U8436 ( .A1(n13478), .A2(n13505), .ZN(n7285) );
  OR2_X1 U8437 ( .A1(n8760), .A2(n11090), .ZN(n8762) );
  NOR2_X1 U8438 ( .A1(n8762), .A2(n8410), .ZN(n8781) );
  NAND2_X1 U8439 ( .A1(n7046), .A2(n7045), .ZN(n11074) );
  AOI21_X1 U8440 ( .B1(n12425), .B2(n7289), .A(n6660), .ZN(n7287) );
  AOI21_X1 U8441 ( .B1(n10861), .B2(n7397), .A(n7398), .ZN(n11018) );
  NOR2_X1 U8442 ( .A1(n7400), .A2(n7404), .ZN(n7397) );
  NAND2_X1 U8443 ( .A1(n6586), .A2(n12239), .ZN(n7405) );
  NOR2_X1 U8444 ( .A1(n8637), .A2(n8636), .ZN(n8660) );
  NAND2_X1 U8445 ( .A1(n10686), .A2(n13313), .ZN(n7419) );
  OAI21_X1 U8446 ( .B1(n10686), .B2(n13313), .A(n10776), .ZN(n7420) );
  OR2_X1 U8447 ( .A1(n10776), .A2(n14934), .ZN(n10521) );
  NAND2_X1 U8448 ( .A1(n7262), .A2(n7261), .ZN(n10523) );
  NAND2_X1 U8449 ( .A1(n10523), .A2(n10524), .ZN(n10688) );
  NOR2_X1 U8450 ( .A1(n15119), .A2(n7048), .ZN(n7047) );
  INV_X1 U8451 ( .A(n7049), .ZN(n7048) );
  NAND2_X1 U8452 ( .A1(n10254), .A2(n10253), .ZN(n7263) );
  NAND2_X1 U8453 ( .A1(n9806), .A2(n7049), .ZN(n10261) );
  NAND2_X1 U8454 ( .A1(n9806), .A2(n12196), .ZN(n10069) );
  AOI21_X1 U8455 ( .B1(n9743), .B2(n9746), .A(n9535), .ZN(n9799) );
  AND3_X1 U8456 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8546) );
  AND4_X1 U8457 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n12192)
         );
  INV_X1 U8458 ( .A(n15084), .ZN(n12179) );
  OR2_X1 U8459 ( .A1(n8466), .A2(n13325), .ZN(n7574) );
  OAI21_X1 U8460 ( .B1(n6930), .B2(n6926), .A(n8466), .ZN(n6928) );
  NOR2_X1 U8461 ( .A1(n11550), .A2(n8916), .ZN(n6930) );
  NAND2_X1 U8462 ( .A1(n12148), .A2(n9128), .ZN(n9904) );
  CLKBUF_X1 U8463 ( .A(n9525), .Z(n12403) );
  AOI21_X1 U8464 ( .B1(n7384), .B2(n7389), .A(n6687), .ZN(n7381) );
  INV_X1 U8465 ( .A(n7384), .ZN(n7382) );
  CLKBUF_X1 U8466 ( .A(n9126), .Z(n9127) );
  NAND2_X1 U8467 ( .A1(n10067), .A2(n12414), .ZN(n10258) );
  NAND2_X1 U8468 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  INV_X1 U8469 ( .A(n15097), .ZN(n15118) );
  OR2_X1 U8470 ( .A1(n15033), .A2(n12457), .ZN(n15097) );
  AND2_X1 U8471 ( .A1(n8272), .A2(n6733), .ZN(n8868) );
  NOR2_X1 U8472 ( .A1(n8373), .A2(n13800), .ZN(n8374) );
  INV_X1 U8473 ( .A(n8383), .ZN(n8376) );
  NAND2_X1 U8474 ( .A1(n8389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8390) );
  AND2_X2 U8475 ( .A1(n8423), .A2(n8255), .ZN(n8481) );
  INV_X1 U8476 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8255) );
  INV_X1 U8477 ( .A(n13833), .ZN(n11700) );
  OR2_X1 U8478 ( .A1(n9699), .A2(n10287), .ZN(n10128) );
  NAND2_X1 U8479 ( .A1(n10370), .A2(n6657), .ZN(n10373) );
  NAND2_X1 U8480 ( .A1(n6776), .A2(n11789), .ZN(n6775) );
  NOR2_X1 U8481 ( .A1(n13909), .A2(n7480), .ZN(n7479) );
  NOR2_X1 U8482 ( .A1(n13842), .A2(n6592), .ZN(n7480) );
  NAND2_X1 U8483 ( .A1(n11173), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11326) );
  OR2_X1 U8484 ( .A1(n11326), .A2(n11316), .ZN(n11318) );
  CLKBUF_X1 U8485 ( .A(n9922), .Z(n7490) );
  INV_X1 U8486 ( .A(n11404), .ZN(n11176) );
  NAND2_X1 U8487 ( .A1(n10421), .A2(n10420), .ZN(n10450) );
  AND2_X1 U8488 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n10420) );
  OR2_X1 U8489 ( .A1(n10141), .A2(n10140), .ZN(n10419) );
  NAND2_X1 U8490 ( .A1(n10675), .A2(n10674), .ZN(n10827) );
  INV_X1 U8491 ( .A(n10677), .ZN(n10674) );
  AOI21_X1 U8493 ( .B1(n7478), .B2(n7476), .A(n7475), .ZN(n7474) );
  INV_X1 U8494 ( .A(n13880), .ZN(n7475) );
  INV_X1 U8495 ( .A(n7479), .ZN(n7476) );
  INV_X1 U8496 ( .A(n7478), .ZN(n7477) );
  AND3_X1 U8497 ( .A1(n11544), .A2(n11543), .A3(n11542), .ZN(n11577) );
  BUF_X1 U8498 ( .A(n9322), .Z(n11541) );
  INV_X1 U8499 ( .A(n11540), .ZN(n11511) );
  INV_X1 U8500 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15477) );
  AOI21_X1 U8501 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n9225) );
  INV_X1 U8502 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10127) );
  OAI21_X1 U8503 ( .B1(n14056), .B2(n14054), .A(n14055), .ZN(n14053) );
  INV_X1 U8504 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8962) );
  NOR2_X1 U8505 ( .A1(n14099), .A2(n7349), .ZN(n7344) );
  NAND2_X1 U8506 ( .A1(n14099), .A2(n7348), .ZN(n7346) );
  NAND2_X1 U8507 ( .A1(n11849), .A2(n14098), .ZN(n14101) );
  OAI21_X1 U8508 ( .B1(n14337), .B2(n11797), .A(n11843), .ZN(n12113) );
  OR2_X1 U8509 ( .A1(n7210), .A2(n6596), .ZN(n7208) );
  NOR2_X1 U8510 ( .A1(n7584), .A2(n6596), .ZN(n7209) );
  NAND2_X1 U8511 ( .A1(n14139), .A2(n14345), .ZN(n14121) );
  INV_X1 U8512 ( .A(n6886), .ZN(n6885) );
  INV_X1 U8513 ( .A(n6888), .ZN(n6887) );
  NOR2_X1 U8514 ( .A1(n14154), .A2(n14137), .ZN(n14139) );
  NAND2_X1 U8515 ( .A1(n14153), .A2(n14158), .ZN(n14154) );
  AOI21_X1 U8516 ( .B1(n7360), .B2(n7359), .A(n6681), .ZN(n7358) );
  INV_X1 U8517 ( .A(n6619), .ZN(n7359) );
  NAND2_X1 U8518 ( .A1(n14282), .A2(n7063), .ZN(n14267) );
  NAND2_X1 U8519 ( .A1(n11824), .A2(n11823), .ZN(n14288) );
  OR2_X1 U8520 ( .A1(n14667), .A2(n10565), .ZN(n10566) );
  NAND2_X1 U8521 ( .A1(n7179), .A2(n7176), .ZN(n7175) );
  INV_X1 U8522 ( .A(n11598), .ZN(n10444) );
  AOI21_X1 U8523 ( .B1(n7355), .B2(n10183), .A(n6626), .ZN(n7353) );
  NAND2_X1 U8524 ( .A1(n9709), .A2(n6597), .ZN(n14758) );
  AND2_X1 U8525 ( .A1(n9370), .A2(n9369), .ZN(n14747) );
  INV_X1 U8526 ( .A(n11592), .ZN(n14746) );
  NAND2_X1 U8527 ( .A1(n11211), .A2(n11209), .ZN(n7339) );
  INV_X1 U8528 ( .A(n11588), .ZN(n14778) );
  INV_X1 U8529 ( .A(n14125), .ZN(n14345) );
  NAND2_X1 U8530 ( .A1(n6616), .A2(n11828), .ZN(n14246) );
  INV_X1 U8531 ( .A(n14899), .ZN(n14876) );
  AND2_X1 U8533 ( .A1(n10316), .A2(n10315), .ZN(n10321) );
  XNOR2_X1 U8534 ( .A(n11518), .B(n11517), .ZN(n12305) );
  AND2_X1 U8535 ( .A1(n8253), .A2(n8969), .ZN(n9054) );
  NAND2_X1 U8536 ( .A1(n7548), .A2(n6614), .ZN(n11481) );
  AND2_X1 U8537 ( .A1(n8963), .A2(n9245), .ZN(n7247) );
  NAND2_X1 U8538 ( .A1(n8349), .A2(n9964), .ZN(n8801) );
  XNOR2_X1 U8539 ( .A(n8415), .B(n8414), .ZN(n11302) );
  OAI21_X1 U8540 ( .B1(n8328), .B2(n7080), .A(n7078), .ZN(n8753) );
  NAND2_X1 U8541 ( .A1(n8232), .A2(n8234), .ZN(n7232) );
  NAND2_X1 U8542 ( .A1(n6892), .A2(n6654), .ZN(n8736) );
  XNOR2_X1 U8543 ( .A(n8712), .B(n8711), .ZN(n11280) );
  AND2_X1 U8544 ( .A1(n9858), .A2(n9450), .ZN(n10576) );
  NAND2_X1 U8545 ( .A1(n8328), .A2(n8327), .ZN(n8672) );
  NOR2_X1 U8546 ( .A1(n9104), .A2(n9103), .ZN(n14704) );
  OR2_X1 U8547 ( .A1(n8987), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9100) );
  OAI21_X1 U8548 ( .B1(n8553), .B2(n7537), .A(n8572), .ZN(n7536) );
  INV_X1 U8549 ( .A(n8309), .ZN(n7537) );
  NAND2_X1 U8550 ( .A1(n8541), .A2(n8306), .ZN(n8554) );
  NAND2_X1 U8551 ( .A1(n8554), .A2(n8553), .ZN(n8555) );
  NAND2_X1 U8552 ( .A1(n8539), .A2(n8538), .ZN(n8541) );
  INV_X1 U8553 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U8554 ( .A1(n14440), .A2(n6907), .ZN(n14490) );
  NAND2_X1 U8555 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6908), .ZN(n6907) );
  INV_X1 U8556 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6908) );
  XNOR2_X1 U8557 ( .A(n14443), .B(n6903), .ZN(n14498) );
  INV_X1 U8558 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n6903) );
  XNOR2_X1 U8559 ( .A(n14486), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14488) );
  INV_X1 U8560 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U8561 ( .A1(n14509), .A2(n14510), .ZN(n14512) );
  INV_X1 U8562 ( .A(n6902), .ZN(n14518) );
  OAI21_X1 U8563 ( .B1(n14549), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6637), .ZN(
        n6902) );
  AOI21_X1 U8564 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14462), .A(n14461), .ZN(
        n14481) );
  AND2_X1 U8565 ( .A1(n7483), .A2(n10943), .ZN(n7482) );
  OR2_X1 U8566 ( .A1(n7884), .A2(n7485), .ZN(n7483) );
  AOI21_X1 U8567 ( .B1(n7513), .B2(n7515), .A(n7511), .ZN(n7510) );
  INV_X1 U8568 ( .A(n7513), .ZN(n7512) );
  INV_X1 U8569 ( .A(n12588), .ZN(n7511) );
  NAND2_X1 U8570 ( .A1(n7509), .A2(n7513), .ZN(n12589) );
  NAND2_X1 U8571 ( .A1(n6813), .A2(n7514), .ZN(n7509) );
  NAND2_X1 U8572 ( .A1(n8034), .A2(n8033), .ZN(n12608) );
  INV_X1 U8573 ( .A(n11121), .ZN(n14597) );
  NAND2_X1 U8574 ( .A1(n7487), .A2(n7884), .ZN(n10974) );
  INV_X1 U8575 ( .A(n10971), .ZN(n7487) );
  AND2_X1 U8576 ( .A1(n8103), .A2(n8102), .ZN(n12972) );
  OAI21_X1 U8577 ( .B1(n9552), .B2(n6765), .A(n6764), .ZN(n9504) );
  NAND2_X1 U8578 ( .A1(n9552), .A2(n13229), .ZN(n6764) );
  NAND2_X1 U8579 ( .A1(n10974), .A2(n7885), .ZN(n10946) );
  NAND2_X1 U8580 ( .A1(n6674), .A2(n8064), .ZN(n11651) );
  INV_X1 U8581 ( .A(n14610), .ZN(n12694) );
  NAND2_X1 U8582 ( .A1(n9915), .A2(n9916), .ZN(n12576) );
  NAND2_X1 U8583 ( .A1(n7517), .A2(n7983), .ZN(n12701) );
  NAND2_X1 U8584 ( .A1(n7514), .A2(n7517), .ZN(n12702) );
  AND2_X1 U8585 ( .A1(n9835), .A2(n8219), .ZN(n12726) );
  AND2_X1 U8586 ( .A1(n8157), .A2(n8156), .ZN(n12923) );
  NAND2_X1 U8587 ( .A1(n9835), .A2(n8218), .ZN(n12729) );
  INV_X1 U8588 ( .A(n12743), .ZN(n13076) );
  OR2_X1 U8589 ( .A1(n12101), .A2(n12100), .ZN(n7139) );
  INV_X1 U8590 ( .A(n12923), .ZN(n12737) );
  NAND2_X1 U8591 ( .A1(n8139), .A2(n8138), .ZN(n12939) );
  INV_X1 U8592 ( .A(n12691), .ZN(n15156) );
  INV_X1 U8593 ( .A(n14602), .ZN(n12746) );
  INV_X1 U8594 ( .A(n10921), .ZN(n12747) );
  INV_X1 U8595 ( .A(n10703), .ZN(n12631) );
  NOR2_X1 U8596 ( .A1(n10493), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10299) );
  NOR2_X1 U8597 ( .A1(n9715), .A2(n10302), .ZN(n9714) );
  NAND2_X1 U8598 ( .A1(n10294), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U8599 ( .A1(n9583), .A2(n9582), .B1(n9581), .B2(n9580), .ZN(n9607)
         );
  AOI21_X1 U8600 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(n10046) );
  AOI21_X1 U8601 ( .B1(n10043), .B2(n10023), .A(n10022), .ZN(n10238) );
  AOI21_X1 U8602 ( .B1(n12766), .B2(n12765), .A(n12764), .ZN(n12769) );
  NOR2_X1 U8603 ( .A1(n10726), .A2(n7311), .ZN(n10725) );
  INV_X1 U8604 ( .A(n10728), .ZN(n6995) );
  INV_X1 U8605 ( .A(n10729), .ZN(n6996) );
  XNOR2_X1 U8606 ( .A(n10978), .B(n7323), .ZN(n10882) );
  XNOR2_X1 U8607 ( .A(n12813), .B(n12814), .ZN(n12780) );
  NOR2_X1 U8608 ( .A1(n12780), .A2(n12781), .ZN(n12815) );
  NOR2_X1 U8609 ( .A1(n12800), .A2(n6814), .ZN(n12840) );
  NOR2_X1 U8610 ( .A1(n6816), .A2(n12814), .ZN(n6814) );
  INV_X1 U8612 ( .A(n12802), .ZN(n6816) );
  INV_X1 U8613 ( .A(n6992), .ZN(n12848) );
  NAND2_X1 U8614 ( .A1(n11899), .A2(n11898), .ZN(n14617) );
  NAND2_X1 U8615 ( .A1(n12525), .A2(n6747), .ZN(n12526) );
  INV_X1 U8616 ( .A(n12907), .ZN(n12904) );
  NAND2_X1 U8617 ( .A1(n7087), .A2(n7088), .ZN(n12903) );
  NAND2_X1 U8618 ( .A1(n7093), .A2(n11873), .ZN(n12919) );
  NAND2_X1 U8619 ( .A1(n12943), .A2(n12064), .ZN(n7093) );
  OR2_X1 U8620 ( .A1(n6590), .A2(n15368), .ZN(n8131) );
  NAND2_X1 U8621 ( .A1(n13021), .A2(n12047), .ZN(n13000) );
  NAND2_X1 U8622 ( .A1(n7024), .A2(n12467), .ZN(n13061) );
  NAND2_X1 U8623 ( .A1(n13073), .A2(n12465), .ZN(n7024) );
  OAI21_X1 U8624 ( .B1(n11122), .B2(n7109), .A(n7106), .ZN(n13078) );
  NAND2_X1 U8625 ( .A1(n7112), .A2(n12007), .ZN(n11865) );
  NAND2_X1 U8626 ( .A1(n11122), .A2(n7113), .ZN(n7112) );
  AND3_X1 U8627 ( .A1(n7732), .A2(n7731), .A3(n7730), .ZN(n12632) );
  NAND2_X1 U8628 ( .A1(n10328), .A2(n10327), .ZN(n10329) );
  OAI21_X1 U8629 ( .B1(n15168), .B2(n15195), .A(n7095), .ZN(n15169) );
  NAND2_X1 U8630 ( .A1(n10354), .A2(n15184), .ZN(n15198) );
  INV_X1 U8631 ( .A(n15184), .ZN(n15178) );
  INV_X1 U8632 ( .A(n11913), .ZN(n13167) );
  NOR2_X1 U8633 ( .A1(n12899), .A2(n12898), .ZN(n14616) );
  INV_X1 U8634 ( .A(n12611), .ZN(n13187) );
  INV_X2 U8635 ( .A(n15223), .ZN(n15225) );
  INV_X1 U8636 ( .A(n9504), .ZN(n10496) );
  OR2_X1 U8637 ( .A1(n15223), .A2(n15183), .ZN(n13212) );
  AND2_X1 U8638 ( .A1(n9550), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13215) );
  XNOR2_X1 U8639 ( .A(n7633), .B(n7120), .ZN(n10941) );
  NAND2_X1 U8640 ( .A1(n7629), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U8641 ( .A1(n7145), .A2(n8059), .ZN(n8075) );
  NAND2_X1 U8642 ( .A1(n8040), .A2(n7149), .ZN(n7145) );
  XNOR2_X1 U8643 ( .A(n8194), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U8644 ( .A1(n6631), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U8645 ( .A1(n8040), .A2(n8039), .ZN(n8058) );
  INV_X1 U8646 ( .A(n11943), .ZN(n10350) );
  INV_X1 U8647 ( .A(SI_20_), .ZN(n9964) );
  INV_X1 U8648 ( .A(n12849), .ZN(n12864) );
  NOR2_X1 U8649 ( .A1(n7950), .A2(n7968), .ZN(n12830) );
  INV_X1 U8650 ( .A(SI_14_), .ZN(n15462) );
  INV_X1 U8651 ( .A(SI_13_), .ZN(n9107) );
  INV_X1 U8652 ( .A(SI_11_), .ZN(n8956) );
  NAND2_X1 U8653 ( .A1(n7167), .A2(n7821), .ZN(n7841) );
  NAND2_X1 U8654 ( .A1(n7173), .A2(n7171), .ZN(n7167) );
  NAND2_X1 U8655 ( .A1(n7173), .A2(n7803), .ZN(n7823) );
  NAND2_X1 U8656 ( .A1(n7156), .A2(n7153), .ZN(n7719) );
  INV_X1 U8657 ( .A(n7154), .ZN(n7153) );
  NAND2_X1 U8658 ( .A1(n7661), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7300) );
  AOI21_X1 U8659 ( .B1(n7662), .B2(n7299), .A(n7298), .ZN(n7297) );
  NAND2_X1 U8660 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7612) );
  OR2_X1 U8661 ( .A1(n8888), .A2(n8285), .ZN(n9008) );
  INV_X1 U8662 ( .A(n13586), .ZN(n13517) );
  NAND2_X1 U8663 ( .A1(n10628), .A2(n6942), .ZN(n10813) );
  AND2_X1 U8664 ( .A1(n10628), .A2(n8694), .ZN(n10815) );
  NOR2_X1 U8665 ( .A1(n13288), .A2(n7460), .ZN(n13245) );
  NAND2_X1 U8666 ( .A1(n8447), .A2(n8446), .ZN(n9117) );
  NAND2_X1 U8667 ( .A1(n7453), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U8668 ( .A1(n11083), .A2(n6956), .ZN(n6955) );
  INV_X1 U8669 ( .A(n13254), .ZN(n6954) );
  AOI21_X1 U8670 ( .B1(n11083), .B2(n6958), .A(n7453), .ZN(n13253) );
  CLKBUF_X1 U8671 ( .A(n14935), .Z(n14936) );
  NOR2_X1 U8672 ( .A1(n6925), .A2(n6924), .ZN(n6923) );
  INV_X1 U8673 ( .A(n13237), .ZN(n6924) );
  NAND2_X1 U8674 ( .A1(n11632), .A2(n11631), .ZN(n11635) );
  NAND2_X1 U8675 ( .A1(n10931), .A2(n8734), .ZN(n11041) );
  AND2_X1 U8676 ( .A1(n8849), .A2(n8848), .ZN(n13596) );
  NAND2_X1 U8677 ( .A1(n7448), .A2(n8853), .ZN(n8876) );
  NAND2_X1 U8678 ( .A1(n6931), .A2(n6935), .ZN(n9269) );
  OAI21_X1 U8679 ( .B1(n13289), .B2(n7457), .A(n7455), .ZN(n13271) );
  NAND2_X1 U8680 ( .A1(n8790), .A2(n8789), .ZN(n13752) );
  NAND2_X1 U8681 ( .A1(n14936), .A2(n7463), .ZN(n10628) );
  NAND2_X1 U8682 ( .A1(n14935), .A2(n8670), .ZN(n10627) );
  INV_X1 U8683 ( .A(n13314), .ZN(n12211) );
  OR2_X1 U8684 ( .A1(n8630), .A2(n8629), .ZN(n8631) );
  NAND2_X1 U8685 ( .A1(n13259), .A2(n8537), .ZN(n9459) );
  INV_X1 U8686 ( .A(n13570), .ZN(n13594) );
  INV_X1 U8687 ( .A(n13596), .ZN(n13483) );
  INV_X1 U8688 ( .A(n13480), .ZN(n13666) );
  OR3_X1 U8689 ( .A1(n8665), .A2(n8664), .A3(n8663), .ZN(n13312) );
  INV_X1 U8690 ( .A(n12187), .ZN(n13318) );
  INV_X1 U8691 ( .A(n9528), .ZN(n13321) );
  OR2_X1 U8692 ( .A1(n11642), .A2(n9020), .ZN(n8453) );
  OR2_X1 U8693 ( .A1(n8451), .A2(n8437), .ZN(n8440) );
  INV_X1 U8694 ( .A(n13470), .ZN(n13471) );
  NAND2_X1 U8695 ( .A1(n13545), .A2(n13544), .ZN(n13546) );
  NAND2_X1 U8696 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  NAND2_X1 U8697 ( .A1(n13570), .A2(n13667), .ZN(n6831) );
  NAND2_X1 U8698 ( .A1(n13591), .A2(n13485), .ZN(n13583) );
  NAND2_X1 U8699 ( .A1(n7422), .A2(n7426), .ZN(n13599) );
  NAND2_X1 U8700 ( .A1(n7430), .A2(n6625), .ZN(n7422) );
  OR2_X1 U8701 ( .A1(n10880), .A2(n8825), .ZN(n8827) );
  OAI21_X1 U8702 ( .B1(n11079), .B2(n7413), .A(n7412), .ZN(n13686) );
  NAND2_X1 U8703 ( .A1(n7415), .A2(n7414), .ZN(n13504) );
  AND2_X1 U8704 ( .A1(n7415), .A2(n6636), .ZN(n11080) );
  NAND2_X1 U8705 ( .A1(n11079), .A2(n11078), .ZN(n7415) );
  NAND2_X1 U8706 ( .A1(n7290), .A2(n7289), .ZN(n11049) );
  NAND2_X1 U8707 ( .A1(n7399), .A2(n7401), .ZN(n11016) );
  NAND2_X1 U8708 ( .A1(n10861), .A2(n7403), .ZN(n7399) );
  NAND2_X1 U8709 ( .A1(n10861), .A2(n7407), .ZN(n10900) );
  NAND2_X1 U8710 ( .A1(n8657), .A2(n8656), .ZN(n14944) );
  INV_X1 U8711 ( .A(n10776), .ZN(n12215) );
  NAND2_X1 U8712 ( .A1(n8500), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U8713 ( .A1(n8484), .A2(n7466), .ZN(n7465) );
  OAI21_X2 U8714 ( .B1(n9330), .B2(n8825), .A(n7575), .ZN(n15070) );
  NAND2_X1 U8715 ( .A1(n15045), .A2(n9492), .ZN(n13677) );
  INV_X1 U8716 ( .A(n13639), .ZN(n13694) );
  NAND2_X1 U8717 ( .A1(n15045), .A2(n13459), .ZN(n13639) );
  AND3_X2 U8718 ( .A1(n9489), .A2(n9142), .A3(n10781), .ZN(n15141) );
  INV_X1 U8719 ( .A(n13714), .ZN(n6811) );
  AND2_X2 U8720 ( .A1(n10782), .A2(n10781), .ZN(n15129) );
  AND2_X1 U8721 ( .A1(n8888), .A2(n8873), .ZN(n15056) );
  AND2_X1 U8722 ( .A1(n8395), .A2(n7434), .ZN(n7433) );
  INV_X1 U8723 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U8724 ( .A1(n8360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U8725 ( .A1(n8360), .A2(n8277), .ZN(n13815) );
  INV_X1 U8726 ( .A(n12436), .ZN(n13459) );
  INV_X1 U8727 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9625) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9938) );
  INV_X1 U8729 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9856) );
  AND2_X1 U8730 ( .A1(n8677), .A2(n8676), .ZN(n15011) );
  INV_X1 U8731 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9279) );
  INV_X1 U8732 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9161) );
  INV_X1 U8733 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8991) );
  INV_X1 U8734 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8961) );
  INV_X1 U8735 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8952) );
  INV_X1 U8736 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8926) );
  INV_X1 U8737 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U8738 ( .A1(n11689), .A2(n11688), .ZN(n13830) );
  OR2_X1 U8739 ( .A1(n11749), .A2(n11748), .ZN(n11750) );
  CLKBUF_X1 U8740 ( .A(n10667), .Z(n10408) );
  AND2_X1 U8741 ( .A1(n13934), .A2(n7507), .ZN(n13850) );
  NAND2_X1 U8742 ( .A1(n13934), .A2(n11731), .ZN(n13851) );
  NAND2_X1 U8743 ( .A1(n11340), .A2(n11339), .ZN(n14388) );
  NAND2_X1 U8744 ( .A1(n10374), .A2(n10373), .ZN(n10376) );
  NAND2_X1 U8745 ( .A1(n9305), .A2(n7488), .ZN(n9386) );
  NAND2_X1 U8746 ( .A1(n10827), .A2(n10826), .ZN(n13873) );
  NAND2_X1 U8747 ( .A1(n7473), .A2(n7478), .ZN(n13879) );
  NAND2_X1 U8748 ( .A1(n13841), .A2(n7479), .ZN(n7473) );
  AOI21_X1 U8749 ( .B1(n13841), .B2(n13842), .A(n6592), .ZN(n13908) );
  INV_X1 U8750 ( .A(n7505), .ZN(n7503) );
  AOI21_X1 U8751 ( .B1(n7507), .B2(n7506), .A(n6684), .ZN(n7505) );
  CLKBUF_X1 U8752 ( .A(n11684), .Z(n10838) );
  INV_X1 U8753 ( .A(n13951), .ZN(n13916) );
  NAND2_X1 U8754 ( .A1(n9362), .A2(n11627), .ZN(n13949) );
  OR2_X1 U8755 ( .A1(n9355), .A2(n9373), .ZN(n13955) );
  INV_X1 U8756 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15522) );
  NAND2_X1 U8757 ( .A1(n7518), .A2(n11708), .ZN(n13957) );
  INV_X1 U8758 ( .A(n7519), .ZN(n7518) );
  INV_X1 U8759 ( .A(n13955), .ZN(n13959) );
  NAND2_X1 U8760 ( .A1(n11442), .A2(n11441), .ZN(n14167) );
  OR2_X1 U8761 ( .A1(n11390), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9325) );
  OR2_X1 U8762 ( .A1(n11494), .A2(n9323), .ZN(n9327) );
  OR2_X1 U8763 ( .A1(n9666), .A2(n9237), .ZN(n9242) );
  OR2_X1 U8764 ( .A1(n9322), .A2(n9239), .ZN(n9240) );
  NOR2_X1 U8765 ( .A1(n9078), .A2(n9077), .ZN(n14041) );
  NOR2_X1 U8766 ( .A1(n9465), .A2(n9464), .ZN(n9467) );
  XNOR2_X1 U8767 ( .A(n9859), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11281) );
  NOR2_X1 U8768 ( .A1(n10499), .A2(n14718), .ZN(n10502) );
  INV_X1 U8769 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n11679) );
  AND2_X1 U8770 ( .A1(n9065), .A2(n14426), .ZN(n14738) );
  NAND2_X1 U8771 ( .A1(n11569), .A2(n11568), .ZN(n14314) );
  NAND2_X1 U8772 ( .A1(n11533), .A2(n11532), .ZN(n14091) );
  NAND2_X1 U8773 ( .A1(n11189), .A2(n11188), .ZN(n14113) );
  NAND2_X1 U8774 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  AOI21_X1 U8775 ( .B1(n12120), .B2(n14902), .A(n12119), .ZN(n12121) );
  NAND2_X1 U8776 ( .A1(n14131), .A2(n7211), .ZN(n7207) );
  OR2_X1 U8777 ( .A1(n14148), .A2(n6888), .ZN(n14133) );
  NOR2_X1 U8778 ( .A1(n14148), .A2(n6890), .ZN(n14135) );
  AND2_X1 U8779 ( .A1(n7203), .A2(n7202), .ZN(n14161) );
  NAND2_X1 U8780 ( .A1(n14209), .A2(n7372), .ZN(n14185) );
  NAND2_X1 U8781 ( .A1(n14383), .A2(n11854), .ZN(n14202) );
  NAND2_X1 U8782 ( .A1(n7195), .A2(n11829), .ZN(n14219) );
  NAND2_X1 U8783 ( .A1(n6616), .A2(n7199), .ZN(n7195) );
  NAND2_X1 U8784 ( .A1(n7362), .A2(n7364), .ZN(n14251) );
  AND2_X1 U8785 ( .A1(n6879), .A2(n6600), .ZN(n7364) );
  NAND2_X1 U8786 ( .A1(n14276), .A2(n11806), .ZN(n14262) );
  NAND2_X1 U8787 ( .A1(n10466), .A2(n11598), .ZN(n7178) );
  NAND2_X1 U8788 ( .A1(n7356), .A2(n7355), .ZN(n10443) );
  AND2_X1 U8789 ( .A1(n7356), .A2(n10154), .ZN(n10155) );
  NAND2_X1 U8790 ( .A1(n14762), .A2(n14764), .ZN(n7190) );
  AND2_X1 U8791 ( .A1(n9332), .A2(n6629), .ZN(n7192) );
  INV_X1 U8792 ( .A(n14273), .ZN(n14793) );
  INV_X1 U8793 ( .A(n14786), .ZN(n14303) );
  OR2_X1 U8794 ( .A1(n14797), .A2(n9710), .ZN(n14786) );
  INV_X1 U8795 ( .A(n14292), .ZN(n14306) );
  AND2_X2 U8796 ( .A1(n10321), .A2(n10319), .ZN(n14929) );
  INV_X1 U8797 ( .A(n14432), .ZN(n9058) );
  INV_X1 U8798 ( .A(n9236), .ZN(n11162) );
  CLKBUF_X1 U8799 ( .A(n8977), .Z(n14426) );
  INV_X1 U8800 ( .A(n9054), .ZN(n14431) );
  NAND2_X1 U8801 ( .A1(n8824), .A2(n8356), .ZN(n8838) );
  INV_X1 U8802 ( .A(n9247), .ZN(n11192) );
  INV_X1 U8803 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10393) );
  INV_X1 U8804 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9898) );
  INV_X1 U8805 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9629) );
  INV_X1 U8806 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n15464) );
  INV_X1 U8807 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9860) );
  INV_X1 U8808 ( .A(n11281), .ZN(n10504) );
  INV_X1 U8809 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10574) );
  INV_X1 U8810 ( .A(n10576), .ZN(n9863) );
  INV_X1 U8811 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9158) );
  INV_X1 U8812 ( .A(n10439), .ZN(n9409) );
  INV_X1 U8813 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8990) );
  INV_X1 U8814 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8960) );
  INV_X1 U8815 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8951) );
  INV_X1 U8816 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8947) );
  INV_X1 U8817 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8933) );
  XNOR2_X1 U8818 ( .A(n14488), .B(n7129), .ZN(n15543) );
  INV_X1 U8819 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7129) );
  XNOR2_X1 U8820 ( .A(n14505), .B(n14974), .ZN(n14548) );
  XNOR2_X1 U8821 ( .A(n14512), .B(n7127), .ZN(n15546) );
  INV_X1 U8822 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7127) );
  XNOR2_X1 U8823 ( .A(n14514), .B(n14515), .ZN(n14549) );
  OAI21_X1 U8824 ( .B1(n14521), .B2(n14554), .A(n14551), .ZN(n14683) );
  AOI21_X1 U8825 ( .B1(n15320), .B2(n14536), .A(n14696), .ZN(n14569) );
  INV_X1 U8826 ( .A(n6758), .ZN(n6757) );
  OAI21_X1 U8827 ( .B1(n13094), .B2(n12734), .A(n12557), .ZN(n6758) );
  NAND2_X1 U8828 ( .A1(n7498), .A2(n12724), .ZN(n7495) );
  INV_X1 U8829 ( .A(n6991), .ZN(n10983) );
  OAI211_X1 U8830 ( .C1(n12897), .C2(n12896), .A(n6761), .B(n6760), .ZN(
        P3_U3201) );
  INV_X1 U8831 ( .A(n6762), .ZN(n6761) );
  NAND2_X1 U8832 ( .A1(n12894), .A2(n12895), .ZN(n6760) );
  NAND2_X1 U8833 ( .A1(n15233), .A2(n6820), .ZN(n6819) );
  INV_X1 U8834 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8835 ( .A1(n9110), .A2(n8472), .ZN(n9152) );
  NAND2_X1 U8836 ( .A1(n7439), .A2(n7445), .ZN(n7437) );
  NAND2_X1 U8837 ( .A1(n7540), .A2(n12455), .ZN(n6751) );
  NAND2_X1 U8838 ( .A1(n6669), .A2(n6750), .ZN(n6749) );
  OR2_X1 U8839 ( .A1(n11626), .A2(n11625), .ZN(n6783) );
  OAI21_X1 U8840 ( .B1(n14328), .B2(n14828), .A(n6779), .ZN(n6883) );
  NAND2_X1 U8841 ( .A1(n14909), .A2(n14906), .ZN(n7217) );
  OAI21_X1 U8842 ( .B1(n14327), .B2(n14908), .A(n7213), .ZN(n7216) );
  NOR2_X1 U8843 ( .A1(n6721), .A2(n14687), .ZN(n14686) );
  INV_X1 U8844 ( .A(n14530), .ZN(n14689) );
  NOR2_X1 U8845 ( .A1(n14534), .A2(n14535), .ZN(n14693) );
  AND2_X1 U8846 ( .A1(n14534), .A2(n14535), .ZN(n14694) );
  XNOR2_X1 U8847 ( .A(n6901), .B(n6632), .ZN(SUB_1596_U4) );
  OAI21_X1 U8848 ( .B1(n14571), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6642), .ZN(
        n6901) );
  INV_X2 U8849 ( .A(n12225), .ZN(n12275) );
  OR2_X1 U8850 ( .A1(n8340), .A2(n8737), .ZN(n6591) );
  AND2_X2 U8851 ( .A1(n11545), .A2(n11194), .ZN(n11431) );
  INV_X1 U8852 ( .A(n13478), .ZN(n13763) );
  INV_X1 U8853 ( .A(n13555), .ZN(n7390) );
  AND2_X1 U8854 ( .A1(n11756), .A2(n11755), .ZN(n6592) );
  AND2_X1 U8855 ( .A1(n7328), .A2(n7327), .ZN(n6593) );
  INV_X1 U8856 ( .A(n9634), .ZN(n9503) );
  INV_X1 U8857 ( .A(n12226), .ZN(n6866) );
  INV_X1 U8858 ( .A(n12739), .ZN(n7036) );
  NAND2_X1 U8859 ( .A1(n11521), .A2(n11520), .ZN(n14330) );
  INV_X1 U8860 ( .A(n14330), .ZN(n14098) );
  OR2_X1 U8861 ( .A1(n7457), .A2(n6722), .ZN(n6594) );
  AND2_X1 U8862 ( .A1(n8853), .A2(n7447), .ZN(n6595) );
  NAND2_X1 U8863 ( .A1(n11384), .A2(n11383), .ZN(n14374) );
  OAI21_X1 U8864 ( .B1(n7455), .B2(n6722), .A(n7454), .ZN(n7453) );
  INV_X1 U8865 ( .A(n14634), .ZN(n12227) );
  INV_X1 U8866 ( .A(n12931), .ZN(n13175) );
  NAND2_X1 U8867 ( .A1(n8132), .A2(n8131), .ZN(n12931) );
  AND2_X1 U8868 ( .A1(n14125), .A2(n14140), .ZN(n6596) );
  AND2_X1 U8869 ( .A1(n10113), .A2(n7065), .ZN(n6597) );
  AND2_X1 U8870 ( .A1(n7019), .A2(n12468), .ZN(n6598) );
  NAND2_X1 U8871 ( .A1(n12194), .A2(n7309), .ZN(n6599) );
  OR2_X1 U8872 ( .A1(n14647), .A2(n14279), .ZN(n6600) );
  AND2_X1 U8873 ( .A1(n6597), .A2(n7064), .ZN(n6601) );
  AND2_X1 U8874 ( .A1(n15151), .A2(n7015), .ZN(n6602) );
  INV_X1 U8875 ( .A(n11842), .ZN(n14160) );
  AND2_X1 U8876 ( .A1(n13543), .A2(n12307), .ZN(n6603) );
  AND4_X1 U8877 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n13042)
         );
  INV_X1 U8878 ( .A(n13042), .ZN(n6752) );
  AND2_X1 U8879 ( .A1(n7440), .A2(n7438), .ZN(n6604) );
  AND2_X1 U8880 ( .A1(n13715), .A2(n13713), .ZN(n6605) );
  NAND2_X1 U8881 ( .A1(n13768), .A2(n12254), .ZN(n6606) );
  INV_X1 U8882 ( .A(n7389), .ZN(n7388) );
  OAI21_X1 U8883 ( .B1(n6624), .B2(n7390), .A(n7393), .ZN(n7389) );
  AND2_X1 U8884 ( .A1(n12980), .A2(n12738), .ZN(n6607) );
  NAND2_X1 U8885 ( .A1(n12374), .A2(n12373), .ZN(n6608) );
  AND2_X1 U8886 ( .A1(n10832), .A2(n10826), .ZN(n6609) );
  OR2_X1 U8887 ( .A1(n10942), .A2(n7486), .ZN(n7485) );
  AND2_X1 U8888 ( .A1(n7207), .A2(n7210), .ZN(n6610) );
  AND2_X1 U8889 ( .A1(n8330), .A2(n9107), .ZN(n6611) );
  INV_X1 U8890 ( .A(n7101), .ZN(n7100) );
  OAI21_X1 U8891 ( .B1(n12470), .B2(n7102), .A(n12050), .ZN(n7101) );
  INV_X1 U8892 ( .A(n12234), .ZN(n12235) );
  AND2_X1 U8893 ( .A1(n8697), .A2(n8696), .ZN(n12234) );
  AND2_X1 U8894 ( .A1(n7063), .A2(n7062), .ZN(n6612) );
  AND3_X1 U8895 ( .A1(n7573), .A2(n7590), .A3(n6713), .ZN(n6613) );
  INV_X1 U8896 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8363) );
  XNOR2_X1 U8897 ( .A(n14271), .B(n6871), .ZN(n14266) );
  INV_X1 U8898 ( .A(n14266), .ZN(n7183) );
  OR2_X1 U8899 ( .A1(n11155), .A2(SI_25_), .ZN(n6614) );
  INV_X1 U8900 ( .A(n8080), .ZN(n6773) );
  NAND2_X1 U8901 ( .A1(n7802), .A2(n7801), .ZN(n7173) );
  NAND2_X2 U8902 ( .A1(n11172), .A2(n13805), .ZN(n8451) );
  INV_X1 U8903 ( .A(n8671), .ZN(n7082) );
  NAND2_X1 U8904 ( .A1(n7628), .A2(n7629), .ZN(n7636) );
  OR2_X1 U8905 ( .A1(n14304), .A2(n14305), .ZN(n6615) );
  NAND2_X1 U8906 ( .A1(n11161), .A2(n11160), .ZN(n11167) );
  NAND2_X1 U8907 ( .A1(n8148), .A2(n8147), .ZN(n12915) );
  OR2_X1 U8908 ( .A1(n14258), .A2(n11827), .ZN(n6616) );
  NAND2_X1 U8909 ( .A1(n11858), .A2(n7204), .ZN(n7203) );
  AND2_X1 U8910 ( .A1(n13757), .A2(n13668), .ZN(n6617) );
  NAND2_X1 U8911 ( .A1(n15111), .A2(n12204), .ZN(n6618) );
  AND2_X1 U8912 ( .A1(n7183), .A2(n11806), .ZN(n6619) );
  AND2_X1 U8913 ( .A1(n10375), .A2(n10373), .ZN(n6620) );
  NAND2_X1 U8914 ( .A1(n12367), .A2(n12366), .ZN(n6621) );
  NAND4_X1 U8915 ( .A1(n8233), .A2(n7058), .A3(n7059), .A4(n7060), .ZN(n7061)
         );
  OR2_X1 U8916 ( .A1(n12962), .A2(n12972), .ZN(n6622) );
  NOR2_X1 U8917 ( .A1(n12968), .A2(n7031), .ZN(n7030) );
  AND2_X1 U8918 ( .A1(n7761), .A2(n12582), .ZN(n6623) );
  OR2_X1 U8919 ( .A1(n13566), .A2(n13517), .ZN(n6624) );
  AND2_X1 U8920 ( .A1(n7429), .A2(n7431), .ZN(n6625) );
  INV_X1 U8921 ( .A(n12270), .ZN(n7322) );
  AND2_X1 U8922 ( .A1(n11250), .A2(n10442), .ZN(n6626) );
  INV_X1 U8923 ( .A(n12193), .ZN(n7309) );
  INV_X1 U8924 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6905) );
  OR2_X1 U8925 ( .A1(n11413), .A2(n13998), .ZN(n6627) );
  XOR2_X1 U8926 ( .A(n13741), .B(n12513), .Z(n6628) );
  INV_X1 U8927 ( .A(n11548), .ZN(n6974) );
  INV_X1 U8928 ( .A(n9585), .ZN(n9991) );
  OR2_X1 U8929 ( .A1(n11413), .A2(n14012), .ZN(n6629) );
  INV_X1 U8930 ( .A(n7426), .ZN(n7425) );
  NAND2_X1 U8931 ( .A1(n7427), .A2(n7431), .ZN(n7426) );
  OR2_X1 U8932 ( .A1(n13478), .A2(n13505), .ZN(n6630) );
  AOI21_X1 U8933 ( .B1(n8345), .B2(n7562), .A(n7561), .ZN(n8776) );
  NAND2_X1 U8934 ( .A1(n8759), .A2(n8758), .ZN(n13768) );
  INV_X1 U8935 ( .A(n13768), .ZN(n7045) );
  NAND2_X1 U8936 ( .A1(n7621), .A2(n7622), .ZN(n6631) );
  INV_X1 U8937 ( .A(n11631), .ZN(n6925) );
  XOR2_X1 U8938 ( .A(n14581), .B(n14580), .Z(n6632) );
  AND2_X1 U8939 ( .A1(n10028), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6633) );
  INV_X1 U8940 ( .A(n12007), .ZN(n7111) );
  MUX2_X1 U8941 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13821), .S(n8466), .Z(n15035)
         );
  NAND2_X1 U8942 ( .A1(n6777), .A2(n13936), .ZN(n13934) );
  OR3_X1 U8943 ( .A1(n12081), .A2(n12492), .A3(n12080), .ZN(n6634) );
  OR3_X1 U8944 ( .A1(n12145), .A2(n15035), .A3(n12225), .ZN(n6635) );
  INV_X1 U8945 ( .A(n14102), .ZN(n14095) );
  NAND2_X1 U8946 ( .A1(n12502), .A2(n12501), .ZN(n13298) );
  NAND2_X1 U8947 ( .A1(n13768), .A2(n13308), .ZN(n6636) );
  OR2_X1 U8948 ( .A1(n14515), .A2(n14514), .ZN(n6637) );
  AND2_X1 U8949 ( .A1(n7800), .A2(n7820), .ZN(n6638) );
  NAND2_X1 U8950 ( .A1(n12293), .A2(n12292), .ZN(n13706) );
  INV_X1 U8951 ( .A(n13706), .ZN(n7041) );
  AND2_X1 U8952 ( .A1(n6863), .A2(n12220), .ZN(n6639) );
  AND2_X1 U8953 ( .A1(n7430), .A2(n7429), .ZN(n6640) );
  AND2_X1 U8954 ( .A1(n14535), .A2(n6913), .ZN(n6641) );
  MUX2_X1 U8955 ( .A(n14140), .B(n14125), .S(n11504), .Z(n11486) );
  OR2_X1 U8956 ( .A1(n14573), .A2(n14572), .ZN(n6642) );
  AND2_X1 U8957 ( .A1(n12190), .A2(n12191), .ZN(n6643) );
  AOI21_X1 U8958 ( .B1(n7030), .B2(n12484), .A(n6607), .ZN(n7029) );
  NAND2_X1 U8959 ( .A1(n8602), .A2(n8601), .ZN(n15111) );
  INV_X1 U8960 ( .A(n15111), .ZN(n7050) );
  AND2_X1 U8961 ( .A1(n7029), .A2(n7025), .ZN(n6644) );
  NOR2_X1 U8962 ( .A1(n6583), .A2(n13323), .ZN(n6645) );
  AND2_X1 U8963 ( .A1(n8708), .A2(n8707), .ZN(n6646) );
  AND2_X1 U8964 ( .A1(n8552), .A2(n8551), .ZN(n6647) );
  AND2_X1 U8965 ( .A1(n6863), .A2(n12218), .ZN(n6648) );
  AND2_X1 U8966 ( .A1(n10253), .A2(n7264), .ZN(n6649) );
  NOR2_X1 U8967 ( .A1(n11622), .A2(n11621), .ZN(n6650) );
  INV_X1 U8968 ( .A(n11849), .ZN(n12122) );
  NOR2_X1 U8969 ( .A1(n14121), .A2(n14337), .ZN(n11849) );
  INV_X1 U8970 ( .A(n7042), .ZN(n13534) );
  INV_X1 U8971 ( .A(n11507), .ZN(n7251) );
  INV_X1 U8972 ( .A(n7515), .ZN(n7514) );
  NAND2_X1 U8973 ( .A1(n7516), .A2(n7983), .ZN(n7515) );
  NAND2_X1 U8974 ( .A1(n13638), .A2(n7053), .ZN(n7057) );
  OR2_X1 U8975 ( .A1(n7054), .A2(n13594), .ZN(n6651) );
  AND2_X1 U8976 ( .A1(n6852), .A2(n6643), .ZN(n6652) );
  AND2_X1 U8977 ( .A1(n8489), .A2(n8488), .ZN(n6653) );
  INV_X1 U8978 ( .A(n12484), .ZN(n7033) );
  AND2_X1 U8979 ( .A1(n6896), .A2(n8332), .ZN(n6654) );
  OR2_X1 U8980 ( .A1(n13608), .A2(n13516), .ZN(n6655) );
  INV_X1 U8981 ( .A(n14096), .ZN(n7352) );
  AND2_X1 U8982 ( .A1(n15111), .A2(n13315), .ZN(n6656) );
  NAND2_X1 U8983 ( .A1(n10372), .A2(n10371), .ZN(n6657) );
  INV_X1 U8984 ( .A(n7379), .ZN(n7377) );
  NOR2_X1 U8985 ( .A1(n13727), .A2(n13570), .ZN(n7379) );
  AND2_X1 U8986 ( .A1(n7045), .A2(n13308), .ZN(n6658) );
  OAI21_X1 U8987 ( .B1(n12148), .B2(n12331), .A(n7394), .ZN(n7337) );
  INV_X1 U8988 ( .A(n7584), .ZN(n7211) );
  NAND2_X1 U8989 ( .A1(n14586), .A2(n11100), .ZN(n6659) );
  AND2_X1 U8990 ( .A1(n13773), .A2(n12249), .ZN(n6660) );
  AND2_X1 U8991 ( .A1(n12272), .A2(n12273), .ZN(n6661) );
  AND2_X1 U8992 ( .A1(n13624), .A2(n13483), .ZN(n6662) );
  NAND2_X1 U8993 ( .A1(n8166), .A2(n8165), .ZN(n12495) );
  AND2_X1 U8994 ( .A1(n8742), .A2(n8741), .ZN(n12251) );
  INV_X1 U8995 ( .A(n12251), .ZN(n13773) );
  AND2_X1 U8996 ( .A1(n6934), .A2(n6935), .ZN(n6663) );
  OR2_X1 U8997 ( .A1(n12815), .A2(n12816), .ZN(n7296) );
  AND2_X1 U8998 ( .A1(n8092), .A2(n8091), .ZN(n6664) );
  NOR2_X1 U8999 ( .A1(n12271), .A2(n7322), .ZN(n6665) );
  NOR2_X1 U9000 ( .A1(n14388), .A2(n14237), .ZN(n6666) );
  NOR2_X1 U9001 ( .A1(n11770), .A2(n11769), .ZN(n6667) );
  NOR2_X1 U9002 ( .A1(n11103), .A2(n11102), .ZN(n6668) );
  AND2_X1 U9003 ( .A1(n7543), .A2(n12456), .ZN(n6669) );
  NOR2_X1 U9004 ( .A1(n12996), .A2(n7579), .ZN(n6670) );
  MUX2_X1 U9005 ( .A(n13972), .B(n14137), .S(n6799), .Z(n11467) );
  NAND2_X1 U9006 ( .A1(n14305), .A2(n7239), .ZN(n6671) );
  INV_X1 U9007 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8373) );
  INV_X1 U9008 ( .A(n12920), .ZN(n12918) );
  AND2_X1 U9009 ( .A1(n13747), .A2(n13480), .ZN(n6672) );
  OR2_X1 U9010 ( .A1(n8081), .A2(n6778), .ZN(n6673) );
  AND2_X1 U9011 ( .A1(n8072), .A2(n7036), .ZN(n6674) );
  OR2_X1 U9012 ( .A1(n12091), .A2(n11910), .ZN(n6675) );
  INV_X1 U9013 ( .A(n6742), .ZN(n8249) );
  INV_X1 U9014 ( .A(n7349), .ZN(n7348) );
  NAND2_X1 U9015 ( .A1(n7569), .A2(n7350), .ZN(n7349) );
  NOR2_X1 U9016 ( .A1(n12262), .A2(n12261), .ZN(n6676) );
  NOR2_X1 U9017 ( .A1(n11764), .A2(n11763), .ZN(n6677) );
  NAND2_X1 U9018 ( .A1(n7074), .A2(n12307), .ZN(n13712) );
  AND2_X1 U9019 ( .A1(n7348), .A2(n7352), .ZN(n6678) );
  NAND2_X1 U9020 ( .A1(n7660), .A2(n7299), .ZN(n7663) );
  OR2_X1 U9021 ( .A1(n6817), .A2(n7521), .ZN(n6679) );
  INV_X1 U9022 ( .A(n11859), .ZN(n7202) );
  INV_X1 U9023 ( .A(n7404), .ZN(n7403) );
  NAND2_X1 U9024 ( .A1(n7406), .A2(n7407), .ZN(n7404) );
  AND2_X1 U9025 ( .A1(n6862), .A2(n6867), .ZN(n6680) );
  NOR2_X1 U9026 ( .A1(n14397), .A2(n11807), .ZN(n6681) );
  INV_X1 U9027 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7434) );
  AND2_X1 U9028 ( .A1(n8000), .A2(n12742), .ZN(n6682) );
  AND2_X1 U9029 ( .A1(n7099), .A2(n12051), .ZN(n6683) );
  INV_X1 U9030 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8925) );
  AND2_X1 U9031 ( .A1(n11734), .A2(n11735), .ZN(n6684) );
  INV_X1 U9032 ( .A(n7361), .ZN(n7360) );
  NAND2_X1 U9033 ( .A1(n6879), .A2(n6878), .ZN(n7361) );
  OAI21_X1 U9034 ( .B1(n7401), .B2(n7400), .A(n7405), .ZN(n7398) );
  AND2_X1 U9035 ( .A1(n13478), .A2(n13477), .ZN(n6685) );
  NOR2_X1 U9036 ( .A1(n14174), .A2(n14183), .ZN(n6686) );
  AND2_X1 U9037 ( .A1(n13712), .A2(n13543), .ZN(n6687) );
  INV_X1 U9038 ( .A(n7370), .ZN(n7369) );
  OR2_X1 U9039 ( .A1(n14186), .A2(n7371), .ZN(n7370) );
  AND2_X1 U9040 ( .A1(n7582), .A2(n6621), .ZN(n6688) );
  OR2_X1 U9041 ( .A1(n7221), .A2(n14094), .ZN(n6689) );
  NAND2_X1 U9042 ( .A1(n9106), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U9043 ( .A1(n10522), .A2(n6618), .ZN(n6691) );
  NAND2_X1 U9044 ( .A1(n8341), .A2(n7539), .ZN(n6692) );
  INV_X1 U9045 ( .A(n11279), .ZN(n7240) );
  OR2_X1 U9046 ( .A1(n14504), .A2(n14503), .ZN(n6693) );
  AND2_X1 U9047 ( .A1(n7368), .A2(n11840), .ZN(n6694) );
  INV_X1 U9048 ( .A(n13727), .ZN(n7054) );
  AND2_X1 U9049 ( .A1(n7718), .A2(n7577), .ZN(n6695) );
  AND2_X1 U9050 ( .A1(n7527), .A2(n9230), .ZN(n6696) );
  AND2_X1 U9051 ( .A1(n6855), .A2(n6854), .ZN(n6697) );
  OR2_X1 U9052 ( .A1(n12234), .A2(n13311), .ZN(n6698) );
  NAND2_X1 U9053 ( .A1(n11121), .A2(n12745), .ZN(n6699) );
  NOR2_X1 U9054 ( .A1(n14130), .A2(n7584), .ZN(n6700) );
  NOR2_X1 U9055 ( .A1(n7508), .A2(n13852), .ZN(n7507) );
  OR2_X1 U9056 ( .A1(n12946), .A2(n12951), .ZN(n6701) );
  AND2_X1 U9057 ( .A1(n8233), .A2(n8921), .ZN(n6702) );
  NAND4_X1 U9058 ( .A1(n8371), .A2(n8370), .A3(n8373), .A4(n8265), .ZN(n8271)
         );
  AND2_X1 U9059 ( .A1(n11364), .A2(n11363), .ZN(n6703) );
  INV_X1 U9060 ( .A(n10327), .ZN(n7010) );
  AND2_X1 U9061 ( .A1(n11855), .A2(n11854), .ZN(n6704) );
  AND2_X1 U9062 ( .A1(n8064), .A2(n8072), .ZN(n6705) );
  NOR2_X1 U9063 ( .A1(n12223), .A2(n12224), .ZN(n6868) );
  AND2_X1 U9064 ( .A1(n8734), .A2(n7449), .ZN(n6706) );
  INV_X1 U9065 ( .A(n11825), .ZN(n7184) );
  OR2_X1 U9066 ( .A1(n11270), .A2(n11268), .ZN(n6707) );
  OR2_X1 U9067 ( .A1(n11241), .A2(n11239), .ZN(n6708) );
  AND2_X1 U9068 ( .A1(n12503), .A2(n12501), .ZN(n6709) );
  INV_X1 U9069 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8192) );
  AND2_X1 U9070 ( .A1(n7247), .A2(n8964), .ZN(n6710) );
  NAND2_X1 U9071 ( .A1(n12442), .A2(n12445), .ZN(n6711) );
  NAND2_X1 U9072 ( .A1(n12269), .A2(n6847), .ZN(n6712) );
  INV_X1 U9073 ( .A(n14099), .ZN(n7221) );
  AND2_X1 U9074 ( .A1(n7610), .A2(n7120), .ZN(n6713) );
  OR2_X1 U9075 ( .A1(n7308), .A2(n12210), .ZN(n6714) );
  INV_X1 U9076 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9245) );
  AND2_X1 U9077 ( .A1(n11230), .A2(n7224), .ZN(n6715) );
  AND2_X1 U9078 ( .A1(n7292), .A2(n12420), .ZN(n7289) );
  OR2_X1 U9079 ( .A1(n7413), .A2(n6617), .ZN(n6716) );
  INV_X1 U9080 ( .A(n7485), .ZN(n7484) );
  OR2_X1 U9081 ( .A1(n12213), .A2(n12214), .ZN(n6717) );
  INV_X1 U9082 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9657) );
  OR2_X1 U9083 ( .A1(n7274), .A2(n13520), .ZN(n6718) );
  INV_X1 U9084 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9331) );
  INV_X1 U9085 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9312) );
  AND2_X1 U9086 ( .A1(n10154), .A2(n11595), .ZN(n7355) );
  NOR2_X2 U9087 ( .A1(n12137), .A2(n8881), .ZN(n12225) );
  INV_X1 U9088 ( .A(n14279), .ZN(n6871) );
  NAND2_X1 U9089 ( .A1(n10933), .A2(n10932), .ZN(n10931) );
  INV_X1 U9090 ( .A(n13031), .ZN(n6800) );
  NAND2_X1 U9091 ( .A1(n8061), .A2(n8060), .ZN(n12483) );
  INV_X1 U9092 ( .A(n12483), .ZN(n7037) );
  XNOR2_X1 U9093 ( .A(n13778), .B(n12239), .ZN(n12425) );
  INV_X1 U9094 ( .A(n12425), .ZN(n7400) );
  AND2_X1 U9095 ( .A1(n14282), .A2(n6967), .ZN(n6719) );
  INV_X1 U9096 ( .A(n10052), .ZN(n10029) );
  AND2_X1 U9097 ( .A1(n6612), .A2(n14282), .ZN(n6720) );
  INV_X1 U9098 ( .A(n10233), .ZN(n10554) );
  AND2_X1 U9099 ( .A1(n6916), .A2(n6919), .ZN(n6721) );
  NAND2_X1 U9100 ( .A1(n14288), .A2(n11825), .ZN(n14265) );
  INV_X1 U9101 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7120) );
  INV_X1 U9102 ( .A(n8327), .ZN(n6969) );
  INV_X1 U9103 ( .A(n12022), .ZN(n7107) );
  AND2_X1 U9104 ( .A1(n8800), .A2(n8799), .ZN(n6722) );
  AND4_X1 U9105 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n14931)
         );
  INV_X1 U9106 ( .A(n14931), .ZN(n7408) );
  AND4_X1 U9107 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(n12233)
         );
  AND3_X1 U9108 ( .A1(n8233), .A2(n8921), .A3(n8232), .ZN(n8235) );
  INV_X1 U9109 ( .A(n8235), .ZN(n9939) );
  INV_X1 U9110 ( .A(n12252), .ZN(n7318) );
  NAND2_X1 U9111 ( .A1(n7044), .A2(n13478), .ZN(n13691) );
  INV_X1 U9112 ( .A(n13691), .ZN(n7043) );
  INV_X1 U9113 ( .A(n13313), .ZN(n14934) );
  OR3_X1 U9114 ( .A1(n8645), .A2(n8644), .A3(n8643), .ZN(n13313) );
  INV_X1 U9115 ( .A(n13543), .ZN(n13519) );
  OR3_X1 U9116 ( .A1(n12313), .A2(n12312), .A3(n12311), .ZN(n13543) );
  OR2_X1 U9117 ( .A1(n12763), .A2(n10558), .ZN(n6723) );
  NOR2_X1 U9118 ( .A1(n6590), .A2(n15465), .ZN(n6724) );
  AND2_X1 U9119 ( .A1(n6996), .A2(n6995), .ZN(n6725) );
  OR2_X1 U9120 ( .A1(n6817), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n6726) );
  AND2_X1 U9121 ( .A1(n8348), .A2(n9507), .ZN(n6727) );
  AND2_X1 U9122 ( .A1(n10225), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6728) );
  AND2_X1 U9123 ( .A1(n7263), .A2(n6618), .ZN(n6729) );
  AND2_X1 U9124 ( .A1(n11708), .A2(n11707), .ZN(n6730) );
  INV_X1 U9125 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9451) );
  INV_X1 U9126 ( .A(SI_10_), .ZN(n7544) );
  AND2_X1 U9127 ( .A1(n9709), .A2(n10113), .ZN(n6731) );
  INV_X1 U9128 ( .A(n10992), .ZN(n7323) );
  INV_X1 U9129 ( .A(n14397), .ZN(n7062) );
  NAND2_X1 U9130 ( .A1(n10881), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7324) );
  NAND2_X1 U9131 ( .A1(n9659), .A2(n9658), .ZN(n14762) );
  NAND2_X1 U9132 ( .A1(n7178), .A2(n10437), .ZN(n10604) );
  NAND2_X1 U9133 ( .A1(n7190), .A2(n9674), .ZN(n10112) );
  OR2_X1 U9134 ( .A1(n8786), .A2(n8785), .ZN(n6732) );
  XNOR2_X1 U9135 ( .A(n7631), .B(n7630), .ZN(n8176) );
  NAND2_X1 U9136 ( .A1(n7462), .A2(n8571), .ZN(n9942) );
  NAND2_X1 U9137 ( .A1(n6921), .A2(n8274), .ZN(n6733) );
  OR2_X1 U9138 ( .A1(n7235), .A2(n7232), .ZN(n9626) );
  AND2_X1 U9139 ( .A1(n7490), .A2(n7491), .ZN(n9887) );
  OR2_X1 U9140 ( .A1(n11478), .A2(SI_26_), .ZN(n6734) );
  AND2_X1 U9141 ( .A1(n6601), .A2(n9709), .ZN(n6735) );
  INV_X1 U9142 ( .A(n14939), .ZN(n7445) );
  XNOR2_X1 U9143 ( .A(n8362), .B(n8361), .ZN(n9010) );
  NAND2_X1 U9144 ( .A1(n9244), .A2(n11192), .ZN(n9338) );
  AND2_X2 U9145 ( .A1(n10348), .A2(n9853), .ZN(n15235) );
  NAND2_X1 U9146 ( .A1(n8202), .A2(n8201), .ZN(n12724) );
  NAND2_X1 U9147 ( .A1(n10209), .A2(n12076), .ZN(n15193) );
  OR2_X1 U9148 ( .A1(n10209), .A2(n12087), .ZN(n15195) );
  INV_X1 U9149 ( .A(n9555), .ZN(n12884) );
  NAND4_X2 U9150 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n13322)
         );
  INV_X1 U9151 ( .A(n13322), .ZN(n6787) );
  AND2_X1 U9152 ( .A1(n8091), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6736) );
  INV_X1 U9153 ( .A(n14891), .ZN(n7064) );
  INV_X1 U9154 ( .A(n7681), .ZN(n7851) );
  NAND2_X1 U9155 ( .A1(n9111), .A2(n9112), .ZN(n9110) );
  INV_X1 U9156 ( .A(n9650), .ZN(n7338) );
  INV_X1 U9157 ( .A(n10207), .ZN(n7011) );
  INV_X1 U9158 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7160) );
  AND2_X1 U9159 ( .A1(n12135), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U9160 ( .A1(n12818), .A2(n12817), .ZN(n6738) );
  AND2_X2 U9161 ( .A1(n12107), .A2(n11943), .ZN(n12076) );
  NAND2_X1 U9162 ( .A1(n11885), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6739) );
  INV_X1 U9163 ( .A(n12102), .ZN(n7138) );
  INV_X1 U9164 ( .A(n12456), .ZN(n7541) );
  INV_X1 U9165 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14441) );
  INV_X1 U9166 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14442) );
  INV_X1 U9167 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6900) );
  INV_X1 U9168 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6765) );
  AND2_X1 U9169 ( .A1(n11550), .A2(P3_U3151), .ZN(n9400) );
  INV_X1 U9170 ( .A(n10673), .ZN(n10675) );
  OAI21_X2 U9171 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10369) );
  INV_X1 U9172 ( .A(n11745), .ZN(n11758) );
  NAND2_X2 U9173 ( .A1(n11574), .A2(n9251), .ZN(n11745) );
  NAND3_X1 U9174 ( .A1(n6741), .A2(n11277), .A3(n6740), .ZN(n7237) );
  NAND2_X1 U9175 ( .A1(n11272), .A2(n11271), .ZN(n6741) );
  OAI22_X2 U9176 ( .A1(n11523), .A2(n7255), .B1(n11524), .B2(n7254), .ZN(
        n11529) );
  NAND3_X1 U9177 ( .A1(n6702), .A2(n7060), .A3(n7059), .ZN(n6742) );
  NAND3_X1 U9178 ( .A1(n7229), .A2(n7227), .A3(n11588), .ZN(n7226) );
  OR2_X1 U9179 ( .A1(n11448), .A2(n11449), .ZN(n11450) );
  INV_X1 U9180 ( .A(n11229), .ZN(n6796) );
  NAND2_X1 U9181 ( .A1(n6792), .A2(n6791), .ZN(n11273) );
  NAND2_X1 U9182 ( .A1(n6794), .A2(n6793), .ZN(n11244) );
  NAND2_X1 U9183 ( .A1(n11582), .A2(n6745), .ZN(n6744) );
  NOR2_X1 U9184 ( .A1(n11623), .A2(n6743), .ZN(n11628) );
  NAND2_X1 U9185 ( .A1(n11584), .A2(n11504), .ZN(n6966) );
  NAND2_X1 U9186 ( .A1(n11530), .A2(n11531), .ZN(n6976) );
  OAI21_X2 U9187 ( .B1(n7863), .B2(n7862), .A(n7861), .ZN(n7864) );
  OR2_X1 U9188 ( .A1(n13090), .A2(n13112), .ZN(n6808) );
  NAND2_X1 U9189 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  AOI21_X2 U9190 ( .B1(n12491), .B2(n11878), .A(n11877), .ZN(n12537) );
  NAND2_X1 U9191 ( .A1(n7134), .A2(n7920), .ZN(n7941) );
  NAND2_X1 U9192 ( .A1(n7966), .A2(n7965), .ZN(n7986) );
  NAND2_X1 U9193 ( .A1(n7161), .A2(n8021), .ZN(n8035) );
  NAND2_X1 U9194 ( .A1(n6802), .A2(n6801), .ZN(n8004) );
  OAI21_X1 U9195 ( .B1(n7671), .B2(n7576), .A(n7672), .ZN(n7691) );
  NAND2_X1 U9196 ( .A1(n12958), .A2(n12060), .ZN(n12943) );
  NAND2_X1 U9197 ( .A1(n14607), .A2(n11939), .ZN(n14595) );
  NAND2_X1 U9198 ( .A1(n12965), .A2(n12968), .ZN(n12967) );
  NAND2_X1 U9199 ( .A1(n10651), .A2(n11971), .ZN(n10635) );
  NAND2_X1 U9200 ( .A1(n10634), .A2(n11964), .ZN(n10652) );
  NAND2_X1 U9201 ( .A1(n11867), .A2(n12024), .ZN(n13067) );
  NAND2_X1 U9202 ( .A1(n6754), .A2(n11938), .ZN(n14609) );
  NAND2_X1 U9203 ( .A1(n15165), .A2(n11955), .ZN(n10200) );
  OAI21_X2 U9204 ( .B1(n13023), .B2(n7101), .A(n6683), .ZN(n12988) );
  NAND3_X1 U9205 ( .A1(n6751), .A2(n12461), .A3(n6749), .ZN(P2_U3328) );
  NAND2_X2 U9206 ( .A1(n8008), .A2(n8007), .ZN(n13193) );
  NAND2_X1 U9207 ( .A1(n10325), .A2(n11969), .ZN(n10634) );
  NAND2_X1 U9208 ( .A1(n15167), .A2(n15166), .ZN(n15165) );
  NAND2_X1 U9209 ( .A1(n11120), .A2(n11119), .ZN(n6754) );
  NAND2_X1 U9210 ( .A1(n7557), .A2(n7556), .ZN(n8349) );
  XNOR2_X1 U9211 ( .A(n6755), .B(n12436), .ZN(n12435) );
  NAND4_X1 U9212 ( .A1(n7583), .A2(n12434), .A3(n12433), .A4(n13520), .ZN(
        n6755) );
  NAND2_X1 U9213 ( .A1(n12937), .A2(n12942), .ZN(n12936) );
  NAND2_X1 U9214 ( .A1(n7026), .A2(n6771), .ZN(n12953) );
  NOR2_X1 U9215 ( .A1(n12906), .A2(n12907), .ZN(n12905) );
  NAND2_X1 U9216 ( .A1(n12453), .A2(n6711), .ZN(n7542) );
  NAND2_X1 U9217 ( .A1(n9632), .A2(n11950), .ZN(n10198) );
  NAND3_X1 U9218 ( .A1(n6670), .A2(n6598), .A3(n7018), .ZN(n12480) );
  NAND2_X2 U9219 ( .A1(n13568), .A2(n13569), .ZN(n13567) );
  NAND2_X1 U9220 ( .A1(n7286), .A2(n7287), .ZN(n11072) );
  AOI21_X2 U9221 ( .B1(n13614), .B2(n13484), .A(n6662), .ZN(n13592) );
  OAI21_X1 U9222 ( .B1(n12617), .B2(n12619), .A(n12618), .ZN(n12616) );
  OAI21_X2 U9223 ( .B1(n12640), .B2(n7512), .A(n7510), .ZN(n12587) );
  NAND2_X1 U9224 ( .A1(n6759), .A2(n6757), .ZN(P3_U3154) );
  NAND2_X1 U9225 ( .A1(n12554), .A2(n12724), .ZN(n6759) );
  XNOR2_X1 U9226 ( .A(n12802), .B(n12801), .ZN(n12793) );
  NOR2_X1 U9227 ( .A1(n12791), .A2(n12790), .ZN(n12802) );
  NAND2_X1 U9228 ( .A1(n7084), .A2(n11868), .ZN(n13135) );
  AND2_X2 U9229 ( .A1(n11955), .A2(n11953), .ZN(n15166) );
  NAND2_X1 U9230 ( .A1(n15173), .A2(n12752), .ZN(n11953) );
  NAND2_X1 U9231 ( .A1(n13065), .A2(n12023), .ZN(n13055) );
  NAND2_X1 U9232 ( .A1(n13033), .A2(n6800), .ZN(n13032) );
  OR2_X2 U9233 ( .A1(n7632), .A2(n7118), .ZN(n7598) );
  NAND2_X1 U9234 ( .A1(n10198), .A2(n11949), .ZN(n15167) );
  NOR2_X2 U9235 ( .A1(n14101), .A2(n14113), .ZN(n14100) );
  NOR2_X2 U9236 ( .A1(n14374), .A2(n14214), .ZN(n14213) );
  NAND2_X1 U9237 ( .A1(n11550), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U9238 ( .A1(n11684), .A2(n11683), .ZN(n11689) );
  NAND2_X1 U9239 ( .A1(n11779), .A2(n11778), .ZN(n13822) );
  NAND2_X1 U9240 ( .A1(n13898), .A2(n13899), .ZN(n13897) );
  AOI22_X1 U9241 ( .A1(n13822), .A2(n13823), .B1(n11785), .B2(n11784), .ZN(
        n11794) );
  NAND2_X1 U9242 ( .A1(n8460), .A2(n8461), .ZN(n8474) );
  AND2_X2 U9243 ( .A1(n6788), .A2(n8473), .ZN(n8460) );
  NOR2_X1 U9244 ( .A1(n13919), .A2(n6818), .ZN(n13857) );
  NAND2_X1 U9245 ( .A1(n7489), .A2(n9884), .ZN(n9922) );
  NAND2_X1 U9246 ( .A1(n10709), .A2(n11979), .ZN(n11114) );
  INV_X2 U9247 ( .A(n12752), .ZN(n15192) );
  XNOR2_X1 U9248 ( .A(n11775), .B(n11776), .ZN(n13947) );
  NOR2_X1 U9249 ( .A1(n9302), .A2(n9301), .ZN(n9300) );
  XNOR2_X1 U9250 ( .A(n9297), .B(n11692), .ZN(n9302) );
  NAND2_X1 U9251 ( .A1(n12936), .A2(n6701), .ZN(n12921) );
  NAND2_X1 U9252 ( .A1(n10701), .A2(n10700), .ZN(n10702) );
  NAND2_X1 U9253 ( .A1(n7034), .A2(n7029), .ZN(n6771) );
  INV_X1 U9254 ( .A(n10642), .ZN(n7000) );
  INV_X1 U9255 ( .A(n7008), .ZN(n7007) );
  NAND2_X1 U9256 ( .A1(n10640), .A2(n10639), .ZN(n10653) );
  AOI21_X1 U9257 ( .B1(n11130), .B2(n11129), .A(n11105), .ZN(n11106) );
  NOR2_X1 U9258 ( .A1(n12769), .A2(n10542), .ZN(n10544) );
  OAI21_X1 U9259 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10043) );
  NOR3_X1 U9260 ( .A1(n10998), .A2(n10997), .A3(n10999), .ZN(n12791) );
  NOR2_X2 U9261 ( .A1(n12759), .A2(n6767), .ZN(n10548) );
  NAND2_X1 U9262 ( .A1(n9965), .A2(n9569), .ZN(n9570) );
  NAND2_X1 U9263 ( .A1(n7295), .A2(n9581), .ZN(n7294) );
  NOR2_X1 U9264 ( .A1(n12827), .A2(n12828), .ZN(n12850) );
  NOR2_X1 U9265 ( .A1(n10882), .A2(n10883), .ZN(n10979) );
  NAND2_X1 U9266 ( .A1(n7651), .A2(n15168), .ZN(n7654) );
  AOI21_X2 U9267 ( .B1(n7036), .B2(n8064), .A(n6782), .ZN(n8084) );
  OAI21_X1 U9268 ( .B1(n7959), .B2(n7962), .A(n7961), .ZN(n7963) );
  NAND2_X1 U9269 ( .A1(n12606), .A2(n8055), .ZN(n8063) );
  NAND2_X1 U9270 ( .A1(n12670), .A2(n7837), .ZN(n12567) );
  NAND2_X1 U9271 ( .A1(n7525), .A2(n6638), .ZN(n12670) );
  INV_X1 U9272 ( .A(n10201), .ZN(n9633) );
  NAND2_X1 U9273 ( .A1(n7481), .A2(n7482), .ZN(n7959) );
  INV_X1 U9274 ( .A(n6769), .ZN(n11066) );
  NAND2_X1 U9275 ( .A1(n9637), .A2(n7653), .ZN(n9631) );
  NAND2_X1 U9276 ( .A1(n8004), .A2(n8003), .ZN(n8020) );
  INV_X1 U9277 ( .A(n8081), .ZN(n6774) );
  NAND2_X1 U9278 ( .A1(n7005), .A2(n7004), .ZN(n12906) );
  OAI21_X1 U9279 ( .B1(n8040), .B2(n7148), .A(n7146), .ZN(n8078) );
  AND2_X2 U9280 ( .A1(n6772), .A2(n11872), .ZN(n12968) );
  NAND2_X1 U9281 ( .A1(n12921), .A2(n7006), .ZN(n7005) );
  AOI21_X2 U9282 ( .B1(n10489), .B2(n11897), .A(n6724), .ZN(n13111) );
  INV_X1 U9283 ( .A(n12700), .ZN(n7516) );
  INV_X1 U9284 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7002) );
  AOI21_X1 U9285 ( .B1(n7634), .B2(n8176), .A(n10941), .ZN(n8174) );
  NAND2_X1 U9286 ( .A1(n9304), .A2(n6775), .ZN(n9383) );
  INV_X1 U9287 ( .A(n9303), .ZN(n6776) );
  NAND2_X1 U9288 ( .A1(n9357), .A2(n9356), .ZN(n9881) );
  NAND2_X1 U9289 ( .A1(n13897), .A2(n13901), .ZN(n13935) );
  NAND2_X1 U9290 ( .A1(n6938), .A2(n6940), .ZN(n8733) );
  XNOR2_X2 U9291 ( .A(n8852), .B(n8850), .ZN(n13236) );
  AND2_X1 U9292 ( .A1(n9392), .A2(n9321), .ZN(n9357) );
  OAI21_X1 U9293 ( .B1(n8391), .B2(n12388), .A(n13459), .ZN(n9126) );
  NAND2_X1 U9294 ( .A1(n6955), .A2(n6953), .ZN(n13252) );
  INV_X1 U9295 ( .A(n11590), .ZN(n9689) );
  NAND2_X1 U9296 ( .A1(n7366), .A2(n7365), .ZN(n14149) );
  NOR2_X2 U9297 ( .A1(n11810), .A2(n11832), .ZN(n11839) );
  INV_X1 U9298 ( .A(n7216), .ZN(n7215) );
  INV_X1 U9299 ( .A(n8537), .ZN(n6949) );
  INV_X1 U9300 ( .A(n7214), .ZN(n7213) );
  NAND2_X1 U9301 ( .A1(n7354), .A2(n7353), .ZN(n10469) );
  NAND3_X1 U9302 ( .A1(n6945), .A2(n9482), .A3(n6943), .ZN(n7462) );
  INV_X1 U9303 ( .A(n7340), .ZN(n12116) );
  OAI21_X1 U9304 ( .B1(n12093), .B2(n12094), .A(n12095), .ZN(n12096) );
  NAND2_X1 U9305 ( .A1(n6807), .A2(n7905), .ZN(n7889) );
  NAND4_X1 U9306 ( .A1(n12068), .A2(n12918), .A3(n12066), .A4(n12067), .ZN(
        n12072) );
  AOI21_X1 U9307 ( .B1(n12085), .B2(n6780), .A(n12091), .ZN(n6804) );
  NOR2_X1 U9308 ( .A1(n12086), .A2(n12076), .ZN(n6780) );
  OR2_X1 U9309 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  INV_X1 U9310 ( .A(n8002), .ZN(n6802) );
  NOR2_X1 U9311 ( .A1(n12082), .A2(n12083), .ZN(n6806) );
  NAND2_X1 U9312 ( .A1(n11821), .A2(n11820), .ZN(n14304) );
  NAND2_X1 U9313 ( .A1(n7194), .A2(n7193), .ZN(n11834) );
  NAND2_X1 U9314 ( .A1(n8034), .A2(n7524), .ZN(n12606) );
  INV_X2 U9315 ( .A(n7680), .ZN(n7717) );
  NAND2_X1 U9316 ( .A1(n7964), .A2(n7963), .ZN(n12640) );
  OAI21_X1 U9317 ( .B1(n11628), .B2(n11627), .A(n6783), .ZN(P1_U3242) );
  NAND2_X1 U9318 ( .A1(n8652), .A2(n8651), .ZN(n8328) );
  NAND2_X1 U9319 ( .A1(n8594), .A2(n8593), .ZN(n8596) );
  OAI21_X1 U9320 ( .B1(n11550), .B2(n9249), .A(n6784), .ZN(n8289) );
  INV_X1 U9321 ( .A(n11434), .ZN(n7245) );
  NAND2_X1 U9322 ( .A1(n6979), .A2(n6978), .ZN(n6977) );
  NAND2_X1 U9323 ( .A1(n9315), .A2(n9316), .ZN(n9317) );
  NAND2_X1 U9324 ( .A1(n7472), .A2(n7471), .ZN(n13946) );
  NAND3_X1 U9325 ( .A1(n7488), .A2(n9305), .A3(n9383), .ZN(n9384) );
  NAND2_X1 U9326 ( .A1(n9293), .A2(n7247), .ZN(n6789) );
  AND2_X4 U9327 ( .A1(n11195), .A2(n11190), .ZN(n11692) );
  NAND2_X1 U9328 ( .A1(n10403), .A2(n10402), .ZN(n10407) );
  XNOR2_X2 U9329 ( .A(n7611), .B(n7610), .ZN(n9555) );
  OAI21_X2 U9330 ( .B1(n7632), .B2(P3_IR_REG_26__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7611) );
  OR2_X2 U9331 ( .A1(n12943), .A2(n7090), .ZN(n7087) );
  NAND2_X1 U9332 ( .A1(n10652), .A2(n11966), .ZN(n10651) );
  NAND2_X1 U9333 ( .A1(n6811), .A2(n6605), .ZN(n13785) );
  CLKBUF_X1 U9334 ( .A(n9907), .Z(n12400) );
  OAI211_X2 U9335 ( .C1(n8466), .C2(n14954), .A(n8464), .B(n8465), .ZN(n15062)
         );
  OR2_X1 U9336 ( .A1(n10365), .A2(n10366), .ZN(n10370) );
  OR2_X1 U9337 ( .A1(n8292), .A2(SI_2_), .ZN(n6788) );
  NAND2_X1 U9338 ( .A1(n8292), .A2(SI_2_), .ZN(n8473) );
  AOI22_X1 U9339 ( .A1(n11771), .A2(n14831), .B1(n9361), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U9340 ( .A1(n7519), .A2(n11708), .ZN(n13887) );
  NAND3_X1 U9341 ( .A1(n9922), .A2(n7491), .A3(n9888), .ZN(n9923) );
  NAND2_X1 U9342 ( .A1(n12967), .A2(n12062), .ZN(n12958) );
  OR2_X1 U9343 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U9344 ( .A1(n8289), .A2(SI_0_), .ZN(n8420) );
  NAND2_X2 U9345 ( .A1(n9685), .A2(n9684), .ZN(n14875) );
  AND2_X1 U9346 ( .A1(n6973), .A2(n6972), .ZN(n11582) );
  NAND3_X1 U9347 ( .A1(n6873), .A2(n6874), .A3(n7533), .ZN(n8594) );
  NAND2_X1 U9348 ( .A1(n6977), .A2(n6976), .ZN(n6975) );
  NAND2_X1 U9349 ( .A1(n8802), .A2(n8352), .ZN(n8806) );
  NAND2_X1 U9350 ( .A1(n11529), .A2(n11528), .ZN(n6979) );
  NAND3_X1 U9351 ( .A1(n6981), .A2(n6980), .A3(n7251), .ZN(n11508) );
  INV_X1 U9352 ( .A(n9300), .ZN(n7488) );
  OAI21_X1 U9353 ( .B1(n6975), .B2(n6974), .A(n11549), .ZN(n6973) );
  OR2_X1 U9354 ( .A1(n10306), .A2(n11675), .ZN(n11191) );
  NAND3_X1 U9355 ( .A1(n11267), .A2(n11266), .A3(n6707), .ZN(n6792) );
  NAND3_X1 U9356 ( .A1(n11236), .A2(n11237), .A3(n6708), .ZN(n6794) );
  AOI21_X1 U9357 ( .B1(n6796), .B2(n6795), .A(n11233), .ZN(n11234) );
  NAND2_X1 U9358 ( .A1(n6798), .A2(n6797), .ZN(n11205) );
  NAND2_X1 U9359 ( .A1(n11431), .A2(n11202), .ZN(n6797) );
  NAND2_X1 U9360 ( .A1(n12988), .A2(n12054), .ZN(n11870) );
  AOI21_X2 U9361 ( .B1(n10857), .B2(n10856), .A(n10855), .ZN(n10901) );
  NAND2_X1 U9362 ( .A1(n9779), .A2(n9509), .ZN(n9907) );
  NAND2_X1 U9363 ( .A1(n9513), .A2(n12405), .ZN(n9816) );
  NAND2_X1 U9364 ( .A1(n13476), .A2(n7285), .ZN(n7284) );
  INV_X1 U9365 ( .A(n11072), .ZN(n6812) );
  OAI21_X1 U9366 ( .B1(n13681), .B2(n7283), .A(n7282), .ZN(n7281) );
  NAND2_X1 U9367 ( .A1(n13542), .A2(n7568), .ZN(n13547) );
  INV_X1 U9368 ( .A(n7889), .ZN(n7135) );
  NAND2_X1 U9369 ( .A1(n6803), .A2(n12090), .ZN(n12094) );
  NAND2_X1 U9370 ( .A1(n6805), .A2(n6804), .ZN(n6803) );
  NAND2_X1 U9371 ( .A1(n12088), .A2(n12076), .ZN(n6805) );
  NAND2_X1 U9372 ( .A1(n6634), .A2(n6806), .ZN(n12085) );
  NAND2_X1 U9373 ( .A1(n7136), .A2(n7658), .ZN(n7671) );
  NAND2_X1 U9374 ( .A1(n7906), .A2(n7905), .ZN(n7919) );
  INV_X1 U9375 ( .A(n7691), .ZN(n7692) );
  NAND2_X1 U9376 ( .A1(n7152), .A2(n7151), .ZN(n7721) );
  NAND3_X1 U9377 ( .A1(n13089), .A2(n13088), .A3(n6808), .ZN(n13168) );
  INV_X1 U9378 ( .A(n7029), .ZN(n7028) );
  NAND2_X1 U9379 ( .A1(n7919), .A2(n7918), .ZN(n7134) );
  NAND2_X1 U9380 ( .A1(n7135), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U9381 ( .A1(n7164), .A2(n7168), .ZN(n7863) );
  INV_X1 U9382 ( .A(n7027), .ZN(n7026) );
  NAND2_X1 U9383 ( .A1(n6828), .A2(n6698), .ZN(n10903) );
  INV_X1 U9384 ( .A(n7281), .ZN(n13663) );
  NAND2_X1 U9385 ( .A1(n13542), .A2(n7570), .ZN(n13525) );
  OAI21_X2 U9386 ( .B1(n9842), .B2(n12100), .A(n7649), .ZN(n7680) );
  AOI21_X1 U9387 ( .B1(n7106), .B2(n7109), .A(n7105), .ZN(n7104) );
  NAND2_X1 U9388 ( .A1(n7727), .A2(n7590), .ZN(n7870) );
  NOR2_X1 U9389 ( .A1(n7843), .A2(n8939), .ZN(n7016) );
  AND2_X1 U9390 ( .A1(n7139), .A2(n7137), .ZN(n12103) );
  NAND2_X2 U9391 ( .A1(n14595), .A2(n14594), .ZN(n11122) );
  NAND2_X1 U9392 ( .A1(n7085), .A2(n12033), .ZN(n13049) );
  OAI21_X1 U9393 ( .B1(n13169), .B2(n15233), .A(n6819), .ZN(n13093) );
  OAI21_X1 U9394 ( .B1(n12099), .B2(n12098), .A(n7138), .ZN(n7137) );
  INV_X1 U9395 ( .A(n6821), .ZN(P3_U3455) );
  AOI21_X1 U9396 ( .B1(n13169), .B2(n15225), .A(n6822), .ZN(n6821) );
  INV_X1 U9397 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n6823) );
  AOI211_X2 U9398 ( .C1(n13683), .C2(n13602), .A(n13601), .B(n13600), .ZN(
        n13734) );
  NAND2_X1 U9399 ( .A1(n7420), .A2(n7419), .ZN(n10794) );
  OAI21_X1 U9400 ( .B1(n10066), .B2(n10253), .A(n7395), .ZN(n10259) );
  INV_X1 U9401 ( .A(n7409), .ZN(n13661) );
  NAND2_X1 U9402 ( .A1(n7277), .A2(n7275), .ZN(n13568) );
  NAND2_X2 U9403 ( .A1(n13567), .A2(n13488), .ZN(n13541) );
  NAND2_X2 U9404 ( .A1(n10060), .A2(n10059), .ZN(n10254) );
  NAND2_X1 U9405 ( .A1(n9518), .A2(n12409), .ZN(n9748) );
  NAND2_X1 U9406 ( .A1(n10901), .A2(n6829), .ZN(n6828) );
  NAND2_X1 U9407 ( .A1(n12889), .A2(n12888), .ZN(n6825) );
  INV_X1 U9408 ( .A(n12887), .ZN(n6826) );
  NAND2_X1 U9409 ( .A1(n6975), .A2(n6974), .ZN(n6972) );
  NAND2_X1 U9410 ( .A1(n6962), .A2(n6960), .ZN(n11433) );
  NAND2_X1 U9411 ( .A1(n6971), .A2(n11365), .ZN(n6970) );
  NAND2_X1 U9412 ( .A1(n6970), .A2(n6703), .ZN(n11368) );
  NAND2_X1 U9413 ( .A1(n12234), .A2(n13311), .ZN(n6829) );
  OAI21_X1 U9414 ( .B1(n13569), .B2(n13568), .A(n13567), .ZN(n6833) );
  NAND2_X1 U9415 ( .A1(n7133), .A2(n7987), .ZN(n8002) );
  INV_X1 U9416 ( .A(n8109), .ZN(n8108) );
  NAND2_X1 U9417 ( .A1(n7656), .A2(n7657), .ZN(n7136) );
  OAI21_X1 U9418 ( .B1(n12238), .B2(n6840), .A(n6837), .ZN(n12243) );
  INV_X1 U9419 ( .A(n6834), .ZN(n12242) );
  INV_X1 U9420 ( .A(n12267), .ZN(n6844) );
  NAND2_X1 U9421 ( .A1(n12266), .A2(n6712), .ZN(n6843) );
  OAI21_X1 U9422 ( .B1(n6844), .B2(n6843), .A(n6845), .ZN(n7320) );
  INV_X1 U9423 ( .A(n12268), .ZN(n6847) );
  NAND3_X1 U9424 ( .A1(n12258), .A2(n6849), .A3(n6593), .ZN(n6848) );
  NAND4_X1 U9425 ( .A1(n6599), .A2(n12186), .A3(n12185), .A4(n6852), .ZN(n6851) );
  AOI21_X1 U9426 ( .B1(n6599), .B2(n6652), .A(n6853), .ZN(n6850) );
  AOI21_X1 U9427 ( .B1(n12219), .B2(n12218), .A(n6868), .ZN(n6859) );
  NAND2_X1 U9428 ( .A1(n6857), .A2(n6856), .ZN(n12230) );
  NAND2_X1 U9429 ( .A1(n8539), .A2(n6875), .ZN(n6873) );
  AND2_X1 U9430 ( .A1(n11806), .A2(n11805), .ZN(n14291) );
  NAND3_X1 U9431 ( .A1(n7183), .A2(n11806), .A3(n6880), .ZN(n6879) );
  NAND2_X1 U9432 ( .A1(n6882), .A2(n6881), .ZN(P1_U3557) );
  OR2_X1 U9433 ( .A1(n14929), .A2(n11184), .ZN(n6881) );
  NAND2_X1 U9434 ( .A1(n6883), .A2(n14929), .ZN(n6882) );
  NAND2_X1 U9435 ( .A1(n14325), .A2(n14902), .ZN(n14326) );
  NAND2_X1 U9436 ( .A1(n14149), .A2(n6887), .ZN(n6884) );
  NAND2_X1 U9437 ( .A1(n6884), .A2(n6885), .ZN(n14119) );
  NAND2_X1 U9438 ( .A1(n7066), .A2(n6893), .ZN(n6892) );
  NAND2_X1 U9439 ( .A1(n6911), .A2(n6912), .ZN(n14698) );
  AND2_X1 U9440 ( .A1(n6911), .A2(n6909), .ZN(n14696) );
  OAI21_X1 U9441 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(n15544), .A(n6693), .ZN(
        n6914) );
  XNOR2_X1 U9442 ( .A(n14503), .B(n14504), .ZN(n15544) );
  INV_X1 U9443 ( .A(n7125), .ZN(n14690) );
  INV_X1 U9444 ( .A(n14527), .ZN(n6919) );
  NAND2_X1 U9445 ( .A1(n6921), .A2(n8365), .ZN(n8275) );
  NAND2_X1 U9446 ( .A1(n8366), .A2(n6920), .ZN(n13801) );
  AND2_X1 U9447 ( .A1(n6921), .A2(n7433), .ZN(n6920) );
  NAND2_X1 U9448 ( .A1(n8366), .A2(n6921), .ZN(n8394) );
  AND2_X2 U9449 ( .A1(n8576), .A2(n8267), .ZN(n6921) );
  NAND2_X1 U9450 ( .A1(n13236), .A2(n6923), .ZN(n6922) );
  OAI211_X2 U9451 ( .C1(n6595), .C2(n6925), .A(n11636), .B(n6922), .ZN(n12502)
         );
  INV_X1 U9452 ( .A(n6929), .ZN(n12148) );
  NAND2_X2 U9453 ( .A1(n8466), .A2(n7614), .ZN(n12348) );
  NOR2_X1 U9454 ( .A1(n9151), .A2(n6933), .ZN(n6932) );
  NAND2_X1 U9455 ( .A1(n6939), .A2(n6942), .ZN(n6938) );
  INV_X1 U9456 ( .A(n14935), .ZN(n6939) );
  OAI21_X1 U9457 ( .B1(n13258), .B2(n6944), .A(n6946), .ZN(n9481) );
  NAND2_X1 U9458 ( .A1(n6946), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U9459 ( .A1(n13258), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U9460 ( .A1(n6950), .A2(n13235), .ZN(P2_U3186) );
  NAND2_X1 U9461 ( .A1(n6951), .A2(n7445), .ZN(n6950) );
  XNOR2_X1 U9462 ( .A(n13230), .B(n6952), .ZN(n6951) );
  INV_X1 U9463 ( .A(n13231), .ZN(n6952) );
  NAND2_X1 U9464 ( .A1(n6961), .A2(n11419), .ZN(n6960) );
  INV_X1 U9465 ( .A(n6964), .ZN(n6961) );
  NAND2_X1 U9466 ( .A1(n6963), .A2(n11415), .ZN(n6962) );
  NAND2_X1 U9467 ( .A1(n6964), .A2(n11418), .ZN(n6963) );
  NAND2_X1 U9468 ( .A1(n11417), .A2(n11416), .ZN(n6964) );
  AND2_X1 U9469 ( .A1(n11804), .A2(n11806), .ZN(n11584) );
  NAND2_X2 U9470 ( .A1(n11288), .A2(n11287), .ZN(n14402) );
  NAND3_X1 U9471 ( .A1(n7237), .A2(n11301), .A3(n7236), .ZN(n6971) );
  OAI21_X1 U9472 ( .B1(n11466), .B2(n6987), .A(n6986), .ZN(n11485) );
  NAND2_X1 U9473 ( .A1(n11466), .A2(n6984), .ZN(n6980) );
  OAI21_X1 U9474 ( .B1(n6983), .B2(n7253), .A(n7252), .ZN(n6982) );
  NAND2_X1 U9475 ( .A1(n6987), .A2(n6986), .ZN(n6983) );
  NOR2_X1 U9476 ( .A1(n11468), .A2(n11465), .ZN(n6987) );
  OR2_X2 U9477 ( .A1(n10979), .A2(n10980), .ZN(n6991) );
  INV_X1 U9478 ( .A(n7306), .ZN(n9617) );
  INV_X1 U9479 ( .A(n9614), .ZN(n6993) );
  NAND2_X1 U9480 ( .A1(n9615), .A2(n9613), .ZN(n6994) );
  NAND3_X1 U9481 ( .A1(n7311), .A2(n7324), .A3(n6999), .ZN(n6998) );
  INV_X1 U9482 ( .A(n10726), .ZN(n6999) );
  MUX2_X1 U9483 ( .A(n13229), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9484 ( .A(n12883), .B(n10296), .S(n6765), .Z(n10301) );
  NAND2_X1 U9485 ( .A1(n11950), .A2(n11949), .ZN(n15181) );
  AND4_X2 U9486 ( .A1(n7003), .A2(n7299), .A3(n15307), .A4(n7002), .ZN(n7698)
         );
  NAND2_X1 U9487 ( .A1(n10207), .A2(n10327), .ZN(n7009) );
  NAND2_X1 U9488 ( .A1(n7009), .A2(n7007), .ZN(n10638) );
  NAND2_X1 U9489 ( .A1(n11097), .A2(n7014), .ZN(n7012) );
  NAND2_X1 U9490 ( .A1(n7012), .A2(n7013), .ZN(n11130) );
  OAI22_X1 U9491 ( .A1(n7690), .A2(n8940), .B1(n9567), .B2(n9552), .ZN(n7017)
         );
  NAND2_X4 U9492 ( .A1(n12528), .A2(n9555), .ZN(n9552) );
  NAND3_X1 U9493 ( .A1(n7520), .A2(n7728), .A3(n6613), .ZN(n7607) );
  NOR2_X2 U9494 ( .A1(n7870), .A2(n7039), .ZN(n7038) );
  NAND2_X1 U9495 ( .A1(n10530), .A2(n12215), .ZN(n10693) );
  AND2_X2 U9496 ( .A1(n7047), .A2(n9806), .ZN(n10530) );
  NAND2_X1 U9497 ( .A1(n13638), .A2(n7051), .ZN(n13561) );
  INV_X1 U9498 ( .A(n7057), .ZN(n13578) );
  INV_X1 U9499 ( .A(n8246), .ZN(n7059) );
  AND2_X1 U9500 ( .A1(n8921), .A2(n7527), .ZN(n7058) );
  NOR2_X2 U9501 ( .A1(n14194), .A2(n14364), .ZN(n14153) );
  NAND3_X1 U9502 ( .A1(n6612), .A2(n14244), .A3(n14282), .ZN(n14242) );
  NAND3_X1 U9503 ( .A1(n6601), .A2(n10310), .A3(n9709), .ZN(n10467) );
  NAND2_X1 U9504 ( .A1(n11211), .A2(n11771), .ZN(n9315) );
  XNOR2_X1 U9505 ( .A(n11211), .B(n13985), .ZN(n11587) );
  NAND2_X1 U9506 ( .A1(n8619), .A2(n8321), .ZN(n7069) );
  NAND2_X1 U9507 ( .A1(n8619), .A2(n7067), .ZN(n7066) );
  INV_X1 U9508 ( .A(n8632), .ZN(n7068) );
  XNOR2_X1 U9509 ( .A(n7069), .B(n8632), .ZN(n10438) );
  OAI21_X1 U9510 ( .B1(n8356), .B2(n8837), .A(n8358), .ZN(n7073) );
  NAND3_X1 U9511 ( .A1(n7071), .A2(n7070), .A3(n7546), .ZN(n7545) );
  NAND2_X1 U9512 ( .A1(n12305), .A2(n6581), .ZN(n7074) );
  NAND2_X1 U9513 ( .A1(n8328), .A2(n7078), .ZN(n7075) );
  NAND2_X1 U9514 ( .A1(n7075), .A2(n7076), .ZN(n8344) );
  INV_X1 U9515 ( .A(n13049), .ZN(n7084) );
  NAND2_X1 U9516 ( .A1(n13055), .A2(n13054), .ZN(n7085) );
  AND2_X2 U9517 ( .A1(n7087), .A2(n7086), .ZN(n12902) );
  NAND3_X1 U9518 ( .A1(n7098), .A2(n7682), .A3(n12581), .ZN(n11956) );
  INV_X1 U9519 ( .A(n12751), .ZN(n7097) );
  NAND2_X1 U9520 ( .A1(n12751), .A2(n15155), .ZN(n7095) );
  NAND2_X1 U9521 ( .A1(n15154), .A2(n12751), .ZN(n7096) );
  OAI22_X1 U9522 ( .A1(n12685), .A2(n15168), .B1(n7097), .B2(n12729), .ZN(
        n9918) );
  NAND2_X1 U9523 ( .A1(n11122), .A2(n7106), .ZN(n7103) );
  NAND2_X1 U9524 ( .A1(n7103), .A2(n7104), .ZN(n11867) );
  NAND2_X1 U9525 ( .A1(n11122), .A2(n12006), .ZN(n11132) );
  INV_X1 U9526 ( .A(n12006), .ZN(n7114) );
  INV_X1 U9527 ( .A(n7115), .ZN(n7597) );
  NOR2_X2 U9528 ( .A1(n7632), .A2(n7116), .ZN(n7115) );
  NAND3_X1 U9529 ( .A1(n7610), .A2(n7120), .A3(n7119), .ZN(n7118) );
  NOR2_X2 U9530 ( .A1(n7521), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7520) );
  NAND4_X1 U9531 ( .A1(n7121), .A2(n7522), .A3(n7592), .A4(n7593), .ZN(n7521)
         );
  NAND2_X1 U9532 ( .A1(n7125), .A2(n7124), .ZN(n14530) );
  INV_X1 U9533 ( .A(n14691), .ZN(n7124) );
  NAND2_X1 U9534 ( .A1(n8145), .A2(n8144), .ZN(n7131) );
  NAND2_X1 U9535 ( .A1(n8129), .A2(n8128), .ZN(n7132) );
  NAND2_X1 U9536 ( .A1(n7986), .A2(n7985), .ZN(n7133) );
  NAND2_X1 U9537 ( .A1(n7946), .A2(n7945), .ZN(n7966) );
  INV_X1 U9538 ( .A(n8164), .ZN(n7140) );
  NAND2_X1 U9539 ( .A1(n7140), .A2(n11880), .ZN(n7142) );
  NAND2_X1 U9540 ( .A1(n7142), .A2(n7143), .ZN(n11886) );
  NAND2_X1 U9541 ( .A1(n8164), .A2(n8163), .ZN(n11881) );
  NAND2_X1 U9542 ( .A1(n7692), .A2(n6695), .ZN(n7152) );
  NAND2_X1 U9543 ( .A1(n8081), .A2(n6736), .ZN(n7157) );
  NAND3_X1 U9544 ( .A1(n6673), .A2(n7158), .A3(n7157), .ZN(n8109) );
  NAND2_X1 U9545 ( .A1(n8004), .A2(n7162), .ZN(n7161) );
  INV_X1 U9546 ( .A(n8035), .ZN(n8038) );
  NAND2_X1 U9547 ( .A1(n7802), .A2(n7165), .ZN(n7164) );
  NAND3_X1 U9548 ( .A1(n7177), .A2(n7175), .A3(n10605), .ZN(n10610) );
  NAND3_X1 U9549 ( .A1(n7179), .A2(n11597), .A3(n10466), .ZN(n7177) );
  OAI21_X1 U9550 ( .B1(n11824), .B2(n7184), .A(n7181), .ZN(n7182) );
  AOI21_X1 U9551 ( .B1(n14291), .B2(n11825), .A(n7183), .ZN(n7181) );
  NAND2_X1 U9552 ( .A1(n7182), .A2(n11826), .ZN(n14258) );
  OAI21_X1 U9553 ( .B1(n14764), .B2(n7191), .A(n11591), .ZN(n7186) );
  NAND2_X1 U9554 ( .A1(n7187), .A2(n7185), .ZN(n10115) );
  INV_X1 U9555 ( .A(n7186), .ZN(n7185) );
  NOR2_X1 U9556 ( .A1(n7191), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U9557 ( .A1(n14852), .A2(n9650), .ZN(n11214) );
  NAND2_X1 U9558 ( .A1(n14383), .A2(n6704), .ZN(n14204) );
  NAND2_X1 U9559 ( .A1(n6616), .A2(n7196), .ZN(n7194) );
  NAND2_X1 U9560 ( .A1(n11858), .A2(n11857), .ZN(n14176) );
  INV_X1 U9561 ( .A(n7203), .ZN(n14178) );
  NOR2_X1 U9562 ( .A1(n14175), .A2(n7205), .ZN(n7204) );
  INV_X1 U9563 ( .A(n11857), .ZN(n7205) );
  NAND2_X1 U9564 ( .A1(n14131), .A2(n7209), .ZN(n7206) );
  NAND2_X1 U9565 ( .A1(n7206), .A2(n7208), .ZN(n12114) );
  NAND2_X1 U9566 ( .A1(n14335), .A2(n7221), .ZN(n7212) );
  AOI21_X1 U9567 ( .B1(n11229), .B2(n11230), .A(n7224), .ZN(n7222) );
  OAI21_X1 U9568 ( .B1(n11229), .B2(n6715), .A(n7223), .ZN(n7225) );
  NAND2_X1 U9569 ( .A1(n7226), .A2(n11218), .ZN(n11221) );
  NAND2_X1 U9570 ( .A1(n7230), .A2(n7228), .ZN(n7227) );
  NAND2_X1 U9571 ( .A1(n8232), .A2(n7231), .ZN(n7233) );
  NAND2_X1 U9572 ( .A1(n11278), .A2(n7240), .ZN(n7239) );
  OAI21_X1 U9573 ( .B1(n11433), .B2(n7246), .A(n7244), .ZN(n11448) );
  NAND2_X1 U9574 ( .A1(n7243), .A2(n7241), .ZN(n11447) );
  NAND2_X1 U9575 ( .A1(n11433), .A2(n7244), .ZN(n7243) );
  NOR2_X1 U9576 ( .A1(n7245), .A2(n11432), .ZN(n7246) );
  NAND2_X1 U9577 ( .A1(n9293), .A2(n6710), .ZN(n7248) );
  NAND2_X1 U9578 ( .A1(n9293), .A2(n8963), .ZN(n9292) );
  NAND2_X1 U9579 ( .A1(n11485), .A2(n7252), .ZN(n7249) );
  NAND2_X1 U9580 ( .A1(n7249), .A2(n7250), .ZN(n11506) );
  AOI21_X1 U9581 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(n7250) );
  NOR2_X1 U9582 ( .A1(n11484), .A2(n11487), .ZN(n7253) );
  NAND2_X1 U9583 ( .A1(n11191), .A2(n11190), .ZN(n11193) );
  NAND3_X1 U9584 ( .A1(n11191), .A2(n11190), .A3(n11570), .ZN(n11194) );
  NAND2_X1 U9585 ( .A1(n11273), .A2(n11274), .ZN(n11272) );
  NAND2_X1 U9586 ( .A1(n11244), .A2(n11245), .ZN(n11243) );
  NAND2_X1 U9587 ( .A1(n11451), .A2(n11450), .ZN(n11466) );
  NAND2_X1 U9588 ( .A1(n11226), .A2(n11225), .ZN(n11229) );
  OAI21_X1 U9589 ( .B1(n11431), .B2(n11200), .A(n11199), .ZN(n11201) );
  NAND2_X1 U9590 ( .A1(n11509), .A2(n11508), .ZN(n11523) );
  NAND2_X1 U9591 ( .A1(n11252), .A2(n11251), .ZN(n11265) );
  NAND2_X1 U9592 ( .A1(n11937), .A2(n6589), .ZN(n12097) );
  NAND2_X1 U9593 ( .A1(n8111), .A2(n8110), .ZN(n8129) );
  INV_X1 U9594 ( .A(n14291), .ZN(n11823) );
  NAND2_X1 U9595 ( .A1(n12097), .A2(n12096), .ZN(n12105) );
  NAND2_X1 U9596 ( .A1(n7866), .A2(n7867), .ZN(n7887) );
  NAND2_X1 U9597 ( .A1(n8078), .A2(n8077), .ZN(n8081) );
  NAND2_X1 U9598 ( .A1(n12094), .A2(n10351), .ZN(n12095) );
  NOR2_X1 U9599 ( .A1(n9823), .A2(n12179), .ZN(n9762) );
  AND2_X2 U9600 ( .A1(n9753), .A2(n15098), .ZN(n9806) );
  NAND2_X1 U9601 ( .A1(n8555), .A2(n8309), .ZN(n8573) );
  XNOR2_X1 U9602 ( .A(n14891), .B(n14749), .ZN(n11593) );
  OAI21_X2 U9603 ( .B1(n7262), .B2(n12416), .A(n7258), .ZN(n10797) );
  NAND2_X1 U9604 ( .A1(n13541), .A2(n7270), .ZN(n7266) );
  OAI211_X1 U9605 ( .C1(n13541), .C2(n6718), .A(n7266), .B(n7265), .ZN(n13497)
         );
  NAND2_X1 U9606 ( .A1(n13592), .A2(n7278), .ZN(n7277) );
  OAI21_X1 U9607 ( .B1(n13592), .B2(n7280), .A(n7278), .ZN(n13582) );
  INV_X1 U9608 ( .A(n10903), .ZN(n7288) );
  NAND2_X1 U9609 ( .A1(n7289), .A2(n10903), .ZN(n7286) );
  NOR2_X1 U9610 ( .A1(n11012), .A2(n7291), .ZN(n11013) );
  NAND2_X1 U9611 ( .A1(n6586), .A2(n13310), .ZN(n7292) );
  INV_X2 U9612 ( .A(n15103), .ZN(n12196) );
  OAI21_X2 U9613 ( .B1(n10121), .B2(n8825), .A(n8578), .ZN(n15103) );
  MUX2_X1 U9614 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n15180), .S(n9981), .Z(n9967)
         );
  NAND3_X1 U9615 ( .A1(n12209), .A2(n12208), .A3(n6717), .ZN(n7307) );
  NAND2_X1 U9616 ( .A1(n7307), .A2(n6714), .ZN(n12216) );
  OAI21_X1 U9617 ( .B1(n12201), .B2(n12198), .A(n12197), .ZN(n12199) );
  OR2_X1 U9618 ( .A1(n7310), .A2(n10726), .ZN(n10549) );
  INV_X1 U9619 ( .A(n7312), .ZN(n7310) );
  INV_X1 U9620 ( .A(n10559), .ZN(n7313) );
  INV_X1 U9621 ( .A(n10548), .ZN(n7314) );
  NAND4_X1 U9622 ( .A1(n8365), .A2(n8576), .A3(n8363), .A4(n8267), .ZN(n8360)
         );
  INV_X1 U9623 ( .A(n12260), .ZN(n7332) );
  NAND3_X1 U9624 ( .A1(n7334), .A2(n7333), .A3(n7335), .ZN(n12184) );
  NAND2_X1 U9625 ( .A1(n12174), .A2(n7336), .ZN(n7333) );
  NAND2_X1 U9626 ( .A1(n12175), .A2(n7336), .ZN(n7334) );
  INV_X1 U9627 ( .A(n11211), .ZN(n14847) );
  NAND2_X1 U9628 ( .A1(n12115), .A2(n7344), .ZN(n7343) );
  NAND2_X1 U9629 ( .A1(n12115), .A2(n11843), .ZN(n14097) );
  OAI211_X1 U9630 ( .C1(n12115), .C2(n7347), .A(n7345), .B(n7343), .ZN(n14325)
         );
  NAND2_X1 U9631 ( .A1(n10189), .A2(n7355), .ZN(n7354) );
  INV_X1 U9632 ( .A(n10189), .ZN(n7357) );
  INV_X1 U9633 ( .A(n14277), .ZN(n7363) );
  NAND2_X1 U9634 ( .A1(n14209), .A2(n7367), .ZN(n7366) );
  INV_X1 U9635 ( .A(n14374), .ZN(n7373) );
  NAND2_X1 U9636 ( .A1(n8235), .A2(n7374), .ZN(n8969) );
  NAND2_X1 U9637 ( .A1(n7380), .A2(n7376), .ZN(n7383) );
  NAND2_X1 U9638 ( .A1(n10259), .A2(n12415), .ZN(n10526) );
  NAND2_X1 U9639 ( .A1(n7402), .A2(n7406), .ZN(n7401) );
  OAI21_X1 U9640 ( .B1(n11079), .B2(n6716), .A(n7410), .ZN(n7409) );
  NAND2_X1 U9641 ( .A1(n14640), .A2(n10795), .ZN(n7417) );
  AND2_X1 U9642 ( .A1(n14944), .A2(n13312), .ZN(n7418) );
  INV_X1 U9643 ( .A(n13635), .ZN(n7430) );
  NAND2_X1 U9644 ( .A1(n13635), .A2(n7426), .ZN(n7421) );
  NOR2_X1 U9645 ( .A1(n6640), .A2(n7432), .ZN(n13626) );
  NAND2_X1 U9646 ( .A1(n13230), .A2(n7436), .ZN(n7435) );
  OAI211_X1 U9647 ( .C1(n13230), .C2(n7437), .A(n12520), .B(n7435), .ZN(
        P2_U3192) );
  INV_X1 U9648 ( .A(n12515), .ZN(n7446) );
  NAND2_X1 U9649 ( .A1(n10931), .A2(n6706), .ZN(n7452) );
  NAND2_X1 U9650 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  INV_X1 U9651 ( .A(n7452), .ZN(n11086) );
  NAND2_X1 U9652 ( .A1(n7450), .A2(n11084), .ZN(n11083) );
  INV_X1 U9653 ( .A(n11085), .ZN(n7451) );
  AND2_X1 U9654 ( .A1(n8774), .A2(n8775), .ZN(n7460) );
  NAND2_X1 U9655 ( .A1(n12502), .A2(n6709), .ZN(n13299) );
  NAND2_X1 U9656 ( .A1(n7462), .A2(n7461), .ZN(n9943) );
  AND2_X1 U9657 ( .A1(n8591), .A2(n8571), .ZN(n7461) );
  NAND2_X2 U9658 ( .A1(n7613), .A2(n14578), .ZN(n7469) );
  NAND3_X1 U9659 ( .A1(n7613), .A2(n14578), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n7468) );
  NAND2_X4 U9660 ( .A1(n7470), .A2(n7469), .ZN(n11550) );
  NAND2_X2 U9661 ( .A1(n7532), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7470) );
  NAND3_X1 U9662 ( .A1(n7470), .A2(n7469), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7467) );
  NAND2_X1 U9663 ( .A1(n13841), .A2(n7474), .ZN(n7472) );
  NAND2_X1 U9664 ( .A1(n10971), .A2(n7484), .ZN(n7481) );
  NAND2_X1 U9665 ( .A1(n9302), .A2(n9301), .ZN(n9305) );
  NAND2_X1 U9666 ( .A1(n9886), .A2(n9885), .ZN(n7491) );
  INV_X1 U9667 ( .A(n9886), .ZN(n7489) );
  NAND2_X1 U9668 ( .A1(n12551), .A2(n7494), .ZN(n7493) );
  OAI211_X1 U9669 ( .C1(n12551), .C2(n7495), .A(n7493), .B(n8225), .ZN(
        P3_U3160) );
  NOR2_X1 U9670 ( .A1(n8173), .A2(n8159), .ZN(n7499) );
  NAND2_X1 U9671 ( .A1(n8173), .A2(n8159), .ZN(n7500) );
  INV_X1 U9672 ( .A(n8173), .ZN(n7501) );
  AND2_X2 U9673 ( .A1(n13831), .A2(n11701), .ZN(n11706) );
  NAND2_X1 U9674 ( .A1(n11689), .A2(n7502), .ZN(n13831) );
  INV_X1 U9675 ( .A(n13935), .ZN(n7504) );
  NAND2_X1 U9676 ( .A1(n13887), .A2(n13888), .ZN(n13886) );
  INV_X1 U9677 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9678 ( .A1(n12626), .A2(n7793), .ZN(n7525) );
  NAND2_X1 U9679 ( .A1(n7525), .A2(n7800), .ZN(n12669) );
  NAND2_X1 U9680 ( .A1(n8249), .A2(n8248), .ZN(n8252) );
  NAND2_X1 U9681 ( .A1(n7621), .A2(n7530), .ZN(n7625) );
  OAI21_X1 U9682 ( .B1(n8554), .B2(n7537), .A(n7535), .ZN(n8575) );
  NAND2_X1 U9683 ( .A1(n8320), .A2(n8321), .ZN(n8617) );
  NAND2_X1 U9684 ( .A1(n11153), .A2(n11152), .ZN(n7554) );
  NAND2_X1 U9685 ( .A1(n7545), .A2(n7549), .ZN(n11501) );
  NAND2_X1 U9686 ( .A1(n7554), .A2(n11154), .ZN(n11462) );
  NAND2_X1 U9687 ( .A1(n8345), .A2(n7558), .ZN(n7557) );
  XNOR2_X1 U9688 ( .A(n8345), .B(n9479), .ZN(n8415) );
  NAND3_X1 U9689 ( .A1(n11564), .A2(n7564), .A3(n11563), .ZN(n13799) );
  OR2_X1 U9690 ( .A1(n13710), .A2(n15078), .ZN(n13715) );
  INV_X1 U9691 ( .A(n10655), .ZN(n10640) );
  NAND2_X1 U9692 ( .A1(n10638), .A2(n10637), .ZN(n10655) );
  NOR2_X1 U9693 ( .A1(n12105), .A2(n12104), .ZN(n12111) );
  NOR2_X1 U9694 ( .A1(n6589), .A2(n12103), .ZN(n12104) );
  NAND2_X1 U9695 ( .A1(n9766), .A2(n9514), .ZN(n12407) );
  MUX2_X2 U9696 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7599), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7600) );
  OAI21_X1 U9697 ( .B1(n9525), .B2(n9524), .A(n9523), .ZN(n9902) );
  NAND4_X2 U9698 ( .A1(n9243), .A2(n9242), .A3(n9241), .A4(n9240), .ZN(n13987)
         );
  NAND2_X1 U9699 ( .A1(n13661), .A2(n13511), .ZN(n13512) );
  NOR2_X1 U9700 ( .A1(n14789), .A2(n14860), .ZN(n14773) );
  AND2_X1 U9701 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  INV_X1 U9702 ( .A(n7601), .ZN(n12524) );
  NAND2_X1 U9703 ( .A1(n9266), .A2(n8511), .ZN(n13258) );
  AND2_X2 U9704 ( .A1(n8481), .A2(n8258), .ZN(n8576) );
  INV_X1 U9705 ( .A(n14938), .ZN(n8666) );
  NAND2_X1 U9706 ( .A1(n9144), .A2(n8445), .ZN(n9120) );
  NAND2_X1 U9707 ( .A1(n9280), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9283) );
  INV_X1 U9708 ( .A(n12152), .ZN(n12155) );
  NAND2_X1 U9709 ( .A1(n8806), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U9710 ( .A1(n7627), .A2(n7626), .ZN(n7629) );
  OR2_X1 U9711 ( .A1(n13987), .A2(n11196), .ZN(n11200) );
  AOI21_X1 U9712 ( .B1(n12278), .B2(n12277), .A(n12276), .ZN(n12337) );
  AND2_X1 U9713 ( .A1(n12342), .A2(n12334), .ZN(n12335) );
  NOR2_X2 U9714 ( .A1(n12144), .A2(n9128), .ZN(n9129) );
  NAND2_X1 U9715 ( .A1(n8444), .A2(n9128), .ZN(n8445) );
  CLKBUF_X1 U9716 ( .A(n10096), .Z(n9931) );
  AND2_X1 U9717 ( .A1(n12280), .A2(n12279), .ZN(n12336) );
  INV_X1 U9718 ( .A(n7625), .ZN(n7627) );
  AOI21_X1 U9719 ( .B1(n9298), .B2(n10100), .A(n9299), .ZN(n9301) );
  XNOR2_X1 U9720 ( .A(n14834), .B(n9298), .ZN(n9727) );
  NAND4_X2 U9721 ( .A1(n9681), .A2(n9680), .A3(n9679), .A4(n9678), .ZN(n14748)
         );
  XNOR2_X1 U9722 ( .A(n11501), .B(n11500), .ZN(n13811) );
  INV_X1 U9723 ( .A(n9235), .ZN(n9238) );
  OAI21_X1 U9724 ( .B1(SI_1_), .B2(n8288), .A(n8290), .ZN(n8421) );
  NAND2_X2 U9725 ( .A1(n13925), .A2(n11750), .ZN(n13841) );
  OAI21_X1 U9726 ( .B1(n11550), .B2(n9331), .A(n8293), .ZN(n8294) );
  NAND2_X1 U9727 ( .A1(n6575), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U9728 ( .A1(n6576), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8291) );
  NAND2_X2 U9729 ( .A1(n8399), .A2(n13805), .ZN(n11642) );
  NAND2_X1 U9730 ( .A1(n9901), .A2(n9511), .ZN(n9778) );
  OR2_X1 U9731 ( .A1(n13541), .A2(n7390), .ZN(n7568) );
  OR2_X1 U9732 ( .A1(n14098), .A2(n14102), .ZN(n7569) );
  AND2_X1 U9733 ( .A1(n13526), .A2(n13527), .ZN(n7570) );
  AND2_X1 U9734 ( .A1(n8819), .A2(n8818), .ZN(n7572) );
  AND4_X1 U9735 ( .A1(n7594), .A2(n7623), .A3(n8192), .A4(n7622), .ZN(n7573)
         );
  AND2_X1 U9736 ( .A1(n8486), .A2(n8485), .ZN(n7575) );
  AND2_X1 U9737 ( .A1(n8917), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7576) );
  INV_X1 U9738 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U9739 ( .A1(n10204), .A2(n10203), .ZN(n10207) );
  INV_X1 U9740 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U9741 ( .A1(n9331), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7577) );
  INV_X1 U9742 ( .A(n12249), .ZN(n13309) );
  INV_X1 U9743 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9234) );
  INV_X1 U9744 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8361) );
  NOR2_X1 U9745 ( .A1(n12437), .A2(n9130), .ZN(n10902) );
  INV_X1 U9746 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8287) );
  INV_X1 U9747 ( .A(n12738), .ZN(n12986) );
  INV_X1 U9748 ( .A(n6589), .ZN(n11936) );
  INV_X1 U9749 ( .A(n11990), .ZN(n10919) );
  AND2_X1 U9750 ( .A1(n8295), .A2(n8475), .ZN(n7578) );
  NOR2_X1 U9751 ( .A1(n12611), .A2(n13016), .ZN(n7579) );
  AND2_X1 U9752 ( .A1(n13094), .A2(n12923), .ZN(n7580) );
  INV_X1 U9753 ( .A(n13520), .ZN(n13492) );
  INV_X1 U9754 ( .A(n7864), .ZN(n7866) );
  NOR3_X1 U9755 ( .A1(n13489), .A2(n13555), .A3(n12432), .ZN(n7583) );
  AND2_X1 U9756 ( .A1(n14137), .A2(n13972), .ZN(n7584) );
  INV_X1 U9757 ( .A(n11812), .ZN(n14220) );
  NOR2_X1 U9758 ( .A1(n14242), .A2(n14388), .ZN(n11812) );
  INV_X1 U9759 ( .A(n14381), .ZN(n11811) );
  INV_X1 U9760 ( .A(n13752), .ZN(n13510) );
  INV_X1 U9761 ( .A(n11595), .ZN(n10433) );
  NOR2_X1 U9762 ( .A1(n11642), .A2(n9493), .ZN(n7585) );
  NAND2_X2 U9763 ( .A1(n9491), .A2(n15037), .ZN(n15045) );
  NAND2_X1 U9764 ( .A1(n12180), .A2(n12144), .ZN(n12138) );
  OR2_X1 U9765 ( .A1(n12148), .A2(n12275), .ZN(n12149) );
  INV_X1 U9766 ( .A(n12153), .ZN(n12154) );
  MUX2_X1 U9767 ( .A(n14875), .B(n14748), .S(n6799), .Z(n11233) );
  INV_X1 U9768 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U9769 ( .A1(n12166), .A2(n12165), .ZN(n12167) );
  MUX2_X1 U9770 ( .A(n13980), .B(n11258), .S(n11504), .Z(n11261) );
  INV_X1 U9771 ( .A(n11278), .ZN(n11284) );
  INV_X1 U9772 ( .A(n12228), .ZN(n12229) );
  NAND2_X1 U9773 ( .A1(n11399), .A2(n11395), .ZN(n11396) );
  NAND2_X1 U9774 ( .A1(n11403), .A2(n11402), .ZN(n11417) );
  OAI21_X1 U9775 ( .B1(n12265), .B2(n12264), .A(n12263), .ZN(n12267) );
  MUX2_X1 U9776 ( .A(n13971), .B(n14337), .S(n11504), .Z(n11505) );
  INV_X1 U9777 ( .A(n15166), .ZN(n11917) );
  NOR3_X1 U9778 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_24__SCAN_IN), .ZN(n8244) );
  INV_X1 U9779 ( .A(n11966), .ZN(n10639) );
  INV_X1 U9780 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7622) );
  INV_X1 U9781 ( .A(n13874), .ZN(n10832) );
  INV_X1 U9782 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7626) );
  INV_X1 U9783 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8680) );
  INV_X1 U9784 ( .A(n8470), .ZN(n8467) );
  AND2_X1 U9785 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(n8892), .ZN(n11638) );
  NAND2_X1 U9786 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  INV_X1 U9787 ( .A(n12412), .ZN(n9802) );
  INV_X1 U9788 ( .A(n11771), .ZN(n11746) );
  INV_X1 U9789 ( .A(n9885), .ZN(n9884) );
  INV_X1 U9790 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11316) );
  INV_X1 U9791 ( .A(n11324), .ZN(n11173) );
  INV_X1 U9792 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10449) );
  INV_X1 U9793 ( .A(n11318), .ZN(n11174) );
  AND2_X1 U9794 ( .A1(n14364), .A2(n14183), .ZN(n11859) );
  INV_X1 U9795 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8964) );
  INV_X1 U9796 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n15306) );
  INV_X1 U9797 ( .A(n7976), .ZN(n7975) );
  INV_X1 U9798 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7813) );
  INV_X1 U9799 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7927) );
  INV_X1 U9800 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10741) );
  INV_X1 U9801 ( .A(n11919), .ZN(n10643) );
  INV_X1 U9802 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7733) );
  INV_X1 U9803 ( .A(n9945), .ZN(n8591) );
  OR2_X1 U9804 ( .A1(n8810), .A2(n8809), .ZN(n8828) );
  NAND2_X1 U9805 ( .A1(n8841), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8843) );
  OR2_X1 U9806 ( .A1(n8681), .A2(n8680), .ZN(n8699) );
  NOR2_X1 U9807 ( .A1(n8843), .A2(n8886), .ZN(n8892) );
  INV_X1 U9808 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8410) );
  AND2_X1 U9809 ( .A1(n11638), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n12296) );
  AOI21_X1 U9810 ( .B1(n13712), .B2(n15118), .A(n13711), .ZN(n13713) );
  INV_X1 U9811 ( .A(n12351), .ZN(n8880) );
  OR2_X1 U9812 ( .A1(n11730), .A2(n11729), .ZN(n11731) );
  OR2_X1 U9813 ( .A1(n11714), .A2(n11713), .ZN(n11715) );
  NAND2_X1 U9814 ( .A1(n11741), .A2(n11742), .ZN(n11743) );
  OR2_X1 U9815 ( .A1(n11470), .A2(n11469), .ZN(n11489) );
  NAND2_X1 U9816 ( .A1(n11178), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U9817 ( .A1(n11175), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U9818 ( .A1(n11176), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U9819 ( .A1(n11174), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U9820 ( .A1(n10587), .A2(n10586), .ZN(n11290) );
  NAND2_X1 U9821 ( .A1(n11413), .A2(n7614), .ZN(n9329) );
  INV_X1 U9822 ( .A(SI_22_), .ZN(n8354) );
  INV_X1 U9823 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14458) );
  OR2_X1 U9824 ( .A1(n7911), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7929) );
  OR2_X1 U9825 ( .A1(n8086), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9826 ( .A1(n8010), .A2(n8009), .ZN(n8025) );
  NAND2_X1 U9827 ( .A1(n8114), .A2(n15524), .ZN(n8133) );
  NAND2_X1 U9828 ( .A1(n7975), .A2(n7974), .ZN(n7993) );
  NAND2_X1 U9829 ( .A1(n7896), .A2(n7895), .ZN(n7911) );
  OR2_X1 U9830 ( .A1(n8133), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U9831 ( .A1(n7928), .A2(n7927), .ZN(n7953) );
  INV_X1 U9832 ( .A(n15142), .ZN(n12837) );
  OR2_X1 U9833 ( .A1(n8167), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12533) );
  INV_X1 U9834 ( .A(n12740), .ZN(n13030) );
  AND4_X1 U9835 ( .A1(n7981), .A2(n7980), .A3(n7979), .A4(n7978), .ZN(n13041)
         );
  INV_X1 U9836 ( .A(n10351), .ZN(n15186) );
  AND2_X1 U9837 ( .A1(n9848), .A2(n10343), .ZN(n10345) );
  NOR2_X1 U9838 ( .A1(n8199), .A2(n13214), .ZN(n9835) );
  AND2_X1 U9839 ( .A1(n7886), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U9840 ( .A1(n8743), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8760) );
  INV_X1 U9841 ( .A(n10626), .ZN(n8693) );
  INV_X1 U9842 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15436) );
  INV_X1 U9843 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U9844 ( .A1(n9014), .A2(n9013), .ZN(n14996) );
  NAND2_X1 U9845 ( .A1(n13586), .A2(n13667), .ZN(n13544) );
  INV_X1 U9846 ( .A(n13585), .ZN(n13516) );
  INV_X1 U9847 ( .A(n13509), .ZN(n13513) );
  INV_X1 U9848 ( .A(n13667), .ZN(n13595) );
  INV_X1 U9849 ( .A(n12389), .ZN(n12457) );
  INV_X1 U9850 ( .A(n13971), .ZN(n11797) );
  OR2_X1 U9851 ( .A1(n11435), .A2(n13911), .ZN(n11453) );
  OR2_X1 U9852 ( .A1(n11572), .A2(n9359), .ZN(n9372) );
  AND2_X1 U9853 ( .A1(n11489), .A2(n11471), .ZN(n14122) );
  OR2_X1 U9854 ( .A1(n11385), .A2(n13862), .ZN(n11404) );
  INV_X1 U9855 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10287) );
  NAND2_X1 U9856 ( .A1(n13970), .A2(n14750), .ZN(n11846) );
  INV_X1 U9857 ( .A(n14153), .ZN(n14170) );
  NAND2_X1 U9858 ( .A1(n11812), .A2(n11811), .ZN(n14214) );
  INV_X1 U9859 ( .A(n14205), .ZN(n11855) );
  OAI21_X1 U9860 ( .B1(n14339), .B2(n14879), .A(n14338), .ZN(n14340) );
  OR2_X1 U9861 ( .A1(n11692), .A2(n10305), .ZN(n14556) );
  INV_X1 U9862 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14453) );
  NAND2_X2 U9863 ( .A1(n8211), .A2(n8210), .ZN(n12731) );
  AND2_X1 U9864 ( .A1(n11906), .A2(n11905), .ZN(n12530) );
  INV_X1 U9865 ( .A(n11900), .ZN(n8171) );
  AND4_X1 U9866 ( .A1(n7916), .A2(n7915), .A3(n7914), .A4(n7913), .ZN(n13075)
         );
  INV_X1 U9867 ( .A(n12883), .ZN(n12834) );
  INV_X1 U9868 ( .A(n12891), .ZN(n12767) );
  INV_X1 U9869 ( .A(n12896), .ZN(n12819) );
  AND2_X1 U9870 ( .A1(n9556), .A2(n12862), .ZN(n12895) );
  INV_X1 U9871 ( .A(n13041), .ZN(n13063) );
  INV_X1 U9872 ( .A(n15195), .ZN(n15154) );
  INV_X1 U9873 ( .A(n12983), .ZN(n14611) );
  NAND2_X1 U9874 ( .A1(n10349), .A2(n15186), .ZN(n15184) );
  INV_X1 U9875 ( .A(n13112), .ZN(n15221) );
  OR2_X1 U9876 ( .A1(n8174), .A2(n13213), .ZN(n15236) );
  INV_X1 U9877 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7647) );
  INV_X1 U9878 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7923) );
  INV_X1 U9879 ( .A(n12188), .ZN(n15090) );
  OR2_X1 U9880 ( .A1(n6583), .A2(n13551), .ZN(n12324) );
  OR2_X1 U9881 ( .A1(n13605), .A2(n8438), .ZN(n8406) );
  AND4_X1 U9882 ( .A1(n8750), .A2(n8749), .A3(n8748), .A4(n8747), .ZN(n12249)
         );
  AND2_X1 U9883 ( .A1(n9039), .A2(n9010), .ZN(n15002) );
  AND2_X1 U9884 ( .A1(n9014), .A2(n13807), .ZN(n9039) );
  INV_X1 U9885 ( .A(n13489), .ZN(n13526) );
  AND2_X1 U9886 ( .A1(n13479), .A2(n12399), .ZN(n13664) );
  INV_X1 U9887 ( .A(n15039), .ZN(n13665) );
  NOR2_X1 U9888 ( .A1(n9138), .A2(n9137), .ZN(n9489) );
  AND2_X1 U9889 ( .A1(n9127), .A2(n12137), .ZN(n15078) );
  INV_X1 U9890 ( .A(n9127), .ZN(n15126) );
  INV_X1 U9891 ( .A(n12137), .ZN(n15088) );
  AND2_X1 U9892 ( .A1(n11007), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8873) );
  AND2_X1 U9893 ( .A1(n8968), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9055) );
  INV_X1 U9894 ( .A(n9383), .ZN(n9387) );
  OR2_X1 U9895 ( .A1(n13826), .A2(n11491), .ZN(n11497) );
  NAND4_X2 U9896 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9650)
         );
  AND2_X1 U9897 ( .A1(n8976), .A2(n8975), .ZN(n9065) );
  INV_X1 U9898 ( .A(n14723), .ZN(n14733) );
  XNOR2_X1 U9899 ( .A(n14097), .B(n11860), .ZN(n11848) );
  INV_X1 U9900 ( .A(n14189), .ZN(n14750) );
  INV_X1 U9901 ( .A(n11831), .ZN(n14227) );
  NAND2_X1 U9902 ( .A1(n9697), .A2(n9696), .ZN(n14902) );
  XNOR2_X1 U9903 ( .A(n13877), .B(n13978), .ZN(n11599) );
  AOI21_X1 U9904 ( .B1(n9354), .B2(n9341), .A(n9340), .ZN(n10319) );
  INV_X1 U9905 ( .A(n14340), .ZN(n14341) );
  AND2_X1 U9906 ( .A1(n14556), .A2(n14879), .ZN(n14828) );
  INV_X1 U9907 ( .A(n14556), .ZN(n14882) );
  INV_X1 U9908 ( .A(n14828), .ZN(n14906) );
  INV_X1 U9909 ( .A(n9371), .ZN(n9378) );
  INV_X1 U9910 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U9911 ( .A1(n14451), .A2(n14450), .ZN(n14507) );
  AND2_X1 U9912 ( .A1(n9564), .A2(n9563), .ZN(n15142) );
  INV_X1 U9913 ( .A(n12915), .ZN(n13094) );
  INV_X1 U9914 ( .A(n8224), .ZN(n8225) );
  INV_X1 U9915 ( .A(n12724), .ZN(n12699) );
  NAND2_X1 U9916 ( .A1(n8203), .A2(n10349), .ZN(n12734) );
  OR2_X1 U9917 ( .A1(n8286), .A2(n13213), .ZN(n12753) );
  INV_X1 U9918 ( .A(n12895), .ZN(n10243) );
  NAND2_X1 U9919 ( .A1(P3_U3897), .A2(n12528), .ZN(n12891) );
  NAND2_X1 U9920 ( .A1(n15198), .A2(n15197), .ZN(n12983) );
  INV_X1 U9921 ( .A(n14583), .ZN(n13081) );
  INV_X1 U9922 ( .A(n12632), .ZN(n10812) );
  INV_X1 U9923 ( .A(n15235), .ZN(n15233) );
  INV_X1 U9924 ( .A(n12495), .ZN(n13170) );
  INV_X1 U9925 ( .A(n12675), .ZN(n11109) );
  AND2_X1 U9926 ( .A1(n9837), .A2(n9836), .ZN(n15223) );
  INV_X1 U9927 ( .A(n13215), .ZN(n13213) );
  INV_X1 U9928 ( .A(SI_27_), .ZN(n12499) );
  NOR2_X1 U9929 ( .A1(n6575), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13221) );
  INV_X1 U9930 ( .A(SI_17_), .ZN(n9456) );
  INV_X1 U9931 ( .A(SI_12_), .ZN(n8985) );
  NAND2_X1 U9932 ( .A1(n9109), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14947) );
  OR2_X1 U9933 ( .A1(n13238), .A2(n15039), .ZN(n14932) );
  NAND2_X1 U9934 ( .A1(n8884), .A2(n8875), .ZN(n14939) );
  NAND2_X1 U9935 ( .A1(n8406), .A2(n8405), .ZN(n13585) );
  OR2_X1 U9936 ( .A1(n8767), .A2(n8766), .ZN(n13308) );
  INV_X1 U9937 ( .A(n15002), .ZN(n15018) );
  INV_X1 U9938 ( .A(n14949), .ZN(n15032) );
  INV_X1 U9939 ( .A(n13644), .ZN(n13697) );
  INV_X1 U9940 ( .A(n15141), .ZN(n15139) );
  INV_X1 U9941 ( .A(n15129), .ZN(n15127) );
  NOR2_X1 U9942 ( .A1(n15051), .A2(n15048), .ZN(n15049) );
  NAND2_X1 U9943 ( .A1(n8870), .A2(n8869), .ZN(n15053) );
  INV_X1 U9944 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11009) );
  INV_X1 U9945 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9899) );
  INV_X1 U9946 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9106) );
  INV_X1 U9947 ( .A(n14271), .ZN(n14647) );
  INV_X1 U9948 ( .A(n13949), .ZN(n13963) );
  NAND2_X1 U9949 ( .A1(n11516), .A2(n11515), .ZN(n14102) );
  INV_X1 U9950 ( .A(n13861), .ZN(n14168) );
  INV_X1 U9951 ( .A(n14738), .ZN(n14721) );
  INV_X1 U9952 ( .A(n14731), .ZN(n14729) );
  OR2_X1 U9953 ( .A1(n14103), .A2(n11573), .ZN(n14273) );
  AND2_X1 U9954 ( .A1(n14204), .A2(n14203), .ZN(n14377) );
  AND2_X1 U9955 ( .A1(n14103), .A2(n14783), .ZN(n14797) );
  OR2_X1 U9956 ( .A1(n14797), .A2(n9646), .ZN(n14292) );
  INV_X1 U9957 ( .A(n14929), .ZN(n14926) );
  NAND2_X1 U9958 ( .A1(n14342), .A2(n14341), .ZN(n14409) );
  AND3_X1 U9959 ( .A1(n14658), .A2(n14657), .A3(n14656), .ZN(n14676) );
  INV_X1 U9960 ( .A(n14909), .ZN(n14908) );
  AND2_X2 U9961 ( .A1(n10321), .A2(n10320), .ZN(n14909) );
  CLKBUF_X1 U9962 ( .A(n14810), .Z(n14825) );
  INV_X1 U9963 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12135) );
  INV_X1 U9964 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9277) );
  AND2_X2 U9965 ( .A1(n7698), .A2(n7587), .ZN(n7727) );
  NOR2_X1 U9966 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7594) );
  INV_X1 U9967 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7595) );
  XNOR2_X2 U9968 ( .A(n7596), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U9969 ( .A1(n7598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7599) );
  NAND2_X2 U9970 ( .A1(n7600), .A2(n7597), .ZN(n13225) );
  NAND2_X1 U9971 ( .A1(n7758), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7606) );
  AND2_X2 U9972 ( .A1(n7601), .A2(n7602), .ZN(n7761) );
  NAND2_X1 U9973 ( .A1(n7761), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7605) );
  AND2_X4 U9974 ( .A1(n7601), .A2(n13225), .ZN(n11900) );
  NAND2_X1 U9975 ( .A1(n11900), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7604) );
  AND2_X2 U9976 ( .A1(n12524), .A2(n7602), .ZN(n7681) );
  NAND2_X1 U9977 ( .A1(n7681), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9978 ( .A1(n7607), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7608) );
  MUX2_X1 U9979 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7608), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7609) );
  NAND2_X2 U9980 ( .A1(n7598), .A2(n7609), .ZN(n12528) );
  INV_X1 U9981 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n15307) );
  XNOR2_X1 U9982 ( .A(n15307), .B(n7612), .ZN(n9567) );
  INV_X1 U9983 ( .A(n11550), .ZN(n7614) );
  INV_X1 U9984 ( .A(SI_1_), .ZN(n8940) );
  XNOR2_X1 U9985 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7657) );
  XNOR2_X1 U9986 ( .A(n7657), .B(n7655), .ZN(n8939) );
  NAND2_X1 U9987 ( .A1(n7758), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U9988 ( .A1(n7761), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7617) );
  NAND2_X1 U9989 ( .A1(n11900), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7616) );
  NAND2_X1 U9990 ( .A1(n7681), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7615) );
  NAND4_X1 U9991 ( .A1(n7618), .A2(n7617), .A3(n7615), .A4(n7616), .ZN(n12754)
         );
  INV_X1 U9992 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9249) );
  NAND2_X1 U9993 ( .A1(n9249), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U9994 ( .A1(n7655), .A2(n7619), .ZN(n7620) );
  MUX2_X1 U9995 ( .A(n7620), .B(SI_0_), .S(n11550), .Z(n13229) );
  NAND2_X1 U9996 ( .A1(n7625), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7624) );
  XNOR2_X1 U9997 ( .A(n7636), .B(P3_B_REG_SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9998 ( .A1(n7632), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7633) );
  INV_X1 U9999 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7635) );
  NAND2_X1 U10000 ( .A1(n8174), .A2(n7635), .ZN(n7638) );
  NAND2_X1 U10001 ( .A1(n7636), .A2(n10941), .ZN(n7637) );
  NAND2_X2 U10002 ( .A1(n7638), .A2(n7637), .ZN(n9842) );
  NAND2_X1 U10003 ( .A1(n7642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7639) );
  MUX2_X1 U10004 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7639), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7640) );
  NAND2_X1 U10005 ( .A1(n6679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7641) );
  MUX2_X1 U10006 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7641), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7643) );
  NAND2_X1 U10007 ( .A1(n7643), .A2(n7642), .ZN(n10195) );
  INV_X1 U10008 ( .A(n10195), .ZN(n10205) );
  NAND2_X1 U10009 ( .A1(n10350), .A2(n10205), .ZN(n12100) );
  NAND2_X1 U10010 ( .A1(n12754), .A2(n9504), .ZN(n15188) );
  NAND2_X1 U10011 ( .A1(n7717), .A2(n15188), .ZN(n7650) );
  NAND2_X1 U10012 ( .A1(n10198), .A2(n7650), .ZN(n7653) );
  XNOR2_X1 U10013 ( .A(n6585), .B(n9633), .ZN(n7651) );
  NAND3_X1 U10014 ( .A1(n9503), .A2(n7717), .A3(n9633), .ZN(n7652) );
  NAND2_X1 U10015 ( .A1(n9631), .A2(n7654), .ZN(n9915) );
  OR2_X1 U10016 ( .A1(n7690), .A2(SI_2_), .ZN(n7666) );
  INV_X1 U10017 ( .A(n7655), .ZN(n7656) );
  INV_X1 U10018 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U10019 ( .A1(n8916), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7658) );
  XNOR2_X1 U10020 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7659) );
  XNOR2_X1 U10021 ( .A(n7671), .B(n7659), .ZN(n8936) );
  NOR2_X1 U10022 ( .A1(n7660), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U10023 ( .A1(n8005), .A2(n9981), .ZN(n7664) );
  XNOR2_X1 U10024 ( .A(n7680), .B(n10199), .ZN(n7685) );
  NAND2_X1 U10025 ( .A1(n7761), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U10026 ( .A1(n6584), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U10027 ( .A1(n11900), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7668) );
  NAND2_X1 U10028 ( .A1(n7681), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7667) );
  XNOR2_X1 U10029 ( .A(n7685), .B(n12752), .ZN(n9916) );
  OR2_X1 U10030 ( .A1(n7690), .A2(SI_3_), .ZN(n7679) );
  INV_X1 U10031 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U10032 ( .A1(n9312), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7672) );
  XNOR2_X1 U10033 ( .A(n8915), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7673) );
  XNOR2_X1 U10034 ( .A(n7691), .B(n7673), .ZN(n8909) );
  OR2_X1 U10035 ( .A1(n7843), .A2(n8909), .ZN(n7678) );
  NAND2_X1 U10036 ( .A1(n7663), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7674) );
  MUX2_X1 U10037 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7674), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7676) );
  NAND2_X1 U10038 ( .A1(n7676), .A2(n7675), .ZN(n9593) );
  NAND2_X1 U10039 ( .A1(n8005), .A2(n9593), .ZN(n7677) );
  XNOR2_X1 U10040 ( .A(n7680), .B(n12581), .ZN(n7687) );
  NAND2_X1 U10041 ( .A1(n7758), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U10042 ( .A1(n11900), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U10043 ( .A1(n7681), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7682) );
  INV_X1 U10044 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n12582) );
  XNOR2_X1 U10045 ( .A(n7687), .B(n12751), .ZN(n12578) );
  NAND2_X1 U10046 ( .A1(n7685), .A2(n15192), .ZN(n12575) );
  AND2_X1 U10047 ( .A1(n12578), .A2(n12575), .ZN(n7686) );
  NAND2_X1 U10048 ( .A1(n12576), .A2(n7686), .ZN(n12577) );
  INV_X1 U10049 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U10050 ( .A1(n7688), .A2(n12751), .ZN(n7689) );
  NAND2_X1 U10051 ( .A1(n12577), .A2(n7689), .ZN(n12660) );
  INV_X1 U10052 ( .A(n12660), .ZN(n7715) );
  OR2_X1 U10053 ( .A1(n6590), .A2(SI_4_), .ZN(n7705) );
  NAND2_X1 U10054 ( .A1(n8915), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10055 ( .A1(n9657), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U10056 ( .A1(n8925), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U10057 ( .A1(n7718), .A2(n7694), .ZN(n7695) );
  NAND2_X1 U10058 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  AND2_X1 U10059 ( .A1(n7719), .A2(n7697), .ZN(n8911) );
  OR2_X1 U10060 ( .A1(n7843), .A2(n8911), .ZN(n7704) );
  INV_X1 U10061 ( .A(n7699), .ZN(n7702) );
  NAND2_X1 U10062 ( .A1(n7675), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7700) );
  MUX2_X1 U10063 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7700), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7701) );
  NAND2_X1 U10064 ( .A1(n7702), .A2(n7701), .ZN(n9598) );
  NAND2_X1 U10065 ( .A1(n8005), .A2(n9598), .ZN(n7703) );
  AND3_X2 U10066 ( .A1(n7705), .A2(n7704), .A3(n7703), .ZN(n12663) );
  XNOR2_X1 U10067 ( .A(n7752), .B(n12663), .ZN(n7711) );
  NAND2_X1 U10068 ( .A1(n7758), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U10069 ( .A1(n11900), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7709) );
  AND2_X1 U10070 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7706) );
  NOR2_X1 U10071 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7734) );
  OR2_X1 U10072 ( .A1(n7706), .A2(n7734), .ZN(n12664) );
  NAND2_X1 U10073 ( .A1(n6587), .A2(n12664), .ZN(n7708) );
  NAND2_X1 U10074 ( .A1(n7681), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10075 ( .A1(n7711), .A2(n10657), .ZN(n7716) );
  INV_X1 U10076 ( .A(n7711), .ZN(n7712) );
  NAND2_X1 U10077 ( .A1(n7712), .A2(n12750), .ZN(n7713) );
  NAND2_X1 U10078 ( .A1(n7716), .A2(n7713), .ZN(n12659) );
  NAND2_X1 U10079 ( .A1(n7715), .A2(n7714), .ZN(n12657) );
  NAND2_X1 U10080 ( .A1(n12657), .A2(n7716), .ZN(n12627) );
  OR2_X1 U10081 ( .A1(n6590), .A2(SI_5_), .ZN(n7732) );
  NAND2_X1 U10082 ( .A1(n8933), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10083 ( .A1(n8926), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U10084 ( .A1(n7744), .A2(n7720), .ZN(n7722) );
  NAND2_X1 U10085 ( .A1(n7721), .A2(n7722), .ZN(n7725) );
  INV_X1 U10086 ( .A(n7721), .ZN(n7724) );
  INV_X1 U10087 ( .A(n7722), .ZN(n7723) );
  NAND2_X1 U10088 ( .A1(n7724), .A2(n7723), .ZN(n7745) );
  AND2_X1 U10089 ( .A1(n7725), .A2(n7745), .ZN(n8913) );
  OR2_X1 U10090 ( .A1(n7843), .A2(n8913), .ZN(n7731) );
  NOR2_X1 U10091 ( .A1(n7699), .A2(n7662), .ZN(n7726) );
  MUX2_X1 U10092 ( .A(n7662), .B(n7726), .S(P3_IR_REG_5__SCAN_IN), .Z(n7729)
         );
  OR2_X1 U10093 ( .A1(n7729), .A2(n7728), .ZN(n9585) );
  NAND2_X1 U10094 ( .A1(n8005), .A2(n9585), .ZN(n7730) );
  XNOR2_X1 U10095 ( .A(n9635), .B(n12632), .ZN(n7778) );
  NAND2_X1 U10096 ( .A1(n10271), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7739) );
  INV_X2 U10097 ( .A(n6579), .ZN(n11901) );
  NAND2_X1 U10098 ( .A1(n11901), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10099 ( .A1(n7734), .A2(n7733), .ZN(n7785) );
  OR2_X1 U10100 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U10101 ( .A1(n7785), .A2(n7735), .ZN(n12633) );
  NAND2_X1 U10102 ( .A1(n6587), .A2(n12633), .ZN(n7737) );
  NAND2_X1 U10103 ( .A1(n11900), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7736) );
  XNOR2_X1 U10104 ( .A(n7778), .B(n12749), .ZN(n12628) );
  NAND2_X1 U10105 ( .A1(n7728), .A2(n7779), .ZN(n7772) );
  NAND2_X1 U10106 ( .A1(n7742), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7741) );
  MUX2_X1 U10107 ( .A(n7741), .B(P3_IR_REG_31__SCAN_IN), .S(n7740), .Z(n7743)
         );
  NAND2_X1 U10108 ( .A1(n7743), .A2(n7806), .ZN(n10225) );
  NAND2_X1 U10109 ( .A1(n7745), .A2(n7744), .ZN(n7782) );
  INV_X1 U10110 ( .A(n7781), .ZN(n7746) );
  NAND2_X1 U10111 ( .A1(n8951), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10112 ( .A1(n8952), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10113 ( .A1(n7748), .A2(n7747), .ZN(n7768) );
  XNOR2_X1 U10114 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7749) );
  XNOR2_X1 U10115 ( .A(n7802), .B(n7749), .ZN(n8935) );
  OR2_X1 U10116 ( .A1(n7843), .A2(n8935), .ZN(n7751) );
  INV_X1 U10117 ( .A(SI_8_), .ZN(n8934) );
  OR2_X1 U10118 ( .A1(n6590), .A2(n8934), .ZN(n7750) );
  OAI211_X1 U10119 ( .C1(n9552), .C2(n10225), .A(n7751), .B(n7750), .ZN(n12600) );
  XNOR2_X1 U10120 ( .A(n7752), .B(n10916), .ZN(n7797) );
  NAND2_X1 U10121 ( .A1(n11901), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7757) );
  INV_X2 U10122 ( .A(n7851), .ZN(n10271) );
  NAND2_X1 U10123 ( .A1(n10271), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7756) );
  NOR2_X1 U10124 ( .A1(n7762), .A2(n15525), .ZN(n7753) );
  OR2_X1 U10125 ( .A1(n7814), .A2(n7753), .ZN(n12601) );
  NAND2_X1 U10126 ( .A1(n6587), .A2(n12601), .ZN(n7755) );
  NAND2_X1 U10127 ( .A1(n11900), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U10128 ( .A(n7797), .B(n10921), .ZN(n7794) );
  NAND2_X1 U10129 ( .A1(n6584), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U10130 ( .A1(n7681), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7759) );
  AND2_X1 U10131 ( .A1(n7760), .A2(n7759), .ZN(n7767) );
  AND2_X1 U10132 ( .A1(n7787), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7763) );
  OR2_X1 U10133 ( .A1(n7763), .A2(n7762), .ZN(n12546) );
  NAND2_X1 U10134 ( .A1(n6587), .A2(n12546), .ZN(n7765) );
  NAND2_X1 U10135 ( .A1(n11900), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7764) );
  AND2_X1 U10136 ( .A1(n7765), .A2(n7764), .ZN(n7766) );
  OR2_X1 U10137 ( .A1(n6590), .A2(SI_7_), .ZN(n7777) );
  NAND2_X1 U10138 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  AND2_X1 U10139 ( .A1(n7771), .A2(n7770), .ZN(n8918) );
  OR2_X1 U10140 ( .A1(n7843), .A2(n8918), .ZN(n7776) );
  NAND2_X1 U10141 ( .A1(n7772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7774) );
  INV_X1 U10142 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U10143 ( .A(n7774), .B(n7773), .ZN(n10052) );
  NAND2_X1 U10144 ( .A1(n8005), .A2(n10052), .ZN(n7775) );
  NAND2_X1 U10145 ( .A1(n10645), .A2(n15209), .ZN(n11983) );
  INV_X1 U10146 ( .A(n15209), .ZN(n10711) );
  NAND2_X1 U10147 ( .A1(n12748), .A2(n10711), .ZN(n11982) );
  XNOR2_X1 U10148 ( .A(n10708), .B(n6770), .ZN(n7796) );
  NAND2_X1 U10149 ( .A1(n7778), .A2(n10644), .ZN(n12541) );
  OR2_X1 U10150 ( .A1(n7728), .A2(n7662), .ZN(n7780) );
  XNOR2_X1 U10151 ( .A(n7780), .B(n7779), .ZN(n10028) );
  INV_X1 U10152 ( .A(SI_6_), .ZN(n8942) );
  OR2_X1 U10153 ( .A1(n6590), .A2(n8942), .ZN(n7784) );
  XNOR2_X1 U10154 ( .A(n7782), .B(n7781), .ZN(n8941) );
  OR2_X1 U10155 ( .A1(n7843), .A2(n8941), .ZN(n7783) );
  OAI211_X1 U10156 ( .C1(n9552), .C2(n10028), .A(n7784), .B(n7783), .ZN(n12714) );
  XNOR2_X1 U10157 ( .A(n7752), .B(n12714), .ZN(n12542) );
  NAND2_X1 U10158 ( .A1(n10271), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U10159 ( .A1(n11901), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10160 ( .A1(n7785), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10161 ( .A1(n7787), .A2(n7786), .ZN(n12716) );
  NAND2_X1 U10162 ( .A1(n6587), .A2(n12716), .ZN(n7789) );
  NAND2_X1 U10163 ( .A1(n11900), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10164 ( .A1(n12542), .A2(n10703), .ZN(n7792) );
  AND4_X1 U10165 ( .A1(n7794), .A2(n7796), .A3(n12541), .A4(n7792), .ZN(n7793)
         );
  INV_X1 U10166 ( .A(n7794), .ZN(n12596) );
  INV_X1 U10167 ( .A(n12542), .ZN(n7795) );
  NAND2_X1 U10168 ( .A1(n7795), .A2(n12631), .ZN(n12543) );
  OAI21_X1 U10169 ( .B1(n12596), .B2(n12543), .A(n7796), .ZN(n7799) );
  INV_X1 U10170 ( .A(n7796), .ZN(n12594) );
  OAI21_X1 U10171 ( .B1(n12596), .B2(n10645), .A(n12594), .ZN(n7798) );
  AOI22_X1 U10172 ( .A1(n7799), .A2(n7798), .B1(n7797), .B2(n12747), .ZN(n7800) );
  NAND2_X1 U10173 ( .A1(n8961), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10174 ( .A1(n8960), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7803) );
  XNOR2_X1 U10175 ( .A(n8991), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7804) );
  XNOR2_X1 U10176 ( .A(n7823), .B(n7804), .ZN(n8948) );
  OR2_X1 U10177 ( .A1(n7843), .A2(n8948), .ZN(n7812) );
  OR2_X1 U10178 ( .A1(n6590), .A2(SI_9_), .ZN(n7811) );
  NAND2_X1 U10179 ( .A1(n7806), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7805) );
  MUX2_X1 U10180 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7805), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7809) );
  INV_X1 U10181 ( .A(n7806), .ZN(n7808) );
  INV_X1 U10182 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10183 ( .A1(n7808), .A2(n7807), .ZN(n7844) );
  NAND2_X1 U10184 ( .A1(n7809), .A2(n7844), .ZN(n10233) );
  NAND2_X1 U10185 ( .A1(n8005), .A2(n10233), .ZN(n7810) );
  XNOR2_X1 U10186 ( .A(n9635), .B(n12675), .ZN(n7836) );
  NAND2_X1 U10187 ( .A1(n11901), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U10188 ( .A1(n10271), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7818) );
  OR2_X1 U10189 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  NAND2_X1 U10190 ( .A1(n7830), .A2(n7815), .ZN(n12676) );
  NAND2_X1 U10191 ( .A1(n6587), .A2(n12676), .ZN(n7817) );
  NAND2_X1 U10192 ( .A1(n11900), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7816) );
  NAND4_X1 U10193 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n15153) );
  INV_X1 U10194 ( .A(n15153), .ZN(n11111) );
  XNOR2_X1 U10195 ( .A(n7836), .B(n11111), .ZN(n12672) );
  INV_X1 U10196 ( .A(n12672), .ZN(n7820) );
  NAND2_X1 U10197 ( .A1(n8991), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7821) );
  XNOR2_X1 U10198 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7824) );
  XNOR2_X1 U10199 ( .A(n7841), .B(n7824), .ZN(n8953) );
  OR2_X1 U10200 ( .A1(n7843), .A2(n8953), .ZN(n7829) );
  OR2_X1 U10201 ( .A1(n6590), .A2(SI_10_), .ZN(n7828) );
  NAND2_X1 U10202 ( .A1(n7844), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7826) );
  INV_X1 U10203 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7825) );
  XNOR2_X1 U10204 ( .A(n7826), .B(n7825), .ZN(n10557) );
  NAND2_X1 U10205 ( .A1(n8005), .A2(n10557), .ZN(n7827) );
  XNOR2_X1 U10206 ( .A(n9635), .B(n15159), .ZN(n7838) );
  NAND2_X1 U10207 ( .A1(n10271), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U10208 ( .A1(n11901), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10209 ( .A1(n7830), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10210 ( .A1(n7849), .A2(n7831), .ZN(n15160) );
  NAND2_X1 U10211 ( .A1(n6587), .A2(n15160), .ZN(n7833) );
  NAND2_X1 U10212 ( .A1(n11900), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7832) );
  XNOR2_X1 U10213 ( .A(n7838), .B(n12746), .ZN(n12568) );
  NAND2_X1 U10214 ( .A1(n7836), .A2(n11111), .ZN(n12566) );
  AND2_X1 U10215 ( .A1(n12568), .A2(n12566), .ZN(n7837) );
  INV_X1 U10216 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U10217 ( .A1(n7839), .A2(n12746), .ZN(n7840) );
  XNOR2_X1 U10218 ( .A(n9161), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7842) );
  XNOR2_X1 U10219 ( .A(n7863), .B(n7842), .ZN(n8955) );
  NAND2_X1 U10220 ( .A1(n8955), .A2(n11897), .ZN(n7848) );
  OAI21_X1 U10221 ( .B1(n7844), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7845) );
  XNOR2_X1 U10222 ( .A(n7845), .B(P3_IR_REG_11__SCAN_IN), .ZN(n10559) );
  NAND2_X1 U10223 ( .A1(n8005), .A2(n10559), .ZN(n7847) );
  OR2_X1 U10224 ( .A1(n6590), .A2(n8956), .ZN(n7846) );
  XNOR2_X1 U10225 ( .A(n9635), .B(n12694), .ZN(n7856) );
  AND2_X1 U10226 ( .A1(n7849), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7850) );
  OR2_X1 U10227 ( .A1(n7874), .A2(n7850), .ZN(n14604) );
  NAND2_X1 U10228 ( .A1(n6587), .A2(n14604), .ZN(n7855) );
  NAND2_X1 U10229 ( .A1(n11901), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U10230 ( .A1(n11900), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10231 ( .A1(n10271), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10232 ( .A1(n12690), .A2(n15156), .ZN(n7860) );
  INV_X1 U10233 ( .A(n7856), .ZN(n7857) );
  NAND2_X1 U10234 ( .A1(n7858), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U10235 ( .A1(n7860), .A2(n7859), .ZN(n10971) );
  NAND2_X1 U10236 ( .A1(n9161), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U10237 ( .A1(n9277), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10238 ( .A1(n9279), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7865) );
  INV_X1 U10239 ( .A(n7867), .ZN(n7868) );
  NAND2_X1 U10240 ( .A1(n7864), .A2(n7868), .ZN(n7869) );
  NAND2_X1 U10241 ( .A1(n7887), .A2(n7869), .ZN(n8986) );
  NAND2_X1 U10242 ( .A1(n8986), .A2(n11897), .ZN(n7873) );
  NAND2_X1 U10243 ( .A1(n6817), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7871) );
  XNOR2_X1 U10244 ( .A(n7871), .B(n7523), .ZN(n10881) );
  AOI22_X1 U10245 ( .A1(n8006), .A2(n8985), .B1(n8005), .B2(n10881), .ZN(n7872) );
  XNOR2_X1 U10246 ( .A(n14597), .B(n9635), .ZN(n7881) );
  NAND2_X1 U10247 ( .A1(n7874), .A2(n10741), .ZN(n7897) );
  INV_X1 U10248 ( .A(n7874), .ZN(n7875) );
  NAND2_X1 U10249 ( .A1(n7875), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10250 ( .A1(n7897), .A2(n7876), .ZN(n14593) );
  NAND2_X1 U10251 ( .A1(n6587), .A2(n14593), .ZN(n7880) );
  NAND2_X1 U10252 ( .A1(n11901), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10253 ( .A1(n11900), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U10254 ( .A1(n10271), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7877) );
  NAND4_X1 U10255 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n12745) );
  NAND2_X1 U10256 ( .A1(n7881), .A2(n12745), .ZN(n7883) );
  INV_X1 U10257 ( .A(n7881), .ZN(n7882) );
  NAND2_X1 U10258 ( .A1(n7882), .A2(n14603), .ZN(n7885) );
  NAND2_X1 U10259 ( .A1(n7883), .A2(n7885), .ZN(n10972) );
  INV_X1 U10260 ( .A(n10972), .ZN(n7884) );
  NAND2_X1 U10261 ( .A1(n7889), .A2(n9451), .ZN(n7890) );
  NAND2_X1 U10262 ( .A1(n7906), .A2(n7890), .ZN(n9108) );
  NAND2_X1 U10263 ( .A1(n9108), .A2(n11897), .ZN(n7894) );
  NAND2_X1 U10264 ( .A1(n6726), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7891) );
  MUX2_X1 U10265 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7891), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7892) );
  NAND2_X1 U10266 ( .A1(n7892), .A2(n7644), .ZN(n10992) );
  AOI22_X1 U10267 ( .A1(n8006), .A2(n9107), .B1(n8005), .B2(n10992), .ZN(n7893) );
  NAND2_X1 U10268 ( .A1(n7894), .A2(n7893), .ZN(n13211) );
  XNOR2_X1 U10269 ( .A(n13211), .B(n6770), .ZN(n7903) );
  NAND2_X1 U10270 ( .A1(n10271), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10271 ( .A1(n11901), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7901) );
  INV_X1 U10272 ( .A(n7897), .ZN(n7896) );
  INV_X1 U10273 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U10274 ( .A1(n7897), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U10275 ( .A1(n7911), .A2(n7898), .ZN(n11133) );
  NAND2_X1 U10276 ( .A1(n6587), .A2(n11133), .ZN(n7900) );
  NAND2_X1 U10277 ( .A1(n11900), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7899) );
  NAND4_X1 U10278 ( .A1(n7902), .A2(n7901), .A3(n7900), .A4(n7899), .ZN(n14591) );
  INV_X1 U10279 ( .A(n14591), .ZN(n11104) );
  AND2_X1 U10280 ( .A1(n7903), .A2(n11104), .ZN(n10942) );
  INV_X1 U10281 ( .A(n7903), .ZN(n7904) );
  NAND2_X1 U10282 ( .A1(n7904), .A2(n14591), .ZN(n10943) );
  NAND2_X1 U10283 ( .A1(n9860), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10284 ( .A1(n9856), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10285 ( .A1(n7920), .A2(n7907), .ZN(n7917) );
  XNOR2_X1 U10286 ( .A(n7919), .B(n7917), .ZN(n9177) );
  NAND2_X1 U10287 ( .A1(n9177), .A2(n11897), .ZN(n7910) );
  NAND2_X1 U10288 ( .A1(n7644), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7908) );
  XNOR2_X1 U10289 ( .A(n7908), .B(P3_IR_REG_14__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U10290 ( .A1(n8006), .A2(SI_14_), .B1(n8005), .B2(n10987), .ZN(
        n7909) );
  NAND2_X1 U10291 ( .A1(n7910), .A2(n7909), .ZN(n12462) );
  XNOR2_X1 U10292 ( .A(n12462), .B(n9635), .ZN(n7936) );
  NAND2_X1 U10293 ( .A1(n10271), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10294 ( .A1(n11901), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10295 ( .A1(n7911), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U10296 ( .A1(n7929), .A2(n7912), .ZN(n11124) );
  NAND2_X1 U10297 ( .A1(n6587), .A2(n11124), .ZN(n7914) );
  NAND2_X1 U10298 ( .A1(n11900), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7913) );
  XNOR2_X1 U10299 ( .A(n7936), .B(n13075), .ZN(n11138) );
  INV_X1 U10300 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10301 ( .A1(n15464), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10302 ( .A1(n9938), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10303 ( .A1(n7942), .A2(n7921), .ZN(n7939) );
  XNOR2_X1 U10304 ( .A(n7941), .B(n7939), .ZN(n9263) );
  NAND2_X1 U10305 ( .A1(n9263), .A2(n11897), .ZN(n7926) );
  OR2_X1 U10306 ( .A1(n7922), .A2(n7662), .ZN(n7924) );
  XNOR2_X1 U10307 ( .A(n7924), .B(n7923), .ZN(n12814) );
  INV_X1 U10308 ( .A(n12814), .ZN(n12801) );
  AOI22_X1 U10309 ( .A1(n8006), .A2(SI_15_), .B1(n8005), .B2(n12801), .ZN(
        n7925) );
  NAND2_X1 U10310 ( .A1(n7926), .A2(n7925), .ZN(n12466) );
  XNOR2_X1 U10311 ( .A(n12466), .B(n9635), .ZN(n7937) );
  INV_X1 U10312 ( .A(n7937), .ZN(n7935) );
  NAND2_X1 U10313 ( .A1(n10271), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10314 ( .A1(n11901), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7933) );
  NAND2_X1 U10315 ( .A1(n7929), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10316 ( .A1(n7953), .A2(n7930), .ZN(n13079) );
  NAND2_X1 U10317 ( .A1(n6587), .A2(n13079), .ZN(n7932) );
  NAND2_X1 U10318 ( .A1(n11900), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7931) );
  NAND4_X1 U10319 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n13062) );
  AND2_X1 U10320 ( .A1(n7935), .A2(n13062), .ZN(n7938) );
  OR2_X1 U10321 ( .A1(n11138), .A2(n7938), .ZN(n7962) );
  NAND2_X1 U10322 ( .A1(n7936), .A2(n13075), .ZN(n11139) );
  XNOR2_X1 U10323 ( .A(n7937), .B(n13062), .ZN(n11143) );
  AND2_X1 U10324 ( .A1(n11139), .A2(n11143), .ZN(n11140) );
  OR2_X1 U10325 ( .A1(n7938), .A2(n11140), .ZN(n7960) );
  INV_X1 U10326 ( .A(n7939), .ZN(n7940) );
  NAND2_X1 U10327 ( .A1(n7941), .A2(n7940), .ZN(n7943) );
  NAND2_X1 U10328 ( .A1(n7943), .A2(n7942), .ZN(n7946) );
  NAND2_X1 U10329 ( .A1(n9629), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10330 ( .A1(n9625), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7944) );
  OR2_X1 U10331 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  AND2_X1 U10332 ( .A1(n7966), .A2(n7947), .ZN(n9401) );
  NAND2_X1 U10333 ( .A1(n9401), .A2(n11897), .ZN(n7952) );
  NOR2_X1 U10334 ( .A1(n7948), .A2(n7662), .ZN(n7949) );
  MUX2_X1 U10335 ( .A(n7662), .B(n7949), .S(P3_IR_REG_16__SCAN_IN), .Z(n7950)
         );
  AOI22_X1 U10336 ( .A1(n8006), .A2(SI_16_), .B1(n8005), .B2(n12830), .ZN(
        n7951) );
  NAND2_X1 U10337 ( .A1(n7952), .A2(n7951), .ZN(n13147) );
  XNOR2_X1 U10338 ( .A(n13147), .B(n6770), .ZN(n11064) );
  NAND2_X1 U10339 ( .A1(n10271), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U10340 ( .A1(n11901), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10341 ( .A1(n7953), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10342 ( .A1(n7976), .A2(n7954), .ZN(n13068) );
  NAND2_X1 U10343 ( .A1(n6587), .A2(n13068), .ZN(n7956) );
  NAND2_X1 U10344 ( .A1(n11900), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7955) );
  NAND4_X1 U10345 ( .A1(n7958), .A2(n7957), .A3(n7956), .A4(n7955), .ZN(n12743) );
  OAI21_X1 U10346 ( .B1(n11066), .B2(n11064), .A(n12743), .ZN(n7964) );
  AND2_X1 U10347 ( .A1(n7960), .A2(n11064), .ZN(n7961) );
  XNOR2_X1 U10348 ( .A(n9899), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n7967) );
  XNOR2_X1 U10349 ( .A(n7986), .B(n7967), .ZN(n9455) );
  NAND2_X1 U10350 ( .A1(n9455), .A2(n11897), .ZN(n7973) );
  NOR2_X1 U10351 ( .A1(n7968), .A2(n7662), .ZN(n7969) );
  MUX2_X1 U10352 ( .A(n7662), .B(n7969), .S(P3_IR_REG_17__SCAN_IN), .Z(n7970)
         );
  INV_X1 U10353 ( .A(n7970), .ZN(n7971) );
  AND2_X1 U10354 ( .A1(n7971), .A2(n7989), .ZN(n12849) );
  AOI22_X1 U10355 ( .A1(n8006), .A2(SI_17_), .B1(n8005), .B2(n12849), .ZN(
        n7972) );
  NAND2_X1 U10356 ( .A1(n7973), .A2(n7972), .ZN(n12642) );
  XNOR2_X1 U10357 ( .A(n12642), .B(n6770), .ZN(n12638) );
  NAND2_X1 U10358 ( .A1(n10271), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10359 ( .A1(n11901), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7980) );
  INV_X1 U10360 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10361 ( .A1(n7976), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U10362 ( .A1(n7993), .A2(n7977), .ZN(n13056) );
  NAND2_X1 U10363 ( .A1(n6587), .A2(n13056), .ZN(n7979) );
  NAND2_X1 U10364 ( .A1(n11900), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7978) );
  AND2_X1 U10365 ( .A1(n12638), .A2(n13063), .ZN(n7984) );
  INV_X1 U10366 ( .A(n12638), .ZN(n7982) );
  NAND2_X1 U10367 ( .A1(n7982), .A2(n13041), .ZN(n7983) );
  NAND2_X1 U10368 ( .A1(n9899), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U10369 ( .A1(n9898), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7987) );
  INV_X1 U10370 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U10371 ( .A1(n10107), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8003) );
  INV_X1 U10372 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U10373 ( .A1(n10111), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10374 ( .A1(n8003), .A2(n7988), .ZN(n8001) );
  XNOR2_X1 U10375 ( .A(n8002), .B(n8001), .ZN(n9478) );
  NAND2_X1 U10376 ( .A1(n9478), .A2(n11897), .ZN(n7992) );
  NAND2_X1 U10377 ( .A1(n7989), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7990) );
  XNOR2_X1 U10378 ( .A(n7990), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U10379 ( .A1(n8006), .A2(SI_18_), .B1(n8005), .B2(n12888), .ZN(
        n7991) );
  XNOR2_X1 U10380 ( .A(n13136), .B(n7752), .ZN(n7999) );
  NAND2_X1 U10381 ( .A1(n10271), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10382 ( .A1(n11901), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7997) );
  NAND2_X1 U10383 ( .A1(n7993), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10384 ( .A1(n8011), .A2(n7994), .ZN(n13045) );
  NAND2_X1 U10385 ( .A1(n6587), .A2(n13045), .ZN(n7996) );
  NAND2_X1 U10386 ( .A1(n11900), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7995) );
  XNOR2_X1 U10387 ( .A(n7999), .B(n13053), .ZN(n12700) );
  INV_X1 U10388 ( .A(n7999), .ZN(n8000) );
  INV_X1 U10389 ( .A(n13053), .ZN(n12742) );
  XNOR2_X1 U10390 ( .A(n10393), .B(P1_DATAO_REG_19__SCAN_IN), .ZN(n8019) );
  XNOR2_X1 U10391 ( .A(n8020), .B(n8019), .ZN(n9508) );
  NAND2_X1 U10392 ( .A1(n9508), .A2(n11897), .ZN(n8008) );
  INV_X1 U10393 ( .A(SI_19_), .ZN(n9507) );
  AOI22_X1 U10394 ( .A1(n8006), .A2(n9507), .B1(n8005), .B2(n6589), .ZN(n8007)
         );
  XNOR2_X1 U10395 ( .A(n13193), .B(n9635), .ZN(n8017) );
  NAND2_X1 U10396 ( .A1(n10271), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10397 ( .A1(n11901), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8015) );
  INV_X1 U10398 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U10399 ( .A1(n8011), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10400 ( .A1(n8025), .A2(n8012), .ZN(n13034) );
  NAND2_X1 U10401 ( .A1(n6587), .A2(n13034), .ZN(n8014) );
  NAND2_X1 U10402 ( .A1(n11900), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8013) );
  XNOR2_X1 U10403 ( .A(n8017), .B(n13042), .ZN(n12588) );
  NAND2_X1 U10404 ( .A1(n8017), .A2(n6752), .ZN(n8018) );
  NAND2_X1 U10405 ( .A1(n10393), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8021) );
  INV_X1 U10406 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U10407 ( .A1(n10786), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8039) );
  INV_X1 U10408 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U10409 ( .A1(n10748), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U10410 ( .A1(n8039), .A2(n8022), .ZN(n8036) );
  XNOR2_X1 U10411 ( .A(n8035), .B(n8036), .ZN(n9962) );
  NAND2_X1 U10412 ( .A1(n9962), .A2(n11897), .ZN(n8024) );
  OR2_X1 U10413 ( .A1(n6590), .A2(n9964), .ZN(n8023) );
  NAND2_X2 U10414 ( .A1(n8024), .A2(n8023), .ZN(n13020) );
  XNOR2_X1 U10415 ( .A(n13020), .B(n9635), .ZN(n12681) );
  NAND2_X1 U10416 ( .A1(n10271), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U10417 ( .A1(n11901), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10418 ( .A1(n8025), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10419 ( .A1(n8045), .A2(n8026), .ZN(n13019) );
  NAND2_X1 U10420 ( .A1(n6587), .A2(n13019), .ZN(n8028) );
  NAND2_X1 U10421 ( .A1(n11900), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8027) );
  NAND4_X1 U10422 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n12740) );
  NAND2_X1 U10423 ( .A1(n12681), .A2(n13030), .ZN(n8031) );
  NAND2_X1 U10424 ( .A1(n12683), .A2(n8031), .ZN(n8034) );
  INV_X1 U10425 ( .A(n12681), .ZN(n8032) );
  NAND2_X1 U10426 ( .A1(n8032), .A2(n12740), .ZN(n8033) );
  INV_X1 U10427 ( .A(n8036), .ZN(n8037) );
  XNOR2_X1 U10428 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n8056) );
  XNOR2_X1 U10429 ( .A(n8058), .B(n8056), .ZN(n10220) );
  NAND2_X1 U10430 ( .A1(n10220), .A2(n11897), .ZN(n8042) );
  INV_X1 U10431 ( .A(SI_21_), .ZN(n10221) );
  OR2_X1 U10432 ( .A1(n6590), .A2(n10221), .ZN(n8041) );
  XNOR2_X1 U10433 ( .A(n12611), .B(n9635), .ZN(n8051) );
  INV_X1 U10434 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10435 ( .A1(n8045), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U10436 ( .A1(n8065), .A2(n8046), .ZN(n13002) );
  NAND2_X1 U10437 ( .A1(n13002), .A2(n6587), .ZN(n8050) );
  NAND2_X1 U10438 ( .A1(n7758), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10439 ( .A1(n11900), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10440 ( .A1(n10271), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8047) );
  NAND4_X1 U10441 ( .A1(n8050), .A2(n8049), .A3(n8048), .A4(n8047), .ZN(n13016) );
  NAND2_X1 U10442 ( .A1(n8051), .A2(n12987), .ZN(n8055) );
  INV_X1 U10443 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U10444 ( .A1(n8052), .A2(n13016), .ZN(n8053) );
  NAND2_X1 U10445 ( .A1(n8055), .A2(n8053), .ZN(n12609) );
  INV_X1 U10446 ( .A(n12609), .ZN(n8054) );
  INV_X1 U10447 ( .A(n8056), .ZN(n8057) );
  INV_X1 U10448 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U10449 ( .A1(n11149), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8059) );
  INV_X1 U10450 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8076) );
  XNOR2_X1 U10451 ( .A(n8076), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8073) );
  XNOR2_X1 U10452 ( .A(n8075), .B(n8073), .ZN(n10340) );
  NAND2_X1 U10453 ( .A1(n10340), .A2(n11897), .ZN(n8061) );
  OR2_X1 U10454 ( .A1(n6590), .A2(n8354), .ZN(n8060) );
  XNOR2_X1 U10455 ( .A(n12483), .B(n9635), .ZN(n8062) );
  OR2_X2 U10456 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  INV_X1 U10457 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10458 ( .A1(n8065), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U10459 ( .A1(n8086), .A2(n8066), .ZN(n12990) );
  NAND2_X1 U10460 ( .A1(n12990), .A2(n6587), .ZN(n8070) );
  NAND2_X1 U10461 ( .A1(n10271), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10462 ( .A1(n7758), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8067) );
  AND2_X1 U10463 ( .A1(n8068), .A2(n8067), .ZN(n8069) );
  OAI211_X1 U10464 ( .C1(n8171), .C2(n8071), .A(n8070), .B(n8069), .ZN(n12739)
         );
  INV_X1 U10465 ( .A(n8073), .ZN(n8074) );
  NAND2_X1 U10466 ( .A1(n8076), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10467 ( .A1(n11009), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8091) );
  INV_X1 U10468 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U10469 ( .A1(n15419), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U10470 ( .A1(n8091), .A2(n8079), .ZN(n8080) );
  NAND2_X1 U10471 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U10472 ( .A1(n8092), .A2(n8082), .ZN(n10489) );
  INV_X1 U10473 ( .A(SI_23_), .ZN(n15465) );
  XNOR2_X1 U10474 ( .A(n13111), .B(n7752), .ZN(n8083) );
  NOR2_X1 U10475 ( .A1(n8084), .A2(n8083), .ZN(n8090) );
  INV_X1 U10476 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U10477 ( .A1(n8086), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10478 ( .A1(n8096), .A2(n8087), .ZN(n12976) );
  NAND2_X1 U10479 ( .A1(n12976), .A2(n6587), .ZN(n8089) );
  AOI22_X1 U10480 ( .A1(n10271), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n11901), 
        .B2(P3_REG0_REG_23__SCAN_IN), .ZN(n8088) );
  OAI211_X1 U10481 ( .C1(n8171), .C2(n12978), .A(n8089), .B(n8088), .ZN(n12738) );
  INV_X1 U10482 ( .A(n8090), .ZN(n12648) );
  XNOR2_X1 U10483 ( .A(n8108), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U10484 ( .A1(n10851), .A2(n11897), .ZN(n8094) );
  INV_X1 U10485 ( .A(SI_24_), .ZN(n10852) );
  OR2_X1 U10486 ( .A1(n6590), .A2(n10852), .ZN(n8093) );
  XNOR2_X1 U10487 ( .A(n13107), .B(n9635), .ZN(n8104) );
  INV_X1 U10488 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12650) );
  NAND2_X1 U10489 ( .A1(n8096), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10490 ( .A1(n8115), .A2(n8097), .ZN(n12960) );
  NAND2_X1 U10491 ( .A1(n12960), .A2(n6587), .ZN(n8103) );
  INV_X1 U10492 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10493 ( .A1(n7758), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10494 ( .A1(n10271), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8098) );
  OAI211_X1 U10495 ( .C1(n8100), .C2(n8171), .A(n8099), .B(n8098), .ZN(n8101)
         );
  INV_X1 U10496 ( .A(n8101), .ZN(n8102) );
  NAND2_X1 U10497 ( .A1(n8104), .A2(n12972), .ZN(n8107) );
  INV_X1 U10498 ( .A(n8104), .ZN(n8105) );
  INV_X1 U10499 ( .A(n12972), .ZN(n12938) );
  NAND2_X1 U10500 ( .A1(n8105), .A2(n12938), .ZN(n8106) );
  NAND2_X1 U10501 ( .A1(n8107), .A2(n8106), .ZN(n12647) );
  AOI21_X2 U10502 ( .B1(n12558), .B2(n12648), .A(n12647), .ZN(n12617) );
  INV_X1 U10503 ( .A(n8107), .ZN(n12619) );
  NAND2_X1 U10504 ( .A1(n8109), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10505 ( .A1(n6664), .A2(n7160), .ZN(n8110) );
  INV_X1 U10506 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14435) );
  XNOR2_X1 U10507 ( .A(n14435), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n8127) );
  XNOR2_X1 U10508 ( .A(n8129), .B(n8127), .ZN(n10928) );
  NAND2_X1 U10509 ( .A1(n10928), .A2(n11897), .ZN(n8113) );
  INV_X1 U10510 ( .A(SI_25_), .ZN(n10929) );
  OR2_X1 U10511 ( .A1(n6590), .A2(n10929), .ZN(n8112) );
  XNOR2_X1 U10512 ( .A(n13103), .B(n9635), .ZN(n8123) );
  INV_X1 U10513 ( .A(n8115), .ZN(n8114) );
  INV_X1 U10514 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15524) );
  NAND2_X1 U10515 ( .A1(n8115), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8116) );
  NAND2_X1 U10516 ( .A1(n8133), .A2(n8116), .ZN(n12944) );
  NAND2_X1 U10517 ( .A1(n12944), .A2(n6587), .ZN(n8122) );
  INV_X1 U10518 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10519 ( .A1(n10271), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10520 ( .A1(n11900), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8117) );
  OAI211_X1 U10521 ( .C1(n6579), .C2(n8119), .A(n8118), .B(n8117), .ZN(n8120)
         );
  INV_X1 U10522 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U10523 ( .A1(n8123), .A2(n12951), .ZN(n8126) );
  INV_X1 U10524 ( .A(n8123), .ZN(n8124) );
  INV_X1 U10525 ( .A(n12951), .ZN(n12727) );
  NAND2_X1 U10526 ( .A1(n8124), .A2(n12727), .ZN(n8125) );
  NAND2_X1 U10527 ( .A1(n12616), .A2(n8126), .ZN(n12722) );
  INV_X1 U10528 ( .A(n8127), .ZN(n8128) );
  NAND2_X1 U10529 ( .A1(n14435), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8130) );
  INV_X1 U10530 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15333) );
  XNOR2_X1 U10531 ( .A(n15333), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n8143) );
  XNOR2_X1 U10532 ( .A(n8145), .B(n8143), .ZN(n10939) );
  NAND2_X1 U10533 ( .A1(n10939), .A2(n11897), .ZN(n8132) );
  XNOR2_X1 U10534 ( .A(n12931), .B(n6770), .ZN(n8140) );
  NAND2_X1 U10535 ( .A1(n8133), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10536 ( .A1(n8151), .A2(n8134), .ZN(n12927) );
  NAND2_X1 U10537 ( .A1(n12927), .A2(n6587), .ZN(n8139) );
  INV_X1 U10538 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12929) );
  NAND2_X1 U10539 ( .A1(n10271), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10540 ( .A1(n7758), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8135) );
  OAI211_X1 U10541 ( .C1(n12929), .C2(n8171), .A(n8136), .B(n8135), .ZN(n8137)
         );
  INV_X1 U10542 ( .A(n8137), .ZN(n8138) );
  NOR2_X1 U10543 ( .A1(n8140), .A2(n12939), .ZN(n8141) );
  AOI21_X1 U10544 ( .B1(n8140), .B2(n12939), .A(n8141), .ZN(n12723) );
  NAND2_X1 U10545 ( .A1(n12722), .A2(n12723), .ZN(n12721) );
  INV_X1 U10546 ( .A(n8141), .ZN(n8142) );
  INV_X1 U10547 ( .A(n8143), .ZN(n8144) );
  NAND2_X1 U10548 ( .A1(n15333), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8146) );
  INV_X1 U10549 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14429) );
  XNOR2_X1 U10550 ( .A(n14429), .B(P1_DATAO_REG_27__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10551 ( .A(n8162), .B(n8160), .ZN(n12497) );
  NAND2_X1 U10552 ( .A1(n12497), .A2(n11897), .ZN(n8148) );
  XNOR2_X1 U10553 ( .A(n12915), .B(n6770), .ZN(n8158) );
  INV_X1 U10554 ( .A(n8151), .ZN(n8150) );
  INV_X1 U10555 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U10556 ( .A1(n8150), .A2(n8149), .ZN(n8167) );
  NAND2_X1 U10557 ( .A1(n8151), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10558 ( .A1(n8167), .A2(n8152), .ZN(n12911) );
  NAND2_X1 U10559 ( .A1(n12911), .A2(n6587), .ZN(n8157) );
  INV_X1 U10560 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12912) );
  NAND2_X1 U10561 ( .A1(n10271), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U10562 ( .A1(n6584), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8153) );
  OAI211_X1 U10563 ( .C1(n12912), .C2(n8171), .A(n8154), .B(n8153), .ZN(n8155)
         );
  INV_X1 U10564 ( .A(n8155), .ZN(n8156) );
  NOR2_X1 U10565 ( .A1(n8158), .A2(n12737), .ZN(n8159) );
  AOI21_X1 U10566 ( .B1(n8158), .B2(n12737), .A(n8159), .ZN(n12553) );
  INV_X1 U10567 ( .A(n8160), .ZN(n8161) );
  NAND2_X1 U10568 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  NAND2_X1 U10569 ( .A1(n14429), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10570 ( .A(n12135), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n11879) );
  XNOR2_X1 U10571 ( .A(n11881), .B(n11879), .ZN(n11163) );
  NAND2_X1 U10572 ( .A1(n11163), .A2(n11897), .ZN(n8166) );
  INV_X1 U10573 ( .A(SI_28_), .ZN(n11164) );
  OR2_X1 U10574 ( .A1(n6590), .A2(n11164), .ZN(n8165) );
  NAND2_X1 U10575 ( .A1(n8167), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10576 ( .A1(n12533), .A2(n8168), .ZN(n12488) );
  INV_X1 U10577 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U10578 ( .A1(n10271), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U10579 ( .A1(n6584), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8169) );
  OAI211_X1 U10580 ( .C1(n12489), .C2(n8171), .A(n8170), .B(n8169), .ZN(n8172)
         );
  NAND2_X1 U10581 ( .A1(n12495), .A2(n12909), .ZN(n11878) );
  XOR2_X1 U10582 ( .A(n9635), .B(n12492), .Z(n8173) );
  INV_X1 U10583 ( .A(n9842), .ZN(n13216) );
  INV_X1 U10584 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10585 ( .A1(n8174), .A2(n8175), .ZN(n8178) );
  NAND2_X1 U10586 ( .A1(n8176), .A2(n10941), .ZN(n8177) );
  NOR2_X1 U10587 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8182) );
  NOR4_X1 U10588 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8181) );
  NOR4_X1 U10589 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8180) );
  NOR4_X1 U10590 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8179) );
  NAND4_X1 U10591 ( .A1(n8182), .A2(n8181), .A3(n8180), .A4(n8179), .ZN(n8188)
         );
  NOR4_X1 U10592 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8186) );
  NOR4_X1 U10593 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8185) );
  NOR4_X1 U10594 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8184) );
  NOR4_X1 U10595 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n8183) );
  NAND4_X1 U10596 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8187)
         );
  OAI21_X1 U10597 ( .B1(n8188), .B2(n8187), .A(n8174), .ZN(n9844) );
  AND3_X1 U10598 ( .A1(n13216), .A2(n13214), .A3(n9844), .ZN(n9833) );
  NOR2_X1 U10599 ( .A1(n7636), .A2(n10941), .ZN(n8190) );
  INV_X1 U10600 ( .A(n8176), .ZN(n8189) );
  NAND2_X1 U10601 ( .A1(n8190), .A2(n8189), .ZN(n8286) );
  NAND2_X1 U10602 ( .A1(n8191), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10603 ( .A1(n6589), .A2(n10350), .ZN(n8197) );
  NAND2_X1 U10604 ( .A1(n10350), .A2(n10195), .ZN(n8195) );
  XNOR2_X1 U10605 ( .A(n12107), .B(n8195), .ZN(n8196) );
  NAND2_X1 U10606 ( .A1(n8197), .A2(n8196), .ZN(n9834) );
  INV_X1 U10607 ( .A(n12107), .ZN(n9849) );
  AND2_X1 U10608 ( .A1(n9834), .A2(n15183), .ZN(n10196) );
  AND2_X1 U10609 ( .A1(n9843), .A2(n10196), .ZN(n8198) );
  NAND2_X1 U10610 ( .A1(n9833), .A2(n8198), .ZN(n8202) );
  NAND2_X1 U10611 ( .A1(n9842), .A2(n9844), .ZN(n8199) );
  NAND2_X1 U10612 ( .A1(n11936), .A2(n12107), .ZN(n10206) );
  NOR2_X1 U10613 ( .A1(n10206), .A2(n12100), .ZN(n8204) );
  NAND2_X1 U10614 ( .A1(n9843), .A2(n8204), .ZN(n9831) );
  INV_X1 U10615 ( .A(n9831), .ZN(n8200) );
  NAND2_X1 U10616 ( .A1(n9835), .A2(n8200), .ZN(n8201) );
  NAND2_X1 U10617 ( .A1(n11936), .A2(n10195), .ZN(n10351) );
  OR2_X1 U10618 ( .A1(n9833), .A2(n15186), .ZN(n8203) );
  AND2_X1 U10619 ( .A1(n9843), .A2(n15210), .ZN(n10349) );
  INV_X1 U10620 ( .A(n9834), .ZN(n8208) );
  INV_X1 U10621 ( .A(n8204), .ZN(n8205) );
  OR2_X1 U10622 ( .A1(n9835), .A2(n8205), .ZN(n8207) );
  NAND2_X1 U10623 ( .A1(n6589), .A2(n10195), .ZN(n12092) );
  NAND2_X1 U10624 ( .A1(n12092), .A2(n12076), .ZN(n9848) );
  AND3_X1 U10625 ( .A1(n8286), .A2(n9550), .A3(n9848), .ZN(n8206) );
  OAI211_X1 U10626 ( .C1(n9833), .C2(n8208), .A(n8207), .B(n8206), .ZN(n8209)
         );
  NAND2_X1 U10627 ( .A1(n8209), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8211) );
  NOR2_X1 U10628 ( .A1(n12092), .A2(n12087), .ZN(n9838) );
  NAND2_X1 U10629 ( .A1(n9843), .A2(n9838), .ZN(n12106) );
  OR2_X1 U10630 ( .A1(n9835), .A2(n12106), .ZN(n8210) );
  INV_X1 U10631 ( .A(n12533), .ZN(n8212) );
  NAND2_X1 U10632 ( .A1(n8212), .A2(n6587), .ZN(n11906) );
  INV_X1 U10633 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n15379) );
  NAND2_X1 U10634 ( .A1(n10271), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10635 ( .A1(n11900), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8213) );
  OAI211_X1 U10636 ( .C1(n6579), .C2(n15379), .A(n8214), .B(n8213), .ZN(n8215)
         );
  INV_X1 U10637 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U10638 ( .A1(n11906), .A2(n8216), .ZN(n12736) );
  INV_X1 U10639 ( .A(n12736), .ZN(n8221) );
  INV_X1 U10640 ( .A(n12528), .ZN(n9554) );
  NAND2_X1 U10641 ( .A1(n9554), .A2(n12884), .ZN(n9565) );
  NAND2_X1 U10642 ( .A1(n9565), .A2(n9552), .ZN(n10209) );
  INV_X1 U10643 ( .A(n10209), .ZN(n8217) );
  NOR2_X1 U10644 ( .A1(n12106), .A2(n8217), .ZN(n8218) );
  NOR2_X1 U10645 ( .A1(n12106), .A2(n10209), .ZN(n8219) );
  INV_X2 U10646 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AOI22_X1 U10647 ( .A1(n12737), .A2(n12726), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8220) );
  OAI21_X1 U10648 ( .B1(n8221), .B2(n12729), .A(n8220), .ZN(n8222) );
  AOI21_X1 U10649 ( .B1(n12488), .B2(n12731), .A(n8222), .ZN(n8223) );
  OAI21_X1 U10650 ( .B1(n13170), .B2(n12734), .A(n8223), .ZN(n8224) );
  NOR2_X1 U10651 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .ZN(n8229) );
  AND4_X2 U10652 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n8233)
         );
  AND4_X2 U10653 ( .A1(n8920), .A2(n8929), .A3(n8231), .A4(n8230), .ZN(n8232)
         );
  AND2_X2 U10654 ( .A1(n8902), .A2(n8903), .ZN(n8921) );
  NOR2_X1 U10655 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n8238) );
  NOR2_X1 U10656 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n8237) );
  NOR2_X1 U10657 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8236) );
  NAND2_X1 U10658 ( .A1(n9896), .A2(n8245), .ZN(n8240) );
  NAND2_X1 U10659 ( .A1(n8240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8239) );
  MUX2_X1 U10660 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8239), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8241) );
  NAND2_X1 U10661 ( .A1(n8241), .A2(n8242), .ZN(n8968) );
  INV_X1 U10662 ( .A(n9055), .ZN(n8254) );
  NAND2_X1 U10663 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  NAND2_X1 U10664 ( .A1(n6742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8247) );
  MUX2_X1 U10665 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8247), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8250) );
  NAND2_X1 U10666 ( .A1(n8250), .A2(n8252), .ZN(n14432) );
  NAND2_X1 U10667 ( .A1(n8252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8251) );
  MUX2_X1 U10668 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8251), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8253) );
  NAND3_X2 U10669 ( .A1(n9339), .A2(n9058), .A3(n9054), .ZN(n9251) );
  NOR2_X4 U10670 ( .A1(n8254), .A2(n9251), .ZN(P1_U4016) );
  NOR2_X4 U10671 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8423) );
  NOR2_X1 U10672 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8261) );
  NAND4_X1 U10673 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8653), .ZN(n8755)
         );
  NAND3_X1 U10674 ( .A1(n8597), .A2(n8263), .A3(n8262), .ZN(n8264) );
  NOR2_X2 U10675 ( .A1(n8755), .A2(n8264), .ZN(n8267) );
  NAND2_X1 U10676 ( .A1(n8576), .A2(n8267), .ZN(n8416) );
  NAND2_X1 U10677 ( .A1(n8281), .A2(n8268), .ZN(n8283) );
  NAND2_X1 U10678 ( .A1(n8283), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8266) );
  MUX2_X1 U10679 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8266), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8272) );
  NAND3_X1 U10680 ( .A1(n8269), .A2(n8268), .A3(n8384), .ZN(n8270) );
  NOR2_X2 U10681 ( .A1(n8271), .A2(n8270), .ZN(n8274) );
  AND2_X2 U10682 ( .A1(n8274), .A2(n8273), .ZN(n8365) );
  NAND2_X1 U10683 ( .A1(n8275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8276) );
  MUX2_X1 U10684 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8276), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8277) );
  NAND2_X1 U10685 ( .A1(n6733), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8278) );
  MUX2_X1 U10686 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8278), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8279) );
  NAND2_X1 U10687 ( .A1(n8279), .A2(n8275), .ZN(n13817) );
  NOR2_X1 U10688 ( .A1(n13815), .A2(n13817), .ZN(n8280) );
  NAND2_X1 U10689 ( .A1(n8868), .A2(n8280), .ZN(n8888) );
  INV_X1 U10690 ( .A(n8281), .ZN(n8387) );
  NAND2_X1 U10691 ( .A1(n8387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8282) );
  MUX2_X1 U10692 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8282), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n8284) );
  INV_X1 U10693 ( .A(n11007), .ZN(n8285) );
  OAI21_X1 U10694 ( .B1(n11550), .B2(n9312), .A(n8291), .ZN(n8292) );
  AND2_X1 U10695 ( .A1(n8473), .A2(n8295), .ZN(n8296) );
  OAI21_X1 U10696 ( .B1(n8294), .B2(SI_3_), .A(n8295), .ZN(n8475) );
  AOI21_X2 U10697 ( .B1(n8474), .B2(n8296), .A(n7578), .ZN(n8498) );
  OAI21_X1 U10698 ( .B1(n8297), .B2(SI_4_), .A(n8299), .ZN(n8499) );
  INV_X1 U10699 ( .A(n8499), .ZN(n8298) );
  NAND2_X1 U10700 ( .A1(n8498), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U10701 ( .A1(n8300), .A2(n8299), .ZN(n8522) );
  MUX2_X1 U10702 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n11550), .Z(n8301) );
  NAND2_X1 U10703 ( .A1(n8301), .A2(SI_5_), .ZN(n8303) );
  OAI21_X1 U10704 ( .B1(n8301), .B2(SI_5_), .A(n8303), .ZN(n8302) );
  INV_X1 U10705 ( .A(n8302), .ZN(n8521) );
  NAND2_X1 U10706 ( .A1(n8522), .A2(n8521), .ZN(n8520) );
  MUX2_X1 U10707 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11550), .Z(n8304) );
  NAND2_X1 U10708 ( .A1(n8304), .A2(SI_6_), .ZN(n8306) );
  OAI21_X1 U10709 ( .B1(SI_6_), .B2(n8304), .A(n8306), .ZN(n8305) );
  INV_X1 U10710 ( .A(n8305), .ZN(n8538) );
  MUX2_X1 U10711 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11550), .Z(n8307) );
  NAND2_X1 U10712 ( .A1(n8307), .A2(SI_7_), .ZN(n8309) );
  OAI21_X1 U10713 ( .B1(n8307), .B2(SI_7_), .A(n8309), .ZN(n8308) );
  INV_X1 U10714 ( .A(n8308), .ZN(n8553) );
  MUX2_X1 U10715 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11550), .Z(n8310) );
  NAND2_X1 U10716 ( .A1(n8310), .A2(SI_8_), .ZN(n8312) );
  OAI21_X1 U10717 ( .B1(SI_8_), .B2(n8310), .A(n8312), .ZN(n8311) );
  INV_X1 U10718 ( .A(n8311), .ZN(n8572) );
  MUX2_X1 U10719 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6575), .Z(n8313) );
  NAND2_X1 U10720 ( .A1(n8313), .A2(SI_9_), .ZN(n8315) );
  OAI21_X1 U10721 ( .B1(n8313), .B2(SI_9_), .A(n8315), .ZN(n8314) );
  INV_X1 U10722 ( .A(n8314), .ZN(n8593) );
  INV_X1 U10723 ( .A(n8319), .ZN(n8317) );
  MUX2_X1 U10724 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6575), .Z(n8318) );
  INV_X1 U10725 ( .A(n8318), .ZN(n8316) );
  MUX2_X1 U10726 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11550), .Z(n8322) );
  XNOR2_X1 U10727 ( .A(n8322), .B(SI_11_), .ZN(n8632) );
  INV_X1 U10728 ( .A(n8322), .ZN(n8323) );
  NAND2_X1 U10729 ( .A1(n8323), .A2(n8956), .ZN(n8324) );
  MUX2_X1 U10730 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n6576), .Z(n8325) );
  XNOR2_X1 U10731 ( .A(n8325), .B(n8985), .ZN(n8651) );
  INV_X1 U10732 ( .A(n8325), .ZN(n8326) );
  NAND2_X1 U10733 ( .A1(n8326), .A2(n8985), .ZN(n8327) );
  MUX2_X1 U10734 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11550), .Z(n8329) );
  XNOR2_X1 U10735 ( .A(n8329), .B(n9107), .ZN(n8671) );
  INV_X1 U10736 ( .A(n8329), .ZN(n8330) );
  MUX2_X1 U10737 ( .A(n9860), .B(n9856), .S(n6575), .Z(n8711) );
  MUX2_X1 U10738 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6576), .Z(n8713) );
  NAND2_X1 U10739 ( .A1(n8713), .A2(SI_15_), .ZN(n8335) );
  OAI21_X1 U10740 ( .B1(n15462), .B2(n8711), .A(n8335), .ZN(n8331) );
  INV_X1 U10741 ( .A(n8331), .ZN(n8332) );
  INV_X1 U10742 ( .A(n8711), .ZN(n8333) );
  NOR2_X1 U10743 ( .A1(n8333), .A2(SI_14_), .ZN(n8336) );
  INV_X1 U10744 ( .A(SI_15_), .ZN(n9264) );
  INV_X1 U10745 ( .A(n8713), .ZN(n8334) );
  AOI22_X1 U10746 ( .A1(n8336), .A2(n8335), .B1(n9264), .B2(n8334), .ZN(n8735)
         );
  MUX2_X1 U10747 ( .A(n9629), .B(n9625), .S(n11550), .Z(n8339) );
  NAND2_X1 U10748 ( .A1(n8339), .A2(n8337), .ZN(n8338) );
  AND2_X1 U10749 ( .A1(n8735), .A2(n8338), .ZN(n8341) );
  INV_X1 U10750 ( .A(n8338), .ZN(n8340) );
  XNOR2_X1 U10751 ( .A(n8339), .B(SI_16_), .ZN(n8737) );
  MUX2_X1 U10752 ( .A(n9898), .B(n9899), .S(n11550), .Z(n8342) );
  XNOR2_X1 U10753 ( .A(n8342), .B(SI_17_), .ZN(n8754) );
  NAND2_X1 U10754 ( .A1(n8342), .A2(n9456), .ZN(n8343) );
  INV_X1 U10755 ( .A(SI_18_), .ZN(n9479) );
  MUX2_X1 U10756 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6576), .Z(n8414) );
  INV_X1 U10757 ( .A(n8414), .ZN(n8346) );
  MUX2_X1 U10758 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11550), .Z(n8347) );
  XNOR2_X1 U10759 ( .A(n8347), .B(SI_19_), .ZN(n8777) );
  INV_X1 U10760 ( .A(n8347), .ZN(n8348) );
  MUX2_X1 U10761 ( .A(n10748), .B(n10786), .S(n6576), .Z(n8787) );
  NAND2_X1 U10762 ( .A1(n8788), .A2(n8787), .ZN(n8802) );
  MUX2_X1 U10763 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6575), .Z(n8350) );
  NAND2_X1 U10764 ( .A1(n8350), .A2(SI_21_), .ZN(n8353) );
  OAI21_X1 U10765 ( .B1(SI_21_), .B2(n8350), .A(n8353), .ZN(n8803) );
  INV_X1 U10766 ( .A(n8803), .ZN(n8351) );
  XNOR2_X2 U10767 ( .A(n8355), .B(n8354), .ZN(n11411) );
  MUX2_X1 U10768 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n11550), .Z(n8820) );
  NAND2_X1 U10769 ( .A1(n8355), .A2(SI_22_), .ZN(n8356) );
  MUX2_X1 U10770 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11550), .Z(n8357) );
  NAND2_X1 U10771 ( .A1(n8357), .A2(SI_23_), .ZN(n8358) );
  OAI21_X1 U10772 ( .B1(SI_23_), .B2(n8357), .A(n8358), .ZN(n8837) );
  MUX2_X1 U10773 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6576), .Z(n8359) );
  NAND2_X1 U10774 ( .A1(n8359), .A2(SI_24_), .ZN(n11154) );
  OAI21_X1 U10775 ( .B1(SI_24_), .B2(n8359), .A(n11154), .ZN(n11151) );
  XNOR2_X1 U10776 ( .A(n11153), .B(n11151), .ZN(n11443) );
  AND2_X2 U10777 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  XNOR2_X2 U10778 ( .A(n8367), .B(n7434), .ZN(n9012) );
  NAND2_X2 U10779 ( .A1(n9010), .A2(n9012), .ZN(n8466) );
  NAND2_X1 U10780 ( .A1(n11443), .A2(n6581), .ZN(n8369) );
  INV_X1 U10781 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15323) );
  OR2_X1 U10782 ( .A1(n12348), .A2(n15323), .ZN(n8368) );
  NAND2_X1 U10783 ( .A1(n8388), .A2(n8370), .ZN(n8379) );
  INV_X1 U10784 ( .A(n8379), .ZN(n8372) );
  NAND2_X1 U10785 ( .A1(n8372), .A2(n8371), .ZN(n8381) );
  NAND2_X1 U10786 ( .A1(n8379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U10787 ( .A1(n8383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8385) );
  MUX2_X1 U10788 ( .A(n8385), .B(P2_IR_REG_31__SCAN_IN), .S(n8384), .Z(n8386)
         );
  INV_X1 U10789 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U10790 ( .A1(n9126), .A2(n12140), .ZN(n8426) );
  INV_X2 U10791 ( .A(n8426), .ZN(n8444) );
  INV_X2 U10792 ( .A(n8444), .ZN(n12513) );
  XNOR2_X1 U10793 ( .A(n13732), .B(n12513), .ZN(n8409) );
  NAND2_X1 U10794 ( .A1(n8546), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8562) );
  NOR2_X1 U10795 ( .A1(n8562), .A2(n8561), .ZN(n8580) );
  NAND2_X1 U10796 ( .A1(n8580), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10797 ( .A1(n8660), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8681) );
  INV_X1 U10798 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11090) );
  INV_X1 U10799 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8809) );
  INV_X1 U10800 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13282) );
  INV_X1 U10801 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10802 ( .A1(n8843), .A2(n8886), .ZN(n8393) );
  INV_X1 U10803 ( .A(n8892), .ZN(n8392) );
  NAND2_X1 U10804 ( .A1(n8393), .A2(n8392), .ZN(n13605) );
  XNOR2_X2 U10805 ( .A(n8398), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8400) );
  INV_X1 U10806 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10807 ( .A1(n8436), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10808 ( .A1(n8449), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8401) );
  OAI211_X1 U10809 ( .C1(n12357), .C2(n8403), .A(n8402), .B(n8401), .ZN(n8404)
         );
  INV_X1 U10810 ( .A(n8404), .ZN(n8405) );
  NAND2_X1 U10811 ( .A1(n8881), .A2(n12352), .ZN(n15033) );
  INV_X1 U10812 ( .A(n8879), .ZN(n8407) );
  AND2_X1 U10813 ( .A1(n13585), .A2(n8705), .ZN(n8408) );
  NAND2_X1 U10814 ( .A1(n8409), .A2(n8408), .ZN(n11631) );
  OAI21_X1 U10815 ( .B1(n8409), .B2(n8408), .A(n11631), .ZN(n8878) );
  AND2_X1 U10816 ( .A1(n8762), .A2(n8410), .ZN(n8411) );
  OR2_X1 U10817 ( .A1(n8411), .A2(n8781), .ZN(n13292) );
  AOI22_X1 U10818 ( .A1(n12319), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n8449), 
        .B2(P2_REG1_REG_18__SCAN_IN), .ZN(n8413) );
  INV_X1 U10819 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n11075) );
  OR2_X1 U10820 ( .A1(n6569), .A2(n11075), .ZN(n8412) );
  OAI211_X1 U10821 ( .C1(n13292), .C2(n8438), .A(n8413), .B(n8412), .ZN(n13505) );
  NAND2_X1 U10822 ( .A1(n13505), .A2(n8705), .ZN(n8772) );
  INV_X1 U10823 ( .A(n8772), .ZN(n8775) );
  NAND2_X1 U10824 ( .A1(n11302), .A2(n6581), .ZN(n8419) );
  NAND2_X1 U10825 ( .A1(n8416), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10826 ( .A(n8417), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U10827 ( .A1(n8778), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8484), 
        .B2(n13451), .ZN(n8418) );
  XNOR2_X1 U10828 ( .A(n13478), .B(n12513), .ZN(n8773) );
  INV_X1 U10829 ( .A(n8773), .ZN(n8774) );
  XNOR2_X1 U10830 ( .A(n8421), .B(n8420), .ZN(n9286) );
  NAND2_X1 U10831 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8422) );
  MUX2_X1 U10832 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8422), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8425) );
  INV_X1 U10833 ( .A(n8423), .ZN(n8424) );
  NAND2_X1 U10834 ( .A1(n8425), .A2(n8424), .ZN(n13325) );
  INV_X1 U10835 ( .A(n8434), .ZN(n8432) );
  INV_X1 U10836 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8427) );
  INV_X1 U10837 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13323) );
  INV_X1 U10838 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9493) );
  NOR2_X2 U10839 ( .A1(n6645), .A2(n7585), .ZN(n8429) );
  NAND3_X2 U10840 ( .A1(n8430), .A2(n8429), .A3(n8428), .ZN(n12147) );
  NAND2_X1 U10841 ( .A1(n12147), .A2(n8705), .ZN(n8433) );
  INV_X1 U10842 ( .A(n8433), .ZN(n8431) );
  NAND2_X1 U10843 ( .A1(n8432), .A2(n8431), .ZN(n8435) );
  NAND2_X1 U10844 ( .A1(n8434), .A2(n8433), .ZN(n8448) );
  NAND2_X1 U10845 ( .A1(n8435), .A2(n8448), .ZN(n9119) );
  INV_X1 U10846 ( .A(n9119), .ZN(n8447) );
  INV_X1 U10847 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9045) );
  INV_X1 U10848 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U10849 ( .A1(n8512), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10850 ( .A1(n11550), .A2(SI_0_), .ZN(n8443) );
  XNOR2_X1 U10851 ( .A(n8443), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13821) );
  NAND2_X1 U10852 ( .A1(n12144), .A2(n15035), .ZN(n12402) );
  OR2_X1 U10853 ( .A1(n12402), .A2(n6577), .ZN(n9144) );
  INV_X1 U10854 ( .A(n9120), .ZN(n8446) );
  NAND2_X1 U10855 ( .A1(n9117), .A2(n8448), .ZN(n9111) );
  NAND2_X1 U10856 ( .A1(n6580), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8455) );
  INV_X1 U10857 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9116) );
  OR2_X1 U10858 ( .A1(n8438), .A2(n9116), .ZN(n8454) );
  INV_X1 U10859 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9020) );
  INV_X1 U10860 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8450) );
  OR2_X1 U10861 ( .A1(n8451), .A2(n8450), .ZN(n8452) );
  NAND2_X1 U10862 ( .A1(n13322), .A2(n8705), .ZN(n8469) );
  INV_X1 U10863 ( .A(n8469), .ZN(n8468) );
  NOR2_X1 U10864 ( .A1(n8423), .A2(n13800), .ZN(n8456) );
  MUX2_X1 U10865 ( .A(n13800), .B(n8456), .S(P2_IR_REG_2__SCAN_IN), .Z(n8457)
         );
  INV_X1 U10866 ( .A(n8457), .ZN(n8459) );
  INV_X1 U10867 ( .A(n8481), .ZN(n8458) );
  NAND2_X1 U10868 ( .A1(n8459), .A2(n8458), .ZN(n14954) );
  OAI21_X1 U10869 ( .B1(n8461), .B2(n8460), .A(n8474), .ZN(n8905) );
  INV_X1 U10870 ( .A(n8905), .ZN(n8462) );
  NAND2_X1 U10871 ( .A1(n8468), .A2(n8467), .ZN(n8471) );
  NAND2_X1 U10872 ( .A1(n8470), .A2(n8469), .ZN(n8472) );
  NAND2_X1 U10873 ( .A1(n8474), .A2(n8473), .ZN(n8477) );
  INV_X1 U10874 ( .A(n8475), .ZN(n8476) );
  OR2_X1 U10875 ( .A1(n12348), .A2(n8915), .ZN(n8486) );
  NOR2_X1 U10876 ( .A1(n8481), .A2(n13800), .ZN(n8478) );
  MUX2_X1 U10877 ( .A(n13800), .B(n8478), .S(P2_IR_REG_3__SCAN_IN), .Z(n8479)
         );
  INV_X1 U10878 ( .A(n8479), .ZN(n8482) );
  NAND2_X1 U10879 ( .A1(n8481), .A2(n8480), .ZN(n8524) );
  NAND2_X1 U10880 ( .A1(n8482), .A2(n8524), .ZN(n13336) );
  INV_X1 U10881 ( .A(n13336), .ZN(n8483) );
  INV_X1 U10882 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10883 ( .A1(n6583), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8488) );
  INV_X1 U10884 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8995) );
  NOR2_X1 U10885 ( .A1(n8765), .A2(n8995), .ZN(n8492) );
  INV_X1 U10886 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U10887 ( .A1(n12322), .A2(n9785), .ZN(n8491) );
  NOR2_X1 U10888 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  NAND2_X1 U10889 ( .A1(n13321), .A2(n8705), .ZN(n8494) );
  XNOR2_X1 U10890 ( .A(n8495), .B(n8494), .ZN(n9151) );
  NAND2_X1 U10891 ( .A1(n8524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8497) );
  INV_X1 U10892 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8496) );
  XNOR2_X1 U10893 ( .A(n8497), .B(n8496), .ZN(n13352) );
  XNOR2_X1 U10894 ( .A(n8498), .B(n8499), .ZN(n9653) );
  OR2_X1 U10895 ( .A1(n12348), .A2(n8925), .ZN(n8500) );
  NAND2_X1 U10896 ( .A1(n8449), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8505) );
  INV_X1 U10897 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9821) );
  OR2_X1 U10898 ( .A1(n6569), .A2(n9821), .ZN(n8504) );
  XNOR2_X1 U10899 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9825) );
  OR2_X1 U10900 ( .A1(n8438), .A2(n9825), .ZN(n8503) );
  INV_X1 U10901 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8501) );
  OR2_X1 U10902 ( .A1(n8451), .A2(n8501), .ZN(n8502) );
  NAND2_X1 U10903 ( .A1(n13320), .A2(n8705), .ZN(n8506) );
  NAND2_X1 U10904 ( .A1(n8507), .A2(n8506), .ZN(n8511) );
  INV_X1 U10905 ( .A(n8506), .ZN(n8509) );
  INV_X1 U10906 ( .A(n8507), .ZN(n8508) );
  NAND2_X1 U10907 ( .A1(n8509), .A2(n8508), .ZN(n8510) );
  NAND2_X1 U10908 ( .A1(n8511), .A2(n8510), .ZN(n9268) );
  AOI21_X1 U10909 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8513) );
  NOR2_X1 U10910 ( .A1(n8513), .A2(n8546), .ZN(n13264) );
  NAND2_X1 U10911 ( .A1(n8512), .A2(n13264), .ZN(n8519) );
  INV_X1 U10912 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8514) );
  OR2_X1 U10913 ( .A1(n8765), .A2(n8514), .ZN(n8518) );
  INV_X1 U10914 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9025) );
  OR2_X1 U10915 ( .A1(n6569), .A2(n9025), .ZN(n8517) );
  INV_X1 U10916 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8515) );
  OR2_X1 U10917 ( .A1(n12357), .A2(n8515), .ZN(n8516) );
  AND4_X2 U10918 ( .A1(n8519), .A2(n8518), .A3(n8517), .A4(n8516), .ZN(n12181)
         );
  NOR2_X1 U10919 ( .A1(n12181), .A2(n6577), .ZN(n8532) );
  OR2_X1 U10920 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  NAND2_X1 U10921 ( .A1(n8520), .A2(n8523), .ZN(n9671) );
  OR2_X1 U10922 ( .A1(n9671), .A2(n8825), .ZN(n8531) );
  OR2_X1 U10923 ( .A1(n8524), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10924 ( .A1(n8527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8526) );
  MUX2_X1 U10925 ( .A(n8526), .B(P2_IR_REG_31__SCAN_IN), .S(n8525), .Z(n8529)
         );
  INV_X1 U10926 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10927 ( .A1(n8528), .A2(n8525), .ZN(n8556) );
  NAND2_X1 U10928 ( .A1(n8529), .A2(n8556), .ZN(n13365) );
  INV_X1 U10929 ( .A(n13365), .ZN(n9028) );
  AOI22_X1 U10930 ( .A1(n8778), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8484), .B2(
        n9028), .ZN(n8530) );
  XNOR2_X1 U10931 ( .A(n15084), .B(n8444), .ZN(n8533) );
  NAND2_X1 U10932 ( .A1(n8532), .A2(n8533), .ZN(n8536) );
  INV_X1 U10933 ( .A(n8532), .ZN(n8535) );
  INV_X1 U10934 ( .A(n8533), .ZN(n8534) );
  NAND2_X1 U10935 ( .A1(n8535), .A2(n8534), .ZN(n8537) );
  AND2_X1 U10936 ( .A1(n8536), .A2(n8537), .ZN(n13260) );
  NAND2_X1 U10937 ( .A1(n8541), .A2(n8540), .ZN(n9682) );
  OR2_X1 U10938 ( .A1(n9682), .A2(n8825), .ZN(n8544) );
  NAND2_X1 U10939 ( .A1(n8556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8542) );
  XNOR2_X1 U10940 ( .A(n8542), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9030) );
  AOI22_X1 U10941 ( .A1(n8778), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8484), .B2(
        n9030), .ZN(n8543) );
  AND2_X2 U10942 ( .A1(n8544), .A2(n8543), .ZN(n12188) );
  XNOR2_X1 U10943 ( .A(n12188), .B(n8444), .ZN(n8552) );
  NAND2_X1 U10944 ( .A1(n12319), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8550) );
  INV_X1 U10945 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8545) );
  OR2_X1 U10946 ( .A1(n8765), .A2(n8545), .ZN(n8549) );
  OAI21_X1 U10947 ( .B1(n8546), .B2(P2_REG3_REG_6__SCAN_IN), .A(n8562), .ZN(
        n9755) );
  OR2_X1 U10948 ( .A1(n6583), .A2(n9755), .ZN(n8548) );
  INV_X1 U10949 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9752) );
  OR2_X1 U10950 ( .A1(n6569), .A2(n9752), .ZN(n8547) );
  NOR2_X1 U10951 ( .A1(n12187), .A2(n6577), .ZN(n8551) );
  XNOR2_X1 U10952 ( .A(n8552), .B(n8551), .ZN(n9458) );
  OR2_X1 U10953 ( .A1(n10116), .A2(n8825), .ZN(n8559) );
  OAI21_X1 U10954 ( .B1(n8556), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8557) );
  XNOR2_X1 U10955 ( .A(n8557), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U10956 ( .A1(n8778), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8484), .B2(
        n13380), .ZN(n8558) );
  XNOR2_X1 U10957 ( .A(n15098), .B(n12513), .ZN(n8568) );
  NAND2_X1 U10958 ( .A1(n12319), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8567) );
  INV_X1 U10959 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8560) );
  OR2_X1 U10960 ( .A1(n8765), .A2(n8560), .ZN(n8566) );
  AND2_X1 U10961 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  OR2_X1 U10962 ( .A1(n8563), .A2(n8580), .ZN(n9538) );
  OR2_X1 U10963 ( .A1(n6583), .A2(n9538), .ZN(n8565) );
  INV_X1 U10964 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9539) );
  OR2_X1 U10965 ( .A1(n6568), .A2(n9539), .ZN(n8564) );
  NOR2_X1 U10966 ( .A1(n12192), .A2(n6577), .ZN(n8569) );
  XNOR2_X1 U10967 ( .A(n8568), .B(n8569), .ZN(n9482) );
  INV_X1 U10968 ( .A(n8568), .ZN(n8570) );
  NAND2_X1 U10969 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  OR2_X1 U10970 ( .A1(n8573), .A2(n8572), .ZN(n8574) );
  OR2_X1 U10971 ( .A1(n8576), .A2(n13800), .ZN(n8577) );
  XNOR2_X1 U10972 ( .A(n8577), .B(P2_IR_REG_8__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U10973 ( .A1(n8778), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8484), .B2(
        n13394), .ZN(n8578) );
  XNOR2_X1 U10974 ( .A(n12196), .B(n12513), .ZN(n8586) );
  NAND2_X1 U10975 ( .A1(n12319), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8585) );
  INV_X1 U10976 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n8579) );
  OR2_X1 U10977 ( .A1(n8765), .A2(n8579), .ZN(n8584) );
  OR2_X1 U10978 ( .A1(n8580), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10979 ( .A1(n8604), .A2(n8581), .ZN(n9946) );
  OR2_X1 U10980 ( .A1(n8438), .A2(n9946), .ZN(n8583) );
  INV_X1 U10981 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9807) );
  OR2_X1 U10982 ( .A1(n6569), .A2(n9807), .ZN(n8582) );
  OR2_X1 U10983 ( .A1(n12195), .A2(n6577), .ZN(n8587) );
  NAND2_X1 U10984 ( .A1(n8586), .A2(n8587), .ZN(n8592) );
  INV_X1 U10985 ( .A(n8586), .ZN(n8589) );
  INV_X1 U10986 ( .A(n8587), .ZN(n8588) );
  NAND2_X1 U10987 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  NAND2_X1 U10988 ( .A1(n8592), .A2(n8590), .ZN(n9945) );
  NAND2_X1 U10989 ( .A1(n9943), .A2(n8592), .ZN(n10171) );
  OR2_X1 U10990 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U10991 ( .A1(n8596), .A2(n8595), .ZN(n10136) );
  OR2_X1 U10992 ( .A1(n10136), .A2(n8825), .ZN(n8602) );
  NAND2_X1 U10993 ( .A1(n8576), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10994 ( .A1(n8599), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8598) );
  MUX2_X1 U10995 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8598), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8600) );
  AND2_X1 U10996 ( .A1(n8600), .A2(n8756), .ZN(n9036) );
  AOI22_X1 U10997 ( .A1(n8778), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8484), .B2(
        n9036), .ZN(n8601) );
  XNOR2_X1 U10998 ( .A(n15111), .B(n8444), .ZN(n8611) );
  NAND2_X1 U10999 ( .A1(n8436), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8610) );
  INV_X1 U11000 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9431) );
  OR2_X1 U11001 ( .A1(n8765), .A2(n9431), .ZN(n8609) );
  NAND2_X1 U11002 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  NAND2_X1 U11003 ( .A1(n8623), .A2(n8605), .ZN(n10175) );
  OR2_X1 U11004 ( .A1(n8438), .A2(n10175), .ZN(n8608) );
  INV_X1 U11005 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8606) );
  OR2_X1 U11006 ( .A1(n8451), .A2(n8606), .ZN(n8607) );
  NAND4_X1 U11007 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n13315) );
  NAND2_X1 U11008 ( .A1(n13315), .A2(n8705), .ZN(n8612) );
  NAND2_X1 U11009 ( .A1(n8611), .A2(n8612), .ZN(n8616) );
  INV_X1 U11010 ( .A(n8611), .ZN(n8614) );
  INV_X1 U11011 ( .A(n8612), .ZN(n8613) );
  NAND2_X1 U11012 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  AND2_X1 U11013 ( .A1(n8616), .A2(n8615), .ZN(n10173) );
  NAND2_X1 U11014 ( .A1(n10171), .A2(n10173), .ZN(n10172) );
  NAND2_X1 U11015 ( .A1(n10172), .A2(n8616), .ZN(n10245) );
  NAND2_X1 U11016 ( .A1(n8617), .A2(n7544), .ZN(n8618) );
  NAND2_X1 U11017 ( .A1(n8619), .A2(n8618), .ZN(n10409) );
  OR2_X1 U11018 ( .A1(n10409), .A2(n8825), .ZN(n8622) );
  NAND2_X1 U11019 ( .A1(n8756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8620) );
  XNOR2_X1 U11020 ( .A(n8620), .B(P2_IR_REG_10__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U11021 ( .A1(n8778), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8484), 
        .B2(n13411), .ZN(n8621) );
  XNOR2_X1 U11022 ( .A(n15119), .B(n8444), .ZN(n8630) );
  NAND2_X1 U11023 ( .A1(n12319), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8628) );
  INV_X1 U11024 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11025 ( .A1(n8765), .A2(n9435), .ZN(n8627) );
  NAND2_X1 U11026 ( .A1(n8623), .A2(n15436), .ZN(n8624) );
  NAND2_X1 U11027 ( .A1(n8637), .A2(n8624), .ZN(n10264) );
  OR2_X1 U11028 ( .A1(n6583), .A2(n10264), .ZN(n8626) );
  INV_X1 U11029 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n13412) );
  OR2_X1 U11030 ( .A1(n6568), .A2(n13412), .ZN(n8625) );
  NAND4_X1 U11031 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n13314) );
  NAND2_X1 U11032 ( .A1(n13314), .A2(n8705), .ZN(n8629) );
  XNOR2_X1 U11033 ( .A(n8630), .B(n8629), .ZN(n10246) );
  NAND2_X1 U11034 ( .A1(n10438), .A2(n6581), .ZN(n8635) );
  NOR2_X1 U11035 ( .A1(n8756), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n8654) );
  OR2_X1 U11036 ( .A1(n8654), .A2(n13800), .ZN(n8633) );
  XNOR2_X1 U11037 ( .A(n8633), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14981) );
  AOI22_X1 U11038 ( .A1(n8778), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8484), 
        .B2(n14981), .ZN(n8634) );
  XNOR2_X1 U11039 ( .A(n12215), .B(n12513), .ZN(n8646) );
  NAND2_X1 U11040 ( .A1(n8436), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8640) );
  AND2_X1 U11041 ( .A1(n8637), .A2(n8636), .ZN(n8638) );
  OR2_X1 U11042 ( .A1(n8638), .A2(n8660), .ZN(n10532) );
  OR2_X1 U11043 ( .A1(n8438), .A2(n10532), .ZN(n8639) );
  NAND2_X1 U11044 ( .A1(n8640), .A2(n8639), .ZN(n8645) );
  INV_X1 U11045 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8641) );
  NOR2_X1 U11046 ( .A1(n12357), .A2(n8641), .ZN(n8644) );
  INV_X1 U11047 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8642) );
  NOR2_X1 U11048 ( .A1(n8765), .A2(n8642), .ZN(n8643) );
  NAND2_X1 U11049 ( .A1(n13313), .A2(n8705), .ZN(n8647) );
  NAND2_X1 U11050 ( .A1(n8646), .A2(n8647), .ZN(n10386) );
  NAND2_X1 U11051 ( .A1(n10387), .A2(n10386), .ZN(n8650) );
  INV_X1 U11052 ( .A(n8646), .ZN(n8649) );
  INV_X1 U11053 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U11054 ( .A1(n8649), .A2(n8648), .ZN(n10385) );
  NAND2_X1 U11055 ( .A1(n8650), .A2(n10385), .ZN(n14937) );
  INV_X1 U11056 ( .A(n14937), .ZN(n8667) );
  NAND2_X1 U11057 ( .A1(n10568), .A2(n6581), .ZN(n8657) );
  NAND2_X1 U11058 ( .A1(n8654), .A2(n8653), .ZN(n8673) );
  NAND2_X1 U11059 ( .A1(n8673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8655) );
  XNOR2_X1 U11060 ( .A(n8655), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9437) );
  AOI22_X1 U11061 ( .A1(n8778), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8484), 
        .B2(n9437), .ZN(n8656) );
  XNOR2_X1 U11062 ( .A(n14944), .B(n8444), .ZN(n8669) );
  NAND2_X1 U11063 ( .A1(n12319), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8659) );
  INV_X1 U11064 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10692) );
  OR2_X1 U11065 ( .A1(n6569), .A2(n10692), .ZN(n8658) );
  NAND2_X1 U11066 ( .A1(n8659), .A2(n8658), .ZN(n8665) );
  OR2_X1 U11067 ( .A1(n8660), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11068 ( .A1(n8681), .A2(n8661), .ZN(n14946) );
  NOR2_X1 U11069 ( .A1(n6583), .A2(n14946), .ZN(n8664) );
  INV_X1 U11070 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U11071 ( .A1(n8765), .A2(n8662), .ZN(n8663) );
  NAND2_X1 U11072 ( .A1(n13312), .A2(n8705), .ZN(n8668) );
  XNOR2_X1 U11073 ( .A(n8669), .B(n8668), .ZN(n14938) );
  NAND2_X1 U11074 ( .A1(n8667), .A2(n8666), .ZN(n14935) );
  NAND2_X1 U11075 ( .A1(n8669), .A2(n8668), .ZN(n8670) );
  NAND2_X1 U11076 ( .A1(n10573), .A2(n6581), .ZN(n8679) );
  OR2_X1 U11077 ( .A1(n8673), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11078 ( .A1(n8675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8674) );
  MUX2_X1 U11079 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8674), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8677) );
  INV_X1 U11080 ( .A(n8717), .ZN(n8676) );
  AOI22_X1 U11081 ( .A1(n8778), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8484), 
        .B2(n15011), .ZN(n8678) );
  XNOR2_X1 U11082 ( .A(n14634), .B(n8444), .ZN(n8688) );
  NAND2_X1 U11083 ( .A1(n8449), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11084 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  NAND2_X1 U11085 ( .A1(n8699), .A2(n8682), .ZN(n10802) );
  OR2_X1 U11086 ( .A1(n8438), .A2(n10802), .ZN(n8686) );
  INV_X1 U11087 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10803) );
  OR2_X1 U11088 ( .A1(n6569), .A2(n10803), .ZN(n8685) );
  INV_X1 U11089 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8683) );
  OR2_X1 U11090 ( .A1(n8451), .A2(n8683), .ZN(n8684) );
  NOR2_X1 U11091 ( .A1(n14931), .A2(n6577), .ZN(n8689) );
  NAND2_X1 U11092 ( .A1(n8688), .A2(n8689), .ZN(n8694) );
  INV_X1 U11093 ( .A(n8688), .ZN(n8691) );
  INV_X1 U11094 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U11095 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NAND2_X1 U11096 ( .A1(n8694), .A2(n8692), .ZN(n10626) );
  NAND2_X1 U11097 ( .A1(n11280), .A2(n6581), .ZN(n8697) );
  OR2_X1 U11098 ( .A1(n8717), .A2(n13800), .ZN(n8695) );
  XNOR2_X1 U11099 ( .A(n8695), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U11100 ( .A1(n8778), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10762), 
        .B2(n8484), .ZN(n8696) );
  XNOR2_X1 U11101 ( .A(n12234), .B(n12513), .ZN(n8708) );
  NAND2_X1 U11102 ( .A1(n8449), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8704) );
  INV_X1 U11103 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8698) );
  OR2_X1 U11104 ( .A1(n12357), .A2(n8698), .ZN(n8703) );
  AND2_X1 U11105 ( .A1(n8699), .A2(n10818), .ZN(n8700) );
  OR2_X1 U11106 ( .A1(n8700), .A2(n8725), .ZN(n10864) );
  OR2_X1 U11107 ( .A1(n8438), .A2(n10864), .ZN(n8702) );
  INV_X1 U11108 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10865) );
  OR2_X1 U11109 ( .A1(n6568), .A2(n10865), .ZN(n8701) );
  NOR2_X1 U11110 ( .A1(n12233), .A2(n6577), .ZN(n8706) );
  XNOR2_X1 U11111 ( .A(n8708), .B(n8706), .ZN(n10814) );
  INV_X1 U11112 ( .A(n8706), .ZN(n8707) );
  AND2_X1 U11113 ( .A1(n8709), .A2(n15462), .ZN(n8710) );
  XNOR2_X1 U11114 ( .A(n8713), .B(SI_15_), .ZN(n8714) );
  INV_X1 U11115 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8716) );
  AOI21_X1 U11116 ( .B1(n8717), .B2(n8716), .A(n13800), .ZN(n8718) );
  NAND2_X1 U11117 ( .A1(n8718), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8721) );
  INV_X1 U11118 ( .A(n8718), .ZN(n8720) );
  INV_X1 U11119 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11120 ( .A1(n8720), .A2(n8719), .ZN(n8739) );
  AND2_X1 U11121 ( .A1(n8721), .A2(n8739), .ZN(n10766) );
  NAND2_X1 U11122 ( .A1(n10766), .A2(n8484), .ZN(n8722) );
  OAI21_X1 U11123 ( .B1(n12348), .B2(n9938), .A(n8722), .ZN(n8723) );
  AOI21_X1 U11124 ( .B1(n11285), .B2(n6581), .A(n8723), .ZN(n8724) );
  XNOR2_X1 U11125 ( .A(n13778), .B(n12513), .ZN(n8731) );
  XNOR2_X1 U11126 ( .A(n8733), .B(n8731), .ZN(n10933) );
  NAND2_X1 U11127 ( .A1(n12319), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8730) );
  INV_X1 U11128 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10754) );
  OR2_X1 U11129 ( .A1(n8765), .A2(n10754), .ZN(n8729) );
  NOR2_X1 U11130 ( .A1(n8725), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8726) );
  OR2_X1 U11131 ( .A1(n8743), .A2(n8726), .ZN(n10934) );
  OR2_X1 U11132 ( .A1(n10934), .A2(n6583), .ZN(n8728) );
  INV_X1 U11133 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10910) );
  OR2_X1 U11134 ( .A1(n6568), .A2(n10910), .ZN(n8727) );
  NOR2_X1 U11135 ( .A1(n12239), .A2(n6577), .ZN(n10932) );
  INV_X1 U11136 ( .A(n8731), .ZN(n8732) );
  OR2_X2 U11137 ( .A1(n8733), .A2(n8732), .ZN(n8734) );
  NAND2_X1 U11138 ( .A1(n8736), .A2(n8735), .ZN(n8738) );
  XNOR2_X1 U11139 ( .A(n8738), .B(n8737), .ZN(n11331) );
  NAND2_X1 U11140 ( .A1(n11331), .A2(n6581), .ZN(n8742) );
  NAND2_X1 U11141 ( .A1(n8739), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8740) );
  XNOR2_X1 U11142 ( .A(n8740), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U11143 ( .A1(n15024), .A2(n8484), .B1(n8778), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8741) );
  XNOR2_X1 U11144 ( .A(n13773), .B(n12513), .ZN(n8752) );
  OR2_X1 U11145 ( .A1(n8743), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8744) );
  AND2_X1 U11146 ( .A1(n8760), .A2(n8744), .ZN(n11046) );
  NAND2_X1 U11147 ( .A1(n8512), .A2(n11046), .ZN(n8750) );
  INV_X1 U11148 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8745) );
  OR2_X1 U11149 ( .A1(n8451), .A2(n8745), .ZN(n8749) );
  INV_X1 U11150 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8746) );
  OR2_X1 U11151 ( .A1(n8765), .A2(n8746), .ZN(n8748) );
  INV_X1 U11152 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11020) );
  OR2_X1 U11153 ( .A1(n6568), .A2(n11020), .ZN(n8747) );
  NOR2_X1 U11154 ( .A1(n12249), .A2(n6577), .ZN(n8751) );
  XNOR2_X1 U11155 ( .A(n8752), .B(n8751), .ZN(n11042) );
  NOR2_X1 U11156 ( .A1(n8752), .A2(n8751), .ZN(n11085) );
  XNOR2_X1 U11157 ( .A(n8753), .B(n8754), .ZN(n11312) );
  NAND2_X1 U11158 ( .A1(n11312), .A2(n6581), .ZN(n8759) );
  OAI21_X1 U11159 ( .B1(n8756), .B2(n8755), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8757) );
  XNOR2_X1 U11160 ( .A(n8757), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U11161 ( .A1(n8778), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8484), 
        .B2(n13438), .ZN(n8758) );
  XNOR2_X1 U11162 ( .A(n13768), .B(n12513), .ZN(n8770) );
  NAND2_X1 U11163 ( .A1(n8760), .A2(n11090), .ZN(n8761) );
  NAND2_X1 U11164 ( .A1(n8762), .A2(n8761), .ZN(n11089) );
  INV_X1 U11165 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11053) );
  OAI22_X1 U11166 ( .A1(n11089), .A2(n8438), .B1(n6569), .B2(n11053), .ZN(
        n8767) );
  INV_X1 U11167 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11168 ( .A1(n12319), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8763) );
  OAI21_X1 U11169 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8766) );
  NAND2_X1 U11170 ( .A1(n13308), .A2(n8705), .ZN(n8768) );
  XNOR2_X1 U11171 ( .A(n8770), .B(n8768), .ZN(n11084) );
  INV_X1 U11172 ( .A(n8768), .ZN(n8769) );
  XNOR2_X1 U11173 ( .A(n8773), .B(n8772), .ZN(n13290) );
  XNOR2_X1 U11174 ( .A(n8776), .B(n8777), .ZN(n11337) );
  NAND2_X1 U11175 ( .A1(n11337), .A2(n6581), .ZN(n8780) );
  AOI22_X1 U11176 ( .A1(n8778), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8484), 
        .B2(n12436), .ZN(n8779) );
  XNOR2_X1 U11177 ( .A(n13757), .B(n12513), .ZN(n8786) );
  NOR2_X1 U11178 ( .A1(n8781), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8782) );
  OR2_X1 U11179 ( .A1(n8791), .A2(n8782), .ZN(n13687) );
  AOI22_X1 U11180 ( .A1(n8449), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8436), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11181 ( .A1(n12319), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8783) );
  OAI211_X1 U11182 ( .C1(n13687), .C2(n6583), .A(n8784), .B(n8783), .ZN(n13668) );
  AND2_X1 U11183 ( .A1(n13668), .A2(n8705), .ZN(n8785) );
  NAND2_X1 U11184 ( .A1(n8786), .A2(n8785), .ZN(n13243) );
  XNOR2_X1 U11185 ( .A(n8788), .B(n8787), .ZN(n11375) );
  NAND2_X1 U11186 ( .A1(n11375), .A2(n6581), .ZN(n8790) );
  OR2_X1 U11187 ( .A1(n12348), .A2(n10786), .ZN(n8789) );
  XNOR2_X1 U11188 ( .A(n13752), .B(n8444), .ZN(n8800) );
  OR2_X1 U11189 ( .A1(n8791), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8792) );
  AND2_X1 U11190 ( .A1(n8810), .A2(n8792), .ZN(n13674) );
  NAND2_X1 U11191 ( .A1(n13674), .A2(n8512), .ZN(n8798) );
  INV_X1 U11192 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11193 ( .A1(n8436), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11194 ( .A1(n8449), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8793) );
  OAI211_X1 U11195 ( .C1(n12357), .C2(n8795), .A(n8794), .B(n8793), .ZN(n8796)
         );
  INV_X1 U11196 ( .A(n8796), .ZN(n8797) );
  NAND2_X1 U11197 ( .A1(n8798), .A2(n8797), .ZN(n13509) );
  NAND2_X1 U11198 ( .A1(n13509), .A2(n8705), .ZN(n8799) );
  NOR2_X1 U11199 ( .A1(n8800), .A2(n8799), .ZN(n13269) );
  NAND2_X1 U11200 ( .A1(n8802), .A2(n8801), .ZN(n8804) );
  NAND2_X1 U11201 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  NAND2_X1 U11202 ( .A1(n8806), .A2(n8805), .ZN(n11380) );
  OR2_X1 U11203 ( .A1(n11380), .A2(n8825), .ZN(n8808) );
  INV_X1 U11204 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11150) );
  OR2_X1 U11205 ( .A1(n12348), .A2(n11150), .ZN(n8807) );
  XNOR2_X1 U11206 ( .A(n13747), .B(n12513), .ZN(n8819) );
  NAND2_X1 U11207 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND2_X1 U11208 ( .A1(n8828), .A2(n8811), .ZN(n13652) );
  OR2_X1 U11209 ( .A1(n13652), .A2(n8438), .ZN(n8817) );
  INV_X1 U11210 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8814) );
  NAND2_X1 U11211 ( .A1(n12319), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8813) );
  NAND2_X1 U11212 ( .A1(n8449), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8812) );
  OAI211_X1 U11213 ( .C1(n8814), .C2(n6568), .A(n8813), .B(n8812), .ZN(n8815)
         );
  INV_X1 U11214 ( .A(n8815), .ZN(n8816) );
  NOR2_X1 U11215 ( .A1(n13480), .A2(n6577), .ZN(n8818) );
  XNOR2_X1 U11216 ( .A(n8819), .B(n8818), .ZN(n13254) );
  INV_X1 U11217 ( .A(n11411), .ZN(n8822) );
  INV_X1 U11218 ( .A(n8820), .ZN(n8821) );
  NAND2_X1 U11219 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U11220 ( .A1(n8824), .A2(n8823), .ZN(n10880) );
  INV_X1 U11221 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15495) );
  OR2_X1 U11222 ( .A1(n12348), .A2(n15495), .ZN(n8826) );
  XNOR2_X1 U11223 ( .A(n8834), .B(n6628), .ZN(n13280) );
  AND2_X1 U11224 ( .A1(n8828), .A2(n13282), .ZN(n8829) );
  OR2_X1 U11225 ( .A1(n8829), .A2(n8841), .ZN(n13283) );
  INV_X1 U11226 ( .A(n13283), .ZN(n13640) );
  INV_X1 U11227 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11228 ( .A1(n8449), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11229 ( .A1(n8436), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8830) );
  OAI211_X1 U11230 ( .C1(n12357), .C2(n8832), .A(n8831), .B(n8830), .ZN(n8833)
         );
  AOI21_X1 U11231 ( .B1(n13640), .B2(n8512), .A(n8833), .ZN(n13250) );
  INV_X1 U11232 ( .A(n13250), .ZN(n13514) );
  NAND2_X1 U11233 ( .A1(n13514), .A2(n8705), .ZN(n13279) );
  NAND2_X1 U11234 ( .A1(n13280), .A2(n13279), .ZN(n13278) );
  INV_X1 U11235 ( .A(n8834), .ZN(n8835) );
  NAND2_X1 U11236 ( .A1(n11428), .A2(n6581), .ZN(n8840) );
  OR2_X1 U11237 ( .A1(n12348), .A2(n11009), .ZN(n8839) );
  AND2_X2 U11238 ( .A1(n8840), .A2(n8839), .ZN(n13624) );
  XNOR2_X1 U11239 ( .A(n13624), .B(n8444), .ZN(n8850) );
  OR2_X1 U11240 ( .A1(n8841), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8842) );
  NAND2_X1 U11241 ( .A1(n8843), .A2(n8842), .ZN(n13621) );
  OR2_X1 U11242 ( .A1(n13621), .A2(n6583), .ZN(n8849) );
  INV_X1 U11243 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8846) );
  NAND2_X1 U11244 ( .A1(n8449), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U11245 ( .A1(n8436), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8844) );
  OAI211_X1 U11246 ( .C1(n8846), .C2(n12357), .A(n8845), .B(n8844), .ZN(n8847)
         );
  INV_X1 U11247 ( .A(n8847), .ZN(n8848) );
  NAND2_X1 U11248 ( .A1(n13483), .A2(n8705), .ZN(n13237) );
  INV_X1 U11249 ( .A(n8850), .ZN(n8851) );
  NAND2_X1 U11250 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  INV_X1 U11251 ( .A(P2_B_REG_SCAN_IN), .ZN(n13465) );
  XNOR2_X1 U11252 ( .A(n8868), .B(n13465), .ZN(n8854) );
  NAND2_X1 U11253 ( .A1(n8854), .A2(n13817), .ZN(n8856) );
  INV_X1 U11254 ( .A(n13815), .ZN(n8855) );
  NOR2_X1 U11255 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n8860) );
  NOR4_X1 U11256 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8859) );
  NOR4_X1 U11257 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8858) );
  NOR4_X1 U11258 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8857) );
  AND4_X1 U11259 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n8866)
         );
  NOR4_X1 U11260 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8864) );
  NOR4_X1 U11261 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8863) );
  NOR4_X1 U11262 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8862) );
  NOR4_X1 U11263 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8861) );
  AND4_X1 U11264 ( .A1(n8864), .A2(n8863), .A3(n8862), .A4(n8861), .ZN(n8865)
         );
  NAND2_X1 U11265 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  AND2_X1 U11266 ( .A1(n15048), .A2(n8867), .ZN(n9138) );
  INV_X1 U11267 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U11268 ( .A1(n15048), .A2(n15052), .ZN(n8870) );
  INV_X1 U11269 ( .A(n8868), .ZN(n11061) );
  NAND2_X1 U11270 ( .A1(n11061), .A2(n13815), .ZN(n8869) );
  OR2_X1 U11271 ( .A1(n9138), .A2(n15053), .ZN(n8887) );
  INV_X1 U11272 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U11273 ( .A1(n15048), .A2(n15055), .ZN(n8872) );
  NAND2_X1 U11274 ( .A1(n13815), .A2(n13817), .ZN(n8871) );
  NAND2_X1 U11275 ( .A1(n8872), .A2(n8871), .ZN(n9141) );
  INV_X1 U11276 ( .A(n15056), .ZN(n15051) );
  OR2_X1 U11277 ( .A1(n9141), .A2(n15051), .ZN(n15054) );
  NOR2_X1 U11278 ( .A1(n8887), .A2(n15054), .ZN(n8884) );
  INV_X1 U11279 ( .A(n9006), .ZN(n8874) );
  NAND2_X1 U11280 ( .A1(n8879), .A2(n13459), .ZN(n12389) );
  AND2_X1 U11281 ( .A1(n8874), .A2(n15097), .ZN(n8875) );
  INV_X1 U11282 ( .A(n11632), .ZN(n8877) );
  AOI211_X1 U11283 ( .C1(n8878), .C2(n8876), .A(n14939), .B(n8877), .ZN(n8901)
         );
  INV_X1 U11284 ( .A(n13732), .ZN(n13608) );
  NOR2_X1 U11285 ( .A1(n15033), .A2(n8879), .ZN(n9492) );
  NAND2_X1 U11286 ( .A1(n8884), .A2(n9492), .ZN(n8883) );
  NAND2_X2 U11287 ( .A1(n8880), .A2(n12352), .ZN(n12137) );
  NAND2_X1 U11288 ( .A1(n15088), .A2(n8881), .ZN(n9139) );
  INV_X1 U11289 ( .A(n9139), .ZN(n8882) );
  INV_X1 U11290 ( .A(n14943), .ZN(n13297) );
  NOR2_X1 U11291 ( .A1(n13608), .A2(n13297), .ZN(n8900) );
  NAND2_X1 U11292 ( .A1(n8884), .A2(n12457), .ZN(n13238) );
  INV_X1 U11293 ( .A(n9012), .ZN(n8885) );
  OR2_X1 U11294 ( .A1(n13238), .A2(n13595), .ZN(n14933) );
  OAI22_X1 U11295 ( .A1(n13596), .A2(n14933), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8886), .ZN(n8899) );
  OAI21_X1 U11296 ( .B1(n8887), .B2(n9141), .A(n9139), .ZN(n8890) );
  NAND2_X1 U11297 ( .A1(n9006), .A2(n12389), .ZN(n9136) );
  AND3_X1 U11298 ( .A1(n9136), .A2(n8888), .A3(n11007), .ZN(n8889) );
  NAND2_X1 U11299 ( .A1(n8890), .A2(n8889), .ZN(n9109) );
  NAND2_X1 U11300 ( .A1(n8449), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8897) );
  INV_X1 U11301 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8891) );
  OR2_X1 U11302 ( .A1(n6569), .A2(n8891), .ZN(n8896) );
  INV_X1 U11303 ( .A(n11638), .ZN(n11639) );
  OAI21_X1 U11304 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n8892), .A(n11639), .ZN(
        n13579) );
  OR2_X1 U11305 ( .A1(n6583), .A2(n13579), .ZN(n8895) );
  INV_X1 U11306 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8893) );
  OR2_X1 U11307 ( .A1(n8451), .A2(n8893), .ZN(n8894) );
  NAND4_X1 U11308 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n13570) );
  NAND2_X1 U11309 ( .A1(n9006), .A2(n9012), .ZN(n15039) );
  OAI22_X1 U11310 ( .A1(n13605), .A2(n14947), .B1(n13594), .B2(n14932), .ZN(
        n8898) );
  OR4_X1 U11311 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(P2_U3201) );
  OR2_X1 U11312 ( .A1(n8902), .A2(n8966), .ZN(n8904) );
  NAND2_X1 U11313 ( .A1(n7614), .A2(P1_U3086), .ZN(n14434) );
  AND2_X1 U11314 ( .A1(n6576), .A2(P1_U3086), .ZN(n14423) );
  INV_X2 U11315 ( .A(n14423), .ZN(n14436) );
  OAI222_X1 U11316 ( .A1(P1_U3086), .A2(n13998), .B1(n14434), .B2(n8905), .C1(
        n9312), .C2(n14436), .ZN(P1_U3353) );
  OR2_X1 U11317 ( .A1(n8921), .A2(n8966), .ZN(n8906) );
  XNOR2_X1 U11318 ( .A(n8906), .B(n8920), .ZN(n14012) );
  OAI222_X1 U11319 ( .A1(n14436), .A2(n9331), .B1(n14434), .B2(n9330), .C1(
        P1_U3086), .C2(n14012), .ZN(P1_U3352) );
  INV_X1 U11320 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8908) );
  NAND2_X1 U11321 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8907) );
  INV_X1 U11322 ( .A(n14434), .ZN(n11010) );
  INV_X1 U11323 ( .A(n11010), .ZN(n14428) );
  OAI222_X1 U11324 ( .A1(P1_U3086), .A2(n6574), .B1(n14428), .B2(n9286), .C1(
        n8287), .C2(n14436), .ZN(P1_U3354) );
  INV_X1 U11325 ( .A(n9593), .ZN(n9581) );
  AOI222_X1 U11326 ( .A1(n8909), .A2(n13221), .B1(n9581), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n9400), .ZN(n8910) );
  INV_X1 U11327 ( .A(n8910), .ZN(P3_U3292) );
  INV_X1 U11328 ( .A(n9598), .ZN(n9622) );
  AOI222_X1 U11329 ( .A1(n8911), .A2(n13221), .B1(n9622), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n9400), .ZN(n8912) );
  INV_X1 U11330 ( .A(n8912), .ZN(P3_U3291) );
  AOI222_X1 U11331 ( .A1(n8913), .A2(n13221), .B1(n9991), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n9400), .ZN(n8914) );
  INV_X1 U11332 ( .A(n8914), .ZN(P3_U3290) );
  AND2_X1 U11333 ( .A1(n7614), .A2(P2_U3088), .ZN(n13808) );
  INV_X2 U11334 ( .A(n13808), .ZN(n13820) );
  AND2_X1 U11335 ( .A1(n11550), .A2(P2_U3088), .ZN(n11006) );
  OAI222_X1 U11336 ( .A1(n13820), .A2(n8915), .B1(n13818), .B2(n9330), .C1(
        P2_U3088), .C2(n13336), .ZN(P2_U3324) );
  INV_X2 U11337 ( .A(n11006), .ZN(n13818) );
  OAI222_X1 U11338 ( .A1(P2_U3088), .A2(n13325), .B1(n13820), .B2(n8916), .C1(
        n13818), .C2(n9286), .ZN(P2_U3326) );
  OAI222_X1 U11339 ( .A1(P2_U3088), .A2(n14954), .B1(n13820), .B2(n8917), .C1(
        n13818), .C2(n8905), .ZN(P2_U3325) );
  AOI222_X1 U11340 ( .A1(n8918), .A2(n13221), .B1(SI_7_), .B2(n9400), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10029), .ZN(n8919) );
  INV_X1 U11341 ( .A(n8919), .ZN(P3_U3288) );
  INV_X1 U11342 ( .A(n9653), .ZN(n8924) );
  NAND2_X1 U11343 ( .A1(n8921), .A2(n8920), .ZN(n8927) );
  NAND2_X1 U11344 ( .A1(n8927), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8922) );
  XNOR2_X1 U11345 ( .A(n8922), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9654) );
  INV_X1 U11346 ( .A(n9654), .ZN(n8923) );
  OAI222_X1 U11347 ( .A1(n14436), .A2(n9657), .B1(n14434), .B2(n8924), .C1(
        P1_U3086), .C2(n8923), .ZN(P1_U3351) );
  OAI222_X1 U11348 ( .A1(n13820), .A2(n8925), .B1(n13818), .B2(n8924), .C1(
        P2_U3088), .C2(n13352), .ZN(P2_U3323) );
  OAI222_X1 U11349 ( .A1(n13820), .A2(n8926), .B1(n13818), .B2(n9671), .C1(
        n13365), .C2(P2_U3088), .ZN(P2_U3322) );
  NOR2_X1 U11350 ( .A1(n8927), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8930) );
  OR2_X1 U11351 ( .A1(n8930), .A2(n8966), .ZN(n8928) );
  MUX2_X1 U11352 ( .A(n8928), .B(P1_IR_REG_31__SCAN_IN), .S(n8929), .Z(n8931)
         );
  NAND2_X1 U11353 ( .A1(n8930), .A2(n8929), .ZN(n8945) );
  AND2_X1 U11354 ( .A1(n8931), .A2(n8945), .ZN(n14027) );
  INV_X1 U11355 ( .A(n14027), .ZN(n8932) );
  OAI222_X1 U11356 ( .A1(n14436), .A2(n8933), .B1(n14434), .B2(n9671), .C1(
        n8932), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U11357 ( .A(n13221), .ZN(n13227) );
  INV_X1 U11358 ( .A(n9400), .ZN(n13228) );
  OAI222_X1 U11359 ( .A1(n13227), .A2(n8935), .B1(n13228), .B2(n8934), .C1(
        n10225), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U11360 ( .A(n8936), .ZN(n8938) );
  INV_X1 U11361 ( .A(SI_2_), .ZN(n8937) );
  OAI222_X1 U11362 ( .A1(n9981), .A2(P3_U3151), .B1(n13227), .B2(n8938), .C1(
        n8937), .C2(n13228), .ZN(P3_U3293) );
  OAI222_X1 U11363 ( .A1(P3_U3151), .A2(n9567), .B1(n13228), .B2(n8940), .C1(
        n13227), .C2(n8939), .ZN(P3_U3294) );
  OAI222_X1 U11364 ( .A1(P3_U3151), .A2(n10028), .B1(n13228), .B2(n8942), .C1(
        n13227), .C2(n8941), .ZN(P3_U3289) );
  INV_X1 U11365 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8943) );
  INV_X1 U11366 ( .A(n9030), .ZN(n14967) );
  OAI222_X1 U11367 ( .A1(n13820), .A2(n8943), .B1(n13818), .B2(n9682), .C1(
        n14967), .C2(P2_U3088), .ZN(P2_U3321) );
  NAND2_X1 U11368 ( .A1(n8945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8944) );
  MUX2_X1 U11369 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8944), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n8946) );
  AND2_X1 U11370 ( .A1(n8946), .A2(n8958), .ZN(n9683) );
  INV_X1 U11371 ( .A(n9683), .ZN(n9162) );
  OAI222_X1 U11372 ( .A1(n14436), .A2(n8947), .B1(n14434), .B2(n9682), .C1(
        n9162), .C2(P1_U3086), .ZN(P1_U3349) );
  AOI222_X1 U11373 ( .A1(n8948), .A2(n13221), .B1(SI_9_), .B2(n9400), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10554), .ZN(n8949) );
  INV_X1 U11374 ( .A(n8949), .ZN(P3_U3286) );
  NAND2_X1 U11375 ( .A1(n8958), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8950) );
  XNOR2_X1 U11376 ( .A(n8950), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14044) );
  INV_X1 U11377 ( .A(n14044), .ZN(n14036) );
  OAI222_X1 U11378 ( .A1(n14436), .A2(n8951), .B1(n14434), .B2(n10116), .C1(
        n14036), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U11379 ( .A(n13380), .ZN(n13374) );
  OAI222_X1 U11380 ( .A1(n13820), .A2(n8952), .B1(n13818), .B2(n10116), .C1(
        n13374), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U11381 ( .A(n8953), .ZN(n8954) );
  OAI222_X1 U11382 ( .A1(n10557), .A2(P3_U3151), .B1(n13227), .B2(n8954), .C1(
        n7544), .C2(n13228), .ZN(P3_U3285) );
  INV_X1 U11383 ( .A(n8955), .ZN(n8957) );
  OAI222_X1 U11384 ( .A1(n13227), .A2(n8957), .B1(n7313), .B2(P3_U3151), .C1(
        n8956), .C2(n13228), .ZN(P3_U3284) );
  NAND2_X1 U11385 ( .A1(n8987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U11386 ( .A(n8959), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10122) );
  INV_X1 U11387 ( .A(n10122), .ZN(n9165) );
  OAI222_X1 U11388 ( .A1(n14436), .A2(n8960), .B1(n14434), .B2(n10121), .C1(
        n9165), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U11389 ( .A(n13394), .ZN(n13388) );
  OAI222_X1 U11390 ( .A1(n13820), .A2(n8961), .B1(n13818), .B2(n10121), .C1(
        n13388), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U11391 ( .A1(n9896), .A2(n8962), .ZN(n10108) );
  XNOR2_X2 U11392 ( .A(n8965), .B(P1_IR_REG_22__SCAN_IN), .ZN(n10306) );
  INV_X1 U11393 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U11394 ( .A1(n10306), .A2(n9247), .ZN(n11572) );
  INV_X1 U11395 ( .A(n8968), .ZN(n8973) );
  OR2_X1 U11396 ( .A1(n11572), .A2(n8973), .ZN(n8972) );
  NAND2_X1 U11397 ( .A1(n8969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U11398 ( .A1(n8972), .A2(n11413), .ZN(n8974) );
  NAND2_X1 U11399 ( .A1(n8973), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11627) );
  NAND2_X1 U11400 ( .A1(n9378), .A2(n11627), .ZN(n8975) );
  AND2_X1 U11401 ( .A1(n8974), .A2(n8975), .ZN(n14731) );
  INV_X1 U11402 ( .A(n8974), .ZN(n8976) );
  INV_X1 U11403 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9237) );
  INV_X1 U11404 ( .A(n12134), .ZN(n9369) );
  INV_X1 U11405 ( .A(n14426), .ZN(n8980) );
  INV_X1 U11406 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U11407 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U11408 ( .A1(n9369), .A2(n8981), .ZN(n9259) );
  AOI21_X1 U11409 ( .B1(n14426), .B2(n9237), .A(n9259), .ZN(n8982) );
  INV_X1 U11410 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9258) );
  XNOR2_X1 U11411 ( .A(n8982), .B(n9258), .ZN(n8983) );
  AOI22_X1 U11412 ( .A1(n9065), .A2(n8983), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n8984) );
  OAI21_X1 U11413 ( .B1(n14729), .B2(n6900), .A(n8984), .ZN(P1_U3243) );
  OAI222_X1 U11414 ( .A1(n13227), .A2(n8986), .B1(n13228), .B2(n8985), .C1(
        n10881), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U11415 ( .A1(n9100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8988) );
  XNOR2_X1 U11416 ( .A(n8988), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14061) );
  INV_X1 U11417 ( .A(n14061), .ZN(n8989) );
  OAI222_X1 U11418 ( .A1(n14436), .A2(n8990), .B1(n14434), .B2(n10136), .C1(
        n8989), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U11419 ( .A(n9036), .ZN(n9432) );
  OAI222_X1 U11420 ( .A1(n13820), .A2(n8991), .B1(n13818), .B2(n10136), .C1(
        n9432), .C2(P2_U3088), .ZN(P2_U3318) );
  NOR2_X1 U11421 ( .A1(n14731), .A2(P1_U4016), .ZN(P1_U3085) );
  MUX2_X1 U11422 ( .A(n9431), .B(P2_REG1_REG_9__SCAN_IN), .S(n9036), .Z(n9005)
         );
  XNOR2_X1 U11423 ( .A(n14954), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14952) );
  XNOR2_X1 U11424 ( .A(n13325), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n13332) );
  AND2_X1 U11425 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13331) );
  NAND2_X1 U11426 ( .A1(n13332), .A2(n13331), .ZN(n13330) );
  INV_X1 U11427 ( .A(n13325), .ZN(n9016) );
  NAND2_X1 U11428 ( .A1(n9016), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U11429 ( .A1(n13330), .A2(n8992), .ZN(n14951) );
  NAND2_X1 U11430 ( .A1(n14952), .A2(n14951), .ZN(n14950) );
  INV_X1 U11431 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8993) );
  OR2_X1 U11432 ( .A1(n14954), .A2(n8993), .ZN(n8994) );
  NAND2_X1 U11433 ( .A1(n14950), .A2(n8994), .ZN(n13340) );
  XNOR2_X1 U11434 ( .A(n13336), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U11435 ( .A1(n13340), .A2(n13341), .ZN(n13339) );
  OR2_X1 U11436 ( .A1(n13336), .A2(n8995), .ZN(n8996) );
  NAND2_X1 U11437 ( .A1(n13339), .A2(n8996), .ZN(n13350) );
  XNOR2_X1 U11438 ( .A(n13352), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U11439 ( .A1(n13350), .A2(n13351), .ZN(n13349) );
  INV_X1 U11440 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8997) );
  OR2_X1 U11441 ( .A1(n13352), .A2(n8997), .ZN(n8998) );
  NAND2_X1 U11442 ( .A1(n13349), .A2(n8998), .ZN(n13363) );
  XNOR2_X1 U11443 ( .A(n13365), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n13364) );
  NAND2_X1 U11444 ( .A1(n13363), .A2(n13364), .ZN(n13362) );
  NAND2_X1 U11445 ( .A1(n9028), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11446 ( .A1(n13362), .A2(n8999), .ZN(n14963) );
  MUX2_X1 U11447 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n8545), .S(n9030), .Z(n14964) );
  NAND2_X1 U11448 ( .A1(n14963), .A2(n14964), .ZN(n14962) );
  NAND2_X1 U11449 ( .A1(n9030), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11450 ( .A1(n14962), .A2(n9000), .ZN(n13378) );
  MUX2_X1 U11451 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8560), .S(n13380), .Z(
        n13379) );
  NAND2_X1 U11452 ( .A1(n13378), .A2(n13379), .ZN(n13377) );
  NAND2_X1 U11453 ( .A1(n13380), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11454 ( .A1(n13377), .A2(n9001), .ZN(n13393) );
  MUX2_X1 U11455 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8579), .S(n13394), .Z(
        n13392) );
  NAND2_X1 U11456 ( .A1(n13393), .A2(n13392), .ZN(n13391) );
  NAND2_X1 U11457 ( .A1(n13394), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11458 ( .A1(n13391), .A2(n9002), .ZN(n9004) );
  OR2_X1 U11459 ( .A1(n9004), .A2(n9005), .ZN(n9434) );
  INV_X1 U11460 ( .A(n9434), .ZN(n9003) );
  AOI21_X1 U11461 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9044) );
  NAND2_X1 U11462 ( .A1(n9006), .A2(n11007), .ZN(n9007) );
  NAND2_X1 U11463 ( .A1(n9007), .A2(n6588), .ZN(n9009) );
  AND2_X1 U11464 ( .A1(n9009), .A2(n9008), .ZN(n9011) );
  INV_X1 U11465 ( .A(n9011), .ZN(n9014) );
  NOR2_X1 U11466 ( .A1(n9012), .A2(P2_U3088), .ZN(n13807) );
  AND2_X1 U11467 ( .A1(n9011), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14949) );
  AND2_X1 U11468 ( .A1(n9012), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9013) );
  AND2_X1 U11469 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10178) );
  INV_X1 U11470 ( .A(n10178), .ZN(n9015) );
  OAI21_X1 U11471 ( .B1(n14996), .B2(n9432), .A(n9015), .ZN(n9042) );
  MUX2_X1 U11472 ( .A(n9785), .B(P2_REG2_REG_3__SCAN_IN), .S(n13336), .Z(
        n13343) );
  XNOR2_X1 U11473 ( .A(n14954), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n14957) );
  NAND2_X1 U11474 ( .A1(n9016), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11475 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9017) );
  AOI21_X1 U11476 ( .B1(n13325), .B2(n9493), .A(n9017), .ZN(n9018) );
  NAND2_X1 U11477 ( .A1(n9019), .A2(n9018), .ZN(n13329) );
  NAND2_X1 U11478 ( .A1(n13329), .A2(n9019), .ZN(n14956) );
  NAND2_X1 U11479 ( .A1(n14957), .A2(n14956), .ZN(n9022) );
  OR2_X1 U11480 ( .A1(n14954), .A2(n9020), .ZN(n9021) );
  NAND2_X1 U11481 ( .A1(n9022), .A2(n9021), .ZN(n13342) );
  NAND2_X1 U11482 ( .A1(n13343), .A2(n13342), .ZN(n13355) );
  OR2_X1 U11483 ( .A1(n13336), .A2(n9785), .ZN(n13354) );
  NAND2_X1 U11484 ( .A1(n13355), .A2(n13354), .ZN(n9024) );
  MUX2_X1 U11485 ( .A(n9821), .B(P2_REG2_REG_4__SCAN_IN), .S(n13352), .Z(n9023) );
  NAND2_X1 U11486 ( .A1(n9024), .A2(n9023), .ZN(n13368) );
  OR2_X1 U11487 ( .A1(n13352), .A2(n9821), .ZN(n13367) );
  NAND2_X1 U11488 ( .A1(n13368), .A2(n13367), .ZN(n9027) );
  MUX2_X1 U11489 ( .A(n9025), .B(P2_REG2_REG_5__SCAN_IN), .S(n13365), .Z(n9026) );
  NAND2_X1 U11490 ( .A1(n9027), .A2(n9026), .ZN(n13370) );
  NAND2_X1 U11491 ( .A1(n9028), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11492 ( .A1(n13370), .A2(n9029), .ZN(n14971) );
  MUX2_X1 U11493 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9752), .S(n9030), .Z(n14970) );
  NAND2_X1 U11494 ( .A1(n14971), .A2(n14970), .ZN(n14969) );
  NAND2_X1 U11495 ( .A1(n9030), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U11496 ( .A1(n14969), .A2(n13382), .ZN(n9032) );
  MUX2_X1 U11497 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9539), .S(n13380), .Z(n9031) );
  NAND2_X1 U11498 ( .A1(n9032), .A2(n9031), .ZN(n13397) );
  NAND2_X1 U11499 ( .A1(n13380), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13396) );
  NAND2_X1 U11500 ( .A1(n13397), .A2(n13396), .ZN(n9034) );
  MUX2_X1 U11501 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9807), .S(n13394), .Z(n9033) );
  NAND2_X1 U11502 ( .A1(n9034), .A2(n9033), .ZN(n13399) );
  NAND2_X1 U11503 ( .A1(n13394), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11504 ( .A1(n13399), .A2(n9035), .ZN(n9038) );
  INV_X1 U11505 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10071) );
  MUX2_X1 U11506 ( .A(n10071), .B(P2_REG2_REG_9__SCAN_IN), .S(n9036), .Z(n9037) );
  OR2_X1 U11507 ( .A1(n9038), .A2(n9037), .ZN(n9422) );
  NAND2_X1 U11508 ( .A1(n9038), .A2(n9037), .ZN(n9040) );
  INV_X1 U11509 ( .A(n9010), .ZN(n12458) );
  NAND2_X1 U11510 ( .A1(n9039), .A2(n12458), .ZN(n14998) );
  AOI21_X1 U11511 ( .B1(n9422), .B2(n9040), .A(n14998), .ZN(n9041) );
  AOI211_X1 U11512 ( .C1(n14949), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n9042), .B(
        n9041), .ZN(n9043) );
  OAI21_X1 U11513 ( .B1(n9044), .B2(n15018), .A(n9043), .ZN(P2_U3223) );
  INV_X1 U11514 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n15047) );
  OAI22_X1 U11515 ( .A1(n15018), .A2(n9045), .B1(n15047), .B2(n14998), .ZN(
        n9048) );
  NAND2_X1 U11516 ( .A1(n15002), .A2(n9045), .ZN(n9046) );
  OAI211_X1 U11517 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14998), .A(n9046), .B(
        n14996), .ZN(n9047) );
  MUX2_X1 U11518 ( .A(n9048), .B(n9047), .S(P2_IR_REG_0__SCAN_IN), .Z(n9051)
         );
  INV_X1 U11519 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9049) );
  INV_X1 U11520 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n15038) );
  OAI22_X1 U11521 ( .A1(n15032), .A2(n9049), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15038), .ZN(n9050) );
  OR2_X1 U11522 ( .A1(n9051), .A2(n9050), .ZN(P2_U3214) );
  NAND2_X1 U11523 ( .A1(n14432), .A2(P1_B_REG_SCAN_IN), .ZN(n9052) );
  MUX2_X1 U11524 ( .A(n9052), .B(P1_B_REG_SCAN_IN), .S(n9339), .Z(n9053) );
  NOR2_X2 U11525 ( .A1(n9354), .A2(n9378), .ZN(n14810) );
  NAND2_X1 U11526 ( .A1(n9055), .A2(n14431), .ZN(n9057) );
  OAI22_X1 U11527 ( .A1(n14825), .A2(P1_D_REG_0__SCAN_IN), .B1(n9339), .B2(
        n9057), .ZN(n9056) );
  INV_X1 U11528 ( .A(n9056), .ZN(P1_U3445) );
  OAI22_X1 U11529 ( .A1(n14825), .A2(P1_D_REG_1__SCAN_IN), .B1(n9058), .B2(
        n9057), .ZN(n9059) );
  INV_X1 U11530 ( .A(n9059), .ZN(P1_U3446) );
  NAND2_X1 U11531 ( .A1(n9065), .A2(n12134), .ZN(n14725) );
  AND2_X1 U11532 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9060) );
  INV_X1 U11533 ( .A(n9060), .ZN(n9257) );
  INV_X1 U11534 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9080) );
  MUX2_X1 U11535 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9080), .S(n6574), .Z(n9064)
         );
  MUX2_X1 U11536 ( .A(n9080), .B(P1_REG2_REG_1__SCAN_IN), .S(n6574), .Z(n9061)
         );
  NAND2_X1 U11537 ( .A1(n9061), .A2(n9060), .ZN(n13994) );
  INV_X1 U11538 ( .A(n13994), .ZN(n9063) );
  NOR2_X1 U11539 ( .A1(n12134), .A2(n14426), .ZN(n9062) );
  NAND2_X1 U11540 ( .A1(n9065), .A2(n9062), .ZN(n14723) );
  AOI211_X1 U11541 ( .C1(n9257), .C2(n9064), .A(n9063), .B(n14723), .ZN(n9069)
         );
  INV_X1 U11542 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14911) );
  MUX2_X1 U11543 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14911), .S(n9289), .Z(n9066) );
  NOR3_X1 U11544 ( .A1(n9066), .A2(n9237), .A3(n9258), .ZN(n13990) );
  INV_X1 U11545 ( .A(n13990), .ZN(n9074) );
  OAI21_X1 U11546 ( .B1(n9237), .B2(n9258), .A(n9066), .ZN(n9067) );
  AND3_X1 U11547 ( .A1(n14738), .A2(n9074), .A3(n9067), .ZN(n9068) );
  NOR2_X1 U11548 ( .A1(n9069), .A2(n9068), .ZN(n9071) );
  AOI22_X1 U11549 ( .A1(n14731), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9070) );
  OAI211_X1 U11550 ( .C1(n6574), .C2(n14725), .A(n9071), .B(n9070), .ZN(
        P1_U3244) );
  NOR2_X1 U11551 ( .A1(n6574), .A2(n14911), .ZN(n13989) );
  INV_X1 U11552 ( .A(n13989), .ZN(n9073) );
  INV_X1 U11553 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14913) );
  MUX2_X1 U11554 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14913), .S(n13998), .Z(
        n9072) );
  AOI21_X1 U11555 ( .B1(n9074), .B2(n9073), .A(n9072), .ZN(n13992) );
  INV_X1 U11556 ( .A(n13992), .ZN(n14009) );
  INV_X1 U11557 ( .A(n13998), .ZN(n9083) );
  NAND2_X1 U11558 ( .A1(n9083), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14008) );
  INV_X1 U11559 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14915) );
  MUX2_X1 U11560 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n14915), .S(n14012), .Z(
        n14007) );
  INV_X1 U11561 ( .A(n9225), .ZN(n14011) );
  NOR2_X1 U11562 ( .A1(n14012), .A2(n14915), .ZN(n9224) );
  INV_X1 U11563 ( .A(n9224), .ZN(n9076) );
  INV_X1 U11564 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14917) );
  MUX2_X1 U11565 ( .A(n14917), .B(P1_REG1_REG_4__SCAN_IN), .S(n9654), .Z(n9075) );
  AOI21_X1 U11566 ( .B1(n14011), .B2(n9076), .A(n9075), .ZN(n9227) );
  AOI21_X1 U11567 ( .B1(n9654), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9227), .ZN(
        n14024) );
  INV_X1 U11568 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14919) );
  MUX2_X1 U11569 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14919), .S(n14027), .Z(
        n14025) );
  NAND2_X1 U11570 ( .A1(n14024), .A2(n14025), .ZN(n14023) );
  OAI21_X1 U11571 ( .B1(n14027), .B2(P1_REG1_REG_5__SCAN_IN), .A(n14023), .ZN(
        n9078) );
  INV_X1 U11572 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14921) );
  MUX2_X1 U11573 ( .A(n14921), .B(P1_REG1_REG_6__SCAN_IN), .S(n9683), .Z(n9077) );
  AOI211_X1 U11574 ( .C1(n9078), .C2(n9077), .A(n14041), .B(n14721), .ZN(n9096) );
  INV_X1 U11575 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9661) );
  MUX2_X1 U11576 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9661), .S(n14027), .Z(n9089) );
  INV_X1 U11577 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9079) );
  MUX2_X1 U11578 ( .A(n9079), .B(P1_REG2_REG_2__SCAN_IN), .S(n13998), .Z(n9082) );
  OR2_X1 U11579 ( .A1(n6574), .A2(n9080), .ZN(n13993) );
  NAND2_X1 U11580 ( .A1(n13994), .A2(n13993), .ZN(n9081) );
  NAND2_X1 U11581 ( .A1(n9082), .A2(n9081), .ZN(n14014) );
  NAND2_X1 U11582 ( .A1(n9083), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U11583 ( .A1(n14014), .A2(n14013), .ZN(n9085) );
  INV_X1 U11584 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9323) );
  MUX2_X1 U11585 ( .A(n9323), .B(P1_REG2_REG_3__SCAN_IN), .S(n14012), .Z(n9084) );
  NAND2_X1 U11586 ( .A1(n9085), .A2(n9084), .ZN(n14017) );
  INV_X1 U11587 ( .A(n14012), .ZN(n14006) );
  NAND2_X1 U11588 ( .A1(n14006), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11589 ( .A1(n14017), .A2(n9220), .ZN(n9087) );
  INV_X1 U11590 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9364) );
  MUX2_X1 U11591 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9364), .S(n9654), .Z(n9086)
         );
  NAND2_X1 U11592 ( .A1(n9087), .A2(n9086), .ZN(n14029) );
  NAND2_X1 U11593 ( .A1(n9654), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U11594 ( .A1(n14029), .A2(n14028), .ZN(n9088) );
  NAND2_X1 U11595 ( .A1(n9089), .A2(n9088), .ZN(n14032) );
  NAND2_X1 U11596 ( .A1(n14027), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11597 ( .A1(n14032), .A2(n9093), .ZN(n9091) );
  INV_X1 U11598 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9707) );
  MUX2_X1 U11599 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9707), .S(n9683), .Z(n9090)
         );
  NAND2_X1 U11600 ( .A1(n9091), .A2(n9090), .ZN(n14047) );
  MUX2_X1 U11601 ( .A(n9707), .B(P1_REG2_REG_6__SCAN_IN), .S(n9683), .Z(n9092)
         );
  NAND3_X1 U11602 ( .A1(n14032), .A2(n9093), .A3(n9092), .ZN(n9094) );
  AND3_X1 U11603 ( .A1(n14733), .A2(n14047), .A3(n9094), .ZN(n9095) );
  NOR2_X1 U11604 ( .A1(n9096), .A2(n9095), .ZN(n9099) );
  INV_X1 U11605 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9097) );
  NOR2_X1 U11606 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9097), .ZN(n10103) );
  AOI21_X1 U11607 ( .B1(n14731), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10103), .ZN(
        n9098) );
  OAI211_X1 U11608 ( .C1(n9162), .C2(n14725), .A(n9099), .B(n9098), .ZN(
        P1_U3249) );
  INV_X1 U11609 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9105) );
  NOR2_X1 U11610 ( .A1(n9102), .A2(n8966), .ZN(n9101) );
  MUX2_X1 U11611 ( .A(n8966), .B(n9101), .S(P1_IR_REG_10__SCAN_IN), .Z(n9104)
         );
  NAND2_X1 U11612 ( .A1(n9102), .A2(n15306), .ZN(n9157) );
  INV_X1 U11613 ( .A(n9157), .ZN(n9103) );
  INV_X1 U11614 ( .A(n14704), .ZN(n14712) );
  OAI222_X1 U11615 ( .A1(n14436), .A2(n9105), .B1(n14428), .B2(n10409), .C1(
        n14712), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U11616 ( .A(n13411), .ZN(n13407) );
  OAI222_X1 U11617 ( .A1(n13820), .A2(n9106), .B1(n13818), .B2(n10409), .C1(
        n13407), .C2(P2_U3088), .ZN(P2_U3317) );
  OAI222_X1 U11618 ( .A1(n13227), .A2(n9108), .B1(n13228), .B2(n9107), .C1(
        n10992), .C2(P3_U3151), .ZN(P3_U3282) );
  NOR2_X1 U11619 ( .A1(n9109), .A2(P2_U3088), .ZN(n9146) );
  OAI21_X1 U11620 ( .B1(n9112), .B2(n9111), .A(n9110), .ZN(n9113) );
  NAND2_X1 U11621 ( .A1(n9113), .A2(n7445), .ZN(n9115) );
  INV_X1 U11622 ( .A(n13238), .ZN(n13285) );
  INV_X1 U11623 ( .A(n12147), .ZN(n15040) );
  OAI22_X1 U11624 ( .A1(n15040), .A2(n13595), .B1(n9528), .B2(n15039), .ZN(
        n9910) );
  AOI22_X1 U11625 ( .A1(n13285), .A2(n9910), .B1(n14943), .B2(n15062), .ZN(
        n9114) );
  OAI211_X1 U11626 ( .C1(n9146), .C2(n9116), .A(n9115), .B(n9114), .ZN(
        P2_U3209) );
  INV_X1 U11627 ( .A(n9117), .ZN(n9118) );
  AOI21_X1 U11628 ( .B1(n9120), .B2(n9119), .A(n9118), .ZN(n9124) );
  INV_X1 U11629 ( .A(n14933), .ZN(n13294) );
  NOR2_X1 U11630 ( .A1(n13297), .A2(n12148), .ZN(n9122) );
  OAI22_X1 U11631 ( .A1(n9146), .A2(n13323), .B1(n14932), .B2(n6787), .ZN(
        n9121) );
  AOI211_X1 U11632 ( .C1(n13294), .C2(n12144), .A(n9122), .B(n9121), .ZN(n9123) );
  OAI21_X1 U11633 ( .B1(n9124), .B2(n14939), .A(n9123), .ZN(P2_U3194) );
  XNOR2_X1 U11634 ( .A(n12403), .B(n12402), .ZN(n9134) );
  INV_X1 U11635 ( .A(n9134), .ZN(n9495) );
  AOI21_X1 U11636 ( .B1(n6929), .B2(n15035), .A(n8705), .ZN(n9125) );
  NAND2_X1 U11637 ( .A1(n9125), .A2(n9904), .ZN(n9498) );
  OAI21_X1 U11638 ( .B1(n12148), .B2(n15097), .A(n9498), .ZN(n9135) );
  AOI22_X1 U11639 ( .A1(n13667), .A2(n12144), .B1(n13322), .B2(n13665), .ZN(
        n9133) );
  NAND2_X1 U11640 ( .A1(n9525), .A2(n9129), .ZN(n9510) );
  OAI21_X1 U11641 ( .B1(n9129), .B2(n12403), .A(n9510), .ZN(n9131) );
  NOR2_X1 U11642 ( .A1(n8881), .A2(n8879), .ZN(n12437) );
  NOR2_X1 U11643 ( .A1(n12352), .A2(n13459), .ZN(n9130) );
  NAND2_X1 U11644 ( .A1(n9131), .A2(n13683), .ZN(n9132) );
  OAI211_X1 U11645 ( .C1(n9134), .C2(n9127), .A(n9133), .B(n9132), .ZN(n9500)
         );
  AOI211_X1 U11646 ( .C1(n15088), .C2(n9495), .A(n9135), .B(n9500), .ZN(n15060) );
  INV_X1 U11647 ( .A(n9136), .ZN(n9137) );
  INV_X1 U11648 ( .A(n15053), .ZN(n9142) );
  AND2_X1 U11649 ( .A1(n15056), .A2(n9139), .ZN(n9140) );
  AND2_X1 U11650 ( .A1(n9141), .A2(n9140), .ZN(n10781) );
  NAND2_X1 U11651 ( .A1(n15139), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9143) );
  OAI21_X1 U11652 ( .B1(n15060), .B2(n15139), .A(n9143), .ZN(P2_U3500) );
  INV_X1 U11653 ( .A(n9144), .ZN(n9145) );
  OAI21_X1 U11654 ( .B1(n9145), .B2(n14939), .A(n13297), .ZN(n9148) );
  INV_X1 U11655 ( .A(n9146), .ZN(n9147) );
  AOI22_X1 U11656 ( .A1(n9148), .A2(n15035), .B1(n9147), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9150) );
  NAND4_X1 U11657 ( .A1(n7445), .A2(n8705), .A3(n12144), .A4(n12402), .ZN(
        n9149) );
  OAI211_X1 U11658 ( .C1(n15040), .C2(n14932), .A(n9150), .B(n9149), .ZN(
        P2_U3204) );
  XNOR2_X1 U11659 ( .A(n9152), .B(n9151), .ZN(n9156) );
  INV_X1 U11660 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15314) );
  INV_X1 U11661 ( .A(n14947), .ZN(n13265) );
  AOI22_X1 U11662 ( .A1(n13667), .A2(n13322), .B1(n13320), .B2(n13665), .ZN(
        n9782) );
  OAI22_X1 U11663 ( .A1(n9782), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15314), .ZN(n9154) );
  NOR2_X1 U11664 ( .A1(n13297), .A2(n9536), .ZN(n9153) );
  AOI211_X1 U11665 ( .C1(n15314), .C2(n13265), .A(n9154), .B(n9153), .ZN(n9155) );
  OAI21_X1 U11666 ( .B1(n9156), .B2(n14939), .A(n9155), .ZN(P2_U3190) );
  INV_X1 U11667 ( .A(n10438), .ZN(n9160) );
  NAND2_X1 U11668 ( .A1(n9157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9275) );
  XNOR2_X1 U11669 ( .A(n9275), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10439) );
  OAI222_X1 U11670 ( .A1(n14436), .A2(n9158), .B1(n14428), .B2(n9160), .C1(
        P1_U3086), .C2(n9409), .ZN(P1_U3344) );
  INV_X1 U11671 ( .A(n14981), .ZN(n9159) );
  OAI222_X1 U11672 ( .A1(n13820), .A2(n9161), .B1(n13818), .B2(n9160), .C1(
        P2_U3088), .C2(n9159), .ZN(P2_U3316) );
  INV_X1 U11673 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10126) );
  MUX2_X1 U11674 ( .A(n10126), .B(P1_REG1_REG_8__SCAN_IN), .S(n10122), .Z(
        n9164) );
  INV_X1 U11675 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14923) );
  NOR2_X1 U11676 ( .A1(n9162), .A2(n14921), .ZN(n14040) );
  MUX2_X1 U11677 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14923), .S(n14044), .Z(
        n14039) );
  OAI21_X1 U11678 ( .B1(n14041), .B2(n14040), .A(n14039), .ZN(n14043) );
  OAI21_X1 U11679 ( .B1(n14923), .B2(n14036), .A(n14043), .ZN(n9163) );
  NOR2_X1 U11680 ( .A1(n9163), .A2(n9164), .ZN(n14056) );
  AOI21_X1 U11681 ( .B1(n9164), .B2(n9163), .A(n14056), .ZN(n9176) );
  NOR2_X1 U11682 ( .A1(n10127), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10378) );
  NOR2_X1 U11683 ( .A1(n14725), .A2(n9165), .ZN(n9166) );
  AOI211_X1 U11684 ( .C1(n14731), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10378), .B(
        n9166), .ZN(n9175) );
  NAND2_X1 U11685 ( .A1(n9683), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U11686 ( .A1(n14047), .A2(n14046), .ZN(n9168) );
  INV_X1 U11687 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9698) );
  MUX2_X1 U11688 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9698), .S(n14044), .Z(n9167) );
  NAND2_X1 U11689 ( .A1(n9168), .A2(n9167), .ZN(n14049) );
  NAND2_X1 U11690 ( .A1(n14044), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11691 ( .A1(n14049), .A2(n9172), .ZN(n9170) );
  INV_X1 U11692 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10125) );
  MUX2_X1 U11693 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10125), .S(n10122), .Z(
        n9169) );
  NAND2_X1 U11694 ( .A1(n9170), .A2(n9169), .ZN(n14064) );
  MUX2_X1 U11695 ( .A(n10125), .B(P1_REG2_REG_8__SCAN_IN), .S(n10122), .Z(
        n9171) );
  NAND3_X1 U11696 ( .A1(n14049), .A2(n9172), .A3(n9171), .ZN(n9173) );
  NAND3_X1 U11697 ( .A1(n14733), .A2(n14064), .A3(n9173), .ZN(n9174) );
  OAI211_X1 U11698 ( .C1(n9176), .C2(n14721), .A(n9175), .B(n9174), .ZN(
        P1_U3251) );
  INV_X1 U11699 ( .A(n10987), .ZN(n10991) );
  INV_X1 U11700 ( .A(n9177), .ZN(n9178) );
  OAI222_X1 U11701 ( .A1(n10991), .A2(P3_U3151), .B1(n13227), .B2(n9178), .C1(
        n15462), .C2(n13228), .ZN(P3_U3281) );
  INV_X1 U11702 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14927) );
  NOR2_X1 U11703 ( .A1(n10122), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n14054) );
  INV_X1 U11704 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U11705 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10317), .S(n14061), .Z(
        n14055) );
  OAI21_X1 U11706 ( .B1(n14061), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14053), .ZN(
        n14700) );
  MUX2_X1 U11707 ( .A(n14927), .B(P1_REG1_REG_10__SCAN_IN), .S(n14704), .Z(
        n9179) );
  OR2_X1 U11708 ( .A1(n14700), .A2(n9179), .ZN(n14701) );
  OAI21_X1 U11709 ( .B1(n14927), .B2(n14712), .A(n14701), .ZN(n9181) );
  INV_X1 U11710 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U11711 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n9409), .B1(n10439), 
        .B2(n14673), .ZN(n9180) );
  NOR2_X1 U11712 ( .A1(n9181), .A2(n9180), .ZN(n9404) );
  AOI21_X1 U11713 ( .B1(n9181), .B2(n9180), .A(n9404), .ZN(n9194) );
  NAND2_X1 U11714 ( .A1(n10122), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14063) );
  NAND2_X1 U11715 ( .A1(n14064), .A2(n14063), .ZN(n9183) );
  INV_X1 U11716 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10139) );
  MUX2_X1 U11717 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10139), .S(n14061), .Z(
        n9182) );
  NAND2_X1 U11718 ( .A1(n9183), .A2(n9182), .ZN(n14707) );
  NAND2_X1 U11719 ( .A1(n14061), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U11720 ( .A1(n14707), .A2(n14706), .ZN(n9185) );
  INV_X1 U11721 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10156) );
  MUX2_X1 U11722 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10156), .S(n14704), .Z(
        n9184) );
  NAND2_X1 U11723 ( .A1(n9185), .A2(n9184), .ZN(n14709) );
  NAND2_X1 U11724 ( .A1(n14704), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U11725 ( .A1(n14709), .A2(n9186), .ZN(n9188) );
  INV_X1 U11726 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10460) );
  MUX2_X1 U11727 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10460), .S(n10439), .Z(
        n9187) );
  NAND2_X1 U11728 ( .A1(n9187), .A2(n9188), .ZN(n9408) );
  OAI211_X1 U11729 ( .C1(n9188), .C2(n9187), .A(n14733), .B(n9408), .ZN(n9191)
         );
  NAND2_X1 U11730 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10678)
         );
  INV_X1 U11731 ( .A(n10678), .ZN(n9189) );
  AOI21_X1 U11732 ( .B1(n14731), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9189), .ZN(
        n9190) );
  OAI211_X1 U11733 ( .C1(n14725), .C2(n9409), .A(n9191), .B(n9190), .ZN(n9192)
         );
  INV_X1 U11734 ( .A(n9192), .ZN(n9193) );
  OAI21_X1 U11735 ( .B1(n9194), .B2(n14721), .A(n9193), .ZN(P1_U3254) );
  INV_X1 U11736 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9195) );
  NOR2_X1 U11737 ( .A1(n9218), .A2(n9195), .ZN(P3_U3245) );
  INV_X1 U11738 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15445) );
  NOR2_X1 U11739 ( .A1(n9218), .A2(n15445), .ZN(P3_U3241) );
  INV_X1 U11740 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9196) );
  NOR2_X1 U11741 ( .A1(n9218), .A2(n9196), .ZN(P3_U3240) );
  INV_X1 U11742 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15389) );
  NOR2_X1 U11743 ( .A1(n9218), .A2(n15389), .ZN(P3_U3242) );
  INV_X1 U11744 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9197) );
  NOR2_X1 U11745 ( .A1(n9218), .A2(n9197), .ZN(P3_U3236) );
  INV_X1 U11746 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9198) );
  NOR2_X1 U11747 ( .A1(n9218), .A2(n9198), .ZN(P3_U3244) );
  INV_X1 U11748 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U11749 ( .A1(n9218), .A2(n9199), .ZN(P3_U3237) );
  INV_X1 U11750 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15315) );
  NOR2_X1 U11751 ( .A1(n9218), .A2(n15315), .ZN(P3_U3260) );
  INV_X1 U11752 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9200) );
  NOR2_X1 U11753 ( .A1(n9218), .A2(n9200), .ZN(P3_U3238) );
  INV_X1 U11754 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9201) );
  NOR2_X1 U11755 ( .A1(n9218), .A2(n9201), .ZN(P3_U3262) );
  INV_X1 U11756 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n15492) );
  NOR2_X1 U11757 ( .A1(n9218), .A2(n15492), .ZN(P3_U3243) );
  INV_X1 U11758 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9202) );
  NOR2_X1 U11759 ( .A1(n9218), .A2(n9202), .ZN(P3_U3239) );
  INV_X1 U11760 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9203) );
  NOR2_X1 U11761 ( .A1(n9218), .A2(n9203), .ZN(P3_U3234) );
  INV_X1 U11762 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9204) );
  NOR2_X1 U11763 ( .A1(n9218), .A2(n9204), .ZN(P3_U3235) );
  INV_X2 U11764 ( .A(n15236), .ZN(n9218) );
  INV_X1 U11765 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9205) );
  NOR2_X1 U11766 ( .A1(n9218), .A2(n9205), .ZN(P3_U3263) );
  INV_X1 U11767 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9206) );
  NOR2_X1 U11768 ( .A1(n9218), .A2(n9206), .ZN(P3_U3258) );
  INV_X1 U11769 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9207) );
  NOR2_X1 U11770 ( .A1(n9218), .A2(n9207), .ZN(P3_U3259) );
  INV_X1 U11771 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9208) );
  NOR2_X1 U11772 ( .A1(n9218), .A2(n9208), .ZN(P3_U3250) );
  INV_X1 U11773 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9209) );
  NOR2_X1 U11774 ( .A1(n9218), .A2(n9209), .ZN(P3_U3255) );
  INV_X1 U11775 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9210) );
  NOR2_X1 U11776 ( .A1(n9218), .A2(n9210), .ZN(P3_U3247) );
  INV_X1 U11777 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9211) );
  NOR2_X1 U11778 ( .A1(n9218), .A2(n9211), .ZN(P3_U3251) );
  INV_X1 U11779 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9212) );
  NOR2_X1 U11780 ( .A1(n9218), .A2(n9212), .ZN(P3_U3248) );
  INV_X1 U11781 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9213) );
  NOR2_X1 U11782 ( .A1(n9218), .A2(n9213), .ZN(P3_U3261) );
  INV_X1 U11783 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9214) );
  NOR2_X1 U11784 ( .A1(n9218), .A2(n9214), .ZN(P3_U3253) );
  INV_X1 U11785 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9215) );
  NOR2_X1 U11786 ( .A1(n9218), .A2(n9215), .ZN(P3_U3252) );
  INV_X1 U11787 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U11788 ( .A1(n9218), .A2(n15347), .ZN(P3_U3257) );
  INV_X1 U11789 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9216) );
  NOR2_X1 U11790 ( .A1(n9218), .A2(n9216), .ZN(P3_U3256) );
  INV_X1 U11791 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n15448) );
  NOR2_X1 U11792 ( .A1(n9218), .A2(n15448), .ZN(P3_U3249) );
  INV_X1 U11793 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9217) );
  NOR2_X1 U11794 ( .A1(n9218), .A2(n9217), .ZN(P3_U3254) );
  INV_X1 U11795 ( .A(n14725), .ZN(n14736) );
  INV_X1 U11796 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14487) );
  MUX2_X1 U11797 ( .A(n9364), .B(P1_REG2_REG_4__SCAN_IN), .S(n9654), .Z(n9219)
         );
  NAND3_X1 U11798 ( .A1(n14017), .A2(n9220), .A3(n9219), .ZN(n9221) );
  NAND3_X1 U11799 ( .A1(n14733), .A2(n14029), .A3(n9221), .ZN(n9222) );
  NAND2_X1 U11800 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9892) );
  OAI211_X1 U11801 ( .C1(n14487), .C2(n14729), .A(n9222), .B(n9892), .ZN(n9229) );
  MUX2_X1 U11802 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14917), .S(n9654), .Z(n9223) );
  NOR3_X1 U11803 ( .A1(n9225), .A2(n9224), .A3(n9223), .ZN(n9226) );
  NOR3_X1 U11804 ( .A1(n14721), .A2(n9227), .A3(n9226), .ZN(n9228) );
  AOI211_X1 U11805 ( .C1(n14736), .C2(n9654), .A(n9229), .B(n9228), .ZN(n9262)
         );
  NAND2_X1 U11806 ( .A1(n9233), .A2(n9234), .ZN(n14421) );
  NAND2_X1 U11807 ( .A1(n11181), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11808 ( .A1(n9238), .A2(n9236), .ZN(n9324) );
  INV_X1 U11809 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10088) );
  OR2_X1 U11810 ( .A1(n9324), .A2(n10088), .ZN(n9241) );
  INV_X1 U11811 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9239) );
  INV_X1 U11812 ( .A(n10306), .ZN(n9244) );
  AND2_X2 U11813 ( .A1(n9358), .A2(n11771), .ZN(n10100) );
  NAND2_X1 U11814 ( .A1(n10100), .A2(n13987), .ZN(n9253) );
  INV_X1 U11815 ( .A(SI_0_), .ZN(n9248) );
  NOR2_X1 U11816 ( .A1(n11550), .A2(n9248), .ZN(n9250) );
  XNOR2_X1 U11817 ( .A(n9250), .B(n9249), .ZN(n14438) );
  MUX2_X1 U11818 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14438), .S(n11413), .Z(n14831) );
  INV_X1 U11819 ( .A(n9251), .ZN(n9361) );
  AOI22_X1 U11820 ( .A1(n14831), .A2(n11758), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n9361), .ZN(n9252) );
  AND2_X1 U11821 ( .A1(n9253), .A2(n9252), .ZN(n9256) );
  NAND2_X1 U11822 ( .A1(n13987), .A2(n11758), .ZN(n9255) );
  NAND2_X1 U11823 ( .A1(n9255), .A2(n9254), .ZN(n9303) );
  NAND2_X1 U11824 ( .A1(n9256), .A2(n9303), .ZN(n9304) );
  OAI21_X1 U11825 ( .B1(n9256), .B2(n9303), .A(n9304), .ZN(n9380) );
  MUX2_X1 U11826 ( .A(n9257), .B(n9380), .S(n14426), .Z(n9261) );
  NAND2_X1 U11827 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  OAI211_X1 U11828 ( .C1(n9261), .C2(n12134), .A(P1_U4016), .B(n9260), .ZN(
        n14003) );
  NAND2_X1 U11829 ( .A1(n9262), .A2(n14003), .ZN(P1_U3247) );
  INV_X1 U11830 ( .A(n9263), .ZN(n9265) );
  OAI222_X1 U11831 ( .A1(n12814), .A2(P3_U3151), .B1(n13227), .B2(n9265), .C1(
        n9264), .C2(n13228), .ZN(P3_U3280) );
  INV_X1 U11832 ( .A(n9266), .ZN(n9267) );
  AOI21_X1 U11833 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(n9273) );
  INV_X1 U11834 ( .A(n14932), .ZN(n13262) );
  INV_X1 U11835 ( .A(n12181), .ZN(n13319) );
  AOI22_X1 U11836 ( .A1(n13294), .A2(n13321), .B1(n13262), .B2(n13319), .ZN(
        n9272) );
  AND2_X1 U11837 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13348) );
  NOR2_X1 U11838 ( .A1(n14947), .A2(n9825), .ZN(n9270) );
  AOI211_X1 U11839 ( .C1(n15075), .C2(n14943), .A(n13348), .B(n9270), .ZN(
        n9271) );
  OAI211_X1 U11840 ( .C1(n9273), .C2(n14939), .A(n9272), .B(n9271), .ZN(
        P2_U3202) );
  INV_X1 U11841 ( .A(n10568), .ZN(n9278) );
  INV_X1 U11842 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11843 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U11844 ( .A1(n9276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9446) );
  XNOR2_X1 U11845 ( .A(n9446), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10569) );
  INV_X1 U11846 ( .A(n10569), .ZN(n9415) );
  OAI222_X1 U11847 ( .A1(n14436), .A2(n9277), .B1(n14428), .B2(n9278), .C1(
        n9415), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U11848 ( .A(n9437), .ZN(n14997) );
  OAI222_X1 U11849 ( .A1(n13820), .A2(n9279), .B1(n13818), .B2(n9278), .C1(
        n14997), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U11850 ( .A1(n11181), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9285) );
  INV_X1 U11851 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9731) );
  OR2_X1 U11852 ( .A1(n9324), .A2(n9731), .ZN(n9284) );
  INV_X1 U11853 ( .A(n9666), .ZN(n9280) );
  INV_X1 U11854 ( .A(n9322), .ZN(n9281) );
  NAND2_X1 U11855 ( .A1(n9281), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11856 ( .A1(n9298), .A2(n11758), .ZN(n9291) );
  OR2_X1 U11857 ( .A1(n9329), .A2(n9286), .ZN(n9288) );
  NAND2_X1 U11858 ( .A1(n11413), .A2(n6576), .ZN(n9311) );
  OR2_X1 U11859 ( .A1(n9311), .A2(n8287), .ZN(n9287) );
  NAND2_X1 U11860 ( .A1(n14834), .A2(n11771), .ZN(n9290) );
  NAND2_X1 U11861 ( .A1(n9291), .A2(n9290), .ZN(n9297) );
  INV_X1 U11862 ( .A(n9293), .ZN(n9294) );
  NAND2_X1 U11863 ( .A1(n9294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9295) );
  MUX2_X1 U11864 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9295), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9296) );
  NAND2_X2 U11865 ( .A1(n9292), .A2(n9296), .ZN(n11675) );
  AND2_X1 U11866 ( .A1(n14834), .A2(n11758), .ZN(n9299) );
  NAND2_X1 U11867 ( .A1(n9384), .A2(n9305), .ZN(n9393) );
  NAND2_X1 U11868 ( .A1(n11181), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9310) );
  INV_X1 U11869 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9398) );
  OR2_X1 U11870 ( .A1(n9324), .A2(n9398), .ZN(n9309) );
  OR2_X1 U11871 ( .A1(n9666), .A2(n14913), .ZN(n9308) );
  INV_X1 U11872 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9306) );
  OR2_X1 U11873 ( .A1(n9322), .A2(n9306), .ZN(n9307) );
  NAND2_X1 U11874 ( .A1(n13985), .A2(n11758), .ZN(n9316) );
  OR2_X1 U11875 ( .A1(n11567), .A2(n9312), .ZN(n9314) );
  OR2_X1 U11876 ( .A1(n9329), .A2(n8905), .ZN(n9313) );
  XNOR2_X1 U11877 ( .A(n9317), .B(n11789), .ZN(n9318) );
  INV_X2 U11878 ( .A(n11745), .ZN(n11786) );
  AOI22_X1 U11879 ( .A1(n13985), .A2(n10100), .B1(n11786), .B2(n11211), .ZN(
        n9319) );
  XNOR2_X1 U11880 ( .A(n9318), .B(n9319), .ZN(n9394) );
  NAND2_X1 U11881 ( .A1(n9393), .A2(n9394), .ZN(n9392) );
  INV_X1 U11882 ( .A(n9318), .ZN(n9320) );
  NAND2_X1 U11883 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  NAND2_X1 U11884 ( .A1(n9660), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9328) );
  OR2_X1 U11885 ( .A1(n9666), .A2(n14915), .ZN(n9326) );
  NAND2_X1 U11886 ( .A1(n9650), .A2(n11788), .ZN(n9335) );
  OR2_X1 U11887 ( .A1(n11567), .A2(n9331), .ZN(n9332) );
  NAND2_X1 U11888 ( .A1(n9708), .A2(n6571), .ZN(n9334) );
  NAND2_X1 U11889 ( .A1(n9335), .A2(n9334), .ZN(n9336) );
  XNOR2_X1 U11890 ( .A(n9336), .B(n11789), .ZN(n9879) );
  AND2_X1 U11891 ( .A1(n9708), .A2(n11786), .ZN(n9337) );
  AOI21_X1 U11892 ( .B1(n9650), .B2(n11757), .A(n9337), .ZN(n9877) );
  XNOR2_X1 U11893 ( .A(n9879), .B(n9877), .ZN(n9356) );
  AND2_X1 U11894 ( .A1(n6790), .A2(n11675), .ZN(n9359) );
  NAND3_X1 U11895 ( .A1(n14899), .A2(n9371), .A3(n11572), .ZN(n9355) );
  INV_X1 U11896 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9341) );
  INV_X1 U11897 ( .A(n9339), .ZN(n11062) );
  AND2_X1 U11898 ( .A1(n11062), .A2(n14431), .ZN(n9340) );
  INV_X1 U11899 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9343) );
  AND2_X1 U11900 ( .A1(n14431), .A2(n14432), .ZN(n9342) );
  AOI21_X1 U11901 ( .B1(n9354), .B2(n9343), .A(n9342), .ZN(n9643) );
  NOR4_X1 U11902 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9352) );
  NOR4_X1 U11903 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9351) );
  INV_X1 U11904 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15521) );
  INV_X1 U11905 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15423) );
  INV_X1 U11906 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15305) );
  INV_X1 U11907 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15402) );
  NAND4_X1 U11908 ( .A1(n15521), .A2(n15423), .A3(n15305), .A4(n15402), .ZN(
        n9349) );
  NOR4_X1 U11909 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9347) );
  NOR4_X1 U11910 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9346) );
  NOR4_X1 U11911 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9345) );
  NOR4_X1 U11912 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9344) );
  NAND4_X1 U11913 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9348)
         );
  NOR4_X1 U11914 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9349), .A4(n9348), .ZN(n9350) );
  NAND3_X1 U11915 ( .A1(n9352), .A2(n9351), .A3(n9350), .ZN(n9353) );
  NAND2_X1 U11916 ( .A1(n9354), .A2(n9353), .ZN(n9641) );
  NAND3_X1 U11917 ( .A1(n10319), .A2(n9643), .A3(n9641), .ZN(n9373) );
  OAI211_X1 U11918 ( .C1(n9357), .C2(n9356), .A(n9881), .B(n13959), .ZN(n9377)
         );
  INV_X1 U11919 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14004) );
  NAND2_X1 U11920 ( .A1(n10314), .A2(n9373), .ZN(n9360) );
  NAND2_X1 U11921 ( .A1(n9360), .A2(n9372), .ZN(n9379) );
  OAI21_X1 U11922 ( .B1(n9379), .B2(n9361), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9362) );
  INV_X1 U11923 ( .A(n9338), .ZN(n14832) );
  NAND3_X1 U11924 ( .A1(n14832), .A2(n11570), .A3(n9371), .ZN(n9363) );
  INV_X1 U11925 ( .A(n6564), .ZN(n13969) );
  NAND2_X1 U11926 ( .A1(n9660), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9368) );
  OR2_X1 U11927 ( .A1(n11494), .A2(n9364), .ZN(n9367) );
  NAND2_X1 U11928 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9664) );
  OAI21_X1 U11929 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9664), .ZN(n10081) );
  OR2_X1 U11930 ( .A1(n11390), .A2(n10081), .ZN(n9366) );
  OR2_X1 U11931 ( .A1(n11540), .A2(n14917), .ZN(n9365) );
  INV_X1 U11932 ( .A(n13984), .ZN(n9932) );
  INV_X1 U11933 ( .A(n13985), .ZN(n11209) );
  INV_X1 U11934 ( .A(n11572), .ZN(n9370) );
  OAI22_X1 U11935 ( .A1(n9932), .A2(n14189), .B1(n11209), .B2(n14191), .ZN(
        n14782) );
  NAND2_X1 U11936 ( .A1(n9372), .A2(n9371), .ZN(n11624) );
  OR2_X1 U11937 ( .A1(n11624), .A2(n9373), .ZN(n13951) );
  AOI22_X1 U11938 ( .A1(n14782), .A2(n13916), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9374) );
  OAI21_X1 U11939 ( .B1(n14852), .B2(n13969), .A(n9374), .ZN(n9375) );
  AOI21_X1 U11940 ( .B1(n14004), .B2(n13949), .A(n9375), .ZN(n9376) );
  NAND2_X1 U11941 ( .A1(n9377), .A2(n9376), .ZN(P1_U3218) );
  NOR2_X1 U11942 ( .A1(n9379), .A2(n9378), .ZN(n9399) );
  INV_X1 U11943 ( .A(n9399), .ZN(n9388) );
  AOI22_X1 U11944 ( .A1(n13959), .A2(n9380), .B1(n9388), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U11945 ( .A1(n13951), .A2(n14189), .ZN(n13966) );
  AOI22_X1 U11946 ( .A1(n13966), .A2(n13986), .B1(n6564), .B2(n14831), .ZN(
        n9381) );
  NAND2_X1 U11947 ( .A1(n9382), .A2(n9381), .ZN(P1_U3232) );
  INV_X1 U11948 ( .A(n9384), .ZN(n9385) );
  AOI21_X1 U11949 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n9391) );
  NAND2_X1 U11950 ( .A1(n13916), .A2(n14747), .ZN(n13962) );
  INV_X1 U11951 ( .A(n13962), .ZN(n13939) );
  AOI22_X1 U11952 ( .A1(n13939), .A2(n13987), .B1(n14834), .B2(n6564), .ZN(
        n9390) );
  AOI22_X1 U11953 ( .A1(n9388), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n13966), .B2(
        n13985), .ZN(n9389) );
  OAI211_X1 U11954 ( .C1(n9391), .C2(n13955), .A(n9390), .B(n9389), .ZN(
        P1_U3222) );
  OAI21_X1 U11955 ( .B1(n9394), .B2(n9393), .A(n9392), .ZN(n9395) );
  NAND2_X1 U11956 ( .A1(n9395), .A2(n13959), .ZN(n9397) );
  INV_X1 U11957 ( .A(n9298), .ZN(n11203) );
  OAI22_X1 U11958 ( .A1(n7338), .A2(n14189), .B1(n11203), .B2(n14191), .ZN(
        n9954) );
  AOI22_X1 U11959 ( .A1(n9954), .A2(n13916), .B1(n11211), .B2(n6564), .ZN(
        n9396) );
  OAI211_X1 U11960 ( .C1(n9399), .C2(n9398), .A(n9397), .B(n9396), .ZN(
        P1_U3237) );
  AOI222_X1 U11961 ( .A1(n9401), .A2(n13221), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12830), .C1(SI_16_), .C2(n9400), .ZN(n9402) );
  INV_X1 U11962 ( .A(n9402), .ZN(P3_U3279) );
  INV_X2 U11963 ( .A(n12753), .ZN(P3_U3897) );
  INV_X1 U11964 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15405) );
  NAND2_X1 U11965 ( .A1(n13063), .A2(P3_U3897), .ZN(n9403) );
  OAI21_X1 U11966 ( .B1(P3_U3897), .B2(n15405), .A(n9403), .ZN(P3_U3508) );
  INV_X1 U11967 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14565) );
  AOI22_X1 U11968 ( .A1(n10569), .A2(n14565), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n9415), .ZN(n9405) );
  NOR2_X1 U11969 ( .A1(n9406), .A2(n9405), .ZN(n9465) );
  AOI21_X1 U11970 ( .B1(n9406), .B2(n9405), .A(n9465), .ZN(n9419) );
  INV_X1 U11971 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9407) );
  AOI22_X1 U11972 ( .A1(n10569), .A2(n9407), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9415), .ZN(n9411) );
  OAI21_X1 U11973 ( .B1(n9409), .B2(n10460), .A(n9408), .ZN(n9410) );
  NOR2_X1 U11974 ( .A1(n9411), .A2(n9410), .ZN(n9468) );
  AOI21_X1 U11975 ( .B1(n9411), .B2(n9410), .A(n9468), .ZN(n9412) );
  NOR2_X1 U11976 ( .A1(n9412), .A2(n14723), .ZN(n9417) );
  NOR2_X1 U11977 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10449), .ZN(n9413) );
  AOI21_X1 U11978 ( .B1(n14731), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9413), .ZN(
        n9414) );
  OAI21_X1 U11979 ( .B1(n14725), .B2(n9415), .A(n9414), .ZN(n9416) );
  NOR2_X1 U11980 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  OAI21_X1 U11981 ( .B1(n9419), .B2(n14721), .A(n9418), .ZN(P1_U3255) );
  NAND2_X1 U11982 ( .A1(n15011), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9428) );
  MUX2_X1 U11983 ( .A(n10803), .B(P2_REG2_REG_13__SCAN_IN), .S(n15011), .Z(
        n9420) );
  INV_X1 U11984 ( .A(n9420), .ZN(n15013) );
  NOR2_X1 U11985 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n9437), .ZN(n9427) );
  NOR2_X1 U11986 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n14981), .ZN(n9426) );
  NAND2_X1 U11987 ( .A1(n9432), .A2(n10071), .ZN(n9421) );
  NAND2_X1 U11988 ( .A1(n9422), .A2(n9421), .ZN(n13410) );
  MUX2_X1 U11989 ( .A(n13412), .B(P2_REG2_REG_10__SCAN_IN), .S(n13411), .Z(
        n9423) );
  OR2_X1 U11990 ( .A1(n13410), .A2(n9423), .ZN(n13413) );
  NAND2_X1 U11991 ( .A1(n13411), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9424) );
  AND2_X1 U11992 ( .A1(n13413), .A2(n9424), .ZN(n14978) );
  INV_X1 U11993 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9425) );
  MUX2_X1 U11994 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9425), .S(n14981), .Z(
        n14977) );
  AND2_X1 U11995 ( .A1(n14978), .A2(n14977), .ZN(n14980) );
  NOR2_X1 U11996 ( .A1(n9426), .A2(n14980), .ZN(n14995) );
  AOI22_X1 U11997 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n14997), .B1(n9437), 
        .B2(n10692), .ZN(n14994) );
  NOR2_X1 U11998 ( .A1(n14995), .A2(n14994), .ZN(n14993) );
  NOR2_X1 U11999 ( .A1(n9427), .A2(n14993), .ZN(n15014) );
  NAND2_X1 U12000 ( .A1(n15013), .A2(n15014), .ZN(n15012) );
  NAND2_X1 U12001 ( .A1(n9428), .A2(n15012), .ZN(n10761) );
  XNOR2_X1 U12002 ( .A(n10761), .B(n10762), .ZN(n10763) );
  XNOR2_X1 U12003 ( .A(n10763), .B(n10865), .ZN(n9444) );
  NOR2_X1 U12004 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10818), .ZN(n9430) );
  INV_X1 U12005 ( .A(n10762), .ZN(n9857) );
  NOR2_X1 U12006 ( .A1(n14996), .A2(n9857), .ZN(n9429) );
  AOI211_X1 U12007 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n14949), .A(n9430), .B(
        n9429), .ZN(n9443) );
  INV_X1 U12008 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10877) );
  MUX2_X1 U12009 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n10877), .S(n10762), .Z(
        n9441) );
  AOI22_X1 U12010 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9437), .B1(n14997), 
        .B2(n8662), .ZN(n14992) );
  NAND2_X1 U12011 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  NAND2_X1 U12012 ( .A1(n9434), .A2(n9433), .ZN(n13404) );
  MUX2_X1 U12013 ( .A(n9435), .B(P2_REG1_REG_10__SCAN_IN), .S(n13411), .Z(
        n13403) );
  OR2_X1 U12014 ( .A1(n13404), .A2(n13403), .ZN(n13405) );
  NAND2_X1 U12015 ( .A1(n13411), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U12016 ( .A1(n13405), .A2(n9436), .ZN(n14976) );
  MUX2_X1 U12017 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8642), .S(n14981), .Z(
        n14975) );
  AND2_X1 U12018 ( .A1(n14976), .A2(n14975), .ZN(n14985) );
  AOI21_X1 U12019 ( .B1(n14981), .B2(P2_REG1_REG_11__SCAN_IN), .A(n14985), 
        .ZN(n14991) );
  NAND2_X1 U12020 ( .A1(n14992), .A2(n14991), .ZN(n14990) );
  OAI21_X1 U12021 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n9437), .A(n14990), .ZN(
        n15008) );
  INV_X1 U12022 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U12023 ( .A(n9438), .B(P2_REG1_REG_13__SCAN_IN), .S(n15011), .Z(
        n15007) );
  NOR2_X1 U12024 ( .A1(n15008), .A2(n15007), .ZN(n15006) );
  AOI21_X1 U12025 ( .B1(n15011), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15006), 
        .ZN(n9439) );
  INV_X1 U12026 ( .A(n9439), .ZN(n9440) );
  NAND2_X1 U12027 ( .A1(n9441), .A2(n9440), .ZN(n10751) );
  OAI211_X1 U12028 ( .C1(n9441), .C2(n9440), .A(n15002), .B(n10751), .ZN(n9442) );
  OAI211_X1 U12029 ( .C1(n9444), .C2(n14998), .A(n9443), .B(n9442), .ZN(
        P2_U3228) );
  INV_X1 U12030 ( .A(n10573), .ZN(n9452) );
  INV_X1 U12031 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U12032 ( .A1(n9446), .A2(n9445), .ZN(n9447) );
  NAND2_X1 U12033 ( .A1(n9447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9449) );
  INV_X1 U12034 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U12035 ( .A1(n9449), .A2(n9448), .ZN(n9858) );
  OR2_X1 U12036 ( .A1(n9449), .A2(n9448), .ZN(n9450) );
  OAI222_X1 U12037 ( .A1(n14436), .A2(n10574), .B1(n14428), .B2(n9452), .C1(
        n9863), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12038 ( .A(n15011), .ZN(n9453) );
  OAI222_X1 U12039 ( .A1(P2_U3088), .A2(n9453), .B1(n13818), .B2(n9452), .C1(
        n9451), .C2(n13820), .ZN(P2_U3314) );
  INV_X1 U12040 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n15353) );
  NAND2_X1 U12041 ( .A1(n12631), .A2(P3_U3897), .ZN(n9454) );
  OAI21_X1 U12042 ( .B1(P3_U3897), .B2(n15353), .A(n9454), .ZN(P3_U3497) );
  INV_X1 U12043 ( .A(n9455), .ZN(n9457) );
  OAI222_X1 U12044 ( .A1(n13227), .A2(n9457), .B1(n12864), .B2(P3_U3151), .C1(
        n9456), .C2(n13228), .ZN(P3_U3278) );
  XNOR2_X1 U12045 ( .A(n9459), .B(n9458), .ZN(n9463) );
  NAND2_X1 U12046 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n14965) );
  OAI21_X1 U12047 ( .B1(n14933), .B2(n12181), .A(n14965), .ZN(n9461) );
  OAI22_X1 U12048 ( .A1(n14932), .A2(n12192), .B1(n14947), .B2(n9755), .ZN(
        n9460) );
  AOI211_X1 U12049 ( .C1(n15090), .C2(n14943), .A(n9461), .B(n9460), .ZN(n9462) );
  OAI21_X1 U12050 ( .B1(n9463), .B2(n14939), .A(n9462), .ZN(P2_U3211) );
  NOR2_X1 U12051 ( .A1(n10569), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9464) );
  INV_X1 U12052 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10579) );
  MUX2_X1 U12053 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10579), .S(n10576), .Z(
        n9466) );
  NAND2_X1 U12054 ( .A1(n9467), .A2(n9466), .ZN(n9862) );
  OAI211_X1 U12055 ( .C1(n9467), .C2(n9466), .A(n14738), .B(n9862), .ZN(n9477)
         );
  NAND2_X1 U12056 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n10843)
         );
  NOR2_X1 U12057 ( .A1(n10569), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9469) );
  NOR2_X1 U12058 ( .A1(n9469), .A2(n9468), .ZN(n9473) );
  INV_X1 U12059 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9470) );
  MUX2_X1 U12060 ( .A(n9470), .B(P1_REG2_REG_13__SCAN_IN), .S(n10576), .Z(
        n9471) );
  INV_X1 U12061 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U12062 ( .A1(n9472), .A2(n9473), .ZN(n9867) );
  OAI211_X1 U12063 ( .C1(n9473), .C2(n9472), .A(n14733), .B(n9867), .ZN(n9474)
         );
  NAND2_X1 U12064 ( .A1(n10843), .A2(n9474), .ZN(n9475) );
  AOI21_X1 U12065 ( .B1(n14731), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9475), .ZN(
        n9476) );
  OAI211_X1 U12066 ( .C1(n14725), .C2(n9863), .A(n9477), .B(n9476), .ZN(
        P1_U3256) );
  INV_X1 U12067 ( .A(n12888), .ZN(n12875) );
  INV_X1 U12068 ( .A(n9478), .ZN(n9480) );
  OAI222_X1 U12069 ( .A1(n12875), .A2(P3_U3151), .B1(n13227), .B2(n9480), .C1(
        n9479), .C2(n13228), .ZN(P3_U3277) );
  XNOR2_X1 U12070 ( .A(n9481), .B(n9482), .ZN(n9488) );
  INV_X1 U12071 ( .A(n15098), .ZN(n9541) );
  NOR2_X1 U12072 ( .A1(n14947), .A2(n9538), .ZN(n9486) );
  OR2_X1 U12073 ( .A1(n12195), .A2(n15039), .ZN(n9484) );
  OR2_X1 U12074 ( .A1(n12187), .A2(n13595), .ZN(n9483) );
  AND2_X1 U12075 ( .A1(n9484), .A2(n9483), .ZN(n9521) );
  OAI22_X1 U12076 ( .A1(n9521), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8561), .ZN(n9485) );
  AOI211_X1 U12077 ( .C1(n9541), .C2(n14943), .A(n9486), .B(n9485), .ZN(n9487)
         );
  OAI21_X1 U12078 ( .B1(n9488), .B2(n14939), .A(n9487), .ZN(P2_U3185) );
  AND2_X1 U12079 ( .A1(n9489), .A2(n15053), .ZN(n10782) );
  INV_X1 U12080 ( .A(n15054), .ZN(n9490) );
  NAND2_X1 U12081 ( .A1(n10782), .A2(n9490), .ZN(n9491) );
  INV_X1 U12082 ( .A(n13677), .ZN(n13690) );
  OAI22_X1 U12083 ( .A1(n15045), .A2(n9493), .B1(n13323), .B2(n15037), .ZN(
        n9494) );
  AOI21_X1 U12084 ( .B1(n13690), .B2(n6929), .A(n9494), .ZN(n9497) );
  NOR2_X1 U12085 ( .A1(n12140), .A2(n13459), .ZN(n15044) );
  NAND2_X1 U12086 ( .A1(n15045), .A2(n15044), .ZN(n13609) );
  INV_X1 U12087 ( .A(n13609), .ZN(n9774) );
  NAND2_X1 U12088 ( .A1(n9495), .A2(n9774), .ZN(n9496) );
  OAI211_X1 U12089 ( .C1(n9498), .C2(n13639), .A(n9497), .B(n9496), .ZN(n9499)
         );
  AOI21_X1 U12090 ( .B1(n15045), .B2(n9500), .A(n9499), .ZN(n9501) );
  INV_X1 U12091 ( .A(n9501), .ZN(P2_U3264) );
  AND2_X1 U12092 ( .A1(n12754), .A2(n10496), .ZN(n11942) );
  NOR2_X1 U12093 ( .A1(n9632), .A2(n11942), .ZN(n11921) );
  NOR2_X1 U12094 ( .A1(n12731), .A2(P3_U3151), .ZN(n9921) );
  INV_X1 U12095 ( .A(n9921), .ZN(n9502) );
  NAND2_X1 U12096 ( .A1(n9502), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9506) );
  INV_X1 U12097 ( .A(n12734), .ZN(n12715) );
  INV_X1 U12098 ( .A(n12729), .ZN(n12713) );
  AOI22_X1 U12099 ( .A1(n12715), .A2(n9504), .B1(n12713), .B2(n9503), .ZN(
        n9505) );
  OAI211_X1 U12100 ( .C1(n12699), .C2(n11921), .A(n9506), .B(n9505), .ZN(
        P3_U3172) );
  OAI222_X1 U12101 ( .A1(P3_U3151), .A2(n6589), .B1(n13227), .B2(n9508), .C1(
        n9507), .C2(n13228), .ZN(P3_U3276) );
  NAND2_X1 U12102 ( .A1(n13322), .A2(n9906), .ZN(n9509) );
  INV_X1 U12103 ( .A(n9907), .ZN(n9901) );
  OR2_X1 U12104 ( .A1(n12147), .A2(n12148), .ZN(n9908) );
  NAND2_X1 U12105 ( .A1(n9510), .A2(n9908), .ZN(n9511) );
  NAND2_X1 U12106 ( .A1(n9778), .A2(n9779), .ZN(n9513) );
  AND2_X1 U12107 ( .A1(n9815), .A2(n9512), .ZN(n12405) );
  NAND2_X1 U12108 ( .A1(n9816), .A2(n9815), .ZN(n9515) );
  NAND2_X1 U12109 ( .A1(n13320), .A2(n9826), .ZN(n9514) );
  INV_X1 U12110 ( .A(n12407), .ZN(n9814) );
  NAND2_X1 U12111 ( .A1(n9515), .A2(n9814), .ZN(n9765) );
  NAND2_X1 U12112 ( .A1(n9765), .A2(n9766), .ZN(n9517) );
  NAND2_X1 U12113 ( .A1(n12181), .A2(n12179), .ZN(n9745) );
  NAND2_X1 U12114 ( .A1(n13319), .A2(n15084), .ZN(n9516) );
  NAND2_X1 U12115 ( .A1(n9745), .A2(n9516), .ZN(n12406) );
  INV_X1 U12116 ( .A(n12406), .ZN(n9759) );
  NAND2_X1 U12117 ( .A1(n9517), .A2(n9759), .ZN(n9744) );
  NAND2_X1 U12118 ( .A1(n9744), .A2(n9745), .ZN(n9518) );
  XNOR2_X1 U12119 ( .A(n15090), .B(n13318), .ZN(n12409) );
  NAND2_X1 U12120 ( .A1(n15090), .A2(n12187), .ZN(n9519) );
  NAND2_X1 U12121 ( .A1(n9748), .A2(n9519), .ZN(n9791) );
  INV_X1 U12122 ( .A(n12192), .ZN(n13317) );
  XNOR2_X1 U12123 ( .A(n9541), .B(n13317), .ZN(n12410) );
  XNOR2_X1 U12124 ( .A(n9791), .B(n12410), .ZN(n9520) );
  NAND2_X1 U12125 ( .A1(n9520), .A2(n13683), .ZN(n9522) );
  NAND2_X1 U12126 ( .A1(n9522), .A2(n9521), .ZN(n15099) );
  INV_X1 U12127 ( .A(n15099), .ZN(n9545) );
  INV_X1 U12128 ( .A(n12402), .ZN(n9524) );
  OR2_X1 U12129 ( .A1(n12147), .A2(n6929), .ZN(n9523) );
  NAND2_X1 U12130 ( .A1(n9902), .A2(n12400), .ZN(n9527) );
  OR2_X1 U12131 ( .A1(n13322), .A2(n15062), .ZN(n9526) );
  NAND2_X1 U12132 ( .A1(n9527), .A2(n9526), .ZN(n9777) );
  INV_X1 U12133 ( .A(n12405), .ZN(n9780) );
  NAND2_X1 U12134 ( .A1(n9777), .A2(n9780), .ZN(n9530) );
  NAND2_X1 U12135 ( .A1(n9528), .A2(n9536), .ZN(n9529) );
  NAND2_X1 U12136 ( .A1(n9530), .A2(n9529), .ZN(n9813) );
  NAND2_X1 U12137 ( .A1(n9813), .A2(n12407), .ZN(n9532) );
  OR2_X1 U12138 ( .A1(n13320), .A2(n15075), .ZN(n9531) );
  AND2_X1 U12139 ( .A1(n12181), .A2(n15084), .ZN(n9533) );
  OR2_X1 U12140 ( .A1(n15084), .A2(n12181), .ZN(n9534) );
  INV_X1 U12141 ( .A(n12409), .ZN(n9746) );
  NOR2_X1 U12142 ( .A1(n12188), .A2(n12187), .ZN(n9535) );
  XOR2_X1 U12143 ( .A(n9799), .B(n12410), .Z(n15101) );
  NAND2_X1 U12144 ( .A1(n15045), .A2(n15126), .ZN(n9776) );
  NAND2_X1 U12145 ( .A1(n9776), .A2(n13609), .ZN(n13644) );
  NAND2_X1 U12146 ( .A1(n9903), .A2(n9536), .ZN(n9822) );
  OR2_X1 U12147 ( .A1(n9822), .A2(n15075), .ZN(n9823) );
  AND2_X1 U12148 ( .A1(n9762), .A2(n12188), .ZN(n9753) );
  INV_X1 U12149 ( .A(n9806), .ZN(n9537) );
  OAI211_X1 U12150 ( .C1(n15098), .C2(n9753), .A(n9537), .B(n6577), .ZN(n15096) );
  OAI22_X1 U12151 ( .A1(n15045), .A2(n9539), .B1(n9538), .B2(n15037), .ZN(
        n9540) );
  AOI21_X1 U12152 ( .B1(n13690), .B2(n9541), .A(n9540), .ZN(n9542) );
  OAI21_X1 U12153 ( .B1(n15096), .B2(n13639), .A(n9542), .ZN(n9543) );
  AOI21_X1 U12154 ( .B1(n15101), .B2(n13644), .A(n9543), .ZN(n9544) );
  OAI21_X1 U12155 ( .B1(n6578), .B2(n9545), .A(n9544), .ZN(P2_U3258) );
  MUX2_X1 U12156 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12862), .Z(n9579) );
  XOR2_X1 U12157 ( .A(n9593), .B(n9579), .Z(n9582) );
  INV_X1 U12158 ( .A(n9567), .ZN(n9723) );
  INV_X1 U12159 ( .A(n9546), .ZN(n9547) );
  XNOR2_X1 U12160 ( .A(n9546), .B(n9567), .ZN(n9715) );
  INV_X1 U12161 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10493) );
  INV_X1 U12162 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9854) );
  MUX2_X1 U12163 ( .A(n10493), .B(n9854), .S(n9555), .Z(n10294) );
  MUX2_X1 U12164 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12862), .Z(n9548) );
  XNOR2_X1 U12165 ( .A(n9548), .B(n9981), .ZN(n9976) );
  OAI22_X1 U12166 ( .A1(n9977), .A2(n9976), .B1(n9548), .B2(n9981), .ZN(n9583)
         );
  XOR2_X1 U12167 ( .A(n9582), .B(n9583), .Z(n9578) );
  INV_X1 U12168 ( .A(n9843), .ZN(n9549) );
  OR2_X1 U12169 ( .A1(n9550), .A2(P3_U3151), .ZN(n12110) );
  NAND2_X1 U12170 ( .A1(n9549), .A2(n12110), .ZN(n9564) );
  NAND2_X1 U12171 ( .A1(n9550), .A2(n12076), .ZN(n9551) );
  NAND2_X1 U12172 ( .A1(n9552), .A2(n9551), .ZN(n9563) );
  INV_X1 U12173 ( .A(n9563), .ZN(n9553) );
  NAND2_X1 U12174 ( .A1(n9564), .A2(n9553), .ZN(n9566) );
  MUX2_X1 U12175 ( .A(n9566), .B(n12753), .S(n9554), .Z(n12883) );
  INV_X1 U12176 ( .A(n9566), .ZN(n9556) );
  INV_X1 U12177 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9557) );
  OR2_X1 U12178 ( .A1(n9567), .A2(n9558), .ZN(n9559) );
  NAND2_X1 U12179 ( .A1(n7660), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U12180 ( .A1(n9559), .A2(n9560), .ZN(n9716) );
  INV_X1 U12181 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9561) );
  OAI21_X1 U12182 ( .B1(n9716), .B2(n9561), .A(n9560), .ZN(n9969) );
  NAND2_X1 U12183 ( .A1(n9981), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U12184 ( .A1(n9968), .A2(n9562), .ZN(n9594) );
  XNOR2_X1 U12185 ( .A(n9594), .B(n9581), .ZN(n9592) );
  XOR2_X1 U12186 ( .A(n9592), .B(P3_REG1_REG_3__SCAN_IN), .Z(n9575) );
  NOR2_X1 U12187 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12582), .ZN(n12580) );
  AOI21_X1 U12188 ( .B1(n15142), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n12580), .ZN(
        n9574) );
  OR2_X1 U12189 ( .A1(n9566), .A2(n9565), .ZN(n12896) );
  INV_X1 U12190 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15180) );
  NAND2_X1 U12191 ( .A1(n7660), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9568) );
  OAI21_X1 U12192 ( .B1(n9567), .B2(n10299), .A(n9568), .ZN(n9717) );
  INV_X1 U12193 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15200) );
  OR2_X1 U12194 ( .A1(n9717), .A2(n15200), .ZN(n9719) );
  NAND2_X1 U12195 ( .A1(n9719), .A2(n9568), .ZN(n9966) );
  NAND2_X1 U12196 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  NAND2_X1 U12197 ( .A1(n9981), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U12198 ( .A1(n9570), .A2(n9593), .ZN(n9613) );
  OAI21_X1 U12199 ( .B1(n9571), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9615), .ZN(
        n9572) );
  NAND2_X1 U12200 ( .A1(n12819), .A2(n9572), .ZN(n9573) );
  OAI211_X1 U12201 ( .C1(n10243), .C2(n9575), .A(n9574), .B(n9573), .ZN(n9576)
         );
  AOI21_X1 U12202 ( .B1(n9581), .B2(n12834), .A(n9576), .ZN(n9577) );
  OAI21_X1 U12203 ( .B1(n9578), .B2(n12891), .A(n9577), .ZN(P3_U3185) );
  INV_X1 U12204 ( .A(n9579), .ZN(n9580) );
  MUX2_X1 U12205 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12862), .Z(n9584) );
  XNOR2_X1 U12206 ( .A(n9584), .B(n9598), .ZN(n9608) );
  MUX2_X1 U12207 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12862), .Z(n9586) );
  NAND2_X1 U12208 ( .A1(n9586), .A2(n9585), .ZN(n9589) );
  NAND2_X1 U12209 ( .A1(n9588), .A2(n9589), .ZN(n9987) );
  INV_X1 U12210 ( .A(n9987), .ZN(n9591) );
  INV_X1 U12211 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U12212 ( .A1(n9587), .A2(n9991), .ZN(n9986) );
  AOI21_X1 U12213 ( .B1(n9986), .B2(n9589), .A(n9588), .ZN(n9590) );
  AOI21_X1 U12214 ( .B1(n9591), .B2(n9986), .A(n9590), .ZN(n9606) );
  NAND2_X1 U12215 ( .A1(n9592), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12216 ( .A1(n9594), .A2(n9593), .ZN(n9595) );
  NAND2_X1 U12217 ( .A1(n9596), .A2(n9595), .ZN(n9610) );
  INV_X1 U12218 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9597) );
  MUX2_X1 U12219 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n9597), .S(n9598), .Z(n9609)
         );
  AND2_X1 U12220 ( .A1(n9610), .A2(n9609), .ZN(n9612) );
  XNOR2_X1 U12221 ( .A(n9990), .B(n9991), .ZN(n9992) );
  XNOR2_X1 U12222 ( .A(n9992), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n9603) );
  AND2_X1 U12223 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n12630) );
  AOI21_X1 U12224 ( .B1(n15142), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n12630), .ZN(
        n9602) );
  XNOR2_X1 U12225 ( .A(n9598), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n9614) );
  OAI21_X1 U12226 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n9599), .A(n9998), .ZN(
        n9600) );
  NAND2_X1 U12227 ( .A1(n12819), .A2(n9600), .ZN(n9601) );
  OAI211_X1 U12228 ( .C1(n10243), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9604)
         );
  AOI21_X1 U12229 ( .B1(n9991), .B2(n12834), .A(n9604), .ZN(n9605) );
  OAI21_X1 U12230 ( .B1(n9606), .B2(n12891), .A(n9605), .ZN(P3_U3187) );
  XOR2_X1 U12231 ( .A(n9608), .B(n9607), .Z(n9624) );
  NOR2_X1 U12232 ( .A1(n9610), .A2(n9609), .ZN(n9611) );
  OAI21_X1 U12233 ( .B1(n9612), .B2(n9611), .A(n12895), .ZN(n9620) );
  AND3_X1 U12234 ( .A1(n9615), .A2(n9614), .A3(n9613), .ZN(n9616) );
  OAI21_X1 U12235 ( .B1(n9617), .B2(n9616), .A(n12819), .ZN(n9619) );
  AND2_X1 U12236 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n12662) );
  AOI21_X1 U12237 ( .B1(n15142), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n12662), .ZN(
        n9618) );
  NAND3_X1 U12238 ( .A1(n9620), .A2(n9619), .A3(n9618), .ZN(n9621) );
  AOI21_X1 U12239 ( .B1(n9622), .B2(n12834), .A(n9621), .ZN(n9623) );
  OAI21_X1 U12240 ( .B1(n9624), .B2(n12891), .A(n9623), .ZN(P3_U3186) );
  INV_X1 U12241 ( .A(n15024), .ZN(n10769) );
  INV_X1 U12242 ( .A(n11331), .ZN(n9628) );
  OAI222_X1 U12243 ( .A1(P2_U3088), .A2(n10769), .B1(n13818), .B2(n9628), .C1(
        n9625), .C2(n13820), .ZN(P2_U3311) );
  NAND2_X1 U12244 ( .A1(n9626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9627) );
  XNOR2_X1 U12245 ( .A(n9627), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11332) );
  INV_X1 U12246 ( .A(n11332), .ZN(n11666) );
  OAI222_X1 U12247 ( .A1(n14436), .A2(n9629), .B1(n14428), .B2(n9628), .C1(
        n11666), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12248 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15185) );
  INV_X1 U12249 ( .A(n12726), .ZN(n12685) );
  INV_X1 U12250 ( .A(n12754), .ZN(n15194) );
  OAI22_X1 U12251 ( .A1(n12685), .A2(n15194), .B1(n15192), .B2(n12729), .ZN(
        n9630) );
  AOI21_X1 U12252 ( .B1(n12715), .B2(n9633), .A(n9630), .ZN(n9640) );
  INV_X1 U12253 ( .A(n9632), .ZN(n15182) );
  NAND3_X1 U12254 ( .A1(n15182), .A2(n15181), .A3(n7752), .ZN(n9636) );
  OAI211_X1 U12255 ( .C1(n9637), .C2(n15188), .A(n9631), .B(n9636), .ZN(n9638)
         );
  NAND2_X1 U12256 ( .A1(n9638), .A2(n12724), .ZN(n9639) );
  OAI211_X1 U12257 ( .C1(n9921), .C2(n15185), .A(n9640), .B(n9639), .ZN(
        P3_U3162) );
  INV_X1 U12258 ( .A(n9641), .ZN(n9642) );
  INV_X1 U12259 ( .A(n9643), .ZN(n10313) );
  NOR2_X1 U12260 ( .A1(n10313), .A2(n10319), .ZN(n9644) );
  NAND2_X1 U12261 ( .A1(n10315), .A2(n9644), .ZN(n14103) );
  NOR2_X1 U12262 ( .A1(n11195), .A2(n11190), .ZN(n9645) );
  OR2_X1 U12263 ( .A1(n9645), .A2(n11692), .ZN(n9646) );
  AND2_X1 U12264 ( .A1(n13987), .A2(n14831), .ZN(n9728) );
  OR2_X1 U12265 ( .A1(n9298), .A2(n14834), .ZN(n11204) );
  INV_X1 U12266 ( .A(n11587), .ZN(n9647) );
  NAND2_X1 U12267 ( .A1(n9952), .A2(n9647), .ZN(n9649) );
  OR2_X1 U12268 ( .A1(n13985), .A2(n11211), .ZN(n9648) );
  NAND2_X1 U12269 ( .A1(n9649), .A2(n9648), .ZN(n14777) );
  NAND2_X1 U12270 ( .A1(n14777), .A2(n14778), .ZN(n9652) );
  OR2_X1 U12271 ( .A1(n9650), .A2(n9708), .ZN(n9651) );
  NAND2_X1 U12272 ( .A1(n9652), .A2(n9651), .ZN(n10085) );
  NAND2_X1 U12273 ( .A1(n11565), .A2(n9653), .ZN(n9656) );
  NAND2_X1 U12274 ( .A1(n11338), .A2(n9654), .ZN(n9655) );
  NAND2_X1 U12275 ( .A1(n10085), .A2(n11590), .ZN(n9659) );
  OR2_X1 U12276 ( .A1(n13984), .A2(n14860), .ZN(n9658) );
  NAND2_X1 U12277 ( .A1(n11387), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9670) );
  OR2_X1 U12278 ( .A1(n6573), .A2(n9661), .ZN(n9669) );
  INV_X1 U12279 ( .A(n9664), .ZN(n9662) );
  NAND2_X1 U12280 ( .A1(n9662), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9676) );
  INV_X1 U12281 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12282 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  NAND2_X1 U12283 ( .A1(n9676), .A2(n9665), .ZN(n14768) );
  OR2_X1 U12284 ( .A1(n11390), .A2(n14768), .ZN(n9668) );
  OR2_X1 U12285 ( .A1(n11540), .A2(n14919), .ZN(n9667) );
  NAND4_X2 U12286 ( .A1(n9670), .A2(n9669), .A3(n9668), .A4(n9667), .ZN(n13983) );
  AOI22_X1 U12287 ( .A1(n11519), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11338), 
        .B2(n14027), .ZN(n9673) );
  OR2_X1 U12288 ( .A1(n9671), .A2(n11381), .ZN(n9672) );
  NAND2_X1 U12289 ( .A1(n9673), .A2(n9672), .ZN(n11227) );
  XNOR2_X2 U12290 ( .A(n13983), .B(n14868), .ZN(n14764) );
  INV_X1 U12291 ( .A(n13983), .ZN(n9693) );
  NAND2_X1 U12292 ( .A1(n9693), .A2(n14868), .ZN(n9674) );
  NAND2_X1 U12293 ( .A1(n11387), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9681) );
  OR2_X1 U12294 ( .A1(n6573), .A2(n9707), .ZN(n9680) );
  INV_X1 U12295 ( .A(n9676), .ZN(n9675) );
  NAND2_X1 U12296 ( .A1(n9675), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U12297 ( .A1(n9676), .A2(n9097), .ZN(n9677) );
  NAND2_X1 U12298 ( .A1(n9699), .A2(n9677), .ZN(n10106) );
  OR2_X1 U12299 ( .A1(n11491), .A2(n10106), .ZN(n9679) );
  OR2_X1 U12300 ( .A1(n11540), .A2(n14921), .ZN(n9678) );
  OR2_X1 U12301 ( .A1(n9682), .A2(n11381), .ZN(n9685) );
  AOI22_X1 U12302 ( .A1(n11519), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11338), 
        .B2(n9683), .ZN(n9684) );
  INV_X1 U12303 ( .A(n11591), .ZN(n10147) );
  XNOR2_X1 U12304 ( .A(n10112), .B(n10147), .ZN(n14878) );
  INV_X1 U12305 ( .A(n14834), .ZN(n11202) );
  AND2_X1 U12306 ( .A1(n13986), .A2(n11202), .ZN(n9686) );
  INV_X1 U12307 ( .A(n14831), .ZN(n11196) );
  OAI22_X1 U12308 ( .A1(n9686), .A2(n11200), .B1(n11202), .B2(n13986), .ZN(
        n9953) );
  NAND2_X1 U12309 ( .A1(n9953), .A2(n11587), .ZN(n9687) );
  NAND2_X1 U12310 ( .A1(n9688), .A2(n11213), .ZN(n10079) );
  NAND2_X1 U12311 ( .A1(n9689), .A2(n10079), .ZN(n9691) );
  OR2_X1 U12312 ( .A1(n13984), .A2(n10082), .ZN(n9690) );
  NAND2_X1 U12313 ( .A1(n9691), .A2(n9690), .ZN(n14763) );
  INV_X1 U12314 ( .A(n14764), .ZN(n9692) );
  NAND2_X1 U12315 ( .A1(n14763), .A2(n9692), .ZN(n9695) );
  NAND2_X1 U12316 ( .A1(n9693), .A2(n11227), .ZN(n9694) );
  NAND2_X1 U12317 ( .A1(n9695), .A2(n9694), .ZN(n10148) );
  XNOR2_X1 U12318 ( .A(n10148), .B(n11591), .ZN(n9705) );
  NAND2_X1 U12319 ( .A1(n10306), .A2(n11573), .ZN(n9697) );
  NAND2_X1 U12320 ( .A1(n9247), .A2(n11570), .ZN(n9696) );
  NAND2_X1 U12321 ( .A1(n11387), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9704) );
  OR2_X1 U12322 ( .A1(n6573), .A2(n9698), .ZN(n9703) );
  NAND2_X1 U12323 ( .A1(n9699), .A2(n10287), .ZN(n9700) );
  NAND2_X1 U12324 ( .A1(n10128), .A2(n9700), .ZN(n14754) );
  OR2_X1 U12325 ( .A1(n11390), .A2(n14754), .ZN(n9702) );
  OR2_X1 U12326 ( .A1(n11540), .A2(n14923), .ZN(n9701) );
  NAND4_X1 U12327 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n13982) );
  AOI22_X1 U12328 ( .A1(n14750), .A2(n13982), .B1(n13983), .B2(n14747), .ZN(
        n10101) );
  OAI21_X1 U12329 ( .B1(n9705), .B2(n14863), .A(n10101), .ZN(n14873) );
  INV_X1 U12330 ( .A(n14873), .ZN(n9706) );
  MUX2_X1 U12331 ( .A(n9707), .B(n9706), .S(n14301), .Z(n9713) );
  NOR2_X1 U12332 ( .A1(n14834), .A2(n14831), .ZN(n9956) );
  NAND2_X1 U12333 ( .A1(n9956), .A2(n14847), .ZN(n14788) );
  OR2_X1 U12334 ( .A1(n14788), .A2(n9708), .ZN(n14789) );
  AND2_X1 U12335 ( .A1(n14773), .A2(n14868), .ZN(n9709) );
  INV_X1 U12336 ( .A(n9709), .ZN(n14772) );
  INV_X1 U12337 ( .A(n14875), .ZN(n10113) );
  AOI211_X1 U12338 ( .C1(n14875), .C2(n14772), .A(n14837), .B(n6731), .ZN(
        n14874) );
  OR2_X1 U12339 ( .A1(n9338), .A2(n6790), .ZN(n9710) );
  OAI22_X1 U12340 ( .A1(n14786), .A2(n10113), .B1(n10106), .B2(n14783), .ZN(
        n9711) );
  AOI21_X1 U12341 ( .B1(n14874), .B2(n14793), .A(n9711), .ZN(n9712) );
  OAI211_X1 U12342 ( .C1(n14292), .C2(n14878), .A(n9713), .B(n9712), .ZN(
        P1_U3287) );
  AOI21_X1 U12343 ( .B1(n9715), .B2(n10302), .A(n9714), .ZN(n9726) );
  XOR2_X1 U12344 ( .A(n9716), .B(P3_REG1_REG_1__SCAN_IN), .Z(n9722) );
  OAI22_X1 U12345 ( .A1(n12837), .A2(n14441), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15185), .ZN(n9721) );
  NAND2_X1 U12346 ( .A1(n9717), .A2(n15200), .ZN(n9718) );
  AOI21_X1 U12347 ( .B1(n9719), .B2(n9718), .A(n12896), .ZN(n9720) );
  AOI211_X1 U12348 ( .C1(n12895), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9725)
         );
  NAND2_X1 U12349 ( .A1(n12834), .A2(n9723), .ZN(n9724) );
  OAI211_X1 U12350 ( .C1(n9726), .C2(n12891), .A(n9725), .B(n9724), .ZN(
        P3_U3183) );
  XOR2_X1 U12351 ( .A(n9728), .B(n9727), .Z(n14833) );
  NOR2_X1 U12352 ( .A1(n14273), .A2(n14837), .ZN(n14145) );
  INV_X1 U12353 ( .A(n14145), .ZN(n14087) );
  INV_X1 U12354 ( .A(n9956), .ZN(n9730) );
  NAND2_X1 U12355 ( .A1(n14834), .A2(n14831), .ZN(n9729) );
  NAND2_X1 U12356 ( .A1(n9730), .A2(n9729), .ZN(n14838) );
  OAI22_X1 U12357 ( .A1(n14087), .A2(n14838), .B1(n9731), .B2(n14783), .ZN(
        n9732) );
  AOI21_X1 U12358 ( .B1(n14303), .B2(n14834), .A(n9732), .ZN(n9742) );
  XNOR2_X1 U12359 ( .A(n14838), .B(n13986), .ZN(n9733) );
  NAND2_X1 U12360 ( .A1(n9733), .A2(n14902), .ZN(n9735) );
  INV_X1 U12361 ( .A(n13987), .ZN(n9734) );
  NAND2_X1 U12362 ( .A1(n9735), .A2(n9734), .ZN(n9738) );
  AOI21_X1 U12363 ( .B1(n9727), .B2(n13987), .A(n14863), .ZN(n9736) );
  OR2_X1 U12364 ( .A1(n9736), .A2(n14747), .ZN(n9737) );
  NAND2_X1 U12365 ( .A1(n9738), .A2(n9737), .ZN(n14839) );
  NAND2_X1 U12366 ( .A1(n13985), .A2(n14750), .ZN(n14836) );
  NAND2_X1 U12367 ( .A1(n14839), .A2(n14836), .ZN(n9739) );
  MUX2_X1 U12368 ( .A(n9739), .B(P1_REG2_REG_1__SCAN_IN), .S(n14797), .Z(n9740) );
  INV_X1 U12369 ( .A(n9740), .ZN(n9741) );
  OAI211_X1 U12370 ( .C1(n14292), .C2(n14833), .A(n9742), .B(n9741), .ZN(
        P1_U3292) );
  XNOR2_X1 U12371 ( .A(n9743), .B(n12409), .ZN(n9751) );
  INV_X1 U12372 ( .A(n9751), .ZN(n15093) );
  OAI22_X1 U12373 ( .A1(n12181), .A2(n13595), .B1(n12192), .B2(n15039), .ZN(
        n9750) );
  NAND3_X1 U12374 ( .A1(n9744), .A2(n9746), .A3(n9745), .ZN(n9747) );
  AOI21_X1 U12375 ( .B1(n9748), .B2(n9747), .A(n10902), .ZN(n9749) );
  AOI211_X1 U12376 ( .C1(n15126), .C2(n9751), .A(n9750), .B(n9749), .ZN(n15092) );
  MUX2_X1 U12377 ( .A(n9752), .B(n15092), .S(n15045), .Z(n9758) );
  OAI21_X1 U12378 ( .B1(n9762), .B2(n12188), .A(n6577), .ZN(n9754) );
  NOR2_X1 U12379 ( .A1(n9754), .A2(n9753), .ZN(n15089) );
  OAI22_X1 U12380 ( .A1(n13677), .A2(n12188), .B1(n15037), .B2(n9755), .ZN(
        n9756) );
  AOI21_X1 U12381 ( .B1(n15089), .B2(n13694), .A(n9756), .ZN(n9757) );
  OAI211_X1 U12382 ( .C1(n15093), .C2(n13609), .A(n9758), .B(n9757), .ZN(
        P2_U3259) );
  XNOR2_X1 U12383 ( .A(n9760), .B(n9759), .ZN(n9771) );
  INV_X1 U12384 ( .A(n9771), .ZN(n15087) );
  NAND2_X1 U12385 ( .A1(n9823), .A2(n12179), .ZN(n9761) );
  NAND2_X1 U12386 ( .A1(n9761), .A2(n6577), .ZN(n9763) );
  OR2_X1 U12387 ( .A1(n9763), .A2(n9762), .ZN(n15083) );
  INV_X1 U12388 ( .A(n15037), .ZN(n13673) );
  AOI22_X1 U12389 ( .A1(n13690), .A2(n12179), .B1(n13673), .B2(n13264), .ZN(
        n9764) );
  OAI21_X1 U12390 ( .B1(n13639), .B2(n15083), .A(n9764), .ZN(n9773) );
  INV_X1 U12391 ( .A(n9744), .ZN(n9768) );
  AND3_X1 U12392 ( .A1(n9765), .A2(n9766), .A3(n12406), .ZN(n9767) );
  INV_X2 U12393 ( .A(n10902), .ZN(n13683) );
  OAI21_X1 U12394 ( .B1(n9768), .B2(n9767), .A(n13683), .ZN(n9770) );
  AOI22_X1 U12395 ( .A1(n13318), .A2(n13665), .B1(n13667), .B2(n13320), .ZN(
        n9769) );
  OAI211_X1 U12396 ( .C1(n9771), .C2(n9127), .A(n9770), .B(n9769), .ZN(n15085)
         );
  MUX2_X1 U12397 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15085), .S(n15045), .Z(
        n9772) );
  AOI211_X1 U12398 ( .C1(n9774), .C2(n15087), .A(n9773), .B(n9772), .ZN(n9775)
         );
  INV_X1 U12399 ( .A(n9775), .ZN(P2_U3260) );
  AND2_X1 U12400 ( .A1(n13609), .A2(n9776), .ZN(n13540) );
  XNOR2_X1 U12401 ( .A(n9777), .B(n12405), .ZN(n15072) );
  NAND3_X1 U12402 ( .A1(n9778), .A2(n9780), .A3(n9779), .ZN(n9781) );
  AND2_X1 U12403 ( .A1(n9816), .A2(n9781), .ZN(n9783) );
  OAI21_X1 U12404 ( .B1(n9783), .B2(n10902), .A(n9782), .ZN(n15068) );
  AOI21_X1 U12405 ( .B1(n13673), .B2(n15314), .A(n15068), .ZN(n9784) );
  MUX2_X1 U12406 ( .A(n9785), .B(n9784), .S(n15045), .Z(n9789) );
  INV_X1 U12407 ( .A(n9903), .ZN(n9787) );
  INV_X1 U12408 ( .A(n9822), .ZN(n9786) );
  AOI211_X1 U12409 ( .C1(n15070), .C2(n9787), .A(n8705), .B(n9786), .ZN(n15069) );
  AOI22_X1 U12410 ( .A1(n15069), .A2(n13694), .B1(n13690), .B2(n15070), .ZN(
        n9788) );
  OAI211_X1 U12411 ( .C1(n13540), .C2(n15072), .A(n9789), .B(n9788), .ZN(
        P2_U3262) );
  NAND2_X1 U12412 ( .A1(n15098), .A2(n13317), .ZN(n9790) );
  NAND2_X1 U12413 ( .A1(n9791), .A2(n9790), .ZN(n9793) );
  OR2_X1 U12414 ( .A1(n15098), .A2(n13317), .ZN(n9792) );
  NAND2_X1 U12415 ( .A1(n9793), .A2(n9792), .ZN(n10058) );
  INV_X1 U12416 ( .A(n12195), .ZN(n13316) );
  XNOR2_X1 U12417 ( .A(n15103), .B(n13316), .ZN(n12412) );
  XNOR2_X1 U12418 ( .A(n10058), .B(n12412), .ZN(n9794) );
  NAND2_X1 U12419 ( .A1(n9794), .A2(n13683), .ZN(n9797) );
  OR2_X1 U12420 ( .A1(n12192), .A2(n13595), .ZN(n9796) );
  NAND2_X1 U12421 ( .A1(n13315), .A2(n13665), .ZN(n9795) );
  AND2_X1 U12422 ( .A1(n9796), .A2(n9795), .ZN(n9947) );
  NAND2_X1 U12423 ( .A1(n9797), .A2(n9947), .ZN(n15108) );
  INV_X1 U12424 ( .A(n15108), .ZN(n9812) );
  OR2_X1 U12425 ( .A1(n15098), .A2(n12192), .ZN(n9798) );
  NAND2_X1 U12426 ( .A1(n9799), .A2(n9798), .ZN(n9801) );
  NAND2_X1 U12427 ( .A1(n15098), .A2(n12192), .ZN(n9800) );
  NAND2_X1 U12428 ( .A1(n9801), .A2(n9800), .ZN(n9804) );
  INV_X1 U12429 ( .A(n9804), .ZN(n9803) );
  NAND2_X1 U12430 ( .A1(n9804), .A2(n12412), .ZN(n9805) );
  NAND2_X1 U12431 ( .A1(n10066), .A2(n9805), .ZN(n15106) );
  INV_X1 U12432 ( .A(n15106), .ZN(n15109) );
  INV_X1 U12433 ( .A(n13540), .ZN(n10268) );
  OAI211_X1 U12434 ( .C1(n9806), .C2(n12196), .A(n6577), .B(n10069), .ZN(
        n15105) );
  OAI22_X1 U12435 ( .A1(n15045), .A2(n9807), .B1(n9946), .B2(n15037), .ZN(
        n9808) );
  AOI21_X1 U12436 ( .B1(n15103), .B2(n13690), .A(n9808), .ZN(n9809) );
  OAI21_X1 U12437 ( .B1(n15105), .B2(n13639), .A(n9809), .ZN(n9810) );
  AOI21_X1 U12438 ( .B1(n15109), .B2(n10268), .A(n9810), .ZN(n9811) );
  OAI21_X1 U12439 ( .B1(n9812), .B2(n6578), .A(n9811), .ZN(P2_U3257) );
  XNOR2_X1 U12440 ( .A(n9814), .B(n9813), .ZN(n15079) );
  NAND3_X1 U12441 ( .A1(n9816), .A2(n12407), .A3(n9815), .ZN(n9817) );
  NAND2_X1 U12442 ( .A1(n9765), .A2(n9817), .ZN(n9820) );
  NAND2_X1 U12443 ( .A1(n13321), .A2(n13667), .ZN(n9818) );
  OAI21_X1 U12444 ( .B1(n12181), .B2(n15039), .A(n9818), .ZN(n9819) );
  AOI21_X1 U12445 ( .B1(n9820), .B2(n13683), .A(n9819), .ZN(n15082) );
  MUX2_X1 U12446 ( .A(n9821), .B(n15082), .S(n15045), .Z(n9829) );
  AOI21_X1 U12447 ( .B1(n9822), .B2(n15075), .A(n8705), .ZN(n9824) );
  AND2_X1 U12448 ( .A1(n9824), .A2(n9823), .ZN(n15077) );
  OAI22_X1 U12449 ( .A1(n13677), .A2(n9826), .B1(n15037), .B2(n9825), .ZN(
        n9827) );
  AOI21_X1 U12450 ( .B1(n13694), .B2(n15077), .A(n9827), .ZN(n9828) );
  OAI211_X1 U12451 ( .C1(n13697), .C2(n15079), .A(n9829), .B(n9828), .ZN(
        P2_U3261) );
  INV_X1 U12452 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n15479) );
  NAND2_X1 U12453 ( .A1(n12727), .A2(P3_U3897), .ZN(n9830) );
  OAI21_X1 U12454 ( .B1(P3_U3897), .B2(n15479), .A(n9830), .ZN(P3_U3516) );
  NAND2_X1 U12455 ( .A1(n12106), .A2(n9831), .ZN(n9832) );
  NAND2_X1 U12456 ( .A1(n9833), .A2(n9832), .ZN(n9837) );
  NAND3_X1 U12457 ( .A1(n9835), .A2(n9843), .A3(n9834), .ZN(n9836) );
  OR3_X1 U12458 ( .A1(n11921), .A2(n15210), .A3(n9838), .ZN(n9840) );
  OR2_X1 U12459 ( .A1(n15168), .A2(n15193), .ZN(n9839) );
  AND2_X1 U12460 ( .A1(n9840), .A2(n9839), .ZN(n10491) );
  INV_X1 U12461 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n15338) );
  MUX2_X1 U12462 ( .A(n10491), .B(n15338), .S(n15223), .Z(n9841) );
  OAI21_X1 U12463 ( .B1(n10496), .B2(n13212), .A(n9841), .ZN(P3_U3390) );
  XNOR2_X1 U12464 ( .A(n9842), .B(n13214), .ZN(n9846) );
  AND2_X1 U12465 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  NAND3_X1 U12466 ( .A1(n6589), .A2(n10205), .A3(n12107), .ZN(n9847) );
  NAND2_X1 U12467 ( .A1(n9847), .A2(n12087), .ZN(n10343) );
  OAI22_X1 U12468 ( .A1(n11936), .A2(n9849), .B1(n10205), .B2(n15183), .ZN(
        n9850) );
  AOI21_X1 U12469 ( .B1(n9850), .B2(n12092), .A(n12076), .ZN(n9852) );
  INV_X1 U12470 ( .A(n13214), .ZN(n9851) );
  MUX2_X1 U12471 ( .A(n10345), .B(n9852), .S(n9851), .Z(n9853) );
  NAND2_X1 U12472 ( .A1(n15235), .A2(n15210), .ZN(n13163) );
  MUX2_X1 U12473 ( .A(n10491), .B(n9854), .S(n15233), .Z(n9855) );
  OAI21_X1 U12474 ( .B1(n10496), .B2(n13163), .A(n9855), .ZN(P3_U3459) );
  INV_X1 U12475 ( .A(n11280), .ZN(n9861) );
  OAI222_X1 U12476 ( .A1(P2_U3088), .A2(n9857), .B1(n13818), .B2(n9861), .C1(
        n9856), .C2(n13820), .ZN(P2_U3313) );
  NAND2_X1 U12477 ( .A1(n9858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9859) );
  OAI222_X1 U12478 ( .A1(P1_U3086), .A2(n10504), .B1(n14428), .B2(n9861), .C1(
        n9860), .C2(n14436), .ZN(P1_U3341) );
  INV_X1 U12479 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15332) );
  AOI22_X1 U12480 ( .A1(n11281), .A2(n15332), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10504), .ZN(n9865) );
  OAI21_X1 U12481 ( .B1(n9863), .B2(n10579), .A(n9862), .ZN(n9864) );
  NOR2_X1 U12482 ( .A1(n9865), .A2(n9864), .ZN(n10497) );
  AOI21_X1 U12483 ( .B1(n9865), .B2(n9864), .A(n10497), .ZN(n9873) );
  INV_X1 U12484 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15504) );
  NAND2_X1 U12485 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13837)
         );
  OAI21_X1 U12486 ( .B1(n14729), .B2(n15504), .A(n13837), .ZN(n9866) );
  AOI21_X1 U12487 ( .B1(n11281), .B2(n14736), .A(n9866), .ZN(n9872) );
  NAND2_X1 U12488 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10576), .ZN(n9868) );
  NAND2_X1 U12489 ( .A1(n9868), .A2(n9867), .ZN(n9870) );
  INV_X1 U12490 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14300) );
  MUX2_X1 U12491 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14300), .S(n11281), .Z(
        n9869) );
  NAND2_X1 U12492 ( .A1(n9869), .A2(n9870), .ZN(n10503) );
  OAI211_X1 U12493 ( .C1(n9870), .C2(n9869), .A(n14733), .B(n10503), .ZN(n9871) );
  OAI211_X1 U12494 ( .C1(n9873), .C2(n14721), .A(n9872), .B(n9871), .ZN(
        P1_U3257) );
  NAND2_X1 U12495 ( .A1(n13984), .A2(n11788), .ZN(n9875) );
  NAND2_X1 U12496 ( .A1(n14860), .A2(n11787), .ZN(n9874) );
  NAND2_X1 U12497 ( .A1(n9875), .A2(n9874), .ZN(n9876) );
  XNOR2_X1 U12498 ( .A(n9876), .B(n11692), .ZN(n9888) );
  INV_X1 U12499 ( .A(n9877), .ZN(n9878) );
  NAND2_X1 U12500 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  NAND2_X1 U12501 ( .A1(n9881), .A2(n9880), .ZN(n9886) );
  NAND2_X1 U12502 ( .A1(n13984), .A2(n11757), .ZN(n9883) );
  NAND2_X1 U12503 ( .A1(n14860), .A2(n11788), .ZN(n9882) );
  NAND2_X1 U12504 ( .A1(n9883), .A2(n9882), .ZN(n9885) );
  OAI21_X1 U12505 ( .B1(n9888), .B2(n9887), .A(n9923), .ZN(n9889) );
  NAND2_X1 U12506 ( .A1(n9889), .A2(n13959), .ZN(n9895) );
  NAND2_X1 U12507 ( .A1(n9650), .A2(n14747), .ZN(n9891) );
  NAND2_X1 U12508 ( .A1(n13983), .A2(n14750), .ZN(n9890) );
  AND2_X1 U12509 ( .A1(n9891), .A2(n9890), .ZN(n10080) );
  OAI21_X1 U12510 ( .B1(n10080), .B2(n13951), .A(n9892), .ZN(n9893) );
  AOI21_X1 U12511 ( .B1(n14860), .B2(n6564), .A(n9893), .ZN(n9894) );
  OAI211_X1 U12512 ( .C1(n13963), .C2(n10081), .A(n9895), .B(n9894), .ZN(
        P1_U3230) );
  INV_X1 U12513 ( .A(n11312), .ZN(n9900) );
  OR2_X1 U12514 ( .A1(n9896), .A2(n8966), .ZN(n9897) );
  XNOR2_X1 U12515 ( .A(n9897), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11663) );
  INV_X1 U12516 ( .A(n11663), .ZN(n14080) );
  OAI222_X1 U12517 ( .A1(n14436), .A2(n9898), .B1(n14428), .B2(n9900), .C1(
        n14080), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U12518 ( .A(n13438), .ZN(n13433) );
  OAI222_X1 U12519 ( .A1(P2_U3088), .A2(n13433), .B1(n13818), .B2(n9900), .C1(
        n9899), .C2(n13820), .ZN(P2_U3310) );
  XNOR2_X1 U12520 ( .A(n9902), .B(n9901), .ZN(n15065) );
  AOI211_X1 U12521 ( .C1(n15062), .C2(n9904), .A(n8705), .B(n9903), .ZN(n15061) );
  AOI22_X1 U12522 ( .A1(n6578), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n13673), .ZN(n9905) );
  OAI21_X1 U12523 ( .B1(n9906), .B2(n13677), .A(n9905), .ZN(n9913) );
  NAND3_X1 U12524 ( .A1(n9510), .A2(n12400), .A3(n9908), .ZN(n9909) );
  AOI21_X1 U12525 ( .B1(n9778), .B2(n9909), .A(n10902), .ZN(n9911) );
  NOR2_X1 U12526 ( .A1(n9911), .A2(n9910), .ZN(n15064) );
  NOR2_X1 U12527 ( .A1(n15064), .A2(n6578), .ZN(n9912) );
  AOI211_X1 U12528 ( .C1(n15061), .C2(n13694), .A(n9913), .B(n9912), .ZN(n9914) );
  OAI21_X1 U12529 ( .B1(n13540), .B2(n15065), .A(n9914), .ZN(P2_U3263) );
  INV_X1 U12530 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9972) );
  OAI21_X1 U12531 ( .B1(n9916), .B2(n9915), .A(n12576), .ZN(n9917) );
  NAND2_X1 U12532 ( .A1(n9917), .A2(n12724), .ZN(n9920) );
  AOI21_X1 U12533 ( .B1(n10199), .B2(n12715), .A(n9918), .ZN(n9919) );
  OAI211_X1 U12534 ( .C1(n9921), .C2(n9972), .A(n9920), .B(n9919), .ZN(
        P3_U3177) );
  NAND2_X1 U12535 ( .A1(n9923), .A2(n7490), .ZN(n10096) );
  NAND2_X1 U12536 ( .A1(n13983), .A2(n11788), .ZN(n9925) );
  NAND2_X1 U12537 ( .A1(n11227), .A2(n11787), .ZN(n9924) );
  NAND2_X1 U12538 ( .A1(n9925), .A2(n9924), .ZN(n9926) );
  XNOR2_X1 U12539 ( .A(n9926), .B(n11692), .ZN(n9928) );
  AOI22_X1 U12540 ( .A1(n13983), .A2(n11757), .B1(n11227), .B2(n11788), .ZN(
        n9927) );
  AND2_X1 U12541 ( .A1(n9928), .A2(n9927), .ZN(n10095) );
  INV_X1 U12542 ( .A(n10095), .ZN(n9929) );
  OR2_X1 U12543 ( .A1(n9928), .A2(n9927), .ZN(n10094) );
  NAND2_X1 U12544 ( .A1(n9929), .A2(n10094), .ZN(n9930) );
  XNOR2_X1 U12545 ( .A(n9931), .B(n9930), .ZN(n9937) );
  INV_X1 U12546 ( .A(n14768), .ZN(n9935) );
  OAI22_X1 U12547 ( .A1(n10149), .A2(n14189), .B1(n9932), .B2(n14191), .ZN(
        n14767) );
  AOI22_X1 U12548 ( .A1(n14767), .A2(n13916), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9933) );
  OAI21_X1 U12549 ( .B1(n14868), .B2(n13969), .A(n9933), .ZN(n9934) );
  AOI21_X1 U12550 ( .B1(n9935), .B2(n13949), .A(n9934), .ZN(n9936) );
  OAI21_X1 U12551 ( .B1(n9937), .B2(n13955), .A(n9936), .ZN(P1_U3227) );
  INV_X1 U12552 ( .A(n11285), .ZN(n9941) );
  INV_X1 U12553 ( .A(n10766), .ZN(n13424) );
  OAI222_X1 U12554 ( .A1(n13820), .A2(n9938), .B1(n13818), .B2(n9941), .C1(
        n13424), .C2(P2_U3088), .ZN(P2_U3312) );
  NAND2_X1 U12555 ( .A1(n9939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9940) );
  XNOR2_X1 U12556 ( .A(n9940), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11286) );
  INV_X1 U12557 ( .A(n11286), .ZN(n14724) );
  OAI222_X1 U12558 ( .A1(P1_U3086), .A2(n14724), .B1(n14428), .B2(n9941), .C1(
        n15464), .C2(n14436), .ZN(P1_U3340) );
  INV_X1 U12559 ( .A(n9943), .ZN(n9944) );
  AOI21_X1 U12560 ( .B1(n9942), .B2(n9945), .A(n9944), .ZN(n9951) );
  NOR2_X1 U12561 ( .A1(n14947), .A2(n9946), .ZN(n9949) );
  NAND2_X1 U12562 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n13387) );
  OAI21_X1 U12563 ( .B1(n9947), .B2(n13238), .A(n13387), .ZN(n9948) );
  OAI21_X1 U12564 ( .B1(n9951), .B2(n14939), .A(n9950), .ZN(P2_U3193) );
  XNOR2_X1 U12565 ( .A(n9952), .B(n11587), .ZN(n14844) );
  XNOR2_X1 U12566 ( .A(n11587), .B(n9953), .ZN(n9955) );
  AOI21_X1 U12567 ( .B1(n9955), .B2(n14902), .A(n9954), .ZN(n14846) );
  INV_X1 U12568 ( .A(n14846), .ZN(n9960) );
  INV_X1 U12569 ( .A(n14301), .ZN(n14286) );
  INV_X1 U12570 ( .A(n14783), .ZN(n14284) );
  AOI22_X1 U12571 ( .A1(n14286), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14284), .ZN(n9958) );
  OAI211_X1 U12572 ( .C1(n9956), .C2(n14847), .A(n14788), .B(n14790), .ZN(
        n14845) );
  OR2_X1 U12573 ( .A1(n14273), .A2(n14845), .ZN(n9957) );
  OAI211_X1 U12574 ( .C1(n14786), .C2(n14847), .A(n9958), .B(n9957), .ZN(n9959) );
  AOI21_X1 U12575 ( .B1(n9960), .B2(n14301), .A(n9959), .ZN(n9961) );
  OAI21_X1 U12576 ( .B1(n14292), .B2(n14844), .A(n9961), .ZN(P1_U3291) );
  INV_X1 U12577 ( .A(n9962), .ZN(n9963) );
  OAI222_X1 U12578 ( .A1(n13228), .A2(n9964), .B1(n13227), .B2(n9963), .C1(
        n10195), .C2(P3_U3151), .ZN(P3_U3275) );
  OAI21_X1 U12579 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(n9975) );
  OAI21_X1 U12580 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9971) );
  AND2_X1 U12581 ( .A1(n12895), .A2(n9971), .ZN(n9974) );
  OAI22_X1 U12582 ( .A1(n12837), .A2(n14442), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9972), .ZN(n9973) );
  AOI211_X1 U12583 ( .C1(n12819), .C2(n9975), .A(n9974), .B(n9973), .ZN(n9980)
         );
  XNOR2_X1 U12584 ( .A(n9976), .B(n9977), .ZN(n9978) );
  NAND2_X1 U12585 ( .A1(n9978), .A2(n12767), .ZN(n9979) );
  OAI211_X1 U12586 ( .C1(n12883), .C2(n9981), .A(n9980), .B(n9979), .ZN(
        P3_U3184) );
  INV_X1 U12587 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10648) );
  INV_X1 U12588 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9989) );
  MUX2_X1 U12589 ( .A(n10648), .B(n9989), .S(n12862), .Z(n9982) );
  INV_X1 U12590 ( .A(n10028), .ZN(n10009) );
  NAND2_X1 U12591 ( .A1(n9982), .A2(n10009), .ZN(n10013) );
  INV_X1 U12592 ( .A(n9982), .ZN(n9983) );
  NAND2_X1 U12593 ( .A1(n9983), .A2(n10028), .ZN(n9984) );
  NAND2_X1 U12594 ( .A1(n10013), .A2(n9984), .ZN(n9985) );
  AND3_X1 U12595 ( .A1(n9987), .A2(n9986), .A3(n9985), .ZN(n9988) );
  OAI21_X1 U12596 ( .B1(n10046), .B2(n9988), .A(n12767), .ZN(n10007) );
  MUX2_X1 U12597 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n9989), .S(n10028), .Z(n9994) );
  INV_X1 U12598 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10810) );
  OAI22_X1 U12599 ( .A1(n9992), .A2(n10810), .B1(n9991), .B2(n9990), .ZN(n9993) );
  NAND2_X1 U12600 ( .A1(n9993), .A2(n9994), .ZN(n10008) );
  OAI21_X1 U12601 ( .B1(n9994), .B2(n9993), .A(n10008), .ZN(n10005) );
  INV_X1 U12602 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10003) );
  INV_X1 U12603 ( .A(n9995), .ZN(n9996) );
  MUX2_X1 U12604 ( .A(n10648), .B(P3_REG2_REG_6__SCAN_IN), .S(n10028), .Z(
        n9997) );
  AND3_X1 U12605 ( .A1(n9998), .A2(n9997), .A3(n9996), .ZN(n9999) );
  OAI21_X1 U12606 ( .B1(n10027), .B2(n9999), .A(n12819), .ZN(n10002) );
  INV_X1 U12607 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10000) );
  NOR2_X1 U12608 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10000), .ZN(n12712) );
  INV_X1 U12609 ( .A(n12712), .ZN(n10001) );
  OAI211_X1 U12610 ( .C1(n12837), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10004) );
  AOI21_X1 U12611 ( .B1(n12895), .B2(n10005), .A(n10004), .ZN(n10006) );
  OAI211_X1 U12612 ( .C1(n12883), .C2(n10028), .A(n10007), .B(n10006), .ZN(
        P3_U3188) );
  INV_X1 U12613 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15231) );
  MUX2_X1 U12614 ( .A(n15231), .B(P3_REG1_REG_8__SCAN_IN), .S(n10225), .Z(
        n10012) );
  OAI21_X1 U12615 ( .B1(n10009), .B2(n9989), .A(n10008), .ZN(n10010) );
  XNOR2_X1 U12616 ( .A(n10010), .B(n10029), .ZN(n10042) );
  AOI22_X1 U12617 ( .A1(n10042), .A2(P3_REG1_REG_7__SCAN_IN), .B1(n10052), 
        .B2(n10010), .ZN(n10011) );
  NOR2_X1 U12618 ( .A1(n10011), .A2(n10012), .ZN(n10223) );
  AOI21_X1 U12619 ( .B1(n10012), .B2(n10011), .A(n10223), .ZN(n10040) );
  INV_X1 U12620 ( .A(n10013), .ZN(n10045) );
  INV_X1 U12621 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10014) );
  INV_X1 U12622 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10041) );
  MUX2_X1 U12623 ( .A(n10014), .B(n10041), .S(n12862), .Z(n10015) );
  NAND2_X1 U12624 ( .A1(n10015), .A2(n10029), .ZN(n10023) );
  INV_X1 U12625 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U12626 ( .A1(n10016), .A2(n10052), .ZN(n10017) );
  AND2_X1 U12627 ( .A1(n10023), .A2(n10017), .ZN(n10044) );
  INV_X1 U12628 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10018) );
  MUX2_X1 U12629 ( .A(n10018), .B(n15231), .S(n12862), .Z(n10019) );
  INV_X1 U12630 ( .A(n10225), .ZN(n10037) );
  NAND2_X1 U12631 ( .A1(n10019), .A2(n10037), .ZN(n10230) );
  INV_X1 U12632 ( .A(n10019), .ZN(n10020) );
  NAND2_X1 U12633 ( .A1(n10020), .A2(n10225), .ZN(n10021) );
  NAND2_X1 U12634 ( .A1(n10230), .A2(n10021), .ZN(n10022) );
  AND3_X1 U12635 ( .A1(n10043), .A2(n10023), .A3(n10022), .ZN(n10024) );
  OAI21_X1 U12636 ( .B1(n10238), .B2(n10024), .A(n12767), .ZN(n10039) );
  INV_X1 U12637 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U12638 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15525), .ZN(n12599) );
  INV_X1 U12639 ( .A(n12599), .ZN(n10025) );
  OAI21_X1 U12640 ( .B1(n12837), .B2(n10026), .A(n10025), .ZN(n10036) );
  INV_X1 U12641 ( .A(n10030), .ZN(n10031) );
  XNOR2_X1 U12642 ( .A(n10225), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n10032) );
  INV_X1 U12643 ( .A(n10224), .ZN(n10034) );
  NAND3_X1 U12644 ( .A1(n10049), .A2(n10032), .A3(n10031), .ZN(n10033) );
  AOI21_X1 U12645 ( .B1(n10034), .B2(n10033), .A(n12896), .ZN(n10035) );
  AOI211_X1 U12646 ( .C1(n12834), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10038) );
  OAI211_X1 U12647 ( .C1(n10040), .C2(n10243), .A(n10039), .B(n10038), .ZN(
        P3_U3190) );
  XNOR2_X1 U12648 ( .A(n10042), .B(n10041), .ZN(n10057) );
  INV_X1 U12649 ( .A(n10043), .ZN(n10048) );
  NOR3_X1 U12650 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10047) );
  OAI21_X1 U12651 ( .B1(n10048), .B2(n10047), .A(n12767), .ZN(n10056) );
  OAI21_X1 U12652 ( .B1(n10050), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10049), .ZN(
        n10054) );
  AND2_X1 U12653 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12545) );
  AOI21_X1 U12654 ( .B1(n15142), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12545), .ZN(
        n10051) );
  OAI21_X1 U12655 ( .B1(n12883), .B2(n10052), .A(n10051), .ZN(n10053) );
  AOI21_X1 U12656 ( .B1(n10054), .B2(n12819), .A(n10053), .ZN(n10055) );
  OAI211_X1 U12657 ( .C1(n10057), .C2(n10243), .A(n10056), .B(n10055), .ZN(
        P3_U3189) );
  NAND2_X1 U12658 ( .A1(n10058), .A2(n12412), .ZN(n10060) );
  OR2_X1 U12659 ( .A1(n12196), .A2(n13316), .ZN(n10059) );
  INV_X1 U12660 ( .A(n13315), .ZN(n12204) );
  XNOR2_X1 U12661 ( .A(n15111), .B(n12204), .ZN(n12414) );
  INV_X1 U12662 ( .A(n12414), .ZN(n10253) );
  XNOR2_X1 U12663 ( .A(n10254), .B(n10253), .ZN(n10061) );
  NAND2_X1 U12664 ( .A1(n10061), .A2(n13683), .ZN(n10064) );
  OR2_X1 U12665 ( .A1(n12195), .A2(n13595), .ZN(n10063) );
  NAND2_X1 U12666 ( .A1(n13314), .A2(n13665), .ZN(n10062) );
  AND2_X1 U12667 ( .A1(n10063), .A2(n10062), .ZN(n10176) );
  NAND2_X1 U12668 ( .A1(n10064), .A2(n10176), .ZN(n15115) );
  INV_X1 U12669 ( .A(n15115), .ZN(n10077) );
  OR2_X1 U12670 ( .A1(n12196), .A2(n12195), .ZN(n10065) );
  OR2_X1 U12671 ( .A1(n10067), .A2(n12414), .ZN(n10068) );
  NAND2_X1 U12672 ( .A1(n10258), .A2(n10068), .ZN(n15114) );
  INV_X1 U12673 ( .A(n15114), .ZN(n10075) );
  AOI21_X1 U12674 ( .B1(n10069), .B2(n15111), .A(n8705), .ZN(n10070) );
  NAND2_X1 U12675 ( .A1(n10070), .A2(n10261), .ZN(n15113) );
  OAI22_X1 U12676 ( .A1(n15045), .A2(n10071), .B1(n10175), .B2(n15037), .ZN(
        n10072) );
  AOI21_X1 U12677 ( .B1(n15111), .B2(n13690), .A(n10072), .ZN(n10073) );
  OAI21_X1 U12678 ( .B1(n15113), .B2(n13639), .A(n10073), .ZN(n10074) );
  AOI21_X1 U12679 ( .B1(n10075), .B2(n10268), .A(n10074), .ZN(n10076) );
  OAI21_X1 U12680 ( .B1(n10077), .B2(n6578), .A(n10076), .ZN(P2_U3256) );
  NAND2_X1 U12681 ( .A1(n12753), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10078) );
  OAI21_X1 U12682 ( .B1(n12909), .B2(n12753), .A(n10078), .ZN(P3_U3519) );
  XNOR2_X1 U12683 ( .A(n11590), .B(n10079), .ZN(n14862) );
  NOR2_X1 U12684 ( .A1(n14286), .A2(n14863), .ZN(n14136) );
  INV_X1 U12685 ( .A(n14136), .ZN(n14129) );
  AOI211_X1 U12686 ( .C1(n14860), .C2(n14789), .A(n14837), .B(n14773), .ZN(
        n14858) );
  INV_X1 U12687 ( .A(n10080), .ZN(n14859) );
  MUX2_X1 U12688 ( .A(n14859), .B(P1_REG2_REG_4__SCAN_IN), .S(n14797), .Z(
        n10084) );
  OAI22_X1 U12689 ( .A1(n14786), .A2(n10082), .B1(n10081), .B2(n14783), .ZN(
        n10083) );
  AOI211_X1 U12690 ( .C1(n14858), .C2(n14793), .A(n10084), .B(n10083), .ZN(
        n10087) );
  XNOR2_X1 U12691 ( .A(n10085), .B(n11590), .ZN(n14865) );
  NAND2_X1 U12692 ( .A1(n14865), .A2(n14306), .ZN(n10086) );
  OAI211_X1 U12693 ( .C1(n14862), .C2(n14129), .A(n10087), .B(n10086), .ZN(
        P1_U3289) );
  NAND2_X1 U12694 ( .A1(n13986), .A2(n14750), .ZN(n14826) );
  OAI22_X1 U12695 ( .A1(n14286), .A2(n14826), .B1(n10088), .B2(n14783), .ZN(
        n10090) );
  AOI21_X1 U12696 ( .B1(n14087), .B2(n14786), .A(n11196), .ZN(n10089) );
  AOI211_X1 U12697 ( .C1(n14797), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10090), .B(
        n10089), .ZN(n10093) );
  NAND2_X1 U12698 ( .A1(n13987), .A2(n11196), .ZN(n10091) );
  NAND2_X1 U12699 ( .A1(n11200), .A2(n10091), .ZN(n11586) );
  OAI21_X1 U12700 ( .B1(n14136), .B2(n14306), .A(n11586), .ZN(n10092) );
  NAND2_X1 U12701 ( .A1(n10093), .A2(n10092), .ZN(P1_U3293) );
  NAND2_X1 U12702 ( .A1(n14875), .A2(n11787), .ZN(n10098) );
  NAND2_X1 U12703 ( .A1(n14748), .A2(n11788), .ZN(n10097) );
  NAND2_X1 U12704 ( .A1(n10098), .A2(n10097), .ZN(n10099) );
  XNOR2_X1 U12705 ( .A(n10099), .B(n11789), .ZN(n10277) );
  AOI22_X1 U12706 ( .A1(n14875), .A2(n11786), .B1(n14748), .B2(n11757), .ZN(
        n10278) );
  XNOR2_X1 U12707 ( .A(n10277), .B(n10278), .ZN(n10367) );
  NAND2_X1 U12708 ( .A1(n10369), .A2(n10367), .ZN(n10280) );
  OAI211_X1 U12709 ( .C1(n10369), .C2(n10367), .A(n10280), .B(n13959), .ZN(
        n10105) );
  NOR2_X1 U12710 ( .A1(n10101), .A2(n13951), .ZN(n10102) );
  AOI211_X1 U12711 ( .C1(n14875), .C2(n6564), .A(n10103), .B(n10102), .ZN(
        n10104) );
  OAI211_X1 U12712 ( .C1(n13963), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        P1_U3239) );
  INV_X1 U12713 ( .A(n13451), .ZN(n13445) );
  INV_X1 U12714 ( .A(n11302), .ZN(n10110) );
  OAI222_X1 U12715 ( .A1(P2_U3088), .A2(n13445), .B1(n13818), .B2(n10110), 
        .C1(n10107), .C2(n13820), .ZN(P2_U3309) );
  NAND2_X1 U12716 ( .A1(n10108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10109) );
  XNOR2_X1 U12717 ( .A(n10109), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14735) );
  INV_X1 U12718 ( .A(n14735), .ZN(n11659) );
  OAI222_X1 U12719 ( .A1(n14436), .A2(n10111), .B1(n14428), .B2(n10110), .C1(
        n11659), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X1 U12720 ( .A1(n10113), .A2(n10149), .ZN(n10114) );
  NAND2_X1 U12721 ( .A1(n10115), .A2(n10114), .ZN(n14744) );
  AOI22_X1 U12722 ( .A1(n11519), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11338), 
        .B2(n14044), .ZN(n10117) );
  XNOR2_X1 U12723 ( .A(n11238), .B(n13982), .ZN(n11592) );
  NAND2_X1 U12724 ( .A1(n14744), .A2(n14746), .ZN(n10120) );
  OR2_X1 U12725 ( .A1(n11238), .A2(n13982), .ZN(n10119) );
  NAND2_X1 U12726 ( .A1(n10120), .A2(n10119), .ZN(n10182) );
  OR2_X1 U12727 ( .A1(n10121), .A2(n11381), .ZN(n10124) );
  AOI22_X1 U12728 ( .A1(n11519), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11338), 
        .B2(n10122), .ZN(n10123) );
  NAND2_X1 U12729 ( .A1(n11387), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10133) );
  OR2_X1 U12730 ( .A1(n6573), .A2(n10125), .ZN(n10132) );
  OR2_X1 U12731 ( .A1(n11540), .A2(n10126), .ZN(n10131) );
  NAND2_X1 U12732 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  NAND2_X1 U12733 ( .A1(n10141), .A2(n10129), .ZN(n10381) );
  OR2_X1 U12734 ( .A1(n11491), .A2(n10381), .ZN(n10130) );
  NAND4_X1 U12735 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n14749) );
  INV_X1 U12736 ( .A(n11593), .ZN(n10183) );
  NAND2_X1 U12737 ( .A1(n10182), .A2(n10183), .ZN(n10135) );
  OR2_X1 U12738 ( .A1(n14891), .A2(n14749), .ZN(n10134) );
  NAND2_X1 U12739 ( .A1(n10135), .A2(n10134), .ZN(n10434) );
  OR2_X1 U12740 ( .A1(n10136), .A2(n11381), .ZN(n10138) );
  AOI22_X1 U12741 ( .A1(n11519), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11338), 
        .B2(n14061), .ZN(n10137) );
  NAND2_X1 U12742 ( .A1(n10138), .A2(n10137), .ZN(n11250) );
  NAND2_X1 U12743 ( .A1(n11387), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10146) );
  OR2_X1 U12744 ( .A1(n6573), .A2(n10139), .ZN(n10145) );
  NAND2_X1 U12745 ( .A1(n10141), .A2(n10140), .ZN(n10142) );
  NAND2_X1 U12746 ( .A1(n10419), .A2(n10142), .ZN(n10485) );
  OR2_X1 U12747 ( .A1(n11491), .A2(n10485), .ZN(n10144) );
  OR2_X1 U12748 ( .A1(n11540), .A2(n10317), .ZN(n10143) );
  NAND4_X1 U12749 ( .A1(n10146), .A2(n10145), .A3(n10144), .A4(n10143), .ZN(
        n13981) );
  XNOR2_X1 U12750 ( .A(n11250), .B(n13981), .ZN(n11595) );
  XNOR2_X1 U12751 ( .A(n10434), .B(n10433), .ZN(n10312) );
  INV_X1 U12752 ( .A(n10312), .ZN(n10170) );
  NAND2_X1 U12753 ( .A1(n10148), .A2(n10147), .ZN(n10151) );
  NAND2_X1 U12754 ( .A1(n10149), .A2(n14875), .ZN(n10150) );
  NAND2_X1 U12755 ( .A1(n10151), .A2(n10150), .ZN(n14745) );
  NAND2_X1 U12756 ( .A1(n14745), .A2(n11592), .ZN(n10153) );
  INV_X1 U12757 ( .A(n13982), .ZN(n10190) );
  NAND2_X1 U12758 ( .A1(n11238), .A2(n10190), .ZN(n10152) );
  NAND2_X1 U12759 ( .A1(n10153), .A2(n10152), .ZN(n10189) );
  INV_X1 U12760 ( .A(n14749), .ZN(n10289) );
  OR2_X1 U12761 ( .A1(n14891), .A2(n10289), .ZN(n10154) );
  OAI21_X1 U12762 ( .B1(n10155), .B2(n11595), .A(n10443), .ZN(n10163) );
  NAND2_X1 U12763 ( .A1(n14749), .A2(n14747), .ZN(n10162) );
  NAND2_X1 U12764 ( .A1(n11387), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10160) );
  OR2_X1 U12765 ( .A1(n6573), .A2(n10156), .ZN(n10159) );
  INV_X1 U12766 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10418) );
  XNOR2_X1 U12767 ( .A(n10419), .B(n10418), .ZN(n10470) );
  OR2_X1 U12768 ( .A1(n11491), .A2(n10470), .ZN(n10158) );
  OR2_X1 U12769 ( .A1(n11540), .A2(n14927), .ZN(n10157) );
  NAND4_X1 U12770 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n13980) );
  NAND2_X1 U12771 ( .A1(n13980), .A2(n14750), .ZN(n10161) );
  NAND2_X1 U12772 ( .A1(n10162), .A2(n10161), .ZN(n10483) );
  AOI21_X1 U12773 ( .B1(n10163), .B2(n14902), .A(n10483), .ZN(n10309) );
  INV_X1 U12774 ( .A(n10309), .ZN(n10168) );
  INV_X1 U12775 ( .A(n11250), .ZN(n10310) );
  OAI211_X1 U12776 ( .C1(n6735), .C2(n10310), .A(n10467), .B(n14790), .ZN(
        n10308) );
  NAND2_X1 U12777 ( .A1(n14286), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10164) );
  OAI21_X1 U12778 ( .B1(n14783), .B2(n10485), .A(n10164), .ZN(n10165) );
  AOI21_X1 U12779 ( .B1(n11250), .B2(n14303), .A(n10165), .ZN(n10166) );
  OAI21_X1 U12780 ( .B1(n10308), .B2(n14273), .A(n10166), .ZN(n10167) );
  AOI21_X1 U12781 ( .B1(n10168), .B2(n14301), .A(n10167), .ZN(n10169) );
  OAI21_X1 U12782 ( .B1(n14292), .B2(n10170), .A(n10169), .ZN(P1_U3284) );
  OAI21_X1 U12783 ( .B1(n10173), .B2(n10171), .A(n10172), .ZN(n10174) );
  NAND2_X1 U12784 ( .A1(n10174), .A2(n7445), .ZN(n10181) );
  INV_X1 U12785 ( .A(n10175), .ZN(n10179) );
  NOR2_X1 U12786 ( .A1(n10176), .A2(n13238), .ZN(n10177) );
  AOI211_X1 U12787 ( .C1(n13265), .C2(n10179), .A(n10178), .B(n10177), .ZN(
        n10180) );
  OAI211_X1 U12788 ( .C1(n7050), .C2(n13297), .A(n10181), .B(n10180), .ZN(
        P2_U3203) );
  XNOR2_X1 U12789 ( .A(n10182), .B(n10183), .ZN(n14895) );
  NAND2_X1 U12790 ( .A1(n14758), .A2(n14891), .ZN(n10184) );
  NAND2_X1 U12791 ( .A1(n10184), .A2(n14790), .ZN(n10185) );
  OR2_X1 U12792 ( .A1(n6735), .A2(n10185), .ZN(n14892) );
  NAND2_X1 U12793 ( .A1(n14286), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10186) );
  OAI21_X1 U12794 ( .B1(n14783), .B2(n10381), .A(n10186), .ZN(n10187) );
  AOI21_X1 U12795 ( .B1(n14303), .B2(n14891), .A(n10187), .ZN(n10188) );
  OAI21_X1 U12796 ( .B1(n14892), .B2(n14273), .A(n10188), .ZN(n10193) );
  XNOR2_X1 U12797 ( .A(n10189), .B(n11593), .ZN(n10191) );
  INV_X1 U12798 ( .A(n13981), .ZN(n10442) );
  OAI22_X1 U12799 ( .A1(n10442), .A2(n14189), .B1(n10190), .B2(n14191), .ZN(
        n10379) );
  AOI21_X1 U12800 ( .B1(n10191), .B2(n14902), .A(n10379), .ZN(n14893) );
  NOR2_X1 U12801 ( .A1(n14893), .A2(n14286), .ZN(n10192) );
  AOI211_X1 U12802 ( .C1(n14895), .C2(n14306), .A(n10193), .B(n10192), .ZN(
        n10194) );
  INV_X1 U12803 ( .A(n10194), .ZN(P1_U3285) );
  MUX2_X1 U12804 ( .A(n12107), .B(n10196), .S(n10195), .Z(n10197) );
  NAND2_X1 U12805 ( .A1(n10197), .A2(n6589), .ZN(n12922) );
  OR2_X1 U12806 ( .A1(n10351), .A2(n12107), .ZN(n13098) );
  INV_X1 U12807 ( .A(n12581), .ZN(n10216) );
  NAND2_X1 U12808 ( .A1(n10200), .A2(n11945), .ZN(n10324) );
  OAI21_X1 U12809 ( .B1(n10200), .B2(n11945), .A(n10324), .ZN(n10514) );
  NAND2_X1 U12810 ( .A1(n15168), .A2(n10201), .ZN(n10202) );
  NAND2_X1 U12811 ( .A1(n15164), .A2(n11917), .ZN(n10204) );
  NAND2_X1 U12812 ( .A1(n15192), .A2(n15173), .ZN(n10203) );
  INV_X1 U12813 ( .A(n11945), .ZN(n10208) );
  NAND2_X1 U12814 ( .A1(n11943), .A2(n10205), .ZN(n12102) );
  OAI211_X1 U12815 ( .C1(n7011), .C2(n10208), .A(n15149), .B(n10328), .ZN(
        n10211) );
  INV_X1 U12816 ( .A(n15193), .ZN(n15155) );
  AOI22_X1 U12817 ( .A1(n15154), .A2(n12752), .B1(n12750), .B2(n15155), .ZN(
        n10210) );
  NAND2_X1 U12818 ( .A1(n10211), .A2(n10210), .ZN(n10515) );
  AOI21_X1 U12819 ( .B1(n15221), .B2(n10514), .A(n10515), .ZN(n10219) );
  INV_X1 U12820 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10212) );
  OAI22_X1 U12821 ( .A1(n13163), .A2(n10216), .B1(n15235), .B2(n10212), .ZN(
        n10213) );
  INV_X1 U12822 ( .A(n10213), .ZN(n10214) );
  OAI21_X1 U12823 ( .B1(n10219), .B2(n15233), .A(n10214), .ZN(P3_U3462) );
  INV_X1 U12824 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n10215) );
  OAI22_X1 U12825 ( .A1(n10216), .A2(n13212), .B1(n15225), .B2(n10215), .ZN(
        n10217) );
  INV_X1 U12826 ( .A(n10217), .ZN(n10218) );
  OAI21_X1 U12827 ( .B1(n10219), .B2(n15223), .A(n10218), .ZN(P3_U3399) );
  INV_X1 U12828 ( .A(n10220), .ZN(n10222) );
  OAI222_X1 U12829 ( .A1(P3_U3151), .A2(n10350), .B1(n13227), .B2(n10222), 
        .C1(n10221), .C2(n13228), .ZN(P3_U3274) );
  XNOR2_X1 U12830 ( .A(n10553), .B(n10554), .ZN(n10556) );
  XNOR2_X1 U12831 ( .A(n10556), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n10244) );
  OAI21_X1 U12832 ( .B1(n10226), .B2(P3_REG2_REG_9__SCAN_IN), .A(n12757), .ZN(
        n10229) );
  AND2_X1 U12833 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n12674) );
  AOI21_X1 U12834 ( .B1(n15142), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12674), .ZN(
        n10227) );
  OAI21_X1 U12835 ( .B1(n12883), .B2(n10233), .A(n10227), .ZN(n10228) );
  AOI21_X1 U12836 ( .B1(n10229), .B2(n12819), .A(n10228), .ZN(n10242) );
  INV_X1 U12837 ( .A(n10230), .ZN(n10237) );
  INV_X1 U12838 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10231) );
  INV_X1 U12839 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10555) );
  MUX2_X1 U12840 ( .A(n10231), .B(n10555), .S(n12862), .Z(n10232) );
  NAND2_X1 U12841 ( .A1(n10232), .A2(n10554), .ZN(n12765) );
  INV_X1 U12842 ( .A(n10232), .ZN(n10234) );
  NAND2_X1 U12843 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  AND2_X1 U12844 ( .A1(n12765), .A2(n10235), .ZN(n10236) );
  INV_X1 U12845 ( .A(n12766), .ZN(n10240) );
  NOR3_X1 U12846 ( .A1(n10238), .A2(n10237), .A3(n10236), .ZN(n10239) );
  OAI21_X1 U12847 ( .B1(n10240), .B2(n10239), .A(n12767), .ZN(n10241) );
  OAI211_X1 U12848 ( .C1(n10244), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        P3_U3191) );
  XNOR2_X1 U12849 ( .A(n10245), .B(n10246), .ZN(n10252) );
  NOR2_X1 U12850 ( .A1(n14947), .A2(n10264), .ZN(n10250) );
  NAND2_X1 U12851 ( .A1(n13315), .A2(n13667), .ZN(n10248) );
  NAND2_X1 U12852 ( .A1(n13313), .A2(n13665), .ZN(n10247) );
  AND2_X1 U12853 ( .A1(n10248), .A2(n10247), .ZN(n10256) );
  OAI22_X1 U12854 ( .A1(n13238), .A2(n10256), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15436), .ZN(n10249) );
  AOI211_X1 U12855 ( .C1(n15119), .C2(n14943), .A(n10250), .B(n10249), .ZN(
        n10251) );
  OAI21_X1 U12856 ( .B1(n10252), .B2(n14939), .A(n10251), .ZN(P2_U3189) );
  XNOR2_X1 U12857 ( .A(n15119), .B(n12211), .ZN(n12415) );
  XNOR2_X1 U12858 ( .A(n6729), .B(n12415), .ZN(n10255) );
  NAND2_X1 U12859 ( .A1(n10255), .A2(n13683), .ZN(n10257) );
  NAND2_X1 U12860 ( .A1(n10257), .A2(n10256), .ZN(n15124) );
  INV_X1 U12861 ( .A(n15124), .ZN(n10270) );
  OR2_X1 U12862 ( .A1(n10259), .A2(n12415), .ZN(n10260) );
  NAND2_X1 U12863 ( .A1(n10526), .A2(n10260), .ZN(n15122) );
  INV_X1 U12864 ( .A(n15122), .ZN(n15125) );
  NAND2_X1 U12865 ( .A1(n15119), .A2(n10261), .ZN(n10262) );
  NAND2_X1 U12866 ( .A1(n10262), .A2(n6577), .ZN(n10263) );
  OR2_X1 U12867 ( .A1(n10530), .A2(n10263), .ZN(n15121) );
  OAI22_X1 U12868 ( .A1(n15045), .A2(n13412), .B1(n10264), .B2(n15037), .ZN(
        n10265) );
  AOI21_X1 U12869 ( .B1(n15119), .B2(n13690), .A(n10265), .ZN(n10266) );
  OAI21_X1 U12870 ( .B1(n15121), .B2(n13639), .A(n10266), .ZN(n10267) );
  AOI21_X1 U12871 ( .B1(n15125), .B2(n10268), .A(n10267), .ZN(n10269) );
  OAI21_X1 U12872 ( .B1(n10270), .B2(n6578), .A(n10269), .ZN(P2_U3255) );
  INV_X1 U12873 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15339) );
  NAND2_X1 U12874 ( .A1(n11900), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12875 ( .A1(n10271), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12876 ( .A1(n6584), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10272) );
  AND3_X1 U12877 ( .A1(n10274), .A2(n10273), .A3(n10272), .ZN(n10275) );
  INV_X1 U12878 ( .A(n12899), .ZN(n11909) );
  NAND2_X1 U12879 ( .A1(n11909), .A2(P3_U3897), .ZN(n10276) );
  OAI21_X1 U12880 ( .B1(P3_U3897), .B2(n15339), .A(n10276), .ZN(P3_U3522) );
  INV_X1 U12881 ( .A(n10277), .ZN(n10279) );
  OR2_X1 U12882 ( .A1(n10279), .A2(n10278), .ZN(n10372) );
  NAND2_X1 U12883 ( .A1(n10280), .A2(n10372), .ZN(n10286) );
  NAND2_X1 U12884 ( .A1(n11238), .A2(n6572), .ZN(n10282) );
  NAND2_X1 U12885 ( .A1(n13982), .A2(n11786), .ZN(n10281) );
  NAND2_X1 U12886 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  XNOR2_X1 U12887 ( .A(n10283), .B(n11789), .ZN(n10364) );
  AND2_X1 U12888 ( .A1(n13982), .A2(n11757), .ZN(n10284) );
  AOI21_X1 U12889 ( .B1(n11238), .B2(n11786), .A(n10284), .ZN(n10362) );
  XNOR2_X1 U12890 ( .A(n10364), .B(n10362), .ZN(n10365) );
  NAND2_X1 U12891 ( .A1(n10286), .A2(n10365), .ZN(n10285) );
  OAI211_X1 U12892 ( .C1(n10286), .C2(n10365), .A(n10285), .B(n13959), .ZN(
        n10293) );
  INV_X1 U12893 ( .A(n14754), .ZN(n10291) );
  INV_X1 U12894 ( .A(n13966), .ZN(n13941) );
  NOR2_X1 U12895 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10287), .ZN(n14038) );
  AOI21_X1 U12896 ( .B1(n13939), .B2(n14748), .A(n14038), .ZN(n10288) );
  OAI21_X1 U12897 ( .B1(n10289), .B2(n13941), .A(n10288), .ZN(n10290) );
  AOI21_X1 U12898 ( .B1(n10291), .B2(n13949), .A(n10290), .ZN(n10292) );
  OAI211_X1 U12899 ( .C1(n7065), .C2(n13969), .A(n10293), .B(n10292), .ZN(
        P1_U3213) );
  NOR3_X1 U12900 ( .A1(n12819), .A2(n12895), .A3(n12767), .ZN(n10303) );
  INV_X1 U12901 ( .A(n10294), .ZN(n10295) );
  AOI22_X1 U12902 ( .A1(n12895), .A2(P3_REG1_REG_0__SCAN_IN), .B1(n12767), 
        .B2(n10295), .ZN(n10296) );
  INV_X1 U12903 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10297) );
  OAI22_X1 U12904 ( .A1(n12837), .A2(n14493), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10297), .ZN(n10298) );
  AOI21_X1 U12905 ( .B1(n12819), .B2(n10299), .A(n10298), .ZN(n10300) );
  OAI211_X1 U12906 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        P3_U3182) );
  NAND2_X1 U12907 ( .A1(n6785), .A2(n10306), .ZN(n10304) );
  NAND2_X1 U12908 ( .A1(n10304), .A2(n11675), .ZN(n10305) );
  INV_X1 U12909 ( .A(n11191), .ZN(n10307) );
  NAND2_X1 U12910 ( .A1(n10307), .A2(n6790), .ZN(n14879) );
  OAI211_X1 U12911 ( .C1(n10310), .C2(n14899), .A(n10309), .B(n10308), .ZN(
        n10311) );
  AOI21_X1 U12912 ( .B1(n10312), .B2(n14906), .A(n10311), .ZN(n10323) );
  AND2_X1 U12913 ( .A1(n10314), .A2(n10313), .ZN(n10316) );
  OR2_X1 U12914 ( .A1(n14929), .A2(n10317), .ZN(n10318) );
  OAI21_X1 U12915 ( .B1(n10323), .B2(n14926), .A(n10318), .ZN(P1_U3537) );
  INV_X1 U12916 ( .A(n10319), .ZN(n10320) );
  NAND2_X1 U12917 ( .A1(n14908), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10322) );
  OAI21_X1 U12918 ( .B1(n10323), .B2(n14908), .A(n10322), .ZN(P1_U3486) );
  NAND2_X1 U12919 ( .A1(n10324), .A2(n11956), .ZN(n10325) );
  NAND2_X1 U12920 ( .A1(n10657), .A2(n12663), .ZN(n11964) );
  INV_X1 U12921 ( .A(n12663), .ZN(n10336) );
  NAND2_X1 U12922 ( .A1(n12750), .A2(n10336), .ZN(n11965) );
  NAND2_X1 U12923 ( .A1(n11964), .A2(n11965), .ZN(n11918) );
  INV_X1 U12924 ( .A(n11918), .ZN(n11969) );
  OR2_X1 U12925 ( .A1(n10325), .A2(n11969), .ZN(n10326) );
  AND2_X1 U12926 ( .A1(n10634), .A2(n10326), .ZN(n10357) );
  NAND2_X1 U12927 ( .A1(n12751), .A2(n12581), .ZN(n10327) );
  OAI211_X1 U12928 ( .C1(n10329), .C2(n11918), .A(n10638), .B(n15149), .ZN(
        n10332) );
  INV_X1 U12929 ( .A(n10330), .ZN(n10331) );
  AND2_X1 U12930 ( .A1(n10332), .A2(n10331), .ZN(n10352) );
  OAI21_X1 U12931 ( .B1(n13112), .B2(n10357), .A(n10352), .ZN(n10338) );
  INV_X1 U12932 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10333) );
  OAI22_X1 U12933 ( .A1(n10336), .A2(n13212), .B1(n15225), .B2(n10333), .ZN(
        n10334) );
  AOI21_X1 U12934 ( .B1(n10338), .B2(n15225), .A(n10334), .ZN(n10335) );
  INV_X1 U12935 ( .A(n10335), .ZN(P3_U3402) );
  OAI22_X1 U12936 ( .A1(n13163), .A2(n10336), .B1(n15235), .B2(n9597), .ZN(
        n10337) );
  AOI21_X1 U12937 ( .B1(n10338), .B2(n15235), .A(n10337), .ZN(n10339) );
  INV_X1 U12938 ( .A(n10339), .ZN(P3_U3463) );
  INV_X1 U12939 ( .A(n10340), .ZN(n10342) );
  OAI22_X1 U12940 ( .A1(n12107), .A2(P3_U3151), .B1(SI_22_), .B2(n13228), .ZN(
        n10341) );
  AOI21_X1 U12941 ( .B1(n10342), .B2(n13221), .A(n10341), .ZN(P3_U3273) );
  NAND2_X1 U12942 ( .A1(n13214), .A2(n10343), .ZN(n10344) );
  OAI21_X1 U12943 ( .B1(n13214), .B2(n10345), .A(n10344), .ZN(n10346) );
  INV_X1 U12944 ( .A(n10346), .ZN(n10347) );
  OR2_X1 U12945 ( .A1(n10351), .A2(n10350), .ZN(n15175) );
  NAND2_X1 U12946 ( .A1(n12922), .A2(n15175), .ZN(n15197) );
  INV_X1 U12947 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10353) );
  MUX2_X1 U12948 ( .A(n10353), .B(n10352), .S(n15198), .Z(n10356) );
  OR2_X1 U12949 ( .A1(n10354), .A2(n15186), .ZN(n14596) );
  AOI22_X1 U12950 ( .A1(n14583), .A2(n12663), .B1(n15178), .B2(n12664), .ZN(
        n10355) );
  OAI211_X1 U12951 ( .C1(n10357), .C2(n12983), .A(n10356), .B(n10355), .ZN(
        P3_U3229) );
  NAND2_X1 U12952 ( .A1(n14891), .A2(n11787), .ZN(n10359) );
  NAND2_X1 U12953 ( .A1(n14749), .A2(n11788), .ZN(n10358) );
  NAND2_X1 U12954 ( .A1(n10359), .A2(n10358), .ZN(n10360) );
  XNOR2_X1 U12955 ( .A(n10360), .B(n11692), .ZN(n10401) );
  AND2_X1 U12956 ( .A1(n14749), .A2(n11757), .ZN(n10361) );
  AOI21_X1 U12957 ( .B1(n14891), .B2(n11786), .A(n10361), .ZN(n10400) );
  XNOR2_X1 U12958 ( .A(n10401), .B(n10400), .ZN(n10377) );
  INV_X1 U12959 ( .A(n10362), .ZN(n10363) );
  NAND2_X1 U12960 ( .A1(n10364), .A2(n10363), .ZN(n10371) );
  INV_X1 U12961 ( .A(n10371), .ZN(n10366) );
  AND2_X1 U12962 ( .A1(n10367), .A2(n10370), .ZN(n10368) );
  INV_X1 U12963 ( .A(n10377), .ZN(n10375) );
  INV_X1 U12964 ( .A(n10403), .ZN(n10478) );
  AOI21_X1 U12965 ( .B1(n10377), .B2(n10376), .A(n10478), .ZN(n10384) );
  AOI21_X1 U12966 ( .B1(n10379), .B2(n13916), .A(n10378), .ZN(n10380) );
  OAI21_X1 U12967 ( .B1(n13963), .B2(n10381), .A(n10380), .ZN(n10382) );
  AOI21_X1 U12968 ( .B1(n14891), .B2(n6564), .A(n10382), .ZN(n10383) );
  OAI21_X1 U12969 ( .B1(n10384), .B2(n13955), .A(n10383), .ZN(P1_U3221) );
  NAND2_X1 U12970 ( .A1(n10386), .A2(n10385), .ZN(n10388) );
  XOR2_X1 U12971 ( .A(n10388), .B(n10387), .Z(n10392) );
  NAND2_X1 U12972 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14987)
         );
  OAI21_X1 U12973 ( .B1(n14933), .B2(n12211), .A(n14987), .ZN(n10390) );
  INV_X1 U12974 ( .A(n13312), .ZN(n10795) );
  OAI22_X1 U12975 ( .A1(n14932), .A2(n10795), .B1(n14947), .B2(n10532), .ZN(
        n10389) );
  AOI211_X1 U12976 ( .C1(n10776), .C2(n14943), .A(n10390), .B(n10389), .ZN(
        n10391) );
  OAI21_X1 U12977 ( .B1(n10392), .B2(n14939), .A(n10391), .ZN(P2_U3208) );
  INV_X1 U12978 ( .A(n11337), .ZN(n10394) );
  OAI222_X1 U12979 ( .A1(n14436), .A2(n10393), .B1(n14434), .B2(n10394), .C1(
        P1_U3086), .C2(n11675), .ZN(P1_U3336) );
  INV_X1 U12980 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10395) );
  OAI222_X1 U12981 ( .A1(n13820), .A2(n10395), .B1(n13818), .B2(n10394), .C1(
        n13459), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U12982 ( .A1(n11250), .A2(n11787), .ZN(n10397) );
  NAND2_X1 U12983 ( .A1(n13981), .A2(n11786), .ZN(n10396) );
  NAND2_X1 U12984 ( .A1(n10397), .A2(n10396), .ZN(n10398) );
  XNOR2_X1 U12985 ( .A(n10398), .B(n11692), .ZN(n10480) );
  AND2_X1 U12986 ( .A1(n13981), .A2(n11757), .ZN(n10399) );
  AOI21_X1 U12987 ( .B1(n11250), .B2(n11788), .A(n10399), .ZN(n10404) );
  AND2_X1 U12988 ( .A1(n10401), .A2(n10400), .ZN(n10477) );
  AOI21_X1 U12989 ( .B1(n10480), .B2(n10404), .A(n10477), .ZN(n10402) );
  INV_X1 U12990 ( .A(n10480), .ZN(n10405) );
  INV_X1 U12991 ( .A(n10404), .ZN(n10479) );
  NAND2_X1 U12992 ( .A1(n10405), .A2(n10479), .ZN(n10406) );
  NAND2_X1 U12993 ( .A1(n10407), .A2(n10406), .ZN(n10667) );
  OR2_X1 U12994 ( .A1(n10409), .A2(n11381), .ZN(n10411) );
  AOI22_X1 U12995 ( .A1(n11338), .A2(n14704), .B1(n11519), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12996 ( .A1(n11258), .A2(n11787), .ZN(n10413) );
  NAND2_X1 U12997 ( .A1(n13980), .A2(n11786), .ZN(n10412) );
  NAND2_X1 U12998 ( .A1(n10413), .A2(n10412), .ZN(n10414) );
  XNOR2_X1 U12999 ( .A(n10414), .B(n11692), .ZN(n10668) );
  AND2_X1 U13000 ( .A1(n13980), .A2(n11757), .ZN(n10415) );
  AOI21_X1 U13001 ( .B1(n11258), .B2(n11786), .A(n10415), .ZN(n10665) );
  INV_X1 U13002 ( .A(n10665), .ZN(n10669) );
  XNOR2_X1 U13003 ( .A(n10668), .B(n10669), .ZN(n10416) );
  XNOR2_X1 U13004 ( .A(n10408), .B(n10416), .ZN(n10432) );
  NAND2_X1 U13005 ( .A1(n11387), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10426) );
  OR2_X1 U13006 ( .A1(n6573), .A2(n10460), .ZN(n10425) );
  INV_X1 U13007 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10417) );
  OAI21_X1 U13008 ( .B1(n10419), .B2(n10418), .A(n10417), .ZN(n10422) );
  INV_X1 U13009 ( .A(n10419), .ZN(n10421) );
  NAND2_X1 U13010 ( .A1(n10422), .A2(n10450), .ZN(n10682) );
  OR2_X1 U13011 ( .A1(n11390), .A2(n10682), .ZN(n10424) );
  OR2_X1 U13012 ( .A1(n11540), .A2(n14673), .ZN(n10423) );
  NAND4_X1 U13013 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n13979) );
  AND2_X1 U13014 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n14714) );
  NOR2_X1 U13015 ( .A1(n13962), .A2(n10442), .ZN(n10428) );
  AOI211_X1 U13016 ( .C1(n13966), .C2(n13979), .A(n14714), .B(n10428), .ZN(
        n10429) );
  OAI21_X1 U13017 ( .B1(n13963), .B2(n10470), .A(n10429), .ZN(n10430) );
  AOI21_X1 U13018 ( .B1(n11258), .B2(n6564), .A(n10430), .ZN(n10431) );
  OAI21_X1 U13019 ( .B1(n10432), .B2(n13955), .A(n10431), .ZN(P1_U3217) );
  NAND2_X1 U13020 ( .A1(n10434), .A2(n10433), .ZN(n10436) );
  OR2_X1 U13021 ( .A1(n11250), .A2(n13981), .ZN(n10435) );
  NAND2_X1 U13022 ( .A1(n10436), .A2(n10435), .ZN(n10466) );
  INV_X1 U13023 ( .A(n13980), .ZN(n10679) );
  XNOR2_X1 U13024 ( .A(n11258), .B(n10679), .ZN(n11598) );
  OR2_X1 U13025 ( .A1(n11258), .A2(n13980), .ZN(n10437) );
  NAND2_X1 U13026 ( .A1(n10438), .A2(n11565), .ZN(n10441) );
  AOI22_X1 U13027 ( .A1(n11519), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n10439), 
        .B2(n11338), .ZN(n10440) );
  NAND2_X2 U13028 ( .A1(n10441), .A2(n10440), .ZN(n14667) );
  INV_X1 U13029 ( .A(n13979), .ZN(n10565) );
  XNOR2_X1 U13030 ( .A(n14667), .B(n10565), .ZN(n11597) );
  XNOR2_X1 U13031 ( .A(n10604), .B(n11597), .ZN(n14666) );
  INV_X1 U13032 ( .A(n14666), .ZN(n10465) );
  INV_X1 U13033 ( .A(n10469), .ZN(n10445) );
  NAND2_X1 U13034 ( .A1(n10445), .A2(n10444), .ZN(n14903) );
  OR2_X1 U13035 ( .A1(n11258), .A2(n10679), .ZN(n10446) );
  NAND2_X1 U13036 ( .A1(n14903), .A2(n10446), .ZN(n10448) );
  INV_X1 U13037 ( .A(n11597), .ZN(n10447) );
  NAND2_X1 U13038 ( .A1(n10448), .A2(n10447), .ZN(n10567) );
  OAI211_X1 U13039 ( .C1(n10448), .C2(n10447), .A(n10567), .B(n14902), .ZN(
        n10457) );
  NAND2_X1 U13040 ( .A1(n11387), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U13041 ( .A1(n10450), .A2(n10449), .ZN(n10451) );
  NAND2_X1 U13042 ( .A1(n10590), .A2(n10451), .ZN(n13870) );
  OR2_X1 U13043 ( .A1(n11491), .A2(n13870), .ZN(n10454) );
  OR2_X1 U13044 ( .A1(n6573), .A2(n9407), .ZN(n10453) );
  OR2_X1 U13045 ( .A1(n11540), .A2(n14565), .ZN(n10452) );
  NAND4_X1 U13046 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n13978) );
  AOI22_X1 U13047 ( .A1(n14750), .A2(n13978), .B1(n13980), .B2(n14747), .ZN(
        n10456) );
  NAND2_X1 U13048 ( .A1(n10457), .A2(n10456), .ZN(n14672) );
  INV_X1 U13049 ( .A(n14797), .ZN(n14301) );
  NOR2_X2 U13050 ( .A1(n14667), .A2(n10458), .ZN(n10619) );
  AND2_X1 U13051 ( .A1(n14667), .A2(n10458), .ZN(n10459) );
  OR2_X1 U13052 ( .A1(n10619), .A2(n10459), .ZN(n14669) );
  OAI22_X1 U13053 ( .A1(n14301), .A2(n10460), .B1(n10682), .B2(n14783), .ZN(
        n10461) );
  AOI21_X1 U13054 ( .B1(n14667), .B2(n14303), .A(n10461), .ZN(n10462) );
  OAI21_X1 U13055 ( .B1(n14669), .B2(n14087), .A(n10462), .ZN(n10463) );
  AOI21_X1 U13056 ( .B1(n14672), .B2(n14301), .A(n10463), .ZN(n10464) );
  OAI21_X1 U13057 ( .B1(n14292), .B2(n10465), .A(n10464), .ZN(P1_U3282) );
  XNOR2_X1 U13058 ( .A(n10466), .B(n11598), .ZN(n14907) );
  XOR2_X1 U13059 ( .A(n11258), .B(n10467), .Z(n10468) );
  AOI22_X1 U13060 ( .A1(n10468), .A2(n14790), .B1(n14750), .B2(n13979), .ZN(
        n14898) );
  NAND2_X1 U13061 ( .A1(n10469), .A2(n11598), .ZN(n14901) );
  NAND3_X1 U13062 ( .A1(n14903), .A2(n14901), .A3(n14136), .ZN(n10474) );
  NAND2_X1 U13063 ( .A1(n13981), .A2(n14747), .ZN(n14897) );
  OAI22_X1 U13064 ( .A1(n14286), .A2(n14897), .B1(n10470), .B2(n14783), .ZN(
        n10472) );
  INV_X1 U13065 ( .A(n11258), .ZN(n14900) );
  NOR2_X1 U13066 ( .A1(n14900), .A2(n14786), .ZN(n10471) );
  AOI211_X1 U13067 ( .C1(n14797), .C2(P1_REG2_REG_10__SCAN_IN), .A(n10472), 
        .B(n10471), .ZN(n10473) );
  OAI211_X1 U13068 ( .C1(n14898), .C2(n14273), .A(n10474), .B(n10473), .ZN(
        n10475) );
  AOI21_X1 U13069 ( .B1(n14306), .B2(n14907), .A(n10475), .ZN(n10476) );
  INV_X1 U13070 ( .A(n10476), .ZN(P1_U3283) );
  NOR2_X1 U13071 ( .A1(n10478), .A2(n10477), .ZN(n10482) );
  XNOR2_X1 U13072 ( .A(n10480), .B(n10479), .ZN(n10481) );
  XNOR2_X1 U13073 ( .A(n10482), .B(n10481), .ZN(n10488) );
  AOI22_X1 U13074 ( .A1(n10483), .A2(n13916), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10484) );
  OAI21_X1 U13075 ( .B1(n13963), .B2(n10485), .A(n10484), .ZN(n10486) );
  AOI21_X1 U13076 ( .B1(n11250), .B2(n6564), .A(n10486), .ZN(n10487) );
  OAI21_X1 U13077 ( .B1(n10488), .B2(n13955), .A(n10487), .ZN(P1_U3231) );
  NAND2_X1 U13078 ( .A1(n10489), .A2(n13221), .ZN(n10490) );
  OAI211_X1 U13079 ( .C1(n15465), .C2(n13228), .A(n10490), .B(n12110), .ZN(
        P3_U3272) );
  INV_X1 U13080 ( .A(n10491), .ZN(n10492) );
  AOI21_X1 U13081 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15178), .A(n10492), .ZN(
        n10494) );
  MUX2_X1 U13082 ( .A(n10494), .B(n10493), .S(n14582), .Z(n10495) );
  OAI21_X1 U13083 ( .B1(n10496), .B2(n13081), .A(n10495), .ZN(P3_U3233) );
  NOR2_X1 U13084 ( .A1(n11286), .A2(n10498), .ZN(n10499) );
  XNOR2_X1 U13085 ( .A(n10498), .B(n11286), .ZN(n14719) );
  NOR2_X1 U13086 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14719), .ZN(n14718) );
  INV_X1 U13087 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U13088 ( .A1(n11666), .A2(n14652), .ZN(n10500) );
  AOI21_X1 U13089 ( .B1(n14652), .B2(n11666), .A(n10500), .ZN(n10501) );
  NAND2_X1 U13090 ( .A1(n10501), .A2(n10502), .ZN(n11657) );
  OAI211_X1 U13091 ( .C1(n10502), .C2(n10501), .A(n14738), .B(n11657), .ZN(
        n10513) );
  NAND2_X1 U13092 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13892)
         );
  OAI21_X1 U13093 ( .B1(n14300), .B2(n10504), .A(n10503), .ZN(n10505) );
  NOR2_X1 U13094 ( .A1(n11286), .A2(n10505), .ZN(n10506) );
  XOR2_X1 U13095 ( .A(n10505), .B(n14724), .Z(n14717) );
  NOR2_X1 U13096 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14717), .ZN(n14716) );
  NOR2_X1 U13097 ( .A1(n10506), .A2(n14716), .ZN(n10509) );
  INV_X1 U13098 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14269) );
  NOR2_X1 U13099 ( .A1(n11666), .A2(n14269), .ZN(n10507) );
  AOI21_X1 U13100 ( .B1(n14269), .B2(n11666), .A(n10507), .ZN(n10508) );
  NAND2_X1 U13101 ( .A1(n10508), .A2(n10509), .ZN(n11665) );
  OAI211_X1 U13102 ( .C1(n10509), .C2(n10508), .A(n14733), .B(n11665), .ZN(
        n10510) );
  NAND2_X1 U13103 ( .A1(n13892), .A2(n10510), .ZN(n10511) );
  AOI21_X1 U13104 ( .B1(n14731), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10511), 
        .ZN(n10512) );
  OAI211_X1 U13105 ( .C1(n14725), .C2(n11666), .A(n10513), .B(n10512), .ZN(
        P1_U3259) );
  INV_X1 U13106 ( .A(n10514), .ZN(n10520) );
  INV_X1 U13107 ( .A(n10515), .ZN(n10517) );
  INV_X1 U13108 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10516) );
  MUX2_X1 U13109 ( .A(n10517), .B(n10516), .S(n14582), .Z(n10519) );
  AOI22_X1 U13110 ( .A1(n14583), .A2(n12581), .B1(n15178), .B2(n12582), .ZN(
        n10518) );
  OAI211_X1 U13111 ( .C1(n12983), .C2(n10520), .A(n10519), .B(n10518), .ZN(
        P3_U3230) );
  NAND2_X1 U13112 ( .A1(n10776), .A2(n14934), .ZN(n10687) );
  NAND2_X1 U13113 ( .A1(n10687), .A2(n10521), .ZN(n12416) );
  INV_X1 U13114 ( .A(n12416), .ZN(n10524) );
  NAND2_X1 U13115 ( .A1(n15119), .A2(n12211), .ZN(n10522) );
  INV_X1 U13116 ( .A(n15119), .ZN(n12212) );
  OAI21_X1 U13117 ( .B1(n10524), .B2(n10523), .A(n10688), .ZN(n10529) );
  OAI22_X1 U13118 ( .A1(n12211), .A2(n13595), .B1(n10795), .B2(n15039), .ZN(
        n10528) );
  NAND2_X1 U13119 ( .A1(n15119), .A2(n13314), .ZN(n10525) );
  NAND2_X1 U13120 ( .A1(n10526), .A2(n10525), .ZN(n10686) );
  XNOR2_X1 U13121 ( .A(n10686), .B(n12416), .ZN(n10779) );
  NOR2_X1 U13122 ( .A1(n10779), .A2(n9127), .ZN(n10527) );
  AOI211_X1 U13123 ( .C1(n13683), .C2(n10529), .A(n10528), .B(n10527), .ZN(
        n10778) );
  INV_X1 U13124 ( .A(n10530), .ZN(n10531) );
  INV_X1 U13125 ( .A(n10693), .ZN(n10695) );
  AOI211_X1 U13126 ( .C1(n10776), .C2(n10531), .A(n8705), .B(n10695), .ZN(
        n10775) );
  INV_X1 U13127 ( .A(n10532), .ZN(n10533) );
  AOI22_X1 U13128 ( .A1(n6578), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10533), 
        .B2(n13673), .ZN(n10534) );
  OAI21_X1 U13129 ( .B1(n12215), .B2(n13677), .A(n10534), .ZN(n10536) );
  NOR2_X1 U13130 ( .A1(n10779), .A2(n13609), .ZN(n10535) );
  AOI211_X1 U13131 ( .C1(n10775), .C2(n13694), .A(n10536), .B(n10535), .ZN(
        n10537) );
  OAI21_X1 U13132 ( .B1(n10778), .B2(n6578), .A(n10537), .ZN(P2_U3254) );
  INV_X1 U13133 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10547) );
  INV_X1 U13134 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U13135 ( .A(n10547), .B(n10558), .S(n12862), .Z(n10538) );
  INV_X1 U13136 ( .A(n10557), .ZN(n12763) );
  NAND2_X1 U13137 ( .A1(n10538), .A2(n12763), .ZN(n10541) );
  INV_X1 U13138 ( .A(n10538), .ZN(n10539) );
  NAND2_X1 U13139 ( .A1(n10539), .A2(n10557), .ZN(n10540) );
  NAND2_X1 U13140 ( .A1(n10541), .A2(n10540), .ZN(n12764) );
  INV_X1 U13141 ( .A(n10541), .ZN(n10542) );
  MUX2_X1 U13142 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12862), .Z(n10730) );
  XOR2_X1 U13143 ( .A(n10559), .B(n10730), .Z(n10543) );
  AOI21_X1 U13144 ( .B1(n10544), .B2(n10543), .A(n10733), .ZN(n10564) );
  INV_X1 U13145 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15383) );
  INV_X1 U13146 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15507) );
  NOR2_X1 U13147 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15507), .ZN(n12693) );
  INV_X1 U13148 ( .A(n12693), .ZN(n10545) );
  OAI21_X1 U13149 ( .B1(n12837), .B2(n15383), .A(n10545), .ZN(n10552) );
  INV_X1 U13150 ( .A(n10546), .ZN(n12755) );
  MUX2_X1 U13151 ( .A(n10547), .B(P3_REG2_REG_10__SCAN_IN), .S(n10557), .Z(
        n12756) );
  NOR2_X1 U13152 ( .A1(n10548), .A2(n10559), .ZN(n10726) );
  INV_X1 U13153 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14606) );
  AOI21_X1 U13154 ( .B1(n10549), .B2(n14606), .A(n10725), .ZN(n10550) );
  NOR2_X1 U13155 ( .A1(n10550), .A2(n12896), .ZN(n10551) );
  AOI211_X1 U13156 ( .C1(n12834), .C2(n10559), .A(n10552), .B(n10551), .ZN(
        n10563) );
  OAI22_X1 U13157 ( .A1(n10556), .A2(n10555), .B1(n10554), .B2(n10553), .ZN(
        n12771) );
  MUX2_X1 U13158 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n10558), .S(n10557), .Z(
        n12772) );
  XNOR2_X1 U13159 ( .A(n10736), .B(n10559), .ZN(n10560) );
  NAND2_X1 U13160 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10560), .ZN(n10737) );
  OAI21_X1 U13161 ( .B1(n10560), .B2(P3_REG1_REG_11__SCAN_IN), .A(n10737), 
        .ZN(n10561) );
  NAND2_X1 U13162 ( .A1(n10561), .A2(n12895), .ZN(n10562) );
  OAI211_X1 U13163 ( .C1(n10564), .C2(n12891), .A(n10563), .B(n10562), .ZN(
        P3_U3193) );
  NAND2_X1 U13164 ( .A1(n10567), .A2(n10566), .ZN(n10611) );
  NAND2_X1 U13165 ( .A1(n10568), .A2(n11565), .ZN(n10571) );
  AOI22_X1 U13166 ( .A1(n10569), .A2(n11338), .B1(n11519), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U13167 ( .A1(n10611), .A2(n11599), .ZN(n10616) );
  INV_X1 U13168 ( .A(n13978), .ZN(n10844) );
  NAND2_X1 U13169 ( .A1(n10616), .A2(n10572), .ZN(n10584) );
  NAND2_X1 U13170 ( .A1(n10573), .A2(n11565), .ZN(n10578) );
  NOR2_X1 U13171 ( .A1(n11567), .A2(n10574), .ZN(n10575) );
  AOI21_X1 U13172 ( .B1(n10576), .B2(n11338), .A(n10575), .ZN(n10577) );
  NAND2_X1 U13173 ( .A1(n11387), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10583) );
  OR2_X1 U13174 ( .A1(n6573), .A2(n9470), .ZN(n10582) );
  INV_X1 U13175 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10589) );
  XNOR2_X1 U13176 ( .A(n10590), .B(n10589), .ZN(n10847) );
  OR2_X1 U13177 ( .A1(n11390), .A2(n10847), .ZN(n10581) );
  OR2_X1 U13178 ( .A1(n11540), .A2(n10579), .ZN(n10580) );
  NAND4_X1 U13179 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(
        n13977) );
  XNOR2_X1 U13180 ( .A(n14660), .B(n13977), .ZN(n11600) );
  NAND2_X1 U13181 ( .A1(n10584), .A2(n11600), .ZN(n11803) );
  OAI21_X1 U13182 ( .B1(n10584), .B2(n11600), .A(n11803), .ZN(n14663) );
  INV_X1 U13183 ( .A(n13877), .ZN(n14560) );
  NAND2_X1 U13184 ( .A1(n14560), .A2(n10619), .ZN(n10618) );
  AOI21_X1 U13185 ( .B1(n10618), .B2(n14660), .A(n14837), .ZN(n10585) );
  NAND2_X1 U13186 ( .A1(n10585), .A2(n14308), .ZN(n14661) );
  INV_X1 U13187 ( .A(n14661), .ZN(n10603) );
  NAND2_X1 U13188 ( .A1(n14660), .A2(n14303), .ZN(n10601) );
  NAND2_X1 U13189 ( .A1(n11387), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10595) );
  OR2_X1 U13190 ( .A1(n6573), .A2(n14300), .ZN(n10594) );
  AND2_X1 U13191 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n10586) );
  INV_X1 U13192 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10588) );
  OAI21_X1 U13193 ( .B1(n10590), .B2(n10589), .A(n10588), .ZN(n10591) );
  NAND2_X1 U13194 ( .A1(n11290), .A2(n10591), .ZN(n14299) );
  OR2_X1 U13195 ( .A1(n11491), .A2(n14299), .ZN(n10593) );
  OR2_X1 U13196 ( .A1(n11540), .A2(n15332), .ZN(n10592) );
  NAND4_X1 U13197 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n14278) );
  NAND2_X1 U13198 ( .A1(n14278), .A2(n14750), .ZN(n10597) );
  NAND2_X1 U13199 ( .A1(n13978), .A2(n14747), .ZN(n10596) );
  NAND2_X1 U13200 ( .A1(n10597), .A2(n10596), .ZN(n14659) );
  INV_X1 U13201 ( .A(n14659), .ZN(n10598) );
  OAI22_X1 U13202 ( .A1(n14286), .A2(n10598), .B1(n10847), .B2(n14783), .ZN(
        n10599) );
  INV_X1 U13203 ( .A(n10599), .ZN(n10600) );
  OAI211_X1 U13204 ( .C1(n14301), .C2(n9470), .A(n10601), .B(n10600), .ZN(
        n10602) );
  AOI21_X1 U13205 ( .B1(n10603), .B2(n14793), .A(n10602), .ZN(n10609) );
  OR2_X1 U13206 ( .A1(n14667), .A2(n13979), .ZN(n10605) );
  INV_X1 U13207 ( .A(n11599), .ZN(n10612) );
  NAND2_X1 U13208 ( .A1(n10610), .A2(n10612), .ZN(n10607) );
  OR2_X1 U13209 ( .A1(n13877), .A2(n13978), .ZN(n10606) );
  NAND2_X1 U13210 ( .A1(n10607), .A2(n10606), .ZN(n11819) );
  INV_X1 U13211 ( .A(n11600), .ZN(n11818) );
  XNOR2_X1 U13212 ( .A(n11819), .B(n11818), .ZN(n14665) );
  NAND2_X1 U13213 ( .A1(n14665), .A2(n14306), .ZN(n10608) );
  OAI211_X1 U13214 ( .C1(n14663), .C2(n14129), .A(n10609), .B(n10608), .ZN(
        P1_U3280) );
  XNOR2_X1 U13215 ( .A(n10610), .B(n11599), .ZN(n14557) );
  INV_X1 U13216 ( .A(n10611), .ZN(n10613) );
  AOI21_X1 U13217 ( .B1(n10613), .B2(n10612), .A(n14863), .ZN(n10617) );
  NAND2_X1 U13218 ( .A1(n13979), .A2(n14747), .ZN(n10615) );
  NAND2_X1 U13219 ( .A1(n13977), .A2(n14750), .ZN(n10614) );
  NAND2_X1 U13220 ( .A1(n10615), .A2(n10614), .ZN(n13868) );
  AOI21_X1 U13221 ( .B1(n10617), .B2(n10616), .A(n13868), .ZN(n14559) );
  INV_X1 U13222 ( .A(n14559), .ZN(n10624) );
  OAI211_X1 U13223 ( .C1(n14560), .C2(n10619), .A(n14790), .B(n10618), .ZN(
        n14558) );
  NAND2_X1 U13224 ( .A1(n14286), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10620) );
  OAI21_X1 U13225 ( .B1(n14783), .B2(n13870), .A(n10620), .ZN(n10621) );
  AOI21_X1 U13226 ( .B1(n13877), .B2(n14303), .A(n10621), .ZN(n10622) );
  OAI21_X1 U13227 ( .B1(n14558), .B2(n14273), .A(n10622), .ZN(n10623) );
  AOI21_X1 U13228 ( .B1(n10624), .B2(n14301), .A(n10623), .ZN(n10625) );
  OAI21_X1 U13229 ( .B1(n14292), .B2(n14557), .A(n10625), .ZN(P1_U3281) );
  AOI21_X1 U13230 ( .B1(n10627), .B2(n10626), .A(n14939), .ZN(n10629) );
  NAND2_X1 U13231 ( .A1(n10629), .A2(n10628), .ZN(n10633) );
  INV_X1 U13232 ( .A(n10802), .ZN(n10631) );
  INV_X1 U13233 ( .A(n12233), .ZN(n13311) );
  AOI22_X1 U13234 ( .A1(n13311), .A2(n13665), .B1(n13667), .B2(n13312), .ZN(
        n10798) );
  OAI22_X1 U13235 ( .A1(n10798), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8680), .ZN(n10630) );
  AOI21_X1 U13236 ( .B1(n10631), .B2(n13265), .A(n10630), .ZN(n10632) );
  OAI211_X1 U13237 ( .C1(n14634), .C2(n13297), .A(n10633), .B(n10632), .ZN(
        P2_U3206) );
  NAND2_X1 U13238 ( .A1(n10644), .A2(n12632), .ZN(n11971) );
  NAND2_X1 U13239 ( .A1(n12749), .A2(n10812), .ZN(n11974) );
  NAND2_X1 U13240 ( .A1(n10703), .A2(n12714), .ZN(n11981) );
  INV_X1 U13241 ( .A(n12714), .ZN(n10721) );
  NAND2_X1 U13242 ( .A1(n12631), .A2(n10721), .ZN(n11975) );
  NAND2_X1 U13243 ( .A1(n10635), .A2(n11919), .ZN(n10707) );
  OAI21_X1 U13244 ( .B1(n10635), .B2(n11919), .A(n10707), .ZN(n10636) );
  INV_X1 U13245 ( .A(n10636), .ZN(n10717) );
  NAND2_X1 U13246 ( .A1(n12750), .A2(n12663), .ZN(n10637) );
  NAND2_X1 U13247 ( .A1(n10644), .A2(n10812), .ZN(n10641) );
  AOI21_X1 U13248 ( .B1(n10642), .B2(n11919), .A(n15191), .ZN(n10647) );
  OAI22_X1 U13249 ( .A1(n10645), .A2(n15193), .B1(n10644), .B2(n15195), .ZN(
        n10646) );
  AOI21_X1 U13250 ( .B1(n10647), .B2(n10701), .A(n10646), .ZN(n10716) );
  MUX2_X1 U13251 ( .A(n10716), .B(n10648), .S(n14582), .Z(n10650) );
  AOI22_X1 U13252 ( .A1(n14583), .A2(n12714), .B1(n15178), .B2(n12716), .ZN(
        n10649) );
  OAI211_X1 U13253 ( .C1(n12983), .C2(n10717), .A(n10650), .B(n10649), .ZN(
        P3_U3227) );
  OAI21_X1 U13254 ( .B1(n10652), .B2(n11966), .A(n10651), .ZN(n10787) );
  INV_X1 U13255 ( .A(n10653), .ZN(n10654) );
  AOI21_X1 U13256 ( .B1(n11966), .B2(n10655), .A(n10654), .ZN(n10656) );
  OAI222_X1 U13257 ( .A1(n15195), .A2(n10657), .B1(n15193), .B2(n10703), .C1(
        n15191), .C2(n10656), .ZN(n10788) );
  AOI21_X1 U13258 ( .B1(n15221), .B2(n10787), .A(n10788), .ZN(n10809) );
  INV_X1 U13259 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10658) );
  OAI22_X1 U13260 ( .A1(n10812), .A2(n13212), .B1(n15225), .B2(n10658), .ZN(
        n10659) );
  INV_X1 U13261 ( .A(n10659), .ZN(n10660) );
  OAI21_X1 U13262 ( .B1(n10809), .B2(n15223), .A(n10660), .ZN(P3_U3405) );
  NAND2_X1 U13263 ( .A1(n14667), .A2(n11787), .ZN(n10662) );
  NAND2_X1 U13264 ( .A1(n13979), .A2(n11788), .ZN(n10661) );
  NAND2_X1 U13265 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  XNOR2_X1 U13266 ( .A(n10663), .B(n11692), .ZN(n10825) );
  AND2_X1 U13267 ( .A1(n13979), .A2(n11757), .ZN(n10664) );
  AOI21_X1 U13268 ( .B1(n14667), .B2(n11788), .A(n10664), .ZN(n10824) );
  XNOR2_X1 U13269 ( .A(n10825), .B(n10824), .ZN(n10677) );
  NAND2_X1 U13270 ( .A1(n10668), .A2(n10665), .ZN(n10666) );
  NAND2_X1 U13271 ( .A1(n10667), .A2(n10666), .ZN(n10672) );
  INV_X1 U13272 ( .A(n10668), .ZN(n10670) );
  NAND2_X1 U13273 ( .A1(n10670), .A2(n10669), .ZN(n10671) );
  NAND2_X1 U13274 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  INV_X1 U13275 ( .A(n10827), .ZN(n10676) );
  AOI21_X1 U13276 ( .B1(n10677), .B2(n10673), .A(n10676), .ZN(n10685) );
  OAI21_X1 U13277 ( .B1(n13962), .B2(n10679), .A(n10678), .ZN(n10680) );
  AOI21_X1 U13278 ( .B1(n13966), .B2(n13978), .A(n10680), .ZN(n10681) );
  OAI21_X1 U13279 ( .B1(n13963), .B2(n10682), .A(n10681), .ZN(n10683) );
  AOI21_X1 U13280 ( .B1(n14667), .B2(n6564), .A(n10683), .ZN(n10684) );
  OAI21_X1 U13281 ( .B1(n10685), .B2(n13955), .A(n10684), .ZN(P1_U3236) );
  XNOR2_X1 U13282 ( .A(n14944), .B(n13312), .ZN(n12419) );
  XOR2_X1 U13283 ( .A(n10794), .B(n12419), .Z(n14638) );
  XNOR2_X1 U13284 ( .A(n10797), .B(n12419), .ZN(n10690) );
  OAI22_X1 U13285 ( .A1(n14931), .A2(n15039), .B1(n14934), .B2(n13595), .ZN(
        n10689) );
  AOI21_X1 U13286 ( .B1(n10690), .B2(n13683), .A(n10689), .ZN(n10691) );
  OAI21_X1 U13287 ( .B1(n14638), .B2(n9127), .A(n10691), .ZN(n14641) );
  NAND2_X1 U13288 ( .A1(n14641), .A2(n15045), .ZN(n10699) );
  OAI22_X1 U13289 ( .A1(n15045), .A2(n10692), .B1(n14946), .B2(n15037), .ZN(
        n10697) );
  INV_X1 U13290 ( .A(n14944), .ZN(n14640) );
  INV_X1 U13291 ( .A(n10801), .ZN(n10694) );
  OAI211_X1 U13292 ( .C1(n14640), .C2(n10695), .A(n10694), .B(n6577), .ZN(
        n14639) );
  NOR2_X1 U13293 ( .A1(n14639), .A2(n13639), .ZN(n10696) );
  AOI211_X1 U13294 ( .C1(n13690), .C2(n14944), .A(n10697), .B(n10696), .ZN(
        n10698) );
  OAI211_X1 U13295 ( .C1(n14638), .C2(n13609), .A(n10699), .B(n10698), .ZN(
        P2_U3253) );
  NAND2_X1 U13296 ( .A1(n12631), .A2(n12714), .ZN(n10700) );
  NAND2_X1 U13297 ( .A1(n10702), .A2(n10708), .ZN(n10915) );
  OAI211_X1 U13298 ( .C1(n10702), .C2(n10708), .A(n10915), .B(n15149), .ZN(
        n10706) );
  OAI22_X1 U13299 ( .A1(n10703), .A2(n15195), .B1(n10921), .B2(n15193), .ZN(
        n10704) );
  INV_X1 U13300 ( .A(n10704), .ZN(n10705) );
  AND2_X1 U13301 ( .A1(n10706), .A2(n10705), .ZN(n15213) );
  NAND2_X1 U13302 ( .A1(n10707), .A2(n11981), .ZN(n10709) );
  INV_X1 U13303 ( .A(n10708), .ZN(n11979) );
  OR2_X1 U13304 ( .A1(n10709), .A2(n11979), .ZN(n10710) );
  NAND2_X1 U13305 ( .A1(n11114), .A2(n10710), .ZN(n15211) );
  NOR2_X1 U13306 ( .A1(n13081), .A2(n10711), .ZN(n10714) );
  INV_X1 U13307 ( .A(n12546), .ZN(n10712) );
  OAI22_X1 U13308 ( .A1(n15198), .A2(n10014), .B1(n10712), .B2(n15184), .ZN(
        n10713) );
  AOI211_X1 U13309 ( .C1(n15211), .C2(n14611), .A(n10714), .B(n10713), .ZN(
        n10715) );
  OAI21_X1 U13310 ( .B1(n15213), .B2(n14582), .A(n10715), .ZN(P3_U3226) );
  OAI21_X1 U13311 ( .B1(n10717), .B2(n13112), .A(n10716), .ZN(n10723) );
  OAI22_X1 U13312 ( .A1(n13163), .A2(n10721), .B1(n15235), .B2(n9989), .ZN(
        n10718) );
  AOI21_X1 U13313 ( .B1(n10723), .B2(n15235), .A(n10718), .ZN(n10719) );
  INV_X1 U13314 ( .A(n10719), .ZN(P3_U3465) );
  INV_X1 U13315 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n10720) );
  OAI22_X1 U13316 ( .A1(n10721), .A2(n13212), .B1(n15225), .B2(n10720), .ZN(
        n10722) );
  AOI21_X1 U13317 ( .B1(n10723), .B2(n15225), .A(n10722), .ZN(n10724) );
  INV_X1 U13318 ( .A(n10724), .ZN(P3_U3408) );
  INV_X1 U13319 ( .A(n10881), .ZN(n10888) );
  INV_X1 U13320 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13321 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n10888), .B1(n10881), 
        .B2(n10727), .ZN(n10728) );
  AOI21_X1 U13322 ( .B1(n10729), .B2(n10728), .A(n6725), .ZN(n10747) );
  NOR2_X1 U13323 ( .A1(n10730), .A2(n7313), .ZN(n10732) );
  MUX2_X1 U13324 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12862), .Z(n10887) );
  XNOR2_X1 U13325 ( .A(n10887), .B(n10881), .ZN(n10731) );
  INV_X1 U13326 ( .A(n10892), .ZN(n10735) );
  OAI21_X1 U13327 ( .B1(n10733), .B2(n10732), .A(n10731), .ZN(n10734) );
  NAND3_X1 U13328 ( .A1(n10735), .A2(n12767), .A3(n10734), .ZN(n10746) );
  INV_X1 U13329 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U13330 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10881), .B1(n10888), 
        .B2(n14623), .ZN(n10740) );
  NAND2_X1 U13331 ( .A1(n10736), .A2(n7313), .ZN(n10738) );
  NAND2_X1 U13332 ( .A1(n10738), .A2(n10737), .ZN(n10739) );
  NAND2_X1 U13333 ( .A1(n10740), .A2(n10739), .ZN(n10884) );
  OAI21_X1 U13334 ( .B1(n10740), .B2(n10739), .A(n10884), .ZN(n10744) );
  NOR2_X1 U13335 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10741), .ZN(n10968) );
  AOI21_X1 U13336 ( .B1(n15142), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n10968), 
        .ZN(n10742) );
  OAI21_X1 U13337 ( .B1(n12883), .B2(n10881), .A(n10742), .ZN(n10743) );
  AOI21_X1 U13338 ( .B1(n10744), .B2(n12895), .A(n10743), .ZN(n10745) );
  OAI211_X1 U13339 ( .C1(n10747), .C2(n12896), .A(n10746), .B(n10745), .ZN(
        P3_U3194) );
  INV_X1 U13340 ( .A(n11375), .ZN(n10785) );
  OAI222_X1 U13341 ( .A1(n14436), .A2(n10748), .B1(n14428), .B2(n10785), .C1(
        n6790), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13342 ( .A(n14996), .ZN(n15025) );
  AND2_X1 U13343 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10749) );
  AOI21_X1 U13344 ( .B1(n15025), .B2(n13438), .A(n10749), .ZN(n10750) );
  INV_X1 U13345 ( .A(n10750), .ZN(n10759) );
  INV_X1 U13346 ( .A(n10751), .ZN(n10752) );
  AOI21_X1 U13347 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n10762), .A(n10752), 
        .ZN(n10753) );
  NOR2_X1 U13348 ( .A1(n10753), .A2(n13424), .ZN(n10755) );
  XNOR2_X1 U13349 ( .A(n10753), .B(n13424), .ZN(n13419) );
  NOR2_X1 U13350 ( .A1(n10754), .A2(n13419), .ZN(n13420) );
  NOR2_X1 U13351 ( .A1(n10755), .A2(n13420), .ZN(n15021) );
  XNOR2_X1 U13352 ( .A(n15024), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15020) );
  NOR2_X1 U13353 ( .A1(n15021), .A2(n15020), .ZN(n15019) );
  AOI21_X1 U13354 ( .B1(n15024), .B2(P2_REG1_REG_16__SCAN_IN), .A(n15019), 
        .ZN(n10757) );
  XNOR2_X1 U13355 ( .A(n13438), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n10756) );
  NOR2_X1 U13356 ( .A1(n10757), .A2(n10756), .ZN(n13437) );
  AOI211_X1 U13357 ( .C1(n10757), .C2(n10756), .A(n13437), .B(n15018), .ZN(
        n10758) );
  AOI211_X1 U13358 ( .C1(n14949), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n10759), 
        .B(n10758), .ZN(n10774) );
  NOR2_X1 U13359 ( .A1(n10769), .A2(n11020), .ZN(n10760) );
  AOI21_X1 U13360 ( .B1(n11020), .B2(n10769), .A(n10760), .ZN(n15028) );
  NAND2_X1 U13361 ( .A1(n10762), .A2(n10761), .ZN(n10765) );
  OR2_X1 U13362 ( .A1(n10865), .A2(n10763), .ZN(n10764) );
  NAND2_X1 U13363 ( .A1(n10765), .A2(n10764), .ZN(n10767) );
  NAND2_X1 U13364 ( .A1(n10766), .A2(n10767), .ZN(n10768) );
  XNOR2_X1 U13365 ( .A(n13424), .B(n10767), .ZN(n13428) );
  NAND2_X1 U13366 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13428), .ZN(n13427) );
  NAND2_X1 U13367 ( .A1(n10768), .A2(n13427), .ZN(n15029) );
  NAND2_X1 U13368 ( .A1(n15028), .A2(n15029), .ZN(n15026) );
  OAI21_X1 U13369 ( .B1(n10769), .B2(n11020), .A(n15026), .ZN(n10772) );
  NOR2_X1 U13370 ( .A1(n13433), .A2(n11053), .ZN(n10770) );
  AOI21_X1 U13371 ( .B1(n11053), .B2(n13433), .A(n10770), .ZN(n10771) );
  INV_X1 U13372 ( .A(n14998), .ZN(n15027) );
  NAND2_X1 U13373 ( .A1(n10771), .A2(n10772), .ZN(n13432) );
  OAI211_X1 U13374 ( .C1(n10772), .C2(n10771), .A(n15027), .B(n13432), .ZN(
        n10773) );
  NAND2_X1 U13375 ( .A1(n10774), .A2(n10773), .ZN(P2_U3231) );
  AOI21_X1 U13376 ( .B1(n15118), .B2(n10776), .A(n10775), .ZN(n10777) );
  OAI211_X1 U13377 ( .C1(n12137), .C2(n10779), .A(n10778), .B(n10777), .ZN(
        n10783) );
  NAND2_X1 U13378 ( .A1(n10783), .A2(n15141), .ZN(n10780) );
  OAI21_X1 U13379 ( .B1(n15141), .B2(n8642), .A(n10780), .ZN(P2_U3510) );
  NAND2_X1 U13380 ( .A1(n10783), .A2(n15129), .ZN(n10784) );
  OAI21_X1 U13381 ( .B1(n15129), .B2(n8641), .A(n10784), .ZN(P2_U3463) );
  OAI222_X1 U13382 ( .A1(n13820), .A2(n10786), .B1(P2_U3088), .B2(n8879), .C1(
        n13818), .C2(n10785), .ZN(P2_U3307) );
  INV_X1 U13383 ( .A(n10787), .ZN(n10793) );
  INV_X1 U13384 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10790) );
  INV_X1 U13385 ( .A(n10788), .ZN(n10789) );
  MUX2_X1 U13386 ( .A(n10790), .B(n10789), .S(n15198), .Z(n10792) );
  AOI22_X1 U13387 ( .A1(n14583), .A2(n12632), .B1(n15178), .B2(n12633), .ZN(
        n10791) );
  OAI211_X1 U13388 ( .C1(n10793), .C2(n12983), .A(n10792), .B(n10791), .ZN(
        P3_U3228) );
  OR2_X1 U13389 ( .A1(n12227), .A2(n14931), .ZN(n10854) );
  NAND2_X1 U13390 ( .A1(n12227), .A2(n14931), .ZN(n10856) );
  NAND2_X1 U13391 ( .A1(n10854), .A2(n10856), .ZN(n12418) );
  XOR2_X1 U13392 ( .A(n12418), .B(n10860), .Z(n14637) );
  INV_X1 U13393 ( .A(n14637), .ZN(n10808) );
  NAND2_X1 U13394 ( .A1(n14640), .A2(n13312), .ZN(n10796) );
  XOR2_X1 U13395 ( .A(n10857), .B(n12418), .Z(n10799) );
  OAI21_X1 U13396 ( .B1(n10799), .B2(n10902), .A(n10798), .ZN(n14636) );
  AND2_X1 U13397 ( .A1(n14634), .A2(n10801), .ZN(n10862) );
  INV_X1 U13398 ( .A(n10862), .ZN(n10800) );
  OAI211_X1 U13399 ( .C1(n14634), .C2(n10801), .A(n10800), .B(n6577), .ZN(
        n14633) );
  OAI22_X1 U13400 ( .A1(n15045), .A2(n10803), .B1(n10802), .B2(n15037), .ZN(
        n10804) );
  AOI21_X1 U13401 ( .B1(n12227), .B2(n13690), .A(n10804), .ZN(n10805) );
  OAI21_X1 U13402 ( .B1(n14633), .B2(n13639), .A(n10805), .ZN(n10806) );
  AOI21_X1 U13403 ( .B1(n14636), .B2(n15045), .A(n10806), .ZN(n10807) );
  OAI21_X1 U13404 ( .B1(n10808), .B2(n13697), .A(n10807), .ZN(P2_U3252) );
  MUX2_X1 U13405 ( .A(n10810), .B(n10809), .S(n15235), .Z(n10811) );
  OAI21_X1 U13406 ( .B1(n13163), .B2(n10812), .A(n10811), .ZN(P3_U3464) );
  OAI21_X1 U13407 ( .B1(n10815), .B2(n10814), .A(n10813), .ZN(n10816) );
  NAND2_X1 U13408 ( .A1(n10816), .A2(n7445), .ZN(n10823) );
  INV_X1 U13409 ( .A(n10864), .ZN(n10821) );
  OR2_X1 U13410 ( .A1(n14931), .A2(n13595), .ZN(n10817) );
  OAI21_X1 U13411 ( .B1(n12239), .B2(n15039), .A(n10817), .ZN(n10858) );
  INV_X1 U13412 ( .A(n10858), .ZN(n10819) );
  OAI22_X1 U13413 ( .A1(n10819), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10818), .ZN(n10820) );
  AOI21_X1 U13414 ( .B1(n10821), .B2(n13265), .A(n10820), .ZN(n10822) );
  OAI211_X1 U13415 ( .C1(n12234), .C2(n13297), .A(n10823), .B(n10822), .ZN(
        P2_U3187) );
  NAND2_X1 U13416 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  NAND2_X1 U13417 ( .A1(n13877), .A2(n11787), .ZN(n10829) );
  NAND2_X1 U13418 ( .A1(n13978), .A2(n11786), .ZN(n10828) );
  NAND2_X1 U13419 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  XNOR2_X1 U13420 ( .A(n10830), .B(n11692), .ZN(n10833) );
  AND2_X1 U13421 ( .A1(n13978), .A2(n11757), .ZN(n10831) );
  AOI21_X1 U13422 ( .B1(n13877), .B2(n11788), .A(n10831), .ZN(n10834) );
  XNOR2_X1 U13423 ( .A(n10833), .B(n10834), .ZN(n13874) );
  INV_X1 U13424 ( .A(n10833), .ZN(n10836) );
  INV_X1 U13425 ( .A(n10834), .ZN(n10835) );
  NAND2_X1 U13426 ( .A1(n10836), .A2(n10835), .ZN(n10837) );
  NAND2_X1 U13427 ( .A1(n13871), .A2(n10837), .ZN(n11684) );
  NAND2_X1 U13428 ( .A1(n14660), .A2(n11787), .ZN(n10840) );
  NAND2_X1 U13429 ( .A1(n13977), .A2(n11786), .ZN(n10839) );
  NAND2_X1 U13430 ( .A1(n10840), .A2(n10839), .ZN(n10841) );
  XNOR2_X1 U13431 ( .A(n10841), .B(n11789), .ZN(n11687) );
  AND2_X1 U13432 ( .A1(n13977), .A2(n11757), .ZN(n10842) );
  AOI21_X1 U13433 ( .B1(n14660), .B2(n11788), .A(n10842), .ZN(n11685) );
  XNOR2_X1 U13434 ( .A(n11687), .B(n11685), .ZN(n11683) );
  XNOR2_X1 U13435 ( .A(n10838), .B(n11683), .ZN(n10850) );
  OAI21_X1 U13436 ( .B1(n13962), .B2(n10844), .A(n10843), .ZN(n10845) );
  AOI21_X1 U13437 ( .B1(n13966), .B2(n14278), .A(n10845), .ZN(n10846) );
  OAI21_X1 U13438 ( .B1(n13963), .B2(n10847), .A(n10846), .ZN(n10848) );
  AOI21_X1 U13439 ( .B1(n14660), .B2(n6564), .A(n10848), .ZN(n10849) );
  OAI21_X1 U13440 ( .B1(n10850), .B2(n13955), .A(n10849), .ZN(P1_U3234) );
  INV_X1 U13441 ( .A(n10851), .ZN(n10853) );
  OAI222_X1 U13442 ( .A1(P3_U3151), .A2(n7636), .B1(n13227), .B2(n10853), .C1(
        n10852), .C2(n13228), .ZN(P3_U3271) );
  XNOR2_X1 U13443 ( .A(n12235), .B(n12233), .ZN(n12424) );
  INV_X1 U13444 ( .A(n10854), .ZN(n10855) );
  XOR2_X1 U13445 ( .A(n12424), .B(n10901), .Z(n10859) );
  AOI21_X1 U13446 ( .B1(n10859), .B2(n13683), .A(n10858), .ZN(n10874) );
  XNOR2_X1 U13447 ( .A(n10900), .B(n12424), .ZN(n10875) );
  INV_X1 U13448 ( .A(n10875), .ZN(n10869) );
  AND2_X2 U13449 ( .A1(n12234), .A2(n10862), .ZN(n10907) );
  NOR2_X1 U13450 ( .A1(n12234), .A2(n10862), .ZN(n10863) );
  OR3_X1 U13451 ( .A1(n10907), .A2(n10863), .A3(n8705), .ZN(n10871) );
  OAI22_X1 U13452 ( .A1(n15045), .A2(n10865), .B1(n10864), .B2(n15037), .ZN(
        n10866) );
  AOI21_X1 U13453 ( .B1(n12235), .B2(n13690), .A(n10866), .ZN(n10867) );
  OAI21_X1 U13454 ( .B1(n10871), .B2(n13639), .A(n10867), .ZN(n10868) );
  AOI21_X1 U13455 ( .B1(n10869), .B2(n13644), .A(n10868), .ZN(n10870) );
  OAI21_X1 U13456 ( .B1(n6578), .B2(n10874), .A(n10870), .ZN(P2_U3251) );
  INV_X1 U13457 ( .A(n10871), .ZN(n10872) );
  AOI21_X1 U13458 ( .B1(n15118), .B2(n12235), .A(n10872), .ZN(n10873) );
  OAI211_X1 U13459 ( .C1(n10875), .C2(n15078), .A(n10874), .B(n10873), .ZN(
        n10878) );
  NAND2_X1 U13460 ( .A1(n10878), .A2(n15141), .ZN(n10876) );
  OAI21_X1 U13461 ( .B1(n15141), .B2(n10877), .A(n10876), .ZN(P2_U3513) );
  NAND2_X1 U13462 ( .A1(n10878), .A2(n15129), .ZN(n10879) );
  OAI21_X1 U13463 ( .B1(n15129), .B2(n8698), .A(n10879), .ZN(P2_U3472) );
  OAI222_X1 U13464 ( .A1(n13820), .A2(n15495), .B1(P2_U3088), .B2(n12352), 
        .C1(n13818), .C2(n10880), .ZN(P2_U3305) );
  INV_X1 U13465 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n10883) );
  AOI21_X1 U13466 ( .B1(n10883), .B2(n10882), .A(n10979), .ZN(n10899) );
  XNOR2_X1 U13467 ( .A(n7323), .B(n10984), .ZN(n10885) );
  NAND2_X1 U13468 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n10885), .ZN(n10985) );
  OAI21_X1 U13469 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n10885), .A(n10985), 
        .ZN(n10897) );
  AND2_X1 U13470 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n10947) );
  AOI21_X1 U13471 ( .B1(n15142), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n10947), 
        .ZN(n10886) );
  OAI21_X1 U13472 ( .B1(n12883), .B2(n10992), .A(n10886), .ZN(n10896) );
  INV_X1 U13473 ( .A(n10887), .ZN(n10889) );
  NOR2_X1 U13474 ( .A1(n10889), .A2(n10888), .ZN(n10891) );
  MUX2_X1 U13475 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12862), .Z(n10993) );
  XNOR2_X1 U13476 ( .A(n10993), .B(n10992), .ZN(n10890) );
  INV_X1 U13477 ( .A(n10998), .ZN(n10894) );
  OAI21_X1 U13478 ( .B1(n10892), .B2(n10891), .A(n10890), .ZN(n10893) );
  AOI21_X1 U13479 ( .B1(n10894), .B2(n10893), .A(n12891), .ZN(n10895) );
  AOI211_X1 U13480 ( .C1(n12895), .C2(n10897), .A(n10896), .B(n10895), .ZN(
        n10898) );
  OAI21_X1 U13481 ( .B1(n10899), .B2(n12896), .A(n10898), .ZN(P3_U3195) );
  XOR2_X1 U13482 ( .A(n12425), .B(n11016), .Z(n13781) );
  AOI211_X1 U13483 ( .C1(n12425), .C2(n10903), .A(n10902), .B(n11012), .ZN(
        n10905) );
  OAI22_X1 U13484 ( .A1(n12233), .A2(n13595), .B1(n12249), .B2(n15039), .ZN(
        n10904) );
  NOR2_X1 U13485 ( .A1(n10905), .A2(n10904), .ZN(n13780) );
  OAI21_X1 U13486 ( .B1(n10934), .B2(n15037), .A(n13780), .ZN(n10906) );
  NAND2_X1 U13487 ( .A1(n10906), .A2(n15045), .ZN(n10913) );
  INV_X1 U13488 ( .A(n10907), .ZN(n10909) );
  NAND2_X1 U13489 ( .A1(n6586), .A2(n10907), .ZN(n11022) );
  INV_X1 U13490 ( .A(n11022), .ZN(n10908) );
  AOI211_X1 U13491 ( .C1(n13778), .C2(n10909), .A(n8705), .B(n10908), .ZN(
        n13777) );
  OAI22_X1 U13492 ( .A1(n6586), .A2(n13677), .B1(n15045), .B2(n10910), .ZN(
        n10911) );
  AOI21_X1 U13493 ( .B1(n13777), .B2(n13694), .A(n10911), .ZN(n10912) );
  OAI211_X1 U13494 ( .C1(n13697), .C2(n13781), .A(n10913), .B(n10912), .ZN(
        P2_U3250) );
  NAND2_X1 U13495 ( .A1(n12748), .A2(n15209), .ZN(n10914) );
  NAND2_X1 U13496 ( .A1(n10921), .A2(n12600), .ZN(n11988) );
  NAND2_X1 U13497 ( .A1(n12747), .A2(n10916), .ZN(n11987) );
  NAND2_X1 U13498 ( .A1(n11988), .A2(n11987), .ZN(n10955) );
  NAND2_X1 U13499 ( .A1(n10956), .A2(n10955), .ZN(n10954) );
  NAND2_X1 U13500 ( .A1(n10921), .A2(n10916), .ZN(n10917) );
  NAND2_X1 U13501 ( .A1(n10954), .A2(n10917), .ZN(n10918) );
  XNOR2_X1 U13502 ( .A(n15153), .B(n12675), .ZN(n11990) );
  AOI21_X1 U13503 ( .B1(n10918), .B2(n11990), .A(n15191), .ZN(n10923) );
  INV_X1 U13504 ( .A(n10918), .ZN(n10920) );
  OAI22_X1 U13505 ( .A1(n10921), .A2(n15195), .B1(n14602), .B2(n15193), .ZN(
        n10922) );
  AOI21_X1 U13506 ( .B1(n10923), .B2(n11097), .A(n10922), .ZN(n11030) );
  NAND2_X1 U13507 ( .A1(n11114), .A2(n11983), .ZN(n10953) );
  INV_X1 U13508 ( .A(n10955), .ZN(n11985) );
  NAND2_X1 U13509 ( .A1(n10953), .A2(n11985), .ZN(n15144) );
  NAND2_X1 U13510 ( .A1(n15144), .A2(n11988), .ZN(n10924) );
  XNOR2_X1 U13511 ( .A(n10924), .B(n11990), .ZN(n11028) );
  AOI22_X1 U13512 ( .A1(n14582), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n15178), 
        .B2(n12676), .ZN(n10925) );
  OAI21_X1 U13513 ( .B1(n13081), .B2(n11109), .A(n10925), .ZN(n10926) );
  AOI21_X1 U13514 ( .B1(n11028), .B2(n14611), .A(n10926), .ZN(n10927) );
  OAI21_X1 U13515 ( .B1(n11030), .B2(n14582), .A(n10927), .ZN(P3_U3224) );
  INV_X1 U13516 ( .A(n10928), .ZN(n10930) );
  OAI222_X1 U13517 ( .A1(n13227), .A2(n10930), .B1(P3_U3151), .B2(n8176), .C1(
        n10929), .C2(n13228), .ZN(P3_U3270) );
  OAI211_X1 U13518 ( .C1(n10933), .C2(n10932), .A(n10931), .B(n7445), .ZN(
        n10938) );
  INV_X1 U13519 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13423) );
  OAI22_X1 U13520 ( .A1(n14933), .A2(n12233), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13423), .ZN(n10936) );
  OAI22_X1 U13521 ( .A1(n14932), .A2(n12249), .B1(n14947), .B2(n10934), .ZN(
        n10935) );
  AOI211_X1 U13522 ( .C1(n13778), .C2(n14943), .A(n10936), .B(n10935), .ZN(
        n10937) );
  NAND2_X1 U13523 ( .A1(n10938), .A2(n10937), .ZN(P2_U3213) );
  INV_X1 U13524 ( .A(n10939), .ZN(n10940) );
  OAI222_X1 U13525 ( .A1(n10941), .A2(P3_U3151), .B1(n13228), .B2(n15368), 
        .C1(n13227), .C2(n10940), .ZN(P3_U3269) );
  INV_X1 U13526 ( .A(n10942), .ZN(n10944) );
  NAND2_X1 U13527 ( .A1(n10944), .A2(n10943), .ZN(n10945) );
  XNOR2_X1 U13528 ( .A(n10946), .B(n10945), .ZN(n10952) );
  NOR2_X1 U13529 ( .A1(n12734), .A2(n13211), .ZN(n10950) );
  INV_X1 U13530 ( .A(n13075), .ZN(n12744) );
  AOI21_X1 U13531 ( .B1(n12713), .B2(n12744), .A(n10947), .ZN(n10948) );
  OAI21_X1 U13532 ( .B1(n14603), .B2(n12685), .A(n10948), .ZN(n10949) );
  AOI211_X1 U13533 ( .C1(n11133), .C2(n12731), .A(n10950), .B(n10949), .ZN(
        n10951) );
  OAI21_X1 U13534 ( .B1(n10952), .B2(n12699), .A(n10951), .ZN(P3_U3174) );
  XNOR2_X1 U13535 ( .A(n10953), .B(n10955), .ZN(n10961) );
  OAI21_X1 U13536 ( .B1(n10956), .B2(n10955), .A(n10954), .ZN(n10957) );
  NAND2_X1 U13537 ( .A1(n10957), .A2(n15149), .ZN(n10959) );
  AOI22_X1 U13538 ( .A1(n12748), .A2(n15154), .B1(n15155), .B2(n15153), .ZN(
        n10958) );
  OAI211_X1 U13539 ( .C1(n10961), .C2(n12922), .A(n10959), .B(n10958), .ZN(
        n15215) );
  MUX2_X1 U13540 ( .A(n15215), .B(P3_REG2_REG_8__SCAN_IN), .S(n14582), .Z(
        n10960) );
  INV_X1 U13541 ( .A(n10960), .ZN(n10967) );
  INV_X1 U13542 ( .A(n10961), .ZN(n15218) );
  INV_X1 U13543 ( .A(n15175), .ZN(n10962) );
  NAND2_X1 U13544 ( .A1(n15198), .A2(n10962), .ZN(n12934) );
  INV_X1 U13545 ( .A(n12934), .ZN(n10965) );
  NAND2_X1 U13546 ( .A1(n12600), .A2(n15210), .ZN(n15214) );
  INV_X1 U13547 ( .A(n12601), .ZN(n10963) );
  OAI22_X1 U13548 ( .A1(n14596), .A2(n15214), .B1(n10963), .B2(n15184), .ZN(
        n10964) );
  AOI21_X1 U13549 ( .B1(n15218), .B2(n10965), .A(n10964), .ZN(n10966) );
  NAND2_X1 U13550 ( .A1(n10967), .A2(n10966), .ZN(P3_U3225) );
  AOI21_X1 U13551 ( .B1(n12713), .B2(n14591), .A(n10968), .ZN(n10970) );
  NAND2_X1 U13552 ( .A1(n12726), .A2(n15156), .ZN(n10969) );
  OAI211_X1 U13553 ( .C1(n12734), .C2(n14597), .A(n10970), .B(n10969), .ZN(
        n10976) );
  NAND2_X1 U13554 ( .A1(n10971), .A2(n10972), .ZN(n10973) );
  AOI21_X1 U13555 ( .B1(n10974), .B2(n10973), .A(n12699), .ZN(n10975) );
  AOI211_X1 U13556 ( .C1(n14593), .C2(n12731), .A(n10976), .B(n10975), .ZN(
        n10977) );
  INV_X1 U13557 ( .A(n10977), .ZN(P3_U3164) );
  NOR2_X1 U13558 ( .A1(n7323), .A2(n10978), .ZN(n10980) );
  NAND2_X1 U13559 ( .A1(n10991), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12787) );
  INV_X1 U13560 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U13561 ( .A1(n10987), .A2(n10981), .ZN(n10982) );
  NAND2_X1 U13562 ( .A1(n12787), .A2(n10982), .ZN(n10996) );
  AOI21_X1 U13563 ( .B1(n10983), .B2(n10996), .A(n12778), .ZN(n11005) );
  NAND2_X1 U13564 ( .A1(n10992), .A2(n10984), .ZN(n10986) );
  INV_X1 U13565 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13157) );
  NAND2_X1 U13566 ( .A1(n10991), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12783) );
  INV_X1 U13567 ( .A(n12783), .ZN(n12788) );
  AOI21_X1 U13568 ( .B1(n10987), .B2(n13157), .A(n12788), .ZN(n10994) );
  NAND2_X1 U13569 ( .A1(n10994), .A2(n10988), .ZN(n12782) );
  OAI21_X1 U13570 ( .B1(n10988), .B2(n10994), .A(n12782), .ZN(n11003) );
  INV_X1 U13571 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n10989) );
  NOR2_X1 U13572 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10989), .ZN(n11035) );
  AOI21_X1 U13573 ( .B1(n15142), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11035), 
        .ZN(n10990) );
  OAI21_X1 U13574 ( .B1(n12883), .B2(n10991), .A(n10990), .ZN(n11002) );
  NOR2_X1 U13575 ( .A1(n10993), .A2(n10992), .ZN(n10997) );
  OR2_X1 U13576 ( .A1(n10998), .A2(n10997), .ZN(n11000) );
  INV_X1 U13577 ( .A(n10994), .ZN(n10995) );
  MUX2_X1 U13578 ( .A(n10996), .B(n10995), .S(n12862), .Z(n10999) );
  AOI211_X1 U13579 ( .C1(n11000), .C2(n10999), .A(n12891), .B(n12791), .ZN(
        n11001) );
  AOI211_X1 U13580 ( .C1(n12895), .C2(n11003), .A(n11002), .B(n11001), .ZN(
        n11004) );
  OAI21_X1 U13581 ( .B1(n11005), .B2(n12896), .A(n11004), .ZN(P3_U3196) );
  NAND2_X1 U13582 ( .A1(n11428), .A2(n11006), .ZN(n11008) );
  NOR2_X1 U13583 ( .A1(n11007), .A2(P2_U3088), .ZN(n12456) );
  OAI211_X1 U13584 ( .C1(n11009), .C2(n13820), .A(n11008), .B(n7541), .ZN(
        P2_U3304) );
  NAND2_X1 U13585 ( .A1(n11428), .A2(n11010), .ZN(n11011) );
  OAI211_X1 U13586 ( .C1(n15419), .C2(n14436), .A(n11011), .B(n11627), .ZN(
        P1_U3332) );
  INV_X1 U13587 ( .A(n12239), .ZN(n13310) );
  XNOR2_X1 U13588 ( .A(n13773), .B(n13309), .ZN(n12420) );
  OAI21_X1 U13589 ( .B1(n11013), .B2(n12420), .A(n11049), .ZN(n11015) );
  AOI22_X1 U13590 ( .A1(n13310), .A2(n13667), .B1(n13665), .B2(n13308), .ZN(
        n11043) );
  INV_X1 U13591 ( .A(n11043), .ZN(n11014) );
  AOI21_X1 U13592 ( .B1(n11015), .B2(n13683), .A(n11014), .ZN(n13775) );
  INV_X1 U13593 ( .A(n12420), .ZN(n11017) );
  OAI21_X1 U13594 ( .B1(n11018), .B2(n11017), .A(n11052), .ZN(n13776) );
  INV_X1 U13595 ( .A(n11046), .ZN(n11019) );
  OAI22_X1 U13596 ( .A1(n15045), .A2(n11020), .B1(n11019), .B2(n15037), .ZN(
        n11021) );
  AOI21_X1 U13597 ( .B1(n13773), .B2(n13690), .A(n11021), .ZN(n11025) );
  AOI21_X1 U13598 ( .B1(n11022), .B2(n13773), .A(n8705), .ZN(n11023) );
  AND2_X1 U13599 ( .A1(n11023), .A2(n11055), .ZN(n13772) );
  NAND2_X1 U13600 ( .A1(n13772), .A2(n13694), .ZN(n11024) );
  OAI211_X1 U13601 ( .C1(n13776), .C2(n13697), .A(n11025), .B(n11024), .ZN(
        n11026) );
  INV_X1 U13602 ( .A(n11026), .ZN(n11027) );
  OAI21_X1 U13603 ( .B1(n6578), .B2(n13775), .A(n11027), .ZN(P2_U3249) );
  NAND2_X1 U13604 ( .A1(n11028), .A2(n15221), .ZN(n11029) );
  AND2_X1 U13605 ( .A1(n11030), .A2(n11029), .ZN(n11033) );
  MUX2_X1 U13606 ( .A(n10555), .B(n11033), .S(n15235), .Z(n11031) );
  OAI21_X1 U13607 ( .B1(n13163), .B2(n11109), .A(n11031), .ZN(P3_U3468) );
  INV_X1 U13608 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11032) );
  MUX2_X1 U13609 ( .A(n11033), .B(n11032), .S(n15223), .Z(n11034) );
  OAI21_X1 U13610 ( .B1(n13212), .B2(n11109), .A(n11034), .ZN(P3_U3417) );
  XOR2_X1 U13611 ( .A(n11138), .B(n7959), .Z(n11040) );
  INV_X1 U13612 ( .A(n13062), .ZN(n11866) );
  AOI21_X1 U13613 ( .B1(n12726), .B2(n14591), .A(n11035), .ZN(n11036) );
  OAI21_X1 U13614 ( .B1(n11866), .B2(n12729), .A(n11036), .ZN(n11038) );
  INV_X1 U13615 ( .A(n12462), .ZN(n13208) );
  NOR2_X1 U13616 ( .A1(n13208), .A2(n12734), .ZN(n11037) );
  AOI211_X1 U13617 ( .C1(n11124), .C2(n12731), .A(n11038), .B(n11037), .ZN(
        n11039) );
  OAI21_X1 U13618 ( .B1(n11040), .B2(n12699), .A(n11039), .ZN(P3_U3155) );
  AOI21_X1 U13619 ( .B1(n11042), .B2(n11041), .A(n11086), .ZN(n11048) );
  INV_X1 U13620 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15518) );
  OAI22_X1 U13621 ( .A1(n11043), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15518), .ZN(n11045) );
  NOR2_X1 U13622 ( .A1(n12251), .A2(n13297), .ZN(n11044) );
  AOI211_X1 U13623 ( .C1(n13265), .C2(n11046), .A(n11045), .B(n11044), .ZN(
        n11047) );
  OAI21_X1 U13624 ( .B1(n11048), .B2(n14939), .A(n11047), .ZN(P2_U3198) );
  XNOR2_X1 U13625 ( .A(n13768), .B(n13308), .ZN(n12422) );
  XNOR2_X1 U13626 ( .A(n11072), .B(n12422), .ZN(n11051) );
  AOI22_X1 U13627 ( .A1(n13505), .A2(n13665), .B1(n13309), .B2(n13667), .ZN(
        n11091) );
  INV_X1 U13628 ( .A(n11091), .ZN(n11050) );
  AOI21_X1 U13629 ( .B1(n11051), .B2(n13683), .A(n11050), .ZN(n13770) );
  INV_X1 U13630 ( .A(n12422), .ZN(n11078) );
  XNOR2_X1 U13631 ( .A(n11079), .B(n11078), .ZN(n13771) );
  OAI22_X1 U13632 ( .A1(n15045), .A2(n11053), .B1(n11089), .B2(n15037), .ZN(
        n11054) );
  AOI21_X1 U13633 ( .B1(n13768), .B2(n13690), .A(n11054), .ZN(n11058) );
  AOI21_X1 U13634 ( .B1(n11055), .B2(n13768), .A(n8705), .ZN(n11056) );
  AND2_X1 U13635 ( .A1(n11056), .A2(n11074), .ZN(n13767) );
  NAND2_X1 U13636 ( .A1(n13767), .A2(n13694), .ZN(n11057) );
  OAI211_X1 U13637 ( .C1(n13771), .C2(n13697), .A(n11058), .B(n11057), .ZN(
        n11059) );
  INV_X1 U13638 ( .A(n11059), .ZN(n11060) );
  OAI21_X1 U13639 ( .B1(n6578), .B2(n13770), .A(n11060), .ZN(P2_U3248) );
  INV_X1 U13640 ( .A(n11443), .ZN(n11063) );
  OAI222_X1 U13641 ( .A1(n13820), .A2(n15323), .B1(n13818), .B2(n11063), .C1(
        P2_U3088), .C2(n11061), .ZN(P2_U3303) );
  OAI222_X1 U13642 ( .A1(n14436), .A2(n7160), .B1(n14428), .B2(n11063), .C1(
        n11062), .C2(P1_U3086), .ZN(P1_U3331) );
  XNOR2_X1 U13643 ( .A(n11064), .B(n13076), .ZN(n11065) );
  XNOR2_X1 U13644 ( .A(n11066), .B(n11065), .ZN(n11071) );
  NAND2_X1 U13645 ( .A1(n12726), .A2(n13062), .ZN(n11067) );
  NAND2_X1 U13646 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12809)
         );
  OAI211_X1 U13647 ( .C1(n13041), .C2(n12729), .A(n11067), .B(n12809), .ZN(
        n11069) );
  INV_X1 U13648 ( .A(n13147), .ZN(n13070) );
  NOR2_X1 U13649 ( .A1(n13070), .A2(n12734), .ZN(n11068) );
  AOI211_X1 U13650 ( .C1(n13068), .C2(n12731), .A(n11069), .B(n11068), .ZN(
        n11070) );
  OAI21_X1 U13651 ( .B1(n11071), .B2(n12699), .A(n11070), .ZN(P3_U3166) );
  INV_X1 U13652 ( .A(n13308), .ZN(n12254) );
  INV_X1 U13653 ( .A(n13505), .ZN(n13477) );
  XNOR2_X1 U13654 ( .A(n13763), .B(n13477), .ZN(n12426) );
  XOR2_X1 U13655 ( .A(n13476), .B(n12426), .Z(n11073) );
  AOI222_X1 U13656 ( .A1(n13683), .A2(n11073), .B1(n13308), .B2(n13667), .C1(
        n13668), .C2(n13665), .ZN(n13765) );
  AOI211_X1 U13657 ( .C1(n13763), .C2(n11074), .A(n8705), .B(n7043), .ZN(
        n13762) );
  NOR2_X1 U13658 ( .A1(n13478), .A2(n13677), .ZN(n11077) );
  OAI22_X1 U13659 ( .A1(n15045), .A2(n11075), .B1(n13292), .B2(n15037), .ZN(
        n11076) );
  AOI211_X1 U13660 ( .C1(n13762), .C2(n13694), .A(n11077), .B(n11076), .ZN(
        n11082) );
  OAI21_X1 U13661 ( .B1(n11080), .B2(n12426), .A(n13504), .ZN(n13761) );
  NAND2_X1 U13662 ( .A1(n13761), .A2(n13644), .ZN(n11081) );
  OAI211_X1 U13663 ( .C1(n13765), .C2(n6578), .A(n11082), .B(n11081), .ZN(
        P2_U3247) );
  INV_X1 U13664 ( .A(n11083), .ZN(n11088) );
  NOR3_X1 U13665 ( .A1(n11086), .A2(n11085), .A3(n11084), .ZN(n11087) );
  OAI21_X1 U13666 ( .B1(n11088), .B2(n11087), .A(n7445), .ZN(n11095) );
  INV_X1 U13667 ( .A(n11089), .ZN(n11093) );
  OAI22_X1 U13668 ( .A1(n11091), .A2(n13238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11090), .ZN(n11092) );
  AOI21_X1 U13669 ( .B1(n11093), .B2(n13265), .A(n11092), .ZN(n11094) );
  OAI211_X1 U13670 ( .C1(n7045), .C2(n13297), .A(n11095), .B(n11094), .ZN(
        P2_U3200) );
  NAND2_X1 U13671 ( .A1(n15153), .A2(n12675), .ZN(n11096) );
  NAND2_X1 U13672 ( .A1(n14602), .A2(n15159), .ZN(n11938) );
  INV_X1 U13673 ( .A(n15159), .ZN(n11995) );
  NAND2_X1 U13674 ( .A1(n12746), .A2(n11995), .ZN(n11110) );
  NAND2_X1 U13675 ( .A1(n11938), .A2(n11110), .ZN(n15151) );
  NAND2_X1 U13676 ( .A1(n12746), .A2(n15159), .ZN(n14586) );
  NAND2_X1 U13677 ( .A1(n14603), .A2(n14597), .ZN(n11101) );
  INV_X1 U13678 ( .A(n11101), .ZN(n11099) );
  NAND2_X1 U13679 ( .A1(n15156), .A2(n12694), .ZN(n14588) );
  AND2_X1 U13680 ( .A1(n6699), .A2(n14588), .ZN(n11098) );
  OR2_X1 U13681 ( .A1(n11099), .A2(n11098), .ZN(n11100) );
  INV_X1 U13682 ( .A(n11100), .ZN(n11103) );
  NAND2_X1 U13683 ( .A1(n12691), .A2(n14610), .ZN(n14587) );
  AND2_X1 U13684 ( .A1(n14587), .A2(n11101), .ZN(n11102) );
  OR2_X1 U13685 ( .A1(n13211), .A2(n14591), .ZN(n11123) );
  NAND2_X1 U13686 ( .A1(n13211), .A2(n14591), .ZN(n12007) );
  NAND2_X1 U13687 ( .A1(n11123), .A2(n12007), .ZN(n11129) );
  AND2_X1 U13688 ( .A1(n13211), .A2(n11104), .ZN(n11105) );
  OR2_X1 U13689 ( .A1(n12462), .A2(n13075), .ZN(n12014) );
  NAND2_X1 U13690 ( .A1(n12462), .A2(n13075), .ZN(n12022) );
  NAND2_X1 U13691 ( .A1(n12014), .A2(n12022), .ZN(n12010) );
  NAND2_X1 U13692 ( .A1(n11106), .A2(n12010), .ZN(n12464) );
  OAI211_X1 U13693 ( .C1(n11106), .C2(n12010), .A(n12464), .B(n15149), .ZN(
        n11108) );
  AOI22_X1 U13694 ( .A1(n15154), .A2(n14591), .B1(n13062), .B2(n15155), .ZN(
        n11107) );
  NAND2_X1 U13695 ( .A1(n11108), .A2(n11107), .ZN(n13155) );
  INV_X1 U13696 ( .A(n13155), .ZN(n11128) );
  NAND2_X1 U13697 ( .A1(n15153), .A2(n11109), .ZN(n15145) );
  AND2_X1 U13698 ( .A1(n15145), .A2(n11110), .ZN(n11116) );
  INV_X1 U13699 ( .A(n11116), .ZN(n11112) );
  NAND2_X1 U13700 ( .A1(n11111), .A2(n12675), .ZN(n11992) );
  AND2_X1 U13701 ( .A1(n11988), .A2(n11992), .ZN(n15143) );
  OR2_X1 U13702 ( .A1(n11112), .A2(n15143), .ZN(n11115) );
  AND2_X1 U13703 ( .A1(n11983), .A2(n11115), .ZN(n11113) );
  NAND2_X1 U13704 ( .A1(n11114), .A2(n11113), .ZN(n11120) );
  INV_X1 U13705 ( .A(n11115), .ZN(n11118) );
  AND2_X1 U13706 ( .A1(n11985), .A2(n11116), .ZN(n11117) );
  OR2_X1 U13707 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  NAND2_X1 U13708 ( .A1(n12691), .A2(n12694), .ZN(n11939) );
  NAND2_X1 U13709 ( .A1(n15156), .A2(n14610), .ZN(n12001) );
  NAND2_X1 U13710 ( .A1(n14609), .A2(n14608), .ZN(n14607) );
  NAND2_X1 U13711 ( .A1(n14603), .A2(n11121), .ZN(n12006) );
  NAND2_X1 U13712 ( .A1(n12745), .A2(n14597), .ZN(n12003) );
  INV_X1 U13713 ( .A(n11123), .ZN(n12008) );
  XNOR2_X1 U13714 ( .A(n11865), .B(n12010), .ZN(n13156) );
  AOI22_X1 U13715 ( .A1(n14582), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15178), 
        .B2(n11124), .ZN(n11125) );
  OAI21_X1 U13716 ( .B1(n13081), .B2(n13208), .A(n11125), .ZN(n11126) );
  AOI21_X1 U13717 ( .B1(n13156), .B2(n14611), .A(n11126), .ZN(n11127) );
  OAI21_X1 U13718 ( .B1(n11128), .B2(n14582), .A(n11127), .ZN(P3_U3219) );
  XNOR2_X1 U13719 ( .A(n11130), .B(n12005), .ZN(n11131) );
  OAI222_X1 U13720 ( .A1(n15193), .A2(n13075), .B1(n15195), .B2(n14603), .C1(
        n15191), .C2(n11131), .ZN(n13159) );
  INV_X1 U13721 ( .A(n13159), .ZN(n11137) );
  XNOR2_X1 U13722 ( .A(n11132), .B(n12005), .ZN(n13160) );
  AOI22_X1 U13723 ( .A1(n14582), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15178), 
        .B2(n11133), .ZN(n11134) );
  OAI21_X1 U13724 ( .B1(n13081), .B2(n13211), .A(n11134), .ZN(n11135) );
  AOI21_X1 U13725 ( .B1(n13160), .B2(n14611), .A(n11135), .ZN(n11136) );
  OAI21_X1 U13726 ( .B1(n11137), .B2(n14582), .A(n11136), .ZN(P3_U3220) );
  INV_X1 U13727 ( .A(n12466), .ZN(n13204) );
  OR2_X1 U13728 ( .A1(n7959), .A2(n11138), .ZN(n11141) );
  AND2_X1 U13729 ( .A1(n11141), .A2(n11139), .ZN(n11144) );
  NAND2_X1 U13730 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  OAI211_X1 U13731 ( .C1(n11144), .C2(n11143), .A(n11142), .B(n12724), .ZN(
        n11148) );
  NAND2_X1 U13732 ( .A1(n12726), .A2(n12744), .ZN(n11145) );
  NAND2_X1 U13733 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12785)
         );
  OAI211_X1 U13734 ( .C1(n13076), .C2(n12729), .A(n11145), .B(n12785), .ZN(
        n11146) );
  AOI21_X1 U13735 ( .B1(n13079), .B2(n12731), .A(n11146), .ZN(n11147) );
  OAI211_X1 U13736 ( .C1(n13204), .C2(n12734), .A(n11148), .B(n11147), .ZN(
        P3_U3181) );
  OAI222_X1 U13737 ( .A1(n14436), .A2(n11149), .B1(n14428), .B2(n11380), .C1(
        n11192), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U13738 ( .A1(n13820), .A2(n11150), .B1(P2_U3088), .B2(n8881), .C1(
        n13818), .C2(n11380), .ZN(P2_U3306) );
  INV_X1 U13739 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11885) );
  INV_X1 U13740 ( .A(n11151), .ZN(n11152) );
  MUX2_X1 U13741 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6575), .Z(n11155) );
  XNOR2_X1 U13742 ( .A(n11155), .B(SI_25_), .ZN(n11461) );
  MUX2_X1 U13743 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n11550), .Z(n11478) );
  NAND2_X1 U13744 ( .A1(n11478), .A2(SI_26_), .ZN(n11156) );
  INV_X1 U13745 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13812) );
  MUX2_X1 U13746 ( .A(n14429), .B(n13812), .S(n6576), .Z(n11498) );
  NOR2_X1 U13747 ( .A1(n11498), .A2(n12499), .ZN(n11158) );
  NAND2_X1 U13748 ( .A1(n11498), .A2(n12499), .ZN(n11157) );
  INV_X1 U13749 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12306) );
  MUX2_X1 U13750 ( .A(n12135), .B(n12306), .S(n6575), .Z(n11159) );
  XNOR2_X1 U13751 ( .A(n11159), .B(SI_28_), .ZN(n11517) );
  NAND2_X1 U13752 ( .A1(n11518), .A2(n11517), .ZN(n11161) );
  NAND2_X1 U13753 ( .A1(n11159), .A2(n11164), .ZN(n11160) );
  INV_X1 U13754 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13804) );
  MUX2_X1 U13755 ( .A(n11885), .B(n13804), .S(n6576), .Z(n11168) );
  XNOR2_X1 U13756 ( .A(n11168), .B(SI_29_), .ZN(n11166) );
  INV_X1 U13757 ( .A(n12291), .ZN(n13806) );
  OAI222_X1 U13758 ( .A1(n14436), .A2(n11885), .B1(P1_U3086), .B2(n11162), 
        .C1(n14428), .C2(n13806), .ZN(P1_U3326) );
  INV_X1 U13759 ( .A(n11163), .ZN(n11165) );
  OAI222_X1 U13760 ( .A1(n13227), .A2(n11165), .B1(n12528), .B2(P3_U3151), 
        .C1(n11164), .C2(n13228), .ZN(P3_U3267) );
  INV_X1 U13761 ( .A(SI_29_), .ZN(n15505) );
  NAND2_X1 U13762 ( .A1(n11168), .A2(n15505), .ZN(n11553) );
  NAND2_X1 U13763 ( .A1(n11557), .A2(n11553), .ZN(n11171) );
  INV_X1 U13764 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12133) );
  INV_X1 U13765 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n15406) );
  MUX2_X1 U13766 ( .A(n12133), .B(n15406), .S(n6576), .Z(n11169) );
  INV_X1 U13767 ( .A(SI_30_), .ZN(n12522) );
  NOR2_X1 U13768 ( .A1(n11169), .A2(n12522), .ZN(n11552) );
  INV_X1 U13769 ( .A(n11552), .ZN(n11558) );
  NAND2_X1 U13770 ( .A1(n11169), .A2(n12522), .ZN(n11554) );
  AND2_X1 U13771 ( .A1(n11558), .A2(n11554), .ZN(n11170) );
  INV_X1 U13772 ( .A(n12347), .ZN(n12131) );
  OAI222_X1 U13773 ( .A1(n13818), .A2(n12131), .B1(P2_U3088), .B2(n11172), 
        .C1(n15406), .C2(n13820), .ZN(P2_U3297) );
  INV_X1 U13774 ( .A(n11342), .ZN(n11175) );
  INV_X1 U13775 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11369) );
  INV_X1 U13776 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13862) );
  INV_X1 U13777 ( .A(n11420), .ZN(n11177) );
  INV_X1 U13778 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13911) );
  INV_X1 U13779 ( .A(n11453), .ZN(n11178) );
  INV_X1 U13780 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11469) );
  INV_X1 U13781 ( .A(n11489), .ZN(n11179) );
  NAND2_X1 U13782 ( .A1(n11179), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n14110) );
  NAND2_X1 U13783 ( .A1(n11510), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11180) );
  OR2_X1 U13784 ( .A1(n14110), .A2(n11180), .ZN(n11187) );
  INV_X1 U13785 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U13786 ( .A1(n11387), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U13787 ( .A1(n11538), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11182) );
  OAI211_X1 U13788 ( .C1(n11184), .C2(n11540), .A(n11183), .B(n11182), .ZN(
        n11185) );
  INV_X1 U13789 ( .A(n11185), .ZN(n11186) );
  NAND2_X1 U13790 ( .A1(n11187), .A2(n11186), .ZN(n13970) );
  NAND2_X1 U13791 ( .A1(n12291), .A2(n11565), .ZN(n11189) );
  OR2_X1 U13792 ( .A1(n11567), .A2(n11885), .ZN(n11188) );
  NAND2_X1 U13793 ( .A1(n11193), .A2(n11192), .ZN(n11545) );
  MUX2_X1 U13794 ( .A(n13970), .B(n14113), .S(n6799), .Z(n11528) );
  INV_X1 U13795 ( .A(n11528), .ZN(n11531) );
  OAI21_X1 U13796 ( .B1(n11196), .B2(n11195), .A(n13987), .ZN(n11197) );
  OAI21_X1 U13797 ( .B1(n14831), .B2(n6785), .A(n11197), .ZN(n11198) );
  NAND2_X1 U13798 ( .A1(n11198), .A2(n11431), .ZN(n11199) );
  NAND2_X1 U13799 ( .A1(n11201), .A2(n9727), .ZN(n11207) );
  NAND2_X1 U13800 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  NAND2_X1 U13801 ( .A1(n11351), .A2(n11211), .ZN(n11208) );
  NAND2_X1 U13802 ( .A1(n11209), .A2(n11208), .ZN(n11212) );
  MUX2_X1 U13803 ( .A(n14847), .B(n11209), .S(n6799), .Z(n11210) );
  INV_X1 U13804 ( .A(n11213), .ZN(n11216) );
  INV_X1 U13805 ( .A(n11214), .ZN(n11215) );
  MUX2_X1 U13806 ( .A(n11216), .B(n11215), .S(n11351), .Z(n11217) );
  INV_X1 U13807 ( .A(n11217), .ZN(n11218) );
  MUX2_X1 U13808 ( .A(n14860), .B(n13984), .S(n11351), .Z(n11222) );
  NAND2_X1 U13809 ( .A1(n11221), .A2(n11222), .ZN(n11220) );
  MUX2_X1 U13810 ( .A(n13984), .B(n14860), .S(n11351), .Z(n11219) );
  NAND2_X1 U13811 ( .A1(n11220), .A2(n11219), .ZN(n11226) );
  INV_X1 U13812 ( .A(n11221), .ZN(n11224) );
  INV_X1 U13813 ( .A(n11222), .ZN(n11223) );
  NAND2_X1 U13814 ( .A1(n11224), .A2(n11223), .ZN(n11225) );
  MUX2_X1 U13815 ( .A(n13983), .B(n11227), .S(n11351), .Z(n11230) );
  MUX2_X1 U13816 ( .A(n11227), .B(n13983), .S(n11351), .Z(n11228) );
  MUX2_X1 U13817 ( .A(n14748), .B(n14875), .S(n11351), .Z(n11231) );
  NAND2_X1 U13818 ( .A1(n11232), .A2(n11231), .ZN(n11237) );
  NAND2_X1 U13819 ( .A1(n11235), .A2(n11234), .ZN(n11236) );
  MUX2_X1 U13820 ( .A(n13982), .B(n11238), .S(n6799), .Z(n11240) );
  MUX2_X1 U13821 ( .A(n11238), .B(n13982), .S(n11351), .Z(n11239) );
  INV_X1 U13822 ( .A(n11240), .ZN(n11241) );
  MUX2_X1 U13823 ( .A(n14749), .B(n14891), .S(n11504), .Z(n11245) );
  MUX2_X1 U13824 ( .A(n14749), .B(n14891), .S(n11351), .Z(n11242) );
  NAND2_X1 U13825 ( .A1(n11243), .A2(n11242), .ZN(n11249) );
  INV_X1 U13826 ( .A(n11244), .ZN(n11247) );
  INV_X1 U13827 ( .A(n11245), .ZN(n11246) );
  NAND2_X1 U13828 ( .A1(n11247), .A2(n11246), .ZN(n11248) );
  MUX2_X1 U13829 ( .A(n13981), .B(n11250), .S(n6799), .Z(n11254) );
  NAND2_X1 U13830 ( .A1(n11253), .A2(n11254), .ZN(n11252) );
  MUX2_X1 U13831 ( .A(n13981), .B(n11250), .S(n11504), .Z(n11251) );
  INV_X1 U13832 ( .A(n11253), .ZN(n11256) );
  INV_X1 U13833 ( .A(n11254), .ZN(n11255) );
  NAND2_X1 U13834 ( .A1(n11256), .A2(n11255), .ZN(n11263) );
  NAND2_X1 U13835 ( .A1(n11265), .A2(n11263), .ZN(n11257) );
  NAND2_X1 U13836 ( .A1(n11257), .A2(n11261), .ZN(n11260) );
  MUX2_X1 U13837 ( .A(n13980), .B(n11258), .S(n11351), .Z(n11259) );
  NAND2_X1 U13838 ( .A1(n11260), .A2(n11259), .ZN(n11267) );
  INV_X1 U13839 ( .A(n11261), .ZN(n11262) );
  AND2_X1 U13840 ( .A1(n11263), .A2(n11262), .ZN(n11264) );
  NAND2_X1 U13841 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  MUX2_X1 U13842 ( .A(n13979), .B(n14667), .S(n11351), .Z(n11269) );
  MUX2_X1 U13843 ( .A(n13979), .B(n14667), .S(n11504), .Z(n11268) );
  INV_X1 U13844 ( .A(n11269), .ZN(n11270) );
  MUX2_X1 U13845 ( .A(n13978), .B(n13877), .S(n11504), .Z(n11274) );
  MUX2_X1 U13846 ( .A(n13978), .B(n13877), .S(n6799), .Z(n11271) );
  INV_X1 U13847 ( .A(n11273), .ZN(n11276) );
  INV_X1 U13848 ( .A(n11274), .ZN(n11275) );
  NAND2_X1 U13849 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  MUX2_X1 U13850 ( .A(n13977), .B(n14660), .S(n6799), .Z(n11279) );
  MUX2_X1 U13851 ( .A(n13977), .B(n14660), .S(n11504), .Z(n11278) );
  NAND2_X1 U13852 ( .A1(n11280), .A2(n11565), .ZN(n11283) );
  AOI22_X1 U13853 ( .A1(n11281), .A2(n11338), .B1(n11519), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11282) );
  XNOR2_X1 U13854 ( .A(n11297), .B(n14278), .ZN(n14305) );
  NAND2_X1 U13855 ( .A1(n11285), .A2(n11565), .ZN(n11288) );
  AOI22_X1 U13856 ( .A1(n11519), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11338), 
        .B2(n11286), .ZN(n11287) );
  NAND2_X1 U13857 ( .A1(n11387), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11296) );
  INV_X1 U13858 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11289) );
  OR2_X1 U13859 ( .A1(n6573), .A2(n11289), .ZN(n11295) );
  NAND2_X1 U13860 ( .A1(n11290), .A2(n15522), .ZN(n11291) );
  NAND2_X1 U13861 ( .A1(n11324), .A2(n11291), .ZN(n14283) );
  OR2_X1 U13862 ( .A1(n11390), .A2(n14283), .ZN(n11294) );
  INV_X1 U13863 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11292) );
  OR2_X1 U13864 ( .A1(n11540), .A2(n11292), .ZN(n11293) );
  NAND4_X1 U13865 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n13976) );
  INV_X1 U13866 ( .A(n13976), .ZN(n11299) );
  INV_X1 U13867 ( .A(n14278), .ZN(n13961) );
  NAND2_X1 U13868 ( .A1(n11297), .A2(n13961), .ZN(n11298) );
  OR2_X1 U13869 ( .A1(n11297), .A2(n13961), .ZN(n11804) );
  MUX2_X1 U13870 ( .A(n11805), .B(n11806), .S(n6799), .Z(n11301) );
  NAND2_X1 U13871 ( .A1(n11302), .A2(n11565), .ZN(n11304) );
  AOI22_X1 U13872 ( .A1(n11519), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11338), 
        .B2(n14735), .ZN(n11303) );
  INV_X1 U13873 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U13874 ( .A1(n11318), .A2(n11305), .ZN(n11306) );
  NAND2_X1 U13875 ( .A1(n11342), .A2(n11306), .ZN(n13938) );
  OR2_X1 U13876 ( .A1(n13938), .A2(n11390), .ZN(n11311) );
  INV_X1 U13877 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14243) );
  OR2_X1 U13878 ( .A1(n6573), .A2(n14243), .ZN(n11310) );
  NAND2_X1 U13879 ( .A1(n11387), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11309) );
  INV_X1 U13880 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11307) );
  OR2_X1 U13881 ( .A1(n11540), .A2(n11307), .ZN(n11308) );
  NAND4_X1 U13882 ( .A1(n11311), .A2(n11310), .A3(n11309), .A4(n11308), .ZN(
        n13975) );
  XNOR2_X1 U13883 ( .A(n11350), .B(n13975), .ZN(n14245) );
  NAND2_X1 U13884 ( .A1(n11312), .A2(n11565), .ZN(n11314) );
  AOI22_X1 U13885 ( .A1(n11519), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11338), 
        .B2(n11663), .ZN(n11313) );
  NAND2_X1 U13886 ( .A1(n11387), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11322) );
  INV_X1 U13887 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11315) );
  OR2_X1 U13888 ( .A1(n6573), .A2(n11315), .ZN(n11321) );
  INV_X1 U13889 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11658) );
  OR2_X1 U13890 ( .A1(n11540), .A2(n11658), .ZN(n11320) );
  NAND2_X1 U13891 ( .A1(n11326), .A2(n11316), .ZN(n11317) );
  NAND2_X1 U13892 ( .A1(n11318), .A2(n11317), .ZN(n14254) );
  OR2_X1 U13893 ( .A1(n11491), .A2(n14254), .ZN(n11319) );
  NAND4_X1 U13894 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n14236) );
  XNOR2_X1 U13895 ( .A(n14397), .B(n14236), .ZN(n14257) );
  AND2_X1 U13896 ( .A1(n14245), .A2(n14257), .ZN(n11336) );
  NAND2_X1 U13897 ( .A1(n11387), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11330) );
  OR2_X1 U13898 ( .A1(n6573), .A2(n14269), .ZN(n11329) );
  INV_X1 U13899 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U13900 ( .A1(n11324), .A2(n11323), .ZN(n11325) );
  NAND2_X1 U13901 ( .A1(n11326), .A2(n11325), .ZN(n14268) );
  OR2_X1 U13902 ( .A1(n11390), .A2(n14268), .ZN(n11328) );
  OR2_X1 U13903 ( .A1(n11540), .A2(n14652), .ZN(n11327) );
  NAND4_X1 U13904 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n14279) );
  AOI22_X1 U13905 ( .A1(n11519), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11338), 
        .B2(n11332), .ZN(n11333) );
  MUX2_X1 U13906 ( .A(n6871), .B(n14647), .S(n11351), .Z(n11334) );
  MUX2_X1 U13907 ( .A(n14279), .B(n14271), .S(n11504), .Z(n11335) );
  NAND3_X1 U13908 ( .A1(n11336), .A2(n11335), .A3(n11334), .ZN(n11364) );
  NAND2_X1 U13909 ( .A1(n11337), .A2(n11565), .ZN(n11340) );
  AOI22_X1 U13910 ( .A1(n11519), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11338), 
        .B2(n11573), .ZN(n11339) );
  INV_X1 U13911 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11349) );
  INV_X1 U13912 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U13913 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  NAND2_X1 U13914 ( .A1(n11370), .A2(n11343), .ZN(n14221) );
  OR2_X1 U13915 ( .A1(n14221), .A2(n11390), .ZN(n11348) );
  INV_X1 U13916 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15377) );
  OR2_X1 U13917 ( .A1(n11541), .A2(n15377), .ZN(n11346) );
  INV_X1 U13918 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n11344) );
  OR2_X1 U13919 ( .A1(n6573), .A2(n11344), .ZN(n11345) );
  AND2_X1 U13920 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  OAI211_X1 U13921 ( .C1(n11540), .C2(n11349), .A(n11348), .B(n11347), .ZN(
        n14237) );
  INV_X1 U13922 ( .A(n14237), .ZN(n13942) );
  OR2_X1 U13923 ( .A1(n14388), .A2(n13942), .ZN(n11366) );
  NAND2_X1 U13924 ( .A1(n14388), .A2(n13942), .ZN(n11809) );
  NAND2_X1 U13925 ( .A1(n11366), .A2(n11809), .ZN(n11831) );
  INV_X1 U13926 ( .A(n14236), .ZN(n11807) );
  OR3_X1 U13927 ( .A1(n14397), .A2(n11504), .A3(n11807), .ZN(n11352) );
  NAND2_X1 U13928 ( .A1(n13975), .A2(n11351), .ZN(n11355) );
  AND2_X1 U13929 ( .A1(n11352), .A2(n11355), .ZN(n11361) );
  NAND3_X1 U13930 ( .A1(n14397), .A2(n11504), .A3(n11807), .ZN(n11353) );
  INV_X1 U13931 ( .A(n13975), .ZN(n13903) );
  NAND2_X1 U13932 ( .A1(n13903), .A2(n11504), .ZN(n11356) );
  NAND2_X1 U13933 ( .A1(n11353), .A2(n11356), .ZN(n11354) );
  NAND2_X1 U13934 ( .A1(n11350), .A2(n11354), .ZN(n11360) );
  NOR2_X1 U13935 ( .A1(n11355), .A2(n11807), .ZN(n11358) );
  OAI21_X1 U13936 ( .B1(n14236), .B2(n11356), .A(n14397), .ZN(n11357) );
  OAI21_X1 U13937 ( .B1(n11358), .B2(n14397), .A(n11357), .ZN(n11359) );
  OAI211_X1 U13938 ( .C1(n11350), .C2(n11361), .A(n11360), .B(n11359), .ZN(
        n11362) );
  NOR2_X1 U13939 ( .A1(n11831), .A2(n11362), .ZN(n11363) );
  MUX2_X1 U13940 ( .A(n11809), .B(n11366), .S(n11504), .Z(n11367) );
  INV_X1 U13941 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11374) );
  NAND2_X1 U13942 ( .A1(n11370), .A2(n11369), .ZN(n11371) );
  NAND2_X1 U13943 ( .A1(n11385), .A2(n11371), .ZN(n13918) );
  OR2_X1 U13944 ( .A1(n13918), .A2(n11491), .ZN(n11373) );
  AOI22_X1 U13945 ( .A1(n11387), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n11538), 
        .B2(P1_REG2_REG_20__SCAN_IN), .ZN(n11372) );
  OAI211_X1 U13946 ( .C1(n11540), .C2(n11374), .A(n11373), .B(n11372), .ZN(
        n13974) );
  NAND2_X1 U13947 ( .A1(n11375), .A2(n11565), .ZN(n11377) );
  NAND2_X1 U13948 ( .A1(n11519), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11376) );
  NOR2_X1 U13949 ( .A1(n14381), .A2(n13974), .ZN(n11378) );
  OR2_X1 U13950 ( .A1(n11379), .A2(n11378), .ZN(n11398) );
  NAND2_X1 U13951 ( .A1(n11401), .A2(n11398), .ZN(n11393) );
  NAND2_X1 U13952 ( .A1(n14381), .A2(n13974), .ZN(n11854) );
  NAND2_X1 U13953 ( .A1(n11379), .A2(n11854), .ZN(n11394) );
  INV_X1 U13954 ( .A(n11380), .ZN(n11382) );
  NAND2_X1 U13955 ( .A1(n11519), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U13956 ( .A1(n11385), .A2(n13862), .ZN(n11386) );
  NAND2_X1 U13957 ( .A1(n11404), .A2(n11386), .ZN(n14211) );
  AOI22_X1 U13958 ( .A1(n11387), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n11538), 
        .B2(P1_REG2_REG_21__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U13959 ( .A1(n11511), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11388) );
  OAI211_X1 U13960 ( .C1(n14211), .C2(n11390), .A(n11389), .B(n11388), .ZN(
        n13973) );
  MUX2_X1 U13961 ( .A(n14374), .B(n13973), .S(n11504), .Z(n11399) );
  INV_X1 U13962 ( .A(n11399), .ZN(n11391) );
  AND2_X1 U13963 ( .A1(n11394), .A2(n11391), .ZN(n11392) );
  NAND2_X1 U13964 ( .A1(n11393), .A2(n11392), .ZN(n11416) );
  MUX2_X1 U13965 ( .A(n14374), .B(n13973), .S(n11351), .Z(n11397) );
  INV_X1 U13966 ( .A(n11394), .ZN(n11395) );
  AND2_X1 U13967 ( .A1(n11397), .A2(n11396), .ZN(n11403) );
  AND2_X1 U13968 ( .A1(n11399), .A2(n11398), .ZN(n11400) );
  NAND2_X1 U13969 ( .A1(n11401), .A2(n11400), .ZN(n11402) );
  INV_X1 U13970 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U13971 ( .A1(n11404), .A2(n13929), .ZN(n11405) );
  NAND2_X1 U13972 ( .A1(n11420), .A2(n11405), .ZN(n14192) );
  OR2_X1 U13973 ( .A1(n14192), .A2(n11491), .ZN(n11410) );
  INV_X1 U13974 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15446) );
  NAND2_X1 U13975 ( .A1(n11387), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11407) );
  NAND2_X1 U13976 ( .A1(n11538), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11406) );
  OAI211_X1 U13977 ( .C1(n15446), .C2(n11540), .A(n11407), .B(n11406), .ZN(
        n11408) );
  INV_X1 U13978 ( .A(n11408), .ZN(n11409) );
  NAND2_X1 U13979 ( .A1(n11411), .A2(n7614), .ZN(n11412) );
  XNOR2_X1 U13980 ( .A(n11412), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14437) );
  INV_X1 U13981 ( .A(n14198), .ZN(n14370) );
  MUX2_X1 U13982 ( .A(n13861), .B(n14198), .S(n11351), .Z(n11414) );
  INV_X1 U13983 ( .A(n11414), .ZN(n11415) );
  INV_X1 U13984 ( .A(n11418), .ZN(n11419) );
  INV_X1 U13985 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15519) );
  NAND2_X1 U13986 ( .A1(n11420), .A2(n15519), .ZN(n11421) );
  NAND2_X1 U13987 ( .A1(n11435), .A2(n11421), .ZN(n14171) );
  OR2_X1 U13988 ( .A1(n14171), .A2(n11491), .ZN(n11427) );
  INV_X1 U13989 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U13990 ( .A1(n11387), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U13991 ( .A1(n11538), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11422) );
  OAI211_X1 U13992 ( .C1(n11424), .C2(n11540), .A(n11423), .B(n11422), .ZN(
        n11425) );
  INV_X1 U13993 ( .A(n11425), .ZN(n11426) );
  NAND2_X1 U13994 ( .A1(n11428), .A2(n11565), .ZN(n11430) );
  NAND2_X1 U13995 ( .A1(n11519), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11429) );
  NAND2_X2 U13996 ( .A1(n11430), .A2(n11429), .ZN(n14364) );
  MUX2_X1 U13997 ( .A(n14183), .B(n14364), .S(n6799), .Z(n11434) );
  NAND2_X1 U13998 ( .A1(n11435), .A2(n13911), .ZN(n11436) );
  AND2_X1 U13999 ( .A1(n11453), .A2(n11436), .ZN(n14156) );
  NAND2_X1 U14000 ( .A1(n14156), .A2(n11510), .ZN(n11442) );
  INV_X1 U14001 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11439) );
  NAND2_X1 U14002 ( .A1(n11387), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U14003 ( .A1(n11538), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11437) );
  OAI211_X1 U14004 ( .C1(n11439), .C2(n11540), .A(n11438), .B(n11437), .ZN(
        n11440) );
  INV_X1 U14005 ( .A(n11440), .ZN(n11441) );
  NAND2_X1 U14006 ( .A1(n11443), .A2(n11565), .ZN(n11445) );
  NAND2_X1 U14007 ( .A1(n11519), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11444) );
  NAND2_X2 U14008 ( .A1(n11445), .A2(n11444), .ZN(n14359) );
  MUX2_X1 U14009 ( .A(n14167), .B(n14359), .S(n6799), .Z(n11446) );
  NAND2_X1 U14010 ( .A1(n11447), .A2(n11446), .ZN(n11451) );
  INV_X1 U14011 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U14012 ( .A1(n11453), .A2(n11452), .ZN(n11454) );
  NAND2_X1 U14013 ( .A1(n11470), .A2(n11454), .ZN(n14141) );
  OR2_X1 U14014 ( .A1(n14141), .A2(n11491), .ZN(n11460) );
  INV_X1 U14015 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U14016 ( .A1(n11511), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U14017 ( .A1(n11387), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11455) );
  OAI211_X1 U14018 ( .C1(n6573), .C2(n11457), .A(n11456), .B(n11455), .ZN(
        n11458) );
  INV_X1 U14019 ( .A(n11458), .ZN(n11459) );
  XNOR2_X1 U14020 ( .A(n11462), .B(n11461), .ZN(n13816) );
  NAND2_X1 U14021 ( .A1(n13816), .A2(n11565), .ZN(n11464) );
  NAND2_X1 U14022 ( .A1(n11519), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11463) );
  MUX2_X1 U14023 ( .A(n13972), .B(n14137), .S(n11504), .Z(n11465) );
  INV_X1 U14024 ( .A(n11467), .ZN(n11468) );
  NAND2_X1 U14025 ( .A1(n11470), .A2(n11469), .ZN(n11471) );
  NAND2_X1 U14026 ( .A1(n14122), .A2(n11510), .ZN(n11477) );
  INV_X1 U14027 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11474) );
  NAND2_X1 U14028 ( .A1(n11538), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11473) );
  NAND2_X1 U14029 ( .A1(n11387), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11472) );
  OAI211_X1 U14030 ( .C1(n11540), .C2(n11474), .A(n11473), .B(n11472), .ZN(
        n11475) );
  INV_X1 U14031 ( .A(n11475), .ZN(n11476) );
  INV_X1 U14032 ( .A(n11478), .ZN(n11479) );
  XNOR2_X1 U14033 ( .A(n11479), .B(SI_26_), .ZN(n11480) );
  XNOR2_X1 U14034 ( .A(n11481), .B(n11480), .ZN(n13813) );
  NAND2_X1 U14035 ( .A1(n13813), .A2(n11565), .ZN(n11483) );
  NAND2_X1 U14036 ( .A1(n11519), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11482) );
  MUX2_X1 U14037 ( .A(n14140), .B(n14125), .S(n6799), .Z(n11484) );
  INV_X1 U14038 ( .A(n11486), .ZN(n11487) );
  INV_X1 U14039 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14040 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  NAND2_X1 U14041 ( .A1(n14110), .A2(n11490), .ZN(n13826) );
  INV_X1 U14042 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n12124) );
  NAND2_X1 U14043 ( .A1(n11387), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U14044 ( .A1(n11511), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11492) );
  OAI211_X1 U14045 ( .C1(n6573), .C2(n12124), .A(n11493), .B(n11492), .ZN(
        n11495) );
  INV_X1 U14046 ( .A(n11495), .ZN(n11496) );
  INV_X1 U14047 ( .A(n11498), .ZN(n11499) );
  XNOR2_X1 U14048 ( .A(n11499), .B(SI_27_), .ZN(n11500) );
  NAND2_X1 U14049 ( .A1(n13811), .A2(n11565), .ZN(n11503) );
  NAND2_X1 U14050 ( .A1(n11519), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11502) );
  MUX2_X1 U14051 ( .A(n13971), .B(n14337), .S(n11351), .Z(n11507) );
  NAND2_X1 U14052 ( .A1(n11506), .A2(n11505), .ZN(n11509) );
  XNOR2_X1 U14053 ( .A(n14110), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U14054 ( .A1(n11851), .A2(n11510), .ZN(n11516) );
  INV_X1 U14055 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15400) );
  NAND2_X1 U14056 ( .A1(n11511), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11513) );
  NAND2_X1 U14057 ( .A1(n11538), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11512) );
  OAI211_X1 U14058 ( .C1(n11541), .C2(n15400), .A(n11513), .B(n11512), .ZN(
        n11514) );
  INV_X1 U14059 ( .A(n11514), .ZN(n11515) );
  NAND2_X1 U14060 ( .A1(n12305), .A2(n11565), .ZN(n11521) );
  NAND2_X1 U14061 ( .A1(n11519), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11520) );
  MUX2_X1 U14062 ( .A(n14102), .B(n14330), .S(n6799), .Z(n11522) );
  INV_X1 U14063 ( .A(n11524), .ZN(n11525) );
  INV_X1 U14064 ( .A(n11529), .ZN(n11530) );
  INV_X1 U14065 ( .A(n14113), .ZN(n14322) );
  INV_X1 U14066 ( .A(n13970), .ZN(n11526) );
  MUX2_X1 U14067 ( .A(n14322), .B(n11526), .S(n6799), .Z(n11527) );
  NAND2_X1 U14068 ( .A1(n12347), .A2(n11565), .ZN(n11533) );
  OR2_X1 U14069 ( .A1(n11567), .A2(n12133), .ZN(n11532) );
  INV_X1 U14070 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14071 ( .A1(n11538), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11536) );
  INV_X1 U14072 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n11534) );
  OR2_X1 U14073 ( .A1(n11541), .A2(n11534), .ZN(n11535) );
  OAI211_X1 U14074 ( .C1(n11540), .C2(n11537), .A(n11536), .B(n11535), .ZN(
        n14104) );
  NAND2_X1 U14075 ( .A1(n11538), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11544) );
  INV_X1 U14076 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11539) );
  OR2_X1 U14077 ( .A1(n11540), .A2(n11539), .ZN(n11543) );
  INV_X1 U14078 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15322) );
  OR2_X1 U14079 ( .A1(n11541), .A2(n15322), .ZN(n11542) );
  OAI21_X1 U14080 ( .B1(n11504), .B2(n11577), .A(n11545), .ZN(n11546) );
  AOI22_X1 U14081 ( .A1(n14091), .A2(n11504), .B1(n14104), .B2(n11546), .ZN(
        n11548) );
  INV_X1 U14082 ( .A(n11577), .ZN(n14084) );
  OAI21_X1 U14083 ( .B1(n14084), .B2(n6790), .A(n14104), .ZN(n11547) );
  MUX2_X1 U14084 ( .A(n11547), .B(n14319), .S(n11351), .Z(n11549) );
  MUX2_X1 U14085 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11550), .Z(n11551) );
  XNOR2_X1 U14086 ( .A(n11551), .B(SI_31_), .ZN(n11559) );
  NAND2_X1 U14087 ( .A1(n11554), .A2(n11553), .ZN(n11560) );
  INV_X1 U14088 ( .A(n11559), .ZN(n11555) );
  NOR2_X1 U14089 ( .A1(n11560), .A2(n11555), .ZN(n11556) );
  NAND2_X1 U14090 ( .A1(n11557), .A2(n11556), .ZN(n11564) );
  XNOR2_X1 U14091 ( .A(n11559), .B(n11558), .ZN(n11562) );
  NOR2_X1 U14092 ( .A1(n11560), .A2(n11559), .ZN(n11561) );
  OR2_X1 U14093 ( .A1(n11562), .A2(n11561), .ZN(n11563) );
  NAND2_X1 U14094 ( .A1(n13799), .A2(n11565), .ZN(n11569) );
  INV_X1 U14095 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n11566) );
  OR2_X1 U14096 ( .A1(n11567), .A2(n11566), .ZN(n11568) );
  XNOR2_X1 U14097 ( .A(n14314), .B(n11577), .ZN(n11609) );
  OR2_X1 U14098 ( .A1(n10306), .A2(n11570), .ZN(n11571) );
  NAND2_X1 U14099 ( .A1(n11572), .A2(n11571), .ZN(n11575) );
  NAND2_X1 U14100 ( .A1(n6785), .A2(n11573), .ZN(n12127) );
  NAND2_X1 U14101 ( .A1(n11575), .A2(n12127), .ZN(n11617) );
  NOR3_X1 U14102 ( .A1(n11582), .A2(n11609), .A3(n11617), .ZN(n11623) );
  OR2_X1 U14103 ( .A1(n9247), .A2(n6790), .ZN(n11613) );
  NAND2_X1 U14104 ( .A1(n11617), .A2(n11613), .ZN(n11615) );
  INV_X1 U14105 ( .A(n11615), .ZN(n11581) );
  NOR2_X1 U14106 ( .A1(n14314), .A2(n11577), .ZN(n11579) );
  AND2_X1 U14107 ( .A1(n14314), .A2(n11577), .ZN(n11578) );
  MUX2_X1 U14108 ( .A(n11579), .B(n11578), .S(n11351), .Z(n11618) );
  INV_X1 U14109 ( .A(n11618), .ZN(n11580) );
  NOR2_X1 U14110 ( .A1(n14098), .A2(n14095), .ZN(n14094) );
  AOI21_X1 U14111 ( .B1(n14098), .B2(n14095), .A(n14094), .ZN(n11844) );
  XNOR2_X1 U14112 ( .A(n14125), .B(n12118), .ZN(n14118) );
  NAND2_X1 U14113 ( .A1(n14337), .A2(n11797), .ZN(n11843) );
  XNOR2_X1 U14114 ( .A(n14137), .B(n13972), .ZN(n14134) );
  OR2_X1 U14115 ( .A1(n14198), .A2(n14168), .ZN(n11840) );
  NAND2_X1 U14116 ( .A1(n14198), .A2(n14168), .ZN(n11583) );
  NAND2_X1 U14117 ( .A1(n11840), .A2(n11583), .ZN(n14186) );
  INV_X1 U14118 ( .A(n13974), .ZN(n13860) );
  XNOR2_X1 U14119 ( .A(n14381), .B(n13860), .ZN(n11832) );
  XNOR2_X1 U14120 ( .A(n14374), .B(n13973), .ZN(n14205) );
  INV_X1 U14121 ( .A(n14257), .ZN(n11808) );
  INV_X1 U14122 ( .A(n11584), .ZN(n11604) );
  INV_X1 U14123 ( .A(n11585), .ZN(n11603) );
  INV_X1 U14124 ( .A(n11586), .ZN(n14827) );
  NAND4_X1 U14125 ( .A1(n11588), .A2(n14827), .A3(n9727), .A4(n11587), .ZN(
        n11589) );
  NOR4_X1 U14126 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n14764), .ZN(
        n11594) );
  NAND4_X1 U14127 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  NOR3_X1 U14128 ( .A1(n11598), .A2(n11597), .A3(n11596), .ZN(n11601) );
  NAND4_X1 U14129 ( .A1(n7183), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11602) );
  NOR4_X1 U14130 ( .A1(n11808), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11605) );
  NAND4_X1 U14131 ( .A1(n14205), .A2(n14227), .A3(n11605), .A4(n14245), .ZN(
        n11606) );
  NOR3_X1 U14132 ( .A1(n14186), .A2(n11832), .A3(n11606), .ZN(n11607) );
  XNOR2_X1 U14133 ( .A(n14359), .B(n14167), .ZN(n11842) );
  XNOR2_X1 U14134 ( .A(n14364), .B(n14183), .ZN(n14175) );
  NAND4_X1 U14135 ( .A1(n14134), .A2(n11607), .A3(n11842), .A4(n14175), .ZN(
        n11608) );
  NOR4_X1 U14136 ( .A1(n11844), .A2(n14118), .A3(n12113), .A4(n11608), .ZN(
        n11611) );
  INV_X1 U14137 ( .A(n11609), .ZN(n11616) );
  XNOR2_X1 U14138 ( .A(n14091), .B(n14104), .ZN(n11610) );
  XNOR2_X1 U14139 ( .A(n14113), .B(n13970), .ZN(n14099) );
  NAND4_X1 U14140 ( .A1(n11611), .A2(n11616), .A3(n11610), .A4(n14099), .ZN(
        n11612) );
  XNOR2_X1 U14141 ( .A(n11612), .B(n11675), .ZN(n11614) );
  NOR2_X1 U14142 ( .A1(n11614), .A2(n11613), .ZN(n11622) );
  NOR2_X1 U14143 ( .A1(n11616), .A2(n11615), .ZN(n11620) );
  INV_X1 U14144 ( .A(n11617), .ZN(n11619) );
  MUX2_X1 U14145 ( .A(n11620), .B(n11619), .S(n11618), .Z(n11621) );
  NOR3_X1 U14146 ( .A1(n14191), .A2(n11624), .A3(n14426), .ZN(n11626) );
  OAI21_X1 U14147 ( .B1(n10306), .B2(n11627), .A(P1_B_REG_SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14148 ( .A1(n13816), .A2(n6581), .ZN(n11630) );
  INV_X1 U14149 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13819) );
  OR2_X1 U14150 ( .A1(n12348), .A2(n13819), .ZN(n11629) );
  XNOR2_X1 U14151 ( .A(n13727), .B(n8444), .ZN(n11634) );
  NAND2_X1 U14152 ( .A1(n13570), .A2(n8705), .ZN(n11633) );
  NOR2_X1 U14153 ( .A1(n11634), .A2(n11633), .ZN(n12500) );
  AOI21_X1 U14154 ( .B1(n11634), .B2(n11633), .A(n12500), .ZN(n11636) );
  OAI211_X1 U14155 ( .C1(n11635), .C2(n11636), .A(n12502), .B(n7445), .ZN(
        n11650) );
  NAND2_X1 U14156 ( .A1(n12319), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11646) );
  INV_X1 U14157 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n11637) );
  OR2_X1 U14158 ( .A1(n8765), .A2(n11637), .ZN(n11645) );
  INV_X1 U14159 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13302) );
  NAND2_X1 U14160 ( .A1(n11639), .A2(n13302), .ZN(n11640) );
  NAND2_X1 U14161 ( .A1(n12321), .A2(n11640), .ZN(n13563) );
  OR2_X1 U14162 ( .A1(n6583), .A2(n13563), .ZN(n11644) );
  INV_X1 U14163 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n11641) );
  OR2_X1 U14164 ( .A1(n6569), .A2(n11641), .ZN(n11643) );
  NAND4_X1 U14165 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n13586) );
  NOR2_X1 U14166 ( .A1(n14932), .A2(n13517), .ZN(n11648) );
  OAI22_X1 U14167 ( .A1(n13516), .A2(n14933), .B1(n13579), .B2(n14947), .ZN(
        n11647) );
  AOI211_X1 U14168 ( .C1(P2_REG3_REG_25__SCAN_IN), .C2(P2_U3088), .A(n11648), 
        .B(n11647), .ZN(n11649) );
  OAI211_X1 U14169 ( .C1(n7054), .C2(n13297), .A(n11650), .B(n11649), .ZN(
        P2_U3197) );
  OAI21_X1 U14170 ( .B1(n6705), .B2(n7036), .A(n11651), .ZN(n11652) );
  NAND2_X1 U14171 ( .A1(n11652), .A2(n12724), .ZN(n11656) );
  AOI22_X1 U14172 ( .A1(n12726), .A2(n13016), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11653) );
  OAI21_X1 U14173 ( .B1(n12986), .B2(n12729), .A(n11653), .ZN(n11654) );
  AOI21_X1 U14174 ( .B1(n12990), .B2(n12731), .A(n11654), .ZN(n11655) );
  OAI211_X1 U14175 ( .C1(n7037), .C2(n12734), .A(n11656), .B(n11655), .ZN(
        P3_U3175) );
  XNOR2_X1 U14176 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14080), .ZN(n14074) );
  OAI21_X1 U14177 ( .B1(n14652), .B2(n11666), .A(n11657), .ZN(n14073) );
  NAND2_X1 U14178 ( .A1(n14074), .A2(n14073), .ZN(n14072) );
  OAI21_X1 U14179 ( .B1(n11658), .B2(n14080), .A(n14072), .ZN(n11660) );
  XNOR2_X1 U14180 ( .A(n11659), .B(n11660), .ZN(n14739) );
  NAND2_X1 U14181 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14739), .ZN(n14737) );
  NAND2_X1 U14182 ( .A1(n14735), .A2(n11660), .ZN(n11661) );
  NAND2_X1 U14183 ( .A1(n14737), .A2(n11661), .ZN(n11662) );
  XOR2_X1 U14184 ( .A(n11662), .B(P1_REG1_REG_19__SCAN_IN), .Z(n11674) );
  INV_X1 U14185 ( .A(n11674), .ZN(n11672) );
  NAND2_X1 U14186 ( .A1(n11663), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11667) );
  INV_X1 U14187 ( .A(n11667), .ZN(n11664) );
  AOI21_X1 U14188 ( .B1(n11315), .B2(n14080), .A(n11664), .ZN(n14071) );
  OAI21_X1 U14189 ( .B1(n11666), .B2(n14269), .A(n11665), .ZN(n14070) );
  NAND2_X1 U14190 ( .A1(n14071), .A2(n14070), .ZN(n14069) );
  NAND2_X1 U14191 ( .A1(n11667), .A2(n14069), .ZN(n11668) );
  NAND2_X1 U14192 ( .A1(n14735), .A2(n11668), .ZN(n11669) );
  XOR2_X1 U14193 ( .A(n14735), .B(n11668), .Z(n14734) );
  NAND2_X1 U14194 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14734), .ZN(n14732) );
  NAND2_X1 U14195 ( .A1(n11669), .A2(n14732), .ZN(n11670) );
  XNOR2_X1 U14196 ( .A(n11344), .B(n11670), .ZN(n11673) );
  OAI21_X1 U14197 ( .B1(n11673), .B2(n14723), .A(n14725), .ZN(n11671) );
  AOI21_X1 U14198 ( .B1(n11672), .B2(n14738), .A(n11671), .ZN(n11677) );
  AOI22_X1 U14199 ( .A1(n11674), .A2(n14738), .B1(n14733), .B2(n11673), .ZN(
        n11676) );
  MUX2_X1 U14200 ( .A(n11677), .B(n11676), .S(n11675), .Z(n11678) );
  NAND2_X1 U14201 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13848)
         );
  OAI211_X1 U14202 ( .C1(n11679), .C2(n14729), .A(n11678), .B(n13848), .ZN(
        P1_U3262) );
  AND2_X1 U14203 ( .A1(n13974), .A2(n11757), .ZN(n11680) );
  AOI21_X1 U14204 ( .B1(n14381), .B2(n11786), .A(n11680), .ZN(n11736) );
  INV_X1 U14205 ( .A(n11736), .ZN(n11739) );
  AOI22_X1 U14206 ( .A1(n14381), .A2(n11787), .B1(n11786), .B2(n13974), .ZN(
        n11681) );
  XNOR2_X1 U14207 ( .A(n11681), .B(n11789), .ZN(n11737) );
  INV_X1 U14208 ( .A(n11737), .ZN(n11738) );
  AOI22_X1 U14209 ( .A1(n14388), .A2(n11788), .B1(n11757), .B2(n14237), .ZN(
        n11732) );
  INV_X1 U14210 ( .A(n11732), .ZN(n11735) );
  AOI22_X1 U14211 ( .A1(n14388), .A2(n11787), .B1(n11786), .B2(n14237), .ZN(
        n11682) );
  XNOR2_X1 U14212 ( .A(n11682), .B(n11789), .ZN(n11733) );
  INV_X1 U14213 ( .A(n11733), .ZN(n11734) );
  INV_X1 U14214 ( .A(n11685), .ZN(n11686) );
  NAND2_X1 U14215 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  NAND2_X1 U14216 ( .A1(n11297), .A2(n11787), .ZN(n11691) );
  NAND2_X1 U14217 ( .A1(n14278), .A2(n11786), .ZN(n11690) );
  NAND2_X1 U14218 ( .A1(n11691), .A2(n11690), .ZN(n11693) );
  XNOR2_X1 U14219 ( .A(n11693), .B(n11692), .ZN(n11695) );
  AND2_X1 U14220 ( .A1(n14278), .A2(n11757), .ZN(n11694) );
  AOI21_X1 U14221 ( .B1(n11297), .B2(n11786), .A(n11694), .ZN(n11696) );
  NAND2_X1 U14222 ( .A1(n11695), .A2(n11696), .ZN(n11701) );
  INV_X1 U14223 ( .A(n11695), .ZN(n11698) );
  INV_X1 U14224 ( .A(n11696), .ZN(n11697) );
  NAND2_X1 U14225 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  NAND2_X1 U14226 ( .A1(n11701), .A2(n11699), .ZN(n13833) );
  NAND2_X1 U14227 ( .A1(n14402), .A2(n11787), .ZN(n11703) );
  NAND2_X1 U14228 ( .A1(n13976), .A2(n11786), .ZN(n11702) );
  NAND2_X1 U14229 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  XNOR2_X1 U14230 ( .A(n11704), .B(n11789), .ZN(n11705) );
  OR2_X2 U14231 ( .A1(n11706), .A2(n11705), .ZN(n11708) );
  NAND2_X1 U14232 ( .A1(n11706), .A2(n11705), .ZN(n11707) );
  AOI22_X1 U14233 ( .A1(n14402), .A2(n11788), .B1(n11757), .B2(n13976), .ZN(
        n13958) );
  NAND2_X1 U14234 ( .A1(n14271), .A2(n11787), .ZN(n11710) );
  NAND2_X1 U14235 ( .A1(n14279), .A2(n11788), .ZN(n11709) );
  NAND2_X1 U14236 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  XNOR2_X1 U14237 ( .A(n11711), .B(n11789), .ZN(n11714) );
  AOI22_X1 U14238 ( .A1(n14271), .A2(n11788), .B1(n11757), .B2(n14279), .ZN(
        n11712) );
  XNOR2_X1 U14239 ( .A(n11714), .B(n11712), .ZN(n13888) );
  INV_X1 U14240 ( .A(n11712), .ZN(n11713) );
  NAND2_X1 U14241 ( .A1(n13886), .A2(n11715), .ZN(n13898) );
  NAND2_X1 U14242 ( .A1(n14397), .A2(n11787), .ZN(n11717) );
  NAND2_X1 U14243 ( .A1(n14236), .A2(n11786), .ZN(n11716) );
  NAND2_X1 U14244 ( .A1(n11717), .A2(n11716), .ZN(n11718) );
  XNOR2_X1 U14245 ( .A(n11718), .B(n11789), .ZN(n11721) );
  NAND2_X1 U14246 ( .A1(n14397), .A2(n11786), .ZN(n11720) );
  NAND2_X1 U14247 ( .A1(n14236), .A2(n11757), .ZN(n11719) );
  NAND2_X1 U14248 ( .A1(n11720), .A2(n11719), .ZN(n11722) );
  NAND2_X1 U14249 ( .A1(n11721), .A2(n11722), .ZN(n13899) );
  INV_X1 U14250 ( .A(n11721), .ZN(n11724) );
  INV_X1 U14251 ( .A(n11722), .ZN(n11723) );
  NAND2_X1 U14252 ( .A1(n11724), .A2(n11723), .ZN(n13901) );
  NAND2_X1 U14253 ( .A1(n11350), .A2(n11787), .ZN(n11726) );
  NAND2_X1 U14254 ( .A1(n13975), .A2(n11786), .ZN(n11725) );
  NAND2_X1 U14255 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  XNOR2_X1 U14256 ( .A(n11727), .B(n11789), .ZN(n11730) );
  AOI22_X1 U14257 ( .A1(n11350), .A2(n11788), .B1(n11757), .B2(n13975), .ZN(
        n11728) );
  XNOR2_X1 U14258 ( .A(n11730), .B(n11728), .ZN(n13936) );
  INV_X1 U14259 ( .A(n11728), .ZN(n11729) );
  XNOR2_X1 U14260 ( .A(n11733), .B(n11732), .ZN(n13852) );
  XNOR2_X1 U14261 ( .A(n11737), .B(n11736), .ZN(n13920) );
  AOI22_X1 U14262 ( .A1(n14374), .A2(n11788), .B1(n11757), .B2(n13973), .ZN(
        n11742) );
  AOI22_X1 U14263 ( .A1(n14374), .A2(n11787), .B1(n11786), .B2(n13973), .ZN(
        n11740) );
  XNOR2_X1 U14264 ( .A(n11740), .B(n11789), .ZN(n11741) );
  XOR2_X1 U14265 ( .A(n11742), .B(n11741), .Z(n13858) );
  NAND2_X1 U14266 ( .A1(n13857), .A2(n13858), .ZN(n13856) );
  NAND2_X1 U14267 ( .A1(n13856), .A2(n11743), .ZN(n13926) );
  INV_X1 U14268 ( .A(n11757), .ZN(n11744) );
  OAI22_X1 U14269 ( .A1(n14198), .A2(n11745), .B1(n13861), .B2(n11744), .ZN(
        n11748) );
  OAI22_X1 U14270 ( .A1(n14198), .A2(n11746), .B1(n13861), .B2(n11745), .ZN(
        n11747) );
  XNOR2_X1 U14271 ( .A(n11747), .B(n11789), .ZN(n11749) );
  XOR2_X1 U14272 ( .A(n11748), .B(n11749), .Z(n13927) );
  NAND2_X1 U14273 ( .A1(n14364), .A2(n11787), .ZN(n11752) );
  NAND2_X1 U14274 ( .A1(n14183), .A2(n11788), .ZN(n11751) );
  NAND2_X1 U14275 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  XNOR2_X1 U14276 ( .A(n11753), .B(n11789), .ZN(n11754) );
  AOI22_X1 U14277 ( .A1(n14364), .A2(n11788), .B1(n11757), .B2(n14183), .ZN(
        n11755) );
  XNOR2_X1 U14278 ( .A(n11754), .B(n11755), .ZN(n13842) );
  INV_X1 U14279 ( .A(n11754), .ZN(n11756) );
  AOI22_X1 U14280 ( .A1(n14359), .A2(n11788), .B1(n11757), .B2(n14167), .ZN(
        n11762) );
  NAND2_X1 U14281 ( .A1(n14359), .A2(n6572), .ZN(n11760) );
  NAND2_X1 U14282 ( .A1(n14167), .A2(n11788), .ZN(n11759) );
  NAND2_X1 U14283 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  XNOR2_X1 U14284 ( .A(n11761), .B(n11789), .ZN(n11764) );
  XOR2_X1 U14285 ( .A(n11762), .B(n11764), .Z(n13909) );
  INV_X1 U14286 ( .A(n11762), .ZN(n11763) );
  NAND2_X1 U14287 ( .A1(n14137), .A2(n11787), .ZN(n11766) );
  NAND2_X1 U14288 ( .A1(n13972), .A2(n11786), .ZN(n11765) );
  NAND2_X1 U14289 ( .A1(n11766), .A2(n11765), .ZN(n11767) );
  XNOR2_X1 U14290 ( .A(n11767), .B(n11789), .ZN(n11770) );
  AOI22_X1 U14291 ( .A1(n14137), .A2(n11788), .B1(n11757), .B2(n13972), .ZN(
        n11768) );
  XNOR2_X1 U14292 ( .A(n11770), .B(n11768), .ZN(n13880) );
  INV_X1 U14293 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U14294 ( .A1(n14125), .A2(n6572), .ZN(n11773) );
  NAND2_X1 U14295 ( .A1(n14140), .A2(n11788), .ZN(n11772) );
  NAND2_X1 U14296 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  XNOR2_X1 U14297 ( .A(n11774), .B(n11789), .ZN(n11775) );
  AOI22_X1 U14298 ( .A1(n14125), .A2(n11788), .B1(n11757), .B2(n14140), .ZN(
        n11776) );
  NAND2_X1 U14299 ( .A1(n13946), .A2(n13947), .ZN(n11779) );
  INV_X1 U14300 ( .A(n11775), .ZN(n11777) );
  NAND2_X1 U14301 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  NAND2_X1 U14302 ( .A1(n14337), .A2(n11787), .ZN(n11781) );
  NAND2_X1 U14303 ( .A1(n13971), .A2(n11786), .ZN(n11780) );
  NAND2_X1 U14304 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  XNOR2_X1 U14305 ( .A(n11782), .B(n11789), .ZN(n11783) );
  AOI22_X1 U14306 ( .A1(n14337), .A2(n11788), .B1(n11757), .B2(n13971), .ZN(
        n11784) );
  XNOR2_X1 U14307 ( .A(n11783), .B(n11784), .ZN(n13823) );
  INV_X1 U14308 ( .A(n11783), .ZN(n11785) );
  AOI22_X1 U14309 ( .A1(n14330), .A2(n11787), .B1(n11786), .B2(n14102), .ZN(
        n11792) );
  AOI22_X1 U14310 ( .A1(n14330), .A2(n11788), .B1(n11757), .B2(n14102), .ZN(
        n11790) );
  XNOR2_X1 U14311 ( .A(n11790), .B(n11789), .ZN(n11791) );
  XOR2_X1 U14312 ( .A(n11792), .B(n11791), .Z(n11793) );
  XNOR2_X1 U14313 ( .A(n11794), .B(n11793), .ZN(n11800) );
  AOI22_X1 U14314 ( .A1(n13970), .A2(n13966), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11796) );
  NAND2_X1 U14315 ( .A1(n11851), .A2(n13949), .ZN(n11795) );
  OAI211_X1 U14316 ( .C1(n11797), .C2(n13962), .A(n11796), .B(n11795), .ZN(
        n11798) );
  AOI21_X1 U14317 ( .B1(n14330), .B2(n6564), .A(n11798), .ZN(n11799) );
  OAI21_X1 U14318 ( .B1(n11800), .B2(n13955), .A(n11799), .ZN(P1_U3220) );
  INV_X1 U14319 ( .A(n13977), .ZN(n11801) );
  NAND2_X1 U14320 ( .A1(n11803), .A2(n11802), .ZN(n14297) );
  NAND2_X1 U14321 ( .A1(n14297), .A2(n14305), .ZN(n14296) );
  NAND2_X1 U14322 ( .A1(n14235), .A2(n14245), .ZN(n14234) );
  OR2_X1 U14323 ( .A1(n11350), .A2(n13903), .ZN(n14225) );
  NAND3_X1 U14324 ( .A1(n14234), .A2(n14227), .A3(n14225), .ZN(n14226) );
  NAND2_X1 U14325 ( .A1(n14226), .A2(n11809), .ZN(n11810) );
  NAND2_X1 U14326 ( .A1(n11810), .A2(n11832), .ZN(n14378) );
  NAND2_X1 U14327 ( .A1(n14378), .A2(n14136), .ZN(n11838) );
  INV_X1 U14328 ( .A(n11350), .ZN(n14244) );
  INV_X1 U14329 ( .A(n14214), .ZN(n11813) );
  AOI211_X1 U14330 ( .C1(n14381), .C2(n14220), .A(n14837), .B(n11813), .ZN(
        n14379) );
  INV_X1 U14331 ( .A(n13973), .ZN(n14190) );
  OAI22_X1 U14332 ( .A1(n14190), .A2(n14189), .B1(n13942), .B2(n14191), .ZN(
        n14380) );
  INV_X1 U14333 ( .A(n14380), .ZN(n11814) );
  OAI22_X1 U14334 ( .A1(n11814), .A2(n14286), .B1(n13918), .B2(n14783), .ZN(
        n11815) );
  AOI21_X1 U14335 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(n14286), .A(n11815), 
        .ZN(n11816) );
  OAI21_X1 U14336 ( .B1(n11811), .B2(n14786), .A(n11816), .ZN(n11817) );
  AOI21_X1 U14337 ( .B1(n14379), .B2(n14793), .A(n11817), .ZN(n11837) );
  NAND2_X1 U14338 ( .A1(n11819), .A2(n11818), .ZN(n11821) );
  OR2_X1 U14339 ( .A1(n14660), .A2(n13977), .ZN(n11820) );
  NAND2_X1 U14340 ( .A1(n11297), .A2(n14278), .ZN(n11822) );
  NAND2_X1 U14341 ( .A1(n6615), .A2(n11822), .ZN(n14290) );
  OR2_X1 U14342 ( .A1(n14402), .A2(n13976), .ZN(n11825) );
  OR2_X1 U14343 ( .A1(n14271), .A2(n14279), .ZN(n11826) );
  NOR2_X1 U14344 ( .A1(n14397), .A2(n14236), .ZN(n11827) );
  NAND2_X1 U14345 ( .A1(n14397), .A2(n14236), .ZN(n11828) );
  AND2_X1 U14346 ( .A1(n11350), .A2(n13975), .ZN(n11830) );
  OR2_X1 U14347 ( .A1(n11350), .A2(n13975), .ZN(n11829) );
  INV_X1 U14348 ( .A(n11834), .ZN(n11833) );
  INV_X1 U14349 ( .A(n11832), .ZN(n11835) );
  NAND2_X1 U14350 ( .A1(n11834), .A2(n11835), .ZN(n14382) );
  NAND3_X1 U14351 ( .A1(n14383), .A2(n14382), .A3(n14306), .ZN(n11836) );
  OAI211_X1 U14352 ( .C1(n11839), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        P1_U3273) );
  INV_X1 U14353 ( .A(n14359), .ZN(n14158) );
  NOR2_X1 U14354 ( .A1(n14381), .A2(n13860), .ZN(n14206) );
  OAI21_X2 U14355 ( .B1(n11839), .B2(n14206), .A(n14205), .ZN(n14209) );
  INV_X1 U14356 ( .A(n11840), .ZN(n11841) );
  INV_X1 U14357 ( .A(n14175), .ZN(n14166) );
  INV_X1 U14358 ( .A(n14364), .ZN(n14174) );
  INV_X1 U14359 ( .A(n14137), .ZN(n14353) );
  INV_X1 U14360 ( .A(n12113), .ZN(n12117) );
  NAND2_X1 U14361 ( .A1(n12116), .A2(n12117), .ZN(n12115) );
  INV_X1 U14362 ( .A(n11844), .ZN(n11860) );
  NAND2_X1 U14363 ( .A1(n13971), .A2(n14747), .ZN(n11845) );
  AOI21_X2 U14364 ( .B1(n11848), .B2(n14902), .A(n11847), .ZN(n14333) );
  NAND2_X1 U14365 ( .A1(n14198), .A2(n14213), .ZN(n14194) );
  INV_X1 U14366 ( .A(n14101), .ZN(n11850) );
  AOI21_X1 U14367 ( .B1(n14330), .B2(n12122), .A(n11850), .ZN(n14331) );
  AOI22_X1 U14368 ( .A1(n11851), .A2(n14284), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n14286), .ZN(n11852) );
  OAI21_X1 U14369 ( .B1(n14098), .B2(n14786), .A(n11852), .ZN(n11853) );
  AOI21_X1 U14370 ( .B1(n14331), .B2(n14145), .A(n11853), .ZN(n11864) );
  NAND2_X1 U14371 ( .A1(n7373), .A2(n14190), .ZN(n11856) );
  NAND2_X1 U14372 ( .A1(n14204), .A2(n11856), .ZN(n14182) );
  NAND2_X1 U14373 ( .A1(n14182), .A2(n14186), .ZN(n11858) );
  NAND2_X1 U14374 ( .A1(n14198), .A2(n13861), .ZN(n11857) );
  INV_X1 U14375 ( .A(n14118), .ZN(n14120) );
  INV_X1 U14376 ( .A(n14335), .ZN(n11862) );
  NAND2_X1 U14377 ( .A1(n11861), .A2(n11860), .ZN(n14329) );
  NAND3_X1 U14378 ( .A1(n11862), .A2(n14306), .A3(n14329), .ZN(n11863) );
  OAI211_X1 U14379 ( .C1(n14333), .C2(n14286), .A(n11864), .B(n11863), .ZN(
        P1_U3265) );
  OR2_X1 U14380 ( .A1(n12466), .A2(n11866), .ZN(n12016) );
  NAND2_X1 U14381 ( .A1(n12466), .A2(n11866), .ZN(n12024) );
  XNOR2_X1 U14382 ( .A(n13147), .B(n12743), .ZN(n13066) );
  NAND2_X1 U14383 ( .A1(n13067), .A2(n13066), .ZN(n13065) );
  NAND2_X1 U14384 ( .A1(n13147), .A2(n13076), .ZN(n12023) );
  OR2_X1 U14385 ( .A1(n12642), .A2(n13041), .ZN(n12036) );
  NAND2_X1 U14386 ( .A1(n12642), .A2(n13041), .ZN(n12033) );
  NAND2_X1 U14387 ( .A1(n13136), .A2(n13053), .ZN(n12034) );
  NAND2_X1 U14388 ( .A1(n12035), .A2(n12034), .ZN(n13048) );
  INV_X1 U14389 ( .A(n13048), .ZN(n11868) );
  XNOR2_X1 U14390 ( .A(n13193), .B(n6752), .ZN(n13031) );
  OR2_X1 U14391 ( .A1(n13193), .A2(n6752), .ZN(n12040) );
  NAND2_X1 U14392 ( .A1(n13032), .A2(n12040), .ZN(n13023) );
  INV_X1 U14393 ( .A(n13023), .ZN(n11869) );
  XNOR2_X1 U14394 ( .A(n13020), .B(n12740), .ZN(n12470) );
  OR2_X1 U14395 ( .A1(n13020), .A2(n13030), .ZN(n12047) );
  NAND2_X1 U14396 ( .A1(n12611), .A2(n12987), .ZN(n12050) );
  OR2_X1 U14397 ( .A1(n12611), .A2(n12987), .ZN(n12051) );
  NAND2_X1 U14398 ( .A1(n12483), .A2(n7036), .ZN(n12054) );
  OR2_X1 U14399 ( .A1(n12483), .A2(n7036), .ZN(n12055) );
  NAND2_X1 U14400 ( .A1(n11870), .A2(n12055), .ZN(n12965) );
  NAND2_X1 U14401 ( .A1(n13111), .A2(n12738), .ZN(n11872) );
  INV_X1 U14402 ( .A(n13111), .ZN(n12980) );
  NAND2_X1 U14403 ( .A1(n13107), .A2(n12972), .ZN(n12060) );
  OR2_X1 U14404 ( .A1(n13107), .A2(n12972), .ZN(n11871) );
  INV_X1 U14405 ( .A(n11872), .ZN(n12956) );
  NOR2_X1 U14406 ( .A1(n12955), .A2(n12956), .ZN(n12062) );
  XNOR2_X1 U14407 ( .A(n13103), .B(n12951), .ZN(n12942) );
  INV_X1 U14408 ( .A(n12942), .ZN(n12064) );
  NAND2_X1 U14409 ( .A1(n13103), .A2(n12951), .ZN(n11873) );
  NAND2_X1 U14410 ( .A1(n12931), .A2(n12910), .ZN(n12069) );
  INV_X1 U14411 ( .A(n12069), .ZN(n11874) );
  NAND2_X1 U14412 ( .A1(n12915), .A2(n12923), .ZN(n11876) );
  OR2_X1 U14413 ( .A1(n12915), .A2(n12923), .ZN(n11875) );
  INV_X1 U14414 ( .A(n11876), .ZN(n12080) );
  INV_X1 U14415 ( .A(n12077), .ZN(n11877) );
  INV_X1 U14416 ( .A(n11879), .ZN(n11880) );
  AOI22_X1 U14417 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13804), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n11885), .ZN(n11882) );
  INV_X1 U14418 ( .A(n11882), .ZN(n11883) );
  XNOR2_X1 U14419 ( .A(n11886), .B(n11883), .ZN(n13224) );
  NOR2_X1 U14420 ( .A1(n6590), .A2(n15505), .ZN(n11884) );
  AOI21_X1 U14421 ( .B1(n13224), .B2(n11897), .A(n11884), .ZN(n12534) );
  AND2_X1 U14422 ( .A1(n12534), .A2(n12736), .ZN(n12086) );
  INV_X1 U14423 ( .A(n12086), .ZN(n11911) );
  NAND2_X1 U14424 ( .A1(n13804), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11887) );
  AND2_X1 U14425 ( .A1(n15406), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11889) );
  OAI22_X1 U14426 ( .A1(n11896), .A2(n11889), .B1(P2_DATAO_REG_30__SCAN_IN), 
        .B2(n15406), .ZN(n11891) );
  INV_X1 U14427 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12286) );
  XNOR2_X1 U14428 ( .A(n12286), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n11890) );
  XNOR2_X1 U14429 ( .A(n11891), .B(n11890), .ZN(n13222) );
  NAND2_X1 U14430 ( .A1(n13222), .A2(n11897), .ZN(n11893) );
  INV_X1 U14431 ( .A(SI_31_), .ZN(n13218) );
  OR2_X1 U14432 ( .A1(n6590), .A2(n13218), .ZN(n11892) );
  NAND2_X1 U14433 ( .A1(n11893), .A2(n11892), .ZN(n11913) );
  OR2_X1 U14434 ( .A1(n11913), .A2(n12899), .ZN(n11908) );
  AOI22_X1 U14435 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(
        P2_DATAO_REG_30__SCAN_IN), .B1(n12133), .B2(n15406), .ZN(n11894) );
  INV_X1 U14436 ( .A(n11894), .ZN(n11895) );
  XNOR2_X1 U14437 ( .A(n11896), .B(n11895), .ZN(n12521) );
  NAND2_X1 U14438 ( .A1(n12521), .A2(n11897), .ZN(n11899) );
  OR2_X1 U14439 ( .A1(n6590), .A2(n12522), .ZN(n11898) );
  INV_X1 U14440 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14618) );
  NAND2_X1 U14441 ( .A1(n11900), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U14442 ( .A1(n6584), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n11902) );
  OAI211_X1 U14443 ( .C1(n7851), .C2(n14618), .A(n11903), .B(n11902), .ZN(
        n11904) );
  INV_X1 U14444 ( .A(n11904), .ZN(n11905) );
  NAND2_X1 U14445 ( .A1(n14617), .A2(n12530), .ZN(n11907) );
  NAND2_X1 U14446 ( .A1(n11908), .A2(n11907), .ZN(n12091) );
  INV_X1 U14447 ( .A(n14617), .ZN(n11912) );
  NOR2_X1 U14448 ( .A1(n12534), .A2(n12736), .ZN(n11916) );
  INV_X1 U14449 ( .A(n11916), .ZN(n12084) );
  OAI21_X1 U14450 ( .B1(n11912), .B2(n11909), .A(n12084), .ZN(n11910) );
  INV_X1 U14451 ( .A(n12530), .ZN(n12735) );
  AOI22_X1 U14452 ( .A1(n11913), .A2(n12899), .B1(n11912), .B2(n12735), .ZN(
        n11915) );
  NOR2_X1 U14453 ( .A1(n11915), .A2(n13167), .ZN(n12098) );
  INV_X1 U14454 ( .A(n12098), .ZN(n11914) );
  NAND2_X1 U14455 ( .A1(n11914), .A2(n7138), .ZN(n11935) );
  INV_X1 U14456 ( .A(n11915), .ZN(n12089) );
  INV_X1 U14457 ( .A(n12492), .ZN(n12079) );
  NOR2_X1 U14458 ( .A1(n11918), .A2(n11917), .ZN(n11920) );
  INV_X1 U14459 ( .A(n15181), .ZN(n15189) );
  NAND4_X1 U14460 ( .A1(n11920), .A2(n11919), .A3(n11945), .A4(n15189), .ZN(
        n11923) );
  NAND4_X1 U14461 ( .A1(n11921), .A2(n11985), .A3(n11979), .A4(n11966), .ZN(
        n11922) );
  NOR2_X1 U14462 ( .A1(n11923), .A2(n11922), .ZN(n11926) );
  NOR2_X1 U14463 ( .A1(n10919), .A2(n15151), .ZN(n11925) );
  AND2_X1 U14464 ( .A1(n14594), .A2(n14608), .ZN(n11924) );
  NAND4_X1 U14465 ( .A1(n12005), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11927) );
  NOR2_X1 U14466 ( .A1(n12010), .A2(n11927), .ZN(n11928) );
  NAND4_X1 U14467 ( .A1(n13054), .A2(n13077), .A3(n11928), .A4(n13066), .ZN(
        n11929) );
  NOR4_X1 U14468 ( .A1(n12474), .A2(n13048), .A3(n13031), .A4(n11929), .ZN(
        n11930) );
  XNOR2_X1 U14469 ( .A(n12611), .B(n13016), .ZN(n13001) );
  NAND4_X1 U14470 ( .A1(n12968), .A2(n11930), .A3(n12989), .A4(n13001), .ZN(
        n11931) );
  NOR4_X1 U14471 ( .A1(n12920), .A2(n12942), .A3(n12955), .A4(n11931), .ZN(
        n11932) );
  NAND4_X1 U14472 ( .A1(n12538), .A2(n12079), .A3(n12907), .A4(n11932), .ZN(
        n11933) );
  INV_X1 U14473 ( .A(n12101), .ZN(n11934) );
  OAI22_X1 U14474 ( .A1(n12099), .A2(n11935), .B1(n12100), .B2(n11934), .ZN(
        n11937) );
  INV_X1 U14475 ( .A(n12538), .ZN(n12083) );
  INV_X1 U14476 ( .A(n11938), .ZN(n11941) );
  NAND2_X1 U14477 ( .A1(n12006), .A2(n11939), .ZN(n11940) );
  AOI21_X1 U14478 ( .B1(n14608), .B2(n11941), .A(n11940), .ZN(n12000) );
  INV_X1 U14479 ( .A(n11942), .ZN(n11947) );
  NAND2_X1 U14480 ( .A1(n11947), .A2(n11943), .ZN(n11944) );
  NAND4_X1 U14481 ( .A1(n15182), .A2(n12087), .A3(n11949), .A4(n11944), .ZN(
        n11946) );
  NAND3_X1 U14482 ( .A1(n11946), .A2(n15166), .A3(n11945), .ZN(n11963) );
  NAND2_X1 U14483 ( .A1(n11950), .A2(n11947), .ZN(n11948) );
  NAND2_X1 U14484 ( .A1(n11949), .A2(n11948), .ZN(n11952) );
  INV_X1 U14485 ( .A(n11950), .ZN(n11951) );
  MUX2_X1 U14486 ( .A(n11952), .B(n11951), .S(n12087), .Z(n11962) );
  NAND2_X1 U14487 ( .A1(n11957), .A2(n11953), .ZN(n11954) );
  NAND2_X1 U14488 ( .A1(n11956), .A2(n11954), .ZN(n11960) );
  NAND2_X1 U14489 ( .A1(n11956), .A2(n11955), .ZN(n11958) );
  NAND2_X1 U14490 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  MUX2_X1 U14491 ( .A(n11960), .B(n11959), .S(n12087), .Z(n11961) );
  OAI21_X1 U14492 ( .B1(n11963), .B2(n11962), .A(n11961), .ZN(n11970) );
  MUX2_X1 U14493 ( .A(n11965), .B(n11964), .S(n12087), .Z(n11967) );
  NAND2_X1 U14494 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  AOI21_X1 U14495 ( .B1(n11970), .B2(n11969), .A(n11968), .ZN(n11973) );
  AOI21_X1 U14496 ( .B1(n11981), .B2(n11971), .A(n12087), .ZN(n11972) );
  OAI21_X1 U14497 ( .B1(n11973), .B2(n11972), .A(n11975), .ZN(n11978) );
  NAND2_X1 U14498 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  NAND2_X1 U14499 ( .A1(n11976), .A2(n12087), .ZN(n11977) );
  NAND2_X1 U14500 ( .A1(n11978), .A2(n11977), .ZN(n11980) );
  OAI211_X1 U14501 ( .C1(n12076), .C2(n11981), .A(n11980), .B(n11979), .ZN(
        n11986) );
  MUX2_X1 U14502 ( .A(n11983), .B(n11982), .S(n12087), .Z(n11984) );
  NAND3_X1 U14503 ( .A1(n11986), .A2(n11985), .A3(n11984), .ZN(n11991) );
  MUX2_X1 U14504 ( .A(n11988), .B(n11987), .S(n12076), .Z(n11989) );
  NAND3_X1 U14505 ( .A1(n11991), .A2(n11990), .A3(n11989), .ZN(n11994) );
  INV_X1 U14506 ( .A(n15151), .ZN(n15147) );
  MUX2_X1 U14507 ( .A(n15145), .B(n11992), .S(n12076), .Z(n11993) );
  NAND3_X1 U14508 ( .A1(n11994), .A2(n15147), .A3(n11993), .ZN(n11997) );
  NAND3_X1 U14509 ( .A1(n12746), .A2(n12076), .A3(n11995), .ZN(n11996) );
  NAND2_X1 U14510 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  NAND2_X1 U14511 ( .A1(n11998), .A2(n14608), .ZN(n11999) );
  OAI21_X1 U14512 ( .B1(n12076), .B2(n12000), .A(n11999), .ZN(n12004) );
  AOI21_X1 U14513 ( .B1(n12003), .B2(n12001), .A(n12087), .ZN(n12002) );
  AOI21_X1 U14514 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(n12013) );
  OAI21_X1 U14515 ( .B1(n12087), .B2(n12006), .A(n12005), .ZN(n12012) );
  MUX2_X1 U14516 ( .A(n12008), .B(n7111), .S(n12076), .Z(n12009) );
  NOR2_X1 U14517 ( .A1(n12010), .A2(n12009), .ZN(n12011) );
  OAI211_X1 U14518 ( .C1(n12013), .C2(n12012), .A(n13077), .B(n12011), .ZN(
        n12020) );
  INV_X1 U14519 ( .A(n12014), .ZN(n12015) );
  NAND2_X1 U14520 ( .A1(n13077), .A2(n12015), .ZN(n12017) );
  OAI211_X1 U14521 ( .C1(n13076), .C2(n13147), .A(n12017), .B(n12016), .ZN(
        n12018) );
  NAND2_X1 U14522 ( .A1(n12018), .A2(n12087), .ZN(n12019) );
  NAND2_X1 U14523 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  NAND2_X1 U14524 ( .A1(n12021), .A2(n12023), .ZN(n12028) );
  NAND2_X1 U14525 ( .A1(n13077), .A2(n7107), .ZN(n12025) );
  NAND3_X1 U14526 ( .A1(n12025), .A2(n12024), .A3(n12023), .ZN(n12026) );
  NAND2_X1 U14527 ( .A1(n12026), .A2(n12076), .ZN(n12027) );
  NAND2_X1 U14528 ( .A1(n12028), .A2(n12027), .ZN(n12032) );
  NAND3_X1 U14529 ( .A1(n13070), .A2(n12076), .A3(n12743), .ZN(n12031) );
  INV_X1 U14530 ( .A(n13054), .ZN(n12029) );
  OR2_X1 U14531 ( .A1(n13048), .A2(n12029), .ZN(n12030) );
  AOI21_X1 U14532 ( .B1(n12032), .B2(n12031), .A(n12030), .ZN(n12044) );
  OAI211_X1 U14533 ( .C1(n13048), .C2(n12033), .A(n12040), .B(n12034), .ZN(
        n12039) );
  INV_X1 U14534 ( .A(n12034), .ZN(n12037) );
  NAND2_X1 U14535 ( .A1(n13193), .A2(n6752), .ZN(n12041) );
  OAI211_X1 U14536 ( .C1(n12037), .C2(n12036), .A(n12041), .B(n12035), .ZN(
        n12038) );
  MUX2_X1 U14537 ( .A(n12039), .B(n12038), .S(n12076), .Z(n12043) );
  MUX2_X1 U14538 ( .A(n12041), .B(n12040), .S(n12076), .Z(n12042) );
  OAI21_X1 U14539 ( .B1(n12044), .B2(n12043), .A(n12042), .ZN(n12045) );
  NAND2_X1 U14540 ( .A1(n12045), .A2(n12470), .ZN(n12049) );
  NAND2_X1 U14541 ( .A1(n13020), .A2(n13030), .ZN(n12046) );
  MUX2_X1 U14542 ( .A(n12047), .B(n12046), .S(n12076), .Z(n12048) );
  NAND3_X1 U14543 ( .A1(n12049), .A2(n13001), .A3(n12048), .ZN(n12053) );
  MUX2_X1 U14544 ( .A(n12051), .B(n12050), .S(n12087), .Z(n12052) );
  NAND3_X1 U14545 ( .A1(n12053), .A2(n12989), .A3(n12052), .ZN(n12057) );
  MUX2_X1 U14546 ( .A(n12055), .B(n12054), .S(n12076), .Z(n12056) );
  NAND2_X1 U14547 ( .A1(n12057), .A2(n12056), .ZN(n12059) );
  NOR2_X1 U14548 ( .A1(n12738), .A2(n12087), .ZN(n12058) );
  AOI22_X1 U14549 ( .A1(n12059), .A2(n12968), .B1(n12058), .B2(n12980), .ZN(
        n12065) );
  XNOR2_X1 U14550 ( .A(n12060), .B(n12076), .ZN(n12061) );
  OAI211_X1 U14551 ( .C1(n12065), .C2(n12955), .A(n12064), .B(n12063), .ZN(
        n12068) );
  OR3_X1 U14552 ( .A1(n13103), .A2(n12951), .A3(n12087), .ZN(n12067) );
  NAND3_X1 U14553 ( .A1(n13103), .A2(n12951), .A3(n12087), .ZN(n12066) );
  MUX2_X1 U14554 ( .A(n12070), .B(n12069), .S(n12076), .Z(n12071) );
  NAND2_X1 U14555 ( .A1(n12072), .A2(n12071), .ZN(n12073) );
  NAND2_X1 U14556 ( .A1(n12073), .A2(n12907), .ZN(n12075) );
  OR3_X1 U14557 ( .A1(n12915), .A2(n12923), .A3(n12076), .ZN(n12074) );
  NAND2_X1 U14558 ( .A1(n12075), .A2(n12074), .ZN(n12081) );
  XNOR2_X1 U14559 ( .A(n12077), .B(n12076), .ZN(n12078) );
  AOI21_X1 U14560 ( .B1(n12079), .B2(n12081), .A(n12078), .ZN(n12082) );
  NAND2_X1 U14561 ( .A1(n12085), .A2(n12084), .ZN(n12088) );
  AOI21_X1 U14562 ( .B1(n12899), .B2(n12089), .A(n12098), .ZN(n12090) );
  INV_X1 U14563 ( .A(n12092), .ZN(n12093) );
  NOR3_X1 U14564 ( .A1(n12106), .A2(n12884), .A3(n12528), .ZN(n12109) );
  OAI21_X1 U14565 ( .B1(n12110), .B2(n12107), .A(P3_B_REG_SCAN_IN), .ZN(n12108) );
  OAI22_X1 U14566 ( .A1(n12111), .A2(n12110), .B1(n12109), .B2(n12108), .ZN(
        P3_U3296) );
  OAI21_X1 U14567 ( .B1(n12114), .B2(n12113), .A(n12112), .ZN(n12128) );
  INV_X1 U14568 ( .A(n12128), .ZN(n14339) );
  OAI21_X1 U14569 ( .B1(n12117), .B2(n12116), .A(n12115), .ZN(n12120) );
  OAI22_X1 U14570 ( .A1(n14095), .A2(n14189), .B1(n12118), .B2(n14191), .ZN(
        n12119) );
  AOI211_X1 U14571 ( .C1(n14337), .C2(n14121), .A(n14837), .B(n11849), .ZN(
        n14336) );
  INV_X1 U14572 ( .A(n14337), .ZN(n12123) );
  NOR2_X1 U14573 ( .A1(n12123), .A2(n14786), .ZN(n12126) );
  OAI22_X1 U14574 ( .A1(n13826), .A2(n14783), .B1(n12124), .B2(n14301), .ZN(
        n12125) );
  AOI211_X1 U14575 ( .C1(n14336), .C2(n14793), .A(n12126), .B(n12125), .ZN(
        n12130) );
  NOR2_X1 U14576 ( .A1(n14286), .A2(n12127), .ZN(n14794) );
  NAND2_X1 U14577 ( .A1(n12128), .A2(n14794), .ZN(n12129) );
  OAI211_X1 U14578 ( .C1(n14342), .C2(n14286), .A(n12130), .B(n12129), .ZN(
        P1_U3266) );
  OAI222_X1 U14579 ( .A1(n14436), .A2(n12133), .B1(P1_U3086), .B2(n12132), 
        .C1(n14434), .C2(n12131), .ZN(P1_U3325) );
  INV_X1 U14580 ( .A(n12305), .ZN(n13810) );
  OAI222_X1 U14581 ( .A1(n14436), .A2(n12135), .B1(n14434), .B2(n13810), .C1(
        n12134), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI22_X1 U14582 ( .A1(n12144), .A2(n15035), .B1(n9128), .B2(n12140), .ZN(
        n12136) );
  INV_X1 U14583 ( .A(n12136), .ZN(n12139) );
  NAND2_X1 U14584 ( .A1(n12139), .A2(n12138), .ZN(n12143) );
  INV_X1 U14585 ( .A(n12140), .ZN(n12141) );
  OAI21_X1 U14586 ( .B1(n12460), .B2(n13459), .A(n12141), .ZN(n12142) );
  NAND2_X1 U14587 ( .A1(n12143), .A2(n12142), .ZN(n12146) );
  INV_X1 U14588 ( .A(n12144), .ZN(n12145) );
  NAND2_X1 U14589 ( .A1(n12146), .A2(n6635), .ZN(n12152) );
  NAND2_X1 U14590 ( .A1(n12147), .A2(n12275), .ZN(n12150) );
  NAND2_X1 U14591 ( .A1(n12150), .A2(n12149), .ZN(n12153) );
  NAND2_X1 U14592 ( .A1(n12152), .A2(n12153), .ZN(n12151) );
  NAND2_X1 U14593 ( .A1(n12151), .A2(n7337), .ZN(n12157) );
  NAND2_X1 U14594 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  NAND2_X1 U14595 ( .A1(n12157), .A2(n12156), .ZN(n12163) );
  NAND2_X1 U14596 ( .A1(n13322), .A2(n12225), .ZN(n12159) );
  NAND2_X1 U14597 ( .A1(n15062), .A2(n12275), .ZN(n12158) );
  NAND2_X1 U14598 ( .A1(n12159), .A2(n12158), .ZN(n12164) );
  NAND2_X1 U14599 ( .A1(n12163), .A2(n12164), .ZN(n12162) );
  AOI22_X1 U14600 ( .A1(n13322), .A2(n12275), .B1(n12225), .B2(n15062), .ZN(
        n12160) );
  NAND2_X1 U14601 ( .A1(n12162), .A2(n12161), .ZN(n12168) );
  INV_X1 U14602 ( .A(n12163), .ZN(n12166) );
  INV_X1 U14603 ( .A(n12164), .ZN(n12165) );
  NAND2_X1 U14604 ( .A1(n12168), .A2(n12167), .ZN(n12173) );
  NAND2_X1 U14605 ( .A1(n13321), .A2(n12250), .ZN(n12170) );
  NAND2_X1 U14606 ( .A1(n15070), .A2(n12331), .ZN(n12169) );
  NAND2_X1 U14607 ( .A1(n12170), .A2(n12169), .ZN(n12172) );
  AOI22_X1 U14608 ( .A1(n13321), .A2(n12331), .B1(n15070), .B2(n12275), .ZN(
        n12171) );
  AOI21_X1 U14609 ( .B1(n12173), .B2(n12172), .A(n12171), .ZN(n12175) );
  NOR2_X1 U14610 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NAND2_X1 U14611 ( .A1(n13320), .A2(n12250), .ZN(n12177) );
  NAND2_X1 U14612 ( .A1(n15075), .A2(n12331), .ZN(n12176) );
  NAND2_X1 U14613 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  AOI22_X1 U14614 ( .A1(n13319), .A2(n12275), .B1(n12331), .B2(n12179), .ZN(
        n12183) );
  OAI22_X1 U14615 ( .A1(n12181), .A2(n12180), .B1(n15084), .B2(n12331), .ZN(
        n12182) );
  OAI21_X1 U14616 ( .B1(n12184), .B2(n12183), .A(n12182), .ZN(n12186) );
  NAND2_X1 U14617 ( .A1(n12184), .A2(n12183), .ZN(n12185) );
  OAI22_X1 U14618 ( .A1(n12188), .A2(n12331), .B1(n12187), .B2(n12275), .ZN(
        n12189) );
  OAI22_X1 U14619 ( .A1(n12188), .A2(n12275), .B1(n12187), .B2(n12331), .ZN(
        n12191) );
  INV_X1 U14620 ( .A(n12189), .ZN(n12190) );
  BUF_X1 U14621 ( .A(n12275), .Z(n12250) );
  OAI22_X1 U14622 ( .A1(n15098), .A2(n12250), .B1(n12192), .B2(n12331), .ZN(
        n12193) );
  OAI22_X1 U14623 ( .A1(n15098), .A2(n12331), .B1(n12192), .B2(n12250), .ZN(
        n12194) );
  OAI22_X1 U14624 ( .A1(n12196), .A2(n12331), .B1(n12195), .B2(n12250), .ZN(
        n12200) );
  INV_X1 U14625 ( .A(n12200), .ZN(n12198) );
  OAI22_X1 U14626 ( .A1(n12196), .A2(n12250), .B1(n12195), .B2(n12331), .ZN(
        n12197) );
  INV_X1 U14627 ( .A(n12199), .ZN(n12203) );
  AND2_X1 U14628 ( .A1(n12201), .A2(n12198), .ZN(n12202) );
  NOR2_X1 U14629 ( .A1(n12203), .A2(n12202), .ZN(n12207) );
  AOI22_X1 U14630 ( .A1(n15111), .A2(n12331), .B1(n13315), .B2(n12180), .ZN(
        n12206) );
  OAI22_X1 U14631 ( .A1(n7050), .A2(n12331), .B1(n12204), .B2(n12180), .ZN(
        n12205) );
  OAI21_X1 U14632 ( .B1(n12207), .B2(n12206), .A(n12205), .ZN(n12209) );
  NAND2_X1 U14633 ( .A1(n12207), .A2(n12206), .ZN(n12208) );
  AOI22_X1 U14634 ( .A1(n15119), .A2(n12275), .B1(n12331), .B2(n13314), .ZN(
        n12214) );
  INV_X1 U14635 ( .A(n12214), .ZN(n12210) );
  OAI22_X1 U14636 ( .A1(n12212), .A2(n12275), .B1(n12211), .B2(n12331), .ZN(
        n12213) );
  OAI22_X1 U14637 ( .A1(n12215), .A2(n12250), .B1(n14934), .B2(n12331), .ZN(
        n12217) );
  NAND2_X1 U14638 ( .A1(n12216), .A2(n12217), .ZN(n12221) );
  OAI22_X1 U14639 ( .A1(n12215), .A2(n12331), .B1(n14934), .B2(n12275), .ZN(
        n12220) );
  INV_X1 U14640 ( .A(n12216), .ZN(n12219) );
  INV_X1 U14641 ( .A(n12217), .ZN(n12218) );
  AOI22_X1 U14642 ( .A1(n14944), .A2(n12275), .B1(n12331), .B2(n13312), .ZN(
        n12224) );
  AOI22_X1 U14643 ( .A1(n14944), .A2(n12331), .B1(n13312), .B2(n12275), .ZN(
        n12222) );
  INV_X1 U14644 ( .A(n12222), .ZN(n12223) );
  OAI22_X1 U14645 ( .A1(n14634), .A2(n12250), .B1(n14931), .B2(n12331), .ZN(
        n12226) );
  NAND2_X1 U14646 ( .A1(n6680), .A2(n6866), .ZN(n12232) );
  AOI22_X1 U14647 ( .A1(n12227), .A2(n12275), .B1(n12331), .B2(n7408), .ZN(
        n12228) );
  NAND2_X1 U14648 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U14649 ( .A1(n12232), .A2(n12231), .ZN(n12238) );
  OAI22_X1 U14650 ( .A1(n12234), .A2(n12331), .B1(n12233), .B2(n12180), .ZN(
        n12237) );
  AOI22_X1 U14651 ( .A1(n12235), .A2(n12331), .B1(n13311), .B2(n12275), .ZN(
        n12236) );
  OAI22_X1 U14652 ( .A1(n6586), .A2(n12250), .B1(n12239), .B2(n12331), .ZN(
        n12244) );
  AOI22_X1 U14653 ( .A1(n13778), .A2(n12275), .B1(n12331), .B2(n13310), .ZN(
        n12240) );
  INV_X1 U14654 ( .A(n12240), .ZN(n12241) );
  NAND2_X1 U14655 ( .A1(n12242), .A2(n12241), .ZN(n12248) );
  INV_X1 U14656 ( .A(n12243), .ZN(n12246) );
  INV_X1 U14657 ( .A(n12244), .ZN(n12245) );
  NAND2_X1 U14658 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  OAI22_X1 U14659 ( .A1(n12251), .A2(n12331), .B1(n12249), .B2(n12250), .ZN(
        n12252) );
  OAI22_X1 U14660 ( .A1(n12251), .A2(n12250), .B1(n12249), .B2(n12331), .ZN(
        n12253) );
  AOI22_X1 U14661 ( .A1(n13768), .A2(n12331), .B1(n13308), .B2(n12180), .ZN(
        n12256) );
  OAI22_X1 U14662 ( .A1(n7045), .A2(n12331), .B1(n12254), .B2(n12275), .ZN(
        n12255) );
  NAND2_X1 U14663 ( .A1(n12257), .A2(n12256), .ZN(n12258) );
  OAI22_X1 U14664 ( .A1(n13478), .A2(n12331), .B1(n13477), .B2(n12180), .ZN(
        n12260) );
  AOI22_X1 U14665 ( .A1(n13763), .A2(n12331), .B1(n13505), .B2(n12275), .ZN(
        n12259) );
  AOI22_X1 U14666 ( .A1(n13757), .A2(n12331), .B1(n13668), .B2(n12275), .ZN(
        n12261) );
  INV_X1 U14667 ( .A(n13757), .ZN(n13506) );
  INV_X1 U14668 ( .A(n13668), .ZN(n13507) );
  OAI22_X1 U14669 ( .A1(n13506), .A2(n12331), .B1(n13507), .B2(n12250), .ZN(
        n12262) );
  AOI22_X1 U14670 ( .A1(n13752), .A2(n12275), .B1(n12331), .B2(n13509), .ZN(
        n12264) );
  OAI22_X1 U14671 ( .A1(n13510), .A2(n12250), .B1(n13513), .B2(n12331), .ZN(
        n12263) );
  NAND2_X1 U14672 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  OAI22_X1 U14673 ( .A1(n13655), .A2(n12250), .B1(n13480), .B2(n12331), .ZN(
        n12269) );
  OAI22_X1 U14674 ( .A1(n13655), .A2(n12331), .B1(n13480), .B2(n12250), .ZN(
        n12268) );
  OAI22_X1 U14675 ( .A1(n13741), .A2(n12331), .B1(n13250), .B2(n12250), .ZN(
        n12270) );
  OAI22_X1 U14676 ( .A1(n13741), .A2(n12250), .B1(n13250), .B2(n12331), .ZN(
        n12271) );
  OAI22_X1 U14677 ( .A1(n13624), .A2(n12275), .B1(n13596), .B2(n12331), .ZN(
        n12273) );
  OAI22_X1 U14678 ( .A1(n13624), .A2(n12331), .B1(n13596), .B2(n12250), .ZN(
        n12274) );
  AOI22_X1 U14679 ( .A1(n13732), .A2(n12275), .B1(n12331), .B2(n13585), .ZN(
        n12279) );
  INV_X1 U14680 ( .A(n12279), .ZN(n12277) );
  AOI22_X1 U14681 ( .A1(n13732), .A2(n12331), .B1(n13585), .B2(n12275), .ZN(
        n12276) );
  NAND2_X1 U14682 ( .A1(n13813), .A2(n6581), .ZN(n12282) );
  INV_X1 U14683 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13814) );
  OR2_X1 U14684 ( .A1(n12348), .A2(n13814), .ZN(n12281) );
  AND2_X1 U14685 ( .A1(n13586), .A2(n12180), .ZN(n12283) );
  AOI21_X1 U14686 ( .B1(n13722), .B2(n12331), .A(n12283), .ZN(n12344) );
  NAND2_X1 U14687 ( .A1(n13722), .A2(n12275), .ZN(n12285) );
  NAND2_X1 U14688 ( .A1(n13586), .A2(n12331), .ZN(n12284) );
  NAND2_X1 U14689 ( .A1(n12285), .A2(n12284), .ZN(n12343) );
  OR2_X1 U14690 ( .A1(n12348), .A2(n12286), .ZN(n12287) );
  INV_X1 U14691 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U14692 ( .A1(n8436), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U14693 ( .A1(n8449), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12288) );
  OAI211_X1 U14694 ( .C1(n12357), .C2(n12290), .A(n12289), .B(n12288), .ZN(
        n13307) );
  XNOR2_X1 U14695 ( .A(n12364), .B(n13307), .ZN(n12433) );
  NAND2_X1 U14696 ( .A1(n12291), .A2(n6581), .ZN(n12293) );
  OR2_X1 U14697 ( .A1(n12348), .A2(n13804), .ZN(n12292) );
  NAND2_X1 U14698 ( .A1(n12319), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12300) );
  INV_X1 U14699 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n12294) );
  OR2_X1 U14700 ( .A1(n8765), .A2(n12294), .ZN(n12299) );
  AND2_X1 U14701 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n12295) );
  NAND2_X1 U14702 ( .A1(n12296), .A2(n12295), .ZN(n13500) );
  OR2_X1 U14703 ( .A1(n6583), .A2(n13500), .ZN(n12298) );
  INV_X1 U14704 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13501) );
  OR2_X1 U14705 ( .A1(n6568), .A2(n13501), .ZN(n12297) );
  NAND4_X1 U14706 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n13528) );
  AND2_X1 U14707 ( .A1(n13528), .A2(n12180), .ZN(n12301) );
  AOI21_X1 U14708 ( .B1(n13706), .B2(n12331), .A(n12301), .ZN(n12363) );
  NAND2_X1 U14709 ( .A1(n13706), .A2(n12250), .ZN(n12303) );
  NAND2_X1 U14710 ( .A1(n13528), .A2(n12331), .ZN(n12302) );
  NAND2_X1 U14711 ( .A1(n12303), .A2(n12302), .ZN(n12362) );
  NAND2_X1 U14712 ( .A1(n12363), .A2(n12362), .ZN(n12304) );
  OR2_X1 U14713 ( .A1(n12348), .A2(n12306), .ZN(n12307) );
  NAND2_X1 U14714 ( .A1(n8449), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n12309) );
  INV_X1 U14715 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15494) );
  OR2_X1 U14716 ( .A1(n8451), .A2(n15494), .ZN(n12308) );
  NAND2_X1 U14717 ( .A1(n12309), .A2(n12308), .ZN(n12313) );
  INV_X1 U14718 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13232) );
  INV_X1 U14719 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12516) );
  OAI21_X1 U14720 ( .B1(n12321), .B2(n13232), .A(n12516), .ZN(n12310) );
  NAND2_X1 U14721 ( .A1(n12310), .A2(n13500), .ZN(n13532) );
  NOR2_X1 U14722 ( .A1(n8438), .A2(n13532), .ZN(n12312) );
  INV_X1 U14723 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13535) );
  NOR2_X1 U14724 ( .A1(n6568), .A2(n13535), .ZN(n12311) );
  AND2_X1 U14725 ( .A1(n13543), .A2(n12180), .ZN(n12314) );
  AOI21_X1 U14726 ( .B1(n13712), .B2(n12331), .A(n12314), .ZN(n12367) );
  NAND2_X1 U14727 ( .A1(n13712), .A2(n12275), .ZN(n12316) );
  NAND2_X1 U14728 ( .A1(n13543), .A2(n12331), .ZN(n12315) );
  NAND2_X1 U14729 ( .A1(n12316), .A2(n12315), .ZN(n12366) );
  NAND2_X1 U14730 ( .A1(n13811), .A2(n6581), .ZN(n12318) );
  OR2_X1 U14731 ( .A1(n12348), .A2(n13812), .ZN(n12317) );
  NAND2_X1 U14732 ( .A1(n12319), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n12326) );
  INV_X1 U14733 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n12320) );
  OR2_X1 U14734 ( .A1(n8765), .A2(n12320), .ZN(n12325) );
  XNOR2_X1 U14735 ( .A(n12321), .B(n13232), .ZN(n13551) );
  INV_X1 U14736 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13552) );
  OR2_X1 U14737 ( .A1(n6569), .A2(n13552), .ZN(n12323) );
  NAND4_X1 U14738 ( .A1(n12326), .A2(n12325), .A3(n12324), .A4(n12323), .ZN(
        n13571) );
  AND2_X1 U14739 ( .A1(n13571), .A2(n12275), .ZN(n12327) );
  AOI21_X1 U14740 ( .B1(n13717), .B2(n12331), .A(n12327), .ZN(n12374) );
  NAND2_X1 U14741 ( .A1(n13717), .A2(n12275), .ZN(n12329) );
  NAND2_X1 U14742 ( .A1(n13571), .A2(n12331), .ZN(n12328) );
  NAND2_X1 U14743 ( .A1(n12329), .A2(n12328), .ZN(n12373) );
  AND2_X1 U14744 ( .A1(n13570), .A2(n12180), .ZN(n12330) );
  AOI21_X1 U14745 ( .B1(n13727), .B2(n12331), .A(n12330), .ZN(n12339) );
  NAND2_X1 U14746 ( .A1(n13727), .A2(n12275), .ZN(n12333) );
  NAND2_X1 U14747 ( .A1(n13570), .A2(n12331), .ZN(n12332) );
  NAND2_X1 U14748 ( .A1(n12333), .A2(n12332), .ZN(n12338) );
  NAND2_X1 U14749 ( .A1(n12339), .A2(n12338), .ZN(n12334) );
  OAI21_X1 U14750 ( .B1(n12337), .B2(n12336), .A(n12335), .ZN(n12384) );
  INV_X1 U14751 ( .A(n12338), .ZN(n12341) );
  INV_X1 U14752 ( .A(n12339), .ZN(n12340) );
  INV_X1 U14753 ( .A(n12343), .ZN(n12346) );
  INV_X1 U14754 ( .A(n12344), .ZN(n12345) );
  NAND2_X1 U14755 ( .A1(n12346), .A2(n12345), .ZN(n12380) );
  NAND2_X1 U14756 ( .A1(n12347), .A2(n6581), .ZN(n12350) );
  OR2_X1 U14757 ( .A1(n12348), .A2(n15406), .ZN(n12349) );
  NAND2_X1 U14758 ( .A1(n13307), .A2(n12250), .ZN(n12354) );
  OR2_X1 U14759 ( .A1(n12351), .A2(n12352), .ZN(n12438) );
  NAND4_X1 U14760 ( .A1(n12354), .A2(n12353), .A3(n12438), .A4(n12389), .ZN(
        n12358) );
  INV_X1 U14761 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n15516) );
  NAND2_X1 U14762 ( .A1(n8436), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12356) );
  NAND2_X1 U14763 ( .A1(n8449), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12355) );
  OAI211_X1 U14764 ( .C1(n12357), .C2(n15516), .A(n12356), .B(n12355), .ZN(
        n13493) );
  AND2_X1 U14765 ( .A1(n12358), .A2(n13493), .ZN(n12359) );
  AOI21_X1 U14766 ( .B1(n13469), .B2(n12331), .A(n12359), .ZN(n12441) );
  NAND2_X1 U14767 ( .A1(n13469), .A2(n12275), .ZN(n12361) );
  NAND2_X1 U14768 ( .A1(n13493), .A2(n12331), .ZN(n12360) );
  NAND2_X1 U14769 ( .A1(n12361), .A2(n12360), .ZN(n12440) );
  OAI22_X1 U14770 ( .A1(n12441), .A2(n12440), .B1(n12363), .B2(n12362), .ZN(
        n12372) );
  MUX2_X1 U14771 ( .A(n13307), .B(n12331), .S(n12364), .Z(n12365) );
  NAND2_X1 U14772 ( .A1(n13307), .A2(n12331), .ZN(n12385) );
  NAND2_X1 U14773 ( .A1(n12365), .A2(n12385), .ZN(n12371) );
  INV_X1 U14774 ( .A(n12366), .ZN(n12369) );
  INV_X1 U14775 ( .A(n12367), .ZN(n12368) );
  AND2_X1 U14776 ( .A1(n12369), .A2(n12368), .ZN(n12370) );
  AOI22_X1 U14777 ( .A1(n12372), .A2(n12371), .B1(n7582), .B2(n12370), .ZN(
        n12378) );
  INV_X1 U14778 ( .A(n12373), .ZN(n12376) );
  INV_X1 U14779 ( .A(n12374), .ZN(n12375) );
  NAND3_X1 U14780 ( .A1(n6688), .A2(n12376), .A3(n12375), .ZN(n12377) );
  OAI211_X1 U14781 ( .C1(n12380), .C2(n12379), .A(n12378), .B(n12377), .ZN(
        n12381) );
  NOR2_X1 U14782 ( .A1(n12382), .A2(n12381), .ZN(n12383) );
  NAND2_X1 U14783 ( .A1(n12384), .A2(n12383), .ZN(n12455) );
  OR2_X1 U14784 ( .A1(n12364), .A2(n12385), .ZN(n12387) );
  INV_X1 U14785 ( .A(n13307), .ZN(n13466) );
  NAND3_X1 U14786 ( .A1(n12364), .A2(n13466), .A3(n12275), .ZN(n12386) );
  INV_X1 U14787 ( .A(n12388), .ZN(n12392) );
  OAI21_X1 U14788 ( .B1(n8881), .B2(n12436), .A(n12389), .ZN(n12390) );
  INV_X1 U14789 ( .A(n12390), .ZN(n12391) );
  AND2_X1 U14790 ( .A1(n12392), .A2(n12391), .ZN(n12444) );
  INV_X1 U14791 ( .A(n12444), .ZN(n12393) );
  NAND2_X1 U14792 ( .A1(n12446), .A2(n12393), .ZN(n12454) );
  XNOR2_X1 U14793 ( .A(n13469), .B(n13493), .ZN(n12434) );
  NAND2_X1 U14794 ( .A1(n13712), .A2(n13519), .ZN(n12394) );
  NAND2_X1 U14795 ( .A1(n13491), .A2(n12394), .ZN(n13489) );
  XNOR2_X1 U14796 ( .A(n13717), .B(n13490), .ZN(n13555) );
  NAND2_X1 U14797 ( .A1(n13722), .A2(n13517), .ZN(n13488) );
  OR2_X1 U14798 ( .A1(n13722), .A2(n13517), .ZN(n12395) );
  NAND2_X1 U14799 ( .A1(n13488), .A2(n12395), .ZN(n13487) );
  NAND2_X1 U14800 ( .A1(n13727), .A2(n13594), .ZN(n13486) );
  OR2_X1 U14801 ( .A1(n13727), .A2(n13594), .ZN(n12396) );
  NAND2_X1 U14802 ( .A1(n13732), .A2(n13516), .ZN(n13485) );
  OR2_X1 U14803 ( .A1(n13732), .A2(n13516), .ZN(n12397) );
  NAND2_X1 U14804 ( .A1(n13485), .A2(n12397), .ZN(n13598) );
  NAND2_X1 U14805 ( .A1(n13515), .A2(n13250), .ZN(n12398) );
  NAND2_X1 U14806 ( .A1(n13752), .A2(n13513), .ZN(n13479) );
  OR2_X1 U14807 ( .A1(n13752), .A2(n13513), .ZN(n12399) );
  XNOR2_X1 U14808 ( .A(n13757), .B(n13507), .ZN(n13685) );
  NOR2_X1 U14809 ( .A1(n12400), .A2(n8879), .ZN(n12404) );
  OR2_X1 U14810 ( .A1(n12144), .A2(n15035), .ZN(n12401) );
  NAND2_X1 U14811 ( .A1(n12402), .A2(n12401), .ZN(n15042) );
  NAND4_X1 U14812 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n15042), .ZN(
        n12408) );
  NOR3_X1 U14813 ( .A1(n12408), .A2(n12407), .A3(n12406), .ZN(n12411) );
  NAND4_X1 U14814 ( .A1(n12412), .A2(n12411), .A3(n12410), .A4(n12409), .ZN(
        n12413) );
  OR4_X1 U14815 ( .A1(n12416), .A2(n12415), .A3(n12414), .A4(n12413), .ZN(
        n12417) );
  NOR2_X1 U14816 ( .A1(n12418), .A2(n12417), .ZN(n12421) );
  NAND4_X1 U14817 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12423) );
  OR4_X1 U14818 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        n12427) );
  NOR2_X1 U14819 ( .A1(n13685), .A2(n12427), .ZN(n12428) );
  XNOR2_X1 U14820 ( .A(n13747), .B(n13666), .ZN(n13657) );
  NAND4_X1 U14821 ( .A1(n13636), .A2(n13664), .A3(n12428), .A4(n13657), .ZN(
        n12429) );
  NOR2_X1 U14822 ( .A1(n13598), .A2(n12429), .ZN(n12430) );
  XNOR2_X1 U14823 ( .A(n7056), .B(n13483), .ZN(n13625) );
  NAND3_X1 U14824 ( .A1(n13584), .A2(n12430), .A3(n13625), .ZN(n12431) );
  XNOR2_X1 U14825 ( .A(n13706), .B(n13528), .ZN(n13520) );
  NAND2_X1 U14826 ( .A1(n12435), .A2(n8881), .ZN(n12451) );
  NAND2_X1 U14827 ( .A1(n12437), .A2(n12436), .ZN(n12439) );
  AND2_X1 U14828 ( .A1(n12439), .A2(n12438), .ZN(n12448) );
  NAND2_X1 U14829 ( .A1(n12451), .A2(n12448), .ZN(n12442) );
  NAND2_X1 U14830 ( .A1(n12441), .A2(n12440), .ZN(n12445) );
  INV_X1 U14831 ( .A(n12446), .ZN(n12443) );
  NOR2_X1 U14832 ( .A1(n12443), .A2(n12351), .ZN(n12450) );
  OR2_X1 U14833 ( .A1(n12445), .A2(n12444), .ZN(n12447) );
  MUX2_X1 U14834 ( .A(n12448), .B(n12447), .S(n12446), .Z(n12449) );
  OAI21_X1 U14835 ( .B1(n12451), .B2(n12450), .A(n12449), .ZN(n12452) );
  INV_X1 U14836 ( .A(n12452), .ZN(n12453) );
  NAND4_X1 U14837 ( .A1(n13667), .A2(n12458), .A3(n15056), .A4(n12457), .ZN(
        n12459) );
  OAI211_X1 U14838 ( .C1(n12460), .C2(n7541), .A(n12459), .B(P2_B_REG_SCAN_IN), 
        .ZN(n12461) );
  INV_X1 U14839 ( .A(n13103), .ZN(n12946) );
  NAND2_X1 U14840 ( .A1(n12462), .A2(n12744), .ZN(n12463) );
  NAND2_X1 U14841 ( .A1(n12464), .A2(n12463), .ZN(n13073) );
  OR2_X1 U14842 ( .A1(n12466), .A2(n13062), .ZN(n12465) );
  NAND2_X1 U14843 ( .A1(n12466), .A2(n13062), .ZN(n12467) );
  AND2_X1 U14844 ( .A1(n13147), .A2(n12743), .ZN(n12469) );
  NAND2_X1 U14845 ( .A1(n13070), .A2(n13076), .ZN(n12468) );
  INV_X1 U14846 ( .A(n12475), .ZN(n12473) );
  OR2_X1 U14847 ( .A1(n13136), .A2(n12742), .ZN(n13027) );
  NAND2_X1 U14848 ( .A1(n13193), .A2(n13042), .ZN(n12471) );
  AND2_X1 U14849 ( .A1(n13027), .A2(n12471), .ZN(n12472) );
  NAND2_X1 U14850 ( .A1(n12474), .A2(n13010), .ZN(n12477) );
  NAND2_X1 U14851 ( .A1(n13020), .A2(n12740), .ZN(n12478) );
  AND2_X1 U14852 ( .A1(n13048), .A2(n12475), .ZN(n13009) );
  NAND2_X1 U14853 ( .A1(n12642), .A2(n13063), .ZN(n13007) );
  AND2_X1 U14854 ( .A1(n13009), .A2(n13007), .ZN(n12476) );
  OR2_X1 U14855 ( .A1(n12477), .A2(n12476), .ZN(n13012) );
  AND2_X1 U14856 ( .A1(n12478), .A2(n13012), .ZN(n12997) );
  OR2_X1 U14857 ( .A1(n7579), .A2(n12997), .ZN(n12479) );
  NAND2_X1 U14858 ( .A1(n12611), .A2(n13016), .ZN(n12481) );
  AND2_X1 U14859 ( .A1(n12483), .A2(n12739), .ZN(n12484) );
  INV_X1 U14860 ( .A(n13107), .ZN(n12962) );
  NOR2_X1 U14861 ( .A1(n12905), .A2(n7580), .ZN(n12485) );
  OAI211_X1 U14862 ( .C1(n12485), .C2(n12492), .A(n12525), .B(n15149), .ZN(
        n12487) );
  AOI22_X1 U14863 ( .A1(n12737), .A2(n15154), .B1(n12736), .B2(n15155), .ZN(
        n12486) );
  INV_X1 U14864 ( .A(n12488), .ZN(n12490) );
  OAI22_X1 U14865 ( .A1(n12490), .A2(n15184), .B1(n15198), .B2(n12489), .ZN(
        n12494) );
  XOR2_X1 U14866 ( .A(n12492), .B(n12491), .Z(n13092) );
  NOR2_X1 U14867 ( .A1(n13092), .A2(n12983), .ZN(n12493) );
  AOI211_X1 U14868 ( .C1(n14583), .C2(n12495), .A(n12494), .B(n12493), .ZN(
        n12496) );
  OAI21_X1 U14869 ( .B1(n13091), .B2(n14582), .A(n12496), .ZN(P3_U3205) );
  INV_X1 U14870 ( .A(n12497), .ZN(n12498) );
  OAI222_X1 U14871 ( .A1(P3_U3151), .A2(n12862), .B1(n13228), .B2(n12499), 
        .C1(n13227), .C2(n12498), .ZN(P3_U3268) );
  INV_X1 U14872 ( .A(n12500), .ZN(n12501) );
  XNOR2_X1 U14873 ( .A(n13722), .B(n12513), .ZN(n12504) );
  NOR2_X1 U14874 ( .A1(n13517), .A2(n6577), .ZN(n12505) );
  XNOR2_X1 U14875 ( .A(n12504), .B(n12505), .ZN(n13301) );
  INV_X1 U14876 ( .A(n13301), .ZN(n12503) );
  INV_X1 U14877 ( .A(n12504), .ZN(n12507) );
  INV_X1 U14878 ( .A(n12505), .ZN(n12506) );
  NAND2_X1 U14879 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  XNOR2_X1 U14880 ( .A(n13717), .B(n12513), .ZN(n12510) );
  AND2_X1 U14881 ( .A1(n13571), .A2(n8705), .ZN(n12509) );
  NAND2_X1 U14882 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  OAI21_X1 U14883 ( .B1(n12510), .B2(n12509), .A(n12511), .ZN(n13231) );
  NOR2_X1 U14884 ( .A1(n13519), .A2(n6577), .ZN(n12512) );
  XOR2_X1 U14885 ( .A(n12513), .B(n12512), .Z(n12514) );
  XNOR2_X1 U14886 ( .A(n13712), .B(n12514), .ZN(n12515) );
  INV_X1 U14887 ( .A(n13528), .ZN(n12517) );
  OAI22_X1 U14888 ( .A1(n14932), .A2(n12517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12516), .ZN(n12519) );
  OAI22_X1 U14889 ( .A1(n14933), .A2(n13490), .B1(n14947), .B2(n13532), .ZN(
        n12518) );
  AOI211_X1 U14890 ( .C1(n13712), .C2(n14943), .A(n12519), .B(n12518), .ZN(
        n12520) );
  INV_X1 U14891 ( .A(n12521), .ZN(n12523) );
  OAI222_X1 U14892 ( .A1(n12524), .A2(P3_U3151), .B1(n13227), .B2(n12523), 
        .C1(n12522), .C2(n13228), .ZN(P3_U3265) );
  XNOR2_X1 U14893 ( .A(n12526), .B(n12538), .ZN(n12532) );
  INV_X1 U14894 ( .A(P3_B_REG_SCAN_IN), .ZN(n12527) );
  NOR2_X1 U14895 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  OR2_X1 U14896 ( .A1(n15193), .A2(n12529), .ZN(n12898) );
  OAI22_X1 U14897 ( .A1(n12909), .A2(n15195), .B1(n12530), .B2(n12898), .ZN(
        n12531) );
  AOI21_X2 U14898 ( .B1(n12532), .B2(n15149), .A(n12531), .ZN(n13089) );
  NOR2_X1 U14899 ( .A1(n12533), .A2(n15184), .ZN(n12900) );
  INV_X1 U14900 ( .A(n12534), .ZN(n12535) );
  NAND2_X1 U14901 ( .A1(n12535), .A2(n15210), .ZN(n13088) );
  NOR2_X1 U14902 ( .A1(n13088), .A2(n14596), .ZN(n12536) );
  AOI211_X1 U14903 ( .C1(n14582), .C2(P3_REG2_REG_29__SCAN_IN), .A(n12900), 
        .B(n12536), .ZN(n12540) );
  XOR2_X1 U14904 ( .A(n12538), .B(n12537), .Z(n13090) );
  OR2_X1 U14905 ( .A1(n13090), .A2(n12983), .ZN(n12539) );
  OAI211_X1 U14906 ( .C1(n13089), .C2(n14582), .A(n12540), .B(n12539), .ZN(
        P3_U3204) );
  AND2_X1 U14907 ( .A1(n12626), .A2(n12541), .ZN(n12711) );
  XNOR2_X1 U14908 ( .A(n12542), .B(n12631), .ZN(n12710) );
  NAND2_X1 U14909 ( .A1(n12711), .A2(n12710), .ZN(n12709) );
  NAND2_X1 U14910 ( .A1(n12709), .A2(n12543), .ZN(n12595) );
  XNOR2_X1 U14911 ( .A(n12595), .B(n12594), .ZN(n12544) );
  NAND2_X1 U14912 ( .A1(n12544), .A2(n12724), .ZN(n12550) );
  AOI21_X1 U14913 ( .B1(n12713), .B2(n12747), .A(n12545), .ZN(n12549) );
  AOI22_X1 U14914 ( .A1(n12715), .A2(n15209), .B1(n12726), .B2(n12631), .ZN(
        n12548) );
  NAND2_X1 U14915 ( .A1(n12731), .A2(n12546), .ZN(n12547) );
  NAND4_X1 U14916 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        P3_U3153) );
  OAI21_X1 U14917 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(n12554) );
  AOI22_X1 U14918 ( .A1(n12939), .A2(n12726), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12555) );
  OAI21_X1 U14919 ( .B1(n12909), .B2(n12729), .A(n12555), .ZN(n12556) );
  AOI21_X1 U14920 ( .B1(n12911), .B2(n12731), .A(n12556), .ZN(n12557) );
  OAI21_X1 U14921 ( .B1(n12986), .B2(n12559), .A(n12558), .ZN(n12560) );
  NAND2_X1 U14922 ( .A1(n12560), .A2(n12724), .ZN(n12565) );
  AOI22_X1 U14923 ( .A1(n12726), .A2(n12739), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12562) );
  OAI21_X1 U14924 ( .B1(n12972), .B2(n12729), .A(n12562), .ZN(n12563) );
  AOI21_X1 U14925 ( .B1(n12976), .B2(n12731), .A(n12563), .ZN(n12564) );
  OAI211_X1 U14926 ( .C1(n13111), .C2(n12734), .A(n12565), .B(n12564), .ZN(
        P3_U3156) );
  AND2_X1 U14927 ( .A1(n12670), .A2(n12566), .ZN(n12569) );
  OAI211_X1 U14928 ( .C1(n12569), .C2(n12568), .A(n12724), .B(n12567), .ZN(
        n12574) );
  INV_X1 U14929 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n12570) );
  NOR2_X1 U14930 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12570), .ZN(n12762) );
  AOI21_X1 U14931 ( .B1(n12713), .B2(n15156), .A(n12762), .ZN(n12573) );
  AOI22_X1 U14932 ( .A1(n12715), .A2(n15159), .B1(n12726), .B2(n15153), .ZN(
        n12572) );
  NAND2_X1 U14933 ( .A1(n12731), .A2(n15160), .ZN(n12571) );
  NAND4_X1 U14934 ( .A1(n12574), .A2(n12573), .A3(n12572), .A4(n12571), .ZN(
        P3_U3157) );
  AND2_X1 U14935 ( .A1(n12576), .A2(n12575), .ZN(n12579) );
  OAI211_X1 U14936 ( .C1(n12579), .C2(n12578), .A(n12724), .B(n12577), .ZN(
        n12586) );
  AOI21_X1 U14937 ( .B1(n12713), .B2(n12750), .A(n12580), .ZN(n12585) );
  AOI22_X1 U14938 ( .A1(n12715), .A2(n12581), .B1(n12726), .B2(n12752), .ZN(
        n12584) );
  NAND2_X1 U14939 ( .A1(n12731), .A2(n12582), .ZN(n12583) );
  NAND4_X1 U14940 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        P3_U3158) );
  OAI211_X1 U14941 ( .C1(n12589), .C2(n12588), .A(n12587), .B(n12724), .ZN(
        n12593) );
  NAND2_X1 U14942 ( .A1(n12726), .A2(n12742), .ZN(n12590) );
  NAND2_X1 U14943 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12881)
         );
  OAI211_X1 U14944 ( .C1(n13030), .C2(n12729), .A(n12590), .B(n12881), .ZN(
        n12591) );
  AOI21_X1 U14945 ( .B1(n13034), .B2(n12731), .A(n12591), .ZN(n12592) );
  OAI211_X1 U14946 ( .C1(n12734), .C2(n13193), .A(n12593), .B(n12592), .ZN(
        P3_U3159) );
  MUX2_X1 U14947 ( .A(n12595), .B(n12748), .S(n12594), .Z(n12597) );
  XNOR2_X1 U14948 ( .A(n12597), .B(n12596), .ZN(n12598) );
  NAND2_X1 U14949 ( .A1(n12598), .A2(n12724), .ZN(n12605) );
  AOI21_X1 U14950 ( .B1(n12713), .B2(n15153), .A(n12599), .ZN(n12604) );
  AOI22_X1 U14951 ( .A1(n12715), .A2(n12600), .B1(n12726), .B2(n12748), .ZN(
        n12603) );
  NAND2_X1 U14952 ( .A1(n12731), .A2(n12601), .ZN(n12602) );
  NAND4_X1 U14953 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n12602), .ZN(
        P3_U3161) );
  INV_X1 U14954 ( .A(n12606), .ZN(n12607) );
  AOI21_X1 U14955 ( .B1(n12609), .B2(n12608), .A(n12607), .ZN(n12615) );
  AOI22_X1 U14956 ( .A1(n12726), .A2(n12740), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12610) );
  OAI21_X1 U14957 ( .B1(n7036), .B2(n12729), .A(n12610), .ZN(n12613) );
  NOR2_X1 U14958 ( .A1(n13187), .A2(n12734), .ZN(n12612) );
  AOI211_X1 U14959 ( .C1(n13002), .C2(n12731), .A(n12613), .B(n12612), .ZN(
        n12614) );
  OAI21_X1 U14960 ( .B1(n12615), .B2(n12699), .A(n12614), .ZN(P3_U3163) );
  INV_X1 U14961 ( .A(n12616), .ZN(n12621) );
  NOR3_X1 U14962 ( .A1(n12617), .A2(n12619), .A3(n12618), .ZN(n12620) );
  OAI21_X1 U14963 ( .B1(n12621), .B2(n12620), .A(n12724), .ZN(n12625) );
  NOR2_X1 U14964 ( .A1(n12972), .A2(n12685), .ZN(n12623) );
  OAI22_X1 U14965 ( .A1(n12910), .A2(n12729), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15524), .ZN(n12622) );
  AOI211_X1 U14966 ( .C1(n12944), .C2(n12731), .A(n12623), .B(n12622), .ZN(
        n12624) );
  OAI211_X1 U14967 ( .C1(n12946), .C2(n12734), .A(n12625), .B(n12624), .ZN(
        P3_U3165) );
  OAI21_X1 U14968 ( .B1(n12628), .B2(n12627), .A(n12626), .ZN(n12629) );
  NAND2_X1 U14969 ( .A1(n12629), .A2(n12724), .ZN(n12637) );
  AOI21_X1 U14970 ( .B1(n12713), .B2(n12631), .A(n12630), .ZN(n12636) );
  AOI22_X1 U14971 ( .A1(n12715), .A2(n12632), .B1(n12726), .B2(n12750), .ZN(
        n12635) );
  NAND2_X1 U14972 ( .A1(n12731), .A2(n12633), .ZN(n12634) );
  NAND4_X1 U14973 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        P3_U3167) );
  XNOR2_X1 U14974 ( .A(n12638), .B(n13041), .ZN(n12639) );
  XNOR2_X1 U14975 ( .A(n6813), .B(n12639), .ZN(n12646) );
  NAND2_X1 U14976 ( .A1(n12726), .A2(n12743), .ZN(n12641) );
  NAND2_X1 U14977 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12835)
         );
  OAI211_X1 U14978 ( .C1(n13053), .C2(n12729), .A(n12641), .B(n12835), .ZN(
        n12644) );
  INV_X1 U14979 ( .A(n12642), .ZN(n13199) );
  NOR2_X1 U14980 ( .A1(n13199), .A2(n12734), .ZN(n12643) );
  AOI211_X1 U14981 ( .C1(n13056), .C2(n12731), .A(n12644), .B(n12643), .ZN(
        n12645) );
  OAI21_X1 U14982 ( .B1(n12646), .B2(n12699), .A(n12645), .ZN(P3_U3168) );
  AND3_X1 U14983 ( .A1(n12558), .A2(n12648), .A3(n12647), .ZN(n12649) );
  OAI21_X1 U14984 ( .B1(n12617), .B2(n12649), .A(n12724), .ZN(n12656) );
  OAI22_X1 U14985 ( .A1(n12951), .A2(n12729), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12650), .ZN(n12654) );
  INV_X1 U14986 ( .A(n12731), .ZN(n12652) );
  INV_X1 U14987 ( .A(n12960), .ZN(n12651) );
  NOR2_X1 U14988 ( .A1(n12652), .A2(n12651), .ZN(n12653) );
  AOI211_X1 U14989 ( .C1(n12726), .C2(n12738), .A(n12654), .B(n12653), .ZN(
        n12655) );
  OAI211_X1 U14990 ( .C1(n12962), .C2(n12734), .A(n12656), .B(n12655), .ZN(
        P3_U3169) );
  INV_X1 U14991 ( .A(n12657), .ZN(n12658) );
  AOI21_X1 U14992 ( .B1(n12660), .B2(n12659), .A(n12658), .ZN(n12661) );
  OR2_X1 U14993 ( .A1(n12661), .A2(n12699), .ZN(n12668) );
  AOI21_X1 U14994 ( .B1(n12713), .B2(n12749), .A(n12662), .ZN(n12667) );
  AOI22_X1 U14995 ( .A1(n12715), .A2(n12663), .B1(n12726), .B2(n12751), .ZN(
        n12666) );
  NAND2_X1 U14996 ( .A1(n12731), .A2(n12664), .ZN(n12665) );
  NAND4_X1 U14997 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        P3_U3170) );
  INV_X1 U14998 ( .A(n12670), .ZN(n12671) );
  AOI21_X1 U14999 ( .B1(n12672), .B2(n12669), .A(n12671), .ZN(n12673) );
  OR2_X1 U15000 ( .A1(n12673), .A2(n12699), .ZN(n12680) );
  AOI21_X1 U15001 ( .B1(n12713), .B2(n12746), .A(n12674), .ZN(n12679) );
  AOI22_X1 U15002 ( .A1(n12715), .A2(n12675), .B1(n12726), .B2(n12747), .ZN(
        n12678) );
  NAND2_X1 U15003 ( .A1(n12731), .A2(n12676), .ZN(n12677) );
  NAND4_X1 U15004 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        P3_U3171) );
  XNOR2_X1 U15005 ( .A(n12681), .B(n12740), .ZN(n12682) );
  XNOR2_X1 U15006 ( .A(n12683), .B(n12682), .ZN(n12689) );
  AOI22_X1 U15007 ( .A1(n12713), .A2(n13016), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12684) );
  OAI21_X1 U15008 ( .B1(n13042), .B2(n12685), .A(n12684), .ZN(n12687) );
  INV_X1 U15009 ( .A(n13020), .ZN(n13190) );
  NOR2_X1 U15010 ( .A1(n13190), .A2(n12734), .ZN(n12686) );
  AOI211_X1 U15011 ( .C1(n13019), .C2(n12731), .A(n12687), .B(n12686), .ZN(
        n12688) );
  OAI21_X1 U15012 ( .B1(n12689), .B2(n12699), .A(n12688), .ZN(P3_U3173) );
  XNOR2_X1 U15013 ( .A(n12690), .B(n12691), .ZN(n12692) );
  NAND2_X1 U15014 ( .A1(n12692), .A2(n12724), .ZN(n12698) );
  AOI21_X1 U15015 ( .B1(n12713), .B2(n12745), .A(n12693), .ZN(n12697) );
  AOI22_X1 U15016 ( .A1(n12715), .A2(n12694), .B1(n12726), .B2(n12746), .ZN(
        n12696) );
  NAND2_X1 U15017 ( .A1(n12731), .A2(n14604), .ZN(n12695) );
  NAND4_X1 U15018 ( .A1(n12698), .A2(n12697), .A3(n12696), .A4(n12695), .ZN(
        P3_U3176) );
  INV_X1 U15019 ( .A(n13136), .ZN(n12708) );
  AOI21_X1 U15020 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n12703) );
  NAND2_X1 U15021 ( .A1(n12703), .A2(n12702), .ZN(n12707) );
  NAND2_X1 U15022 ( .A1(n12726), .A2(n13063), .ZN(n12704) );
  NAND2_X1 U15023 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12861)
         );
  OAI211_X1 U15024 ( .C1(n13042), .C2(n12729), .A(n12704), .B(n12861), .ZN(
        n12705) );
  AOI21_X1 U15025 ( .B1(n13045), .B2(n12731), .A(n12705), .ZN(n12706) );
  OAI211_X1 U15026 ( .C1(n12708), .C2(n12734), .A(n12707), .B(n12706), .ZN(
        P3_U3178) );
  OAI211_X1 U15027 ( .C1(n12711), .C2(n12710), .A(n12709), .B(n12724), .ZN(
        n12720) );
  AOI21_X1 U15028 ( .B1(n12713), .B2(n12748), .A(n12712), .ZN(n12719) );
  AOI22_X1 U15029 ( .A1(n12715), .A2(n12714), .B1(n12726), .B2(n12749), .ZN(
        n12718) );
  NAND2_X1 U15030 ( .A1(n12731), .A2(n12716), .ZN(n12717) );
  NAND4_X1 U15031 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        P3_U3179) );
  OAI21_X1 U15032 ( .B1(n12723), .B2(n12722), .A(n12721), .ZN(n12725) );
  NAND2_X1 U15033 ( .A1(n12725), .A2(n12724), .ZN(n12733) );
  AOI22_X1 U15034 ( .A1(n12727), .A2(n12726), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12728) );
  OAI21_X1 U15035 ( .B1(n12923), .B2(n12729), .A(n12728), .ZN(n12730) );
  AOI21_X1 U15036 ( .B1(n12927), .B2(n12731), .A(n12730), .ZN(n12732) );
  OAI211_X1 U15037 ( .C1(n13175), .C2(n12734), .A(n12733), .B(n12732), .ZN(
        P3_U3180) );
  MUX2_X1 U15038 ( .A(n12735), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12753), .Z(
        P3_U3521) );
  MUX2_X1 U15039 ( .A(n12736), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12753), .Z(
        P3_U3520) );
  MUX2_X1 U15040 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12737), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15041 ( .A(n12939), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12753), .Z(
        P3_U3517) );
  MUX2_X1 U15042 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12938), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15043 ( .A(n12738), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12753), .Z(
        P3_U3514) );
  MUX2_X1 U15044 ( .A(n12739), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12753), .Z(
        P3_U3513) );
  MUX2_X1 U15045 ( .A(n13016), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12753), .Z(
        P3_U3512) );
  MUX2_X1 U15046 ( .A(n12740), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12753), .Z(
        P3_U3511) );
  MUX2_X1 U15047 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n6752), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15048 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12742), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15049 ( .A(n12743), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12753), .Z(
        P3_U3507) );
  MUX2_X1 U15050 ( .A(n13062), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12753), .Z(
        P3_U3506) );
  MUX2_X1 U15051 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12744), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15052 ( .A(n14591), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12753), .Z(
        P3_U3504) );
  MUX2_X1 U15053 ( .A(n12745), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12753), .Z(
        P3_U3503) );
  MUX2_X1 U15054 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15156), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15055 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12746), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15056 ( .A(n15153), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12753), .Z(
        P3_U3500) );
  MUX2_X1 U15057 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12747), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15058 ( .A(n12748), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12753), .Z(
        P3_U3498) );
  MUX2_X1 U15059 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12749), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15060 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12750), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15061 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12751), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15062 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12752), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15063 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9503), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15064 ( .A(n12754), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12753), .Z(
        P3_U3491) );
  AND3_X1 U15065 ( .A1(n12757), .A2(n12756), .A3(n12755), .ZN(n12758) );
  OAI21_X1 U15066 ( .B1(n12759), .B2(n12758), .A(n12819), .ZN(n12777) );
  INV_X1 U15067 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n12760) );
  NOR2_X1 U15068 ( .A1(n12837), .A2(n12760), .ZN(n12761) );
  AOI211_X1 U15069 ( .C1(n12834), .C2(n12763), .A(n12762), .B(n12761), .ZN(
        n12776) );
  AND3_X1 U15070 ( .A1(n12766), .A2(n12765), .A3(n12764), .ZN(n12768) );
  OAI21_X1 U15071 ( .B1(n12769), .B2(n12768), .A(n12767), .ZN(n12775) );
  OAI21_X1 U15072 ( .B1(n12772), .B2(n12771), .A(n12770), .ZN(n12773) );
  NAND2_X1 U15073 ( .A1(n12773), .A2(n12895), .ZN(n12774) );
  NAND4_X1 U15074 ( .A1(n12777), .A2(n12776), .A3(n12775), .A4(n12774), .ZN(
        P3_U3192) );
  INV_X1 U15075 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U15076 ( .A1(n12787), .A2(n12779), .ZN(n12813) );
  AOI21_X1 U15077 ( .B1(n12781), .B2(n12780), .A(n12815), .ZN(n12799) );
  NAND2_X1 U15078 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12784), .ZN(n12807) );
  OAI21_X1 U15079 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12784), .A(n12807), 
        .ZN(n12797) );
  INV_X1 U15080 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U15081 ( .A1(n12834), .A2(n12801), .ZN(n12786) );
  OAI211_X1 U15082 ( .C1(n14469), .C2(n12837), .A(n12786), .B(n12785), .ZN(
        n12796) );
  INV_X1 U15083 ( .A(n12787), .ZN(n12789) );
  MUX2_X1 U15084 ( .A(n12789), .B(n12788), .S(n12862), .Z(n12790) );
  MUX2_X1 U15085 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12862), .Z(n12792) );
  AOI21_X1 U15086 ( .B1(n12793), .B2(n12792), .A(n12800), .ZN(n12794) );
  NOR2_X1 U15087 ( .A1(n12794), .A2(n12891), .ZN(n12795) );
  AOI211_X1 U15088 ( .C1(n12895), .C2(n12797), .A(n12796), .B(n12795), .ZN(
        n12798) );
  OAI21_X1 U15089 ( .B1(n12799), .B2(n12896), .A(n12798), .ZN(P3_U3197) );
  INV_X1 U15090 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12824) );
  INV_X1 U15091 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12829) );
  MUX2_X1 U15092 ( .A(n12824), .B(n12829), .S(n12862), .Z(n12803) );
  NOR2_X1 U15093 ( .A1(n12803), .A2(n12830), .ZN(n12839) );
  NAND2_X1 U15094 ( .A1(n12803), .A2(n12830), .ZN(n12838) );
  INV_X1 U15095 ( .A(n12838), .ZN(n12804) );
  NOR2_X1 U15096 ( .A1(n12839), .A2(n12804), .ZN(n12805) );
  XNOR2_X1 U15097 ( .A(n12840), .B(n12805), .ZN(n12823) );
  NAND2_X1 U15098 ( .A1(n12814), .A2(n12806), .ZN(n12808) );
  AND2_X1 U15099 ( .A1(n12808), .A2(n12807), .ZN(n12832) );
  XNOR2_X1 U15100 ( .A(n12830), .B(n12829), .ZN(n12831) );
  XNOR2_X1 U15101 ( .A(n12832), .B(n12831), .ZN(n12812) );
  INV_X1 U15102 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U15103 ( .A1(n12834), .A2(n12830), .ZN(n12810) );
  OAI211_X1 U15104 ( .C1(n15303), .C2(n12837), .A(n12810), .B(n12809), .ZN(
        n12811) );
  AOI21_X1 U15105 ( .B1(n12812), .B2(n12895), .A(n12811), .ZN(n12822) );
  AND2_X1 U15106 ( .A1(n12814), .A2(n12813), .ZN(n12816) );
  OR2_X1 U15107 ( .A1(n12830), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U15108 ( .A1(n12830), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12817) );
  OAI21_X1 U15109 ( .B1(n7296), .B2(n6738), .A(n12826), .ZN(n12820) );
  NAND2_X1 U15110 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  OAI211_X1 U15111 ( .C1(n12823), .C2(n12891), .A(n12822), .B(n12821), .ZN(
        P3_U3198) );
  INV_X1 U15112 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12828) );
  OR2_X1 U15113 ( .A1(n12830), .A2(n12824), .ZN(n12825) );
  AOI21_X1 U15114 ( .B1(n12828), .B2(n12827), .A(n12850), .ZN(n12847) );
  XNOR2_X1 U15115 ( .A(n12855), .B(n12849), .ZN(n12833) );
  NAND2_X1 U15116 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n12833), .ZN(n12856) );
  OAI21_X1 U15117 ( .B1(n12833), .B2(P3_REG1_REG_17__SCAN_IN), .A(n12856), 
        .ZN(n12845) );
  INV_X1 U15118 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U15119 ( .A1(n12834), .A2(n12849), .ZN(n12836) );
  OAI211_X1 U15120 ( .C1(n14538), .C2(n12837), .A(n12836), .B(n12835), .ZN(
        n12844) );
  MUX2_X1 U15121 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12862), .Z(n12865) );
  XNOR2_X1 U15122 ( .A(n12865), .B(n12864), .ZN(n12842) );
  AOI211_X1 U15123 ( .C1(n12842), .C2(n12841), .A(n12891), .B(n12863), .ZN(
        n12843) );
  AOI211_X1 U15124 ( .C1(n12895), .C2(n12845), .A(n12844), .B(n12843), .ZN(
        n12846) );
  OAI21_X1 U15125 ( .B1(n12847), .B2(n12896), .A(n12846), .ZN(P3_U3199) );
  NOR2_X1 U15126 ( .A1(n12849), .A2(n12848), .ZN(n12851) );
  NOR2_X1 U15127 ( .A1(n12851), .A2(n12850), .ZN(n12854) );
  INV_X1 U15128 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15129 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n12888), .B1(n12875), 
        .B2(n12852), .ZN(n12853) );
  NOR2_X1 U15130 ( .A1(n12854), .A2(n12853), .ZN(n12874) );
  AOI21_X1 U15131 ( .B1(n12854), .B2(n12853), .A(n12874), .ZN(n12873) );
  INV_X1 U15132 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U15133 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12875), .B1(n12888), 
        .B2(n13141), .ZN(n12859) );
  NAND2_X1 U15134 ( .A1(n12864), .A2(n12855), .ZN(n12857) );
  NAND2_X1 U15135 ( .A1(n12857), .A2(n12856), .ZN(n12858) );
  OAI21_X1 U15136 ( .B1(n12859), .B2(n12858), .A(n12877), .ZN(n12871) );
  NAND2_X1 U15137 ( .A1(n15142), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12860) );
  OAI211_X1 U15138 ( .C1(n12883), .C2(n12875), .A(n12861), .B(n12860), .ZN(
        n12870) );
  MUX2_X1 U15139 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12862), .Z(n12867) );
  XNOR2_X1 U15140 ( .A(n12889), .B(n12888), .ZN(n12866) );
  AOI21_X1 U15141 ( .B1(n12867), .B2(n12866), .A(n12887), .ZN(n12868) );
  NOR2_X1 U15142 ( .A1(n12868), .A2(n12891), .ZN(n12869) );
  AOI211_X1 U15143 ( .C1(n12895), .C2(n12871), .A(n12870), .B(n12869), .ZN(
        n12872) );
  OAI21_X1 U15144 ( .B1(n12873), .B2(n12896), .A(n12872), .ZN(P3_U3200) );
  XNOR2_X1 U15145 ( .A(n6589), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12885) );
  XOR2_X1 U15146 ( .A(n12885), .B(n12876), .Z(n12897) );
  XNOR2_X1 U15147 ( .A(n6589), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12886) );
  INV_X1 U15148 ( .A(n12886), .ZN(n12878) );
  XNOR2_X1 U15149 ( .A(n12879), .B(n12878), .ZN(n12894) );
  NAND2_X1 U15150 ( .A1(n15142), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12880) );
  OAI211_X1 U15151 ( .C1(n12883), .C2(n6589), .A(n12881), .B(n12880), .ZN(
        n12893) );
  MUX2_X1 U15152 ( .A(n12886), .B(n12885), .S(n12884), .Z(n12890) );
  OAI21_X1 U15153 ( .B1(n14616), .B2(n12900), .A(n15198), .ZN(n14584) );
  NAND2_X1 U15154 ( .A1(n14582), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12901) );
  OAI211_X1 U15155 ( .C1(n13167), .C2(n13081), .A(n14584), .B(n12901), .ZN(
        P3_U3202) );
  AOI21_X1 U15156 ( .B1(n12904), .B2(n12903), .A(n12902), .ZN(n13095) );
  AOI21_X1 U15157 ( .B1(n12907), .B2(n12906), .A(n12905), .ZN(n12908) );
  OAI222_X1 U15158 ( .A1(n15195), .A2(n12910), .B1(n15193), .B2(n12909), .C1(
        n15191), .C2(n12908), .ZN(n13097) );
  NAND2_X1 U15159 ( .A1(n13097), .A2(n15198), .ZN(n12917) );
  INV_X1 U15160 ( .A(n12911), .ZN(n12913) );
  OAI22_X1 U15161 ( .A1(n12913), .A2(n15184), .B1(n15198), .B2(n12912), .ZN(
        n12914) );
  AOI21_X1 U15162 ( .B1(n12915), .B2(n14583), .A(n12914), .ZN(n12916) );
  OAI211_X1 U15163 ( .C1(n13095), .C2(n12983), .A(n12917), .B(n12916), .ZN(
        P3_U3206) );
  XNOR2_X1 U15164 ( .A(n12919), .B(n12918), .ZN(n13100) );
  INV_X1 U15165 ( .A(n13100), .ZN(n12935) );
  XNOR2_X1 U15166 ( .A(n12921), .B(n12920), .ZN(n12926) );
  INV_X1 U15167 ( .A(n12922), .ZN(n15170) );
  OAI22_X1 U15168 ( .A1(n12923), .A2(n15193), .B1(n12951), .B2(n15195), .ZN(
        n12924) );
  AOI21_X1 U15169 ( .B1(n13100), .B2(n15170), .A(n12924), .ZN(n12925) );
  OAI21_X1 U15170 ( .B1(n12926), .B2(n15191), .A(n12925), .ZN(n13099) );
  NAND2_X1 U15171 ( .A1(n13099), .A2(n15198), .ZN(n12933) );
  NAND2_X1 U15172 ( .A1(n12927), .A2(n15178), .ZN(n12928) );
  OAI21_X1 U15173 ( .B1(n15198), .B2(n12929), .A(n12928), .ZN(n12930) );
  AOI21_X1 U15174 ( .B1(n12931), .B2(n14583), .A(n12930), .ZN(n12932) );
  OAI211_X1 U15175 ( .C1(n12935), .C2(n12934), .A(n12933), .B(n12932), .ZN(
        P3_U3207) );
  OAI211_X1 U15176 ( .C1(n12937), .C2(n12942), .A(n12936), .B(n15149), .ZN(
        n12941) );
  AOI22_X1 U15177 ( .A1(n12939), .A2(n15155), .B1(n12938), .B2(n15154), .ZN(
        n12940) );
  AND2_X1 U15178 ( .A1(n12941), .A2(n12940), .ZN(n13105) );
  XNOR2_X1 U15179 ( .A(n12943), .B(n12942), .ZN(n13106) );
  INV_X1 U15180 ( .A(n13106), .ZN(n12948) );
  AOI22_X1 U15181 ( .A1(n14582), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15178), 
        .B2(n12944), .ZN(n12945) );
  OAI21_X1 U15182 ( .B1(n12946), .B2(n13081), .A(n12945), .ZN(n12947) );
  AOI21_X1 U15183 ( .B1(n12948), .B2(n14611), .A(n12947), .ZN(n12949) );
  OAI21_X1 U15184 ( .B1(n13105), .B2(n14582), .A(n12949), .ZN(P3_U3208) );
  INV_X1 U15185 ( .A(n12955), .ZN(n12950) );
  AOI21_X1 U15186 ( .B1(n6644), .B2(n12950), .A(n15191), .ZN(n12954) );
  OAI22_X1 U15187 ( .A1(n12951), .A2(n15193), .B1(n12986), .B2(n15195), .ZN(
        n12952) );
  AOI21_X1 U15188 ( .B1(n12954), .B2(n12953), .A(n12952), .ZN(n13110) );
  INV_X1 U15189 ( .A(n12967), .ZN(n12957) );
  OAI21_X1 U15190 ( .B1(n12957), .B2(n12956), .A(n12955), .ZN(n12959) );
  NAND2_X1 U15191 ( .A1(n12959), .A2(n12958), .ZN(n13108) );
  AOI22_X1 U15192 ( .A1(n14582), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15178), 
        .B2(n12960), .ZN(n12961) );
  OAI21_X1 U15193 ( .B1(n12962), .B2(n13081), .A(n12961), .ZN(n12963) );
  AOI21_X1 U15194 ( .B1(n13108), .B2(n14611), .A(n12963), .ZN(n12964) );
  OAI21_X1 U15195 ( .B1(n13110), .B2(n14582), .A(n12964), .ZN(P3_U3209) );
  OR2_X1 U15196 ( .A1(n12965), .A2(n12968), .ZN(n12966) );
  NAND2_X1 U15197 ( .A1(n12967), .A2(n12966), .ZN(n13113) );
  NAND2_X1 U15198 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  NAND3_X1 U15199 ( .A1(n12971), .A2(n15149), .A3(n12970), .ZN(n12975) );
  OAI22_X1 U15200 ( .A1(n12972), .A2(n15193), .B1(n7036), .B2(n15195), .ZN(
        n12973) );
  INV_X1 U15201 ( .A(n12973), .ZN(n12974) );
  NAND2_X1 U15202 ( .A1(n12975), .A2(n12974), .ZN(n13115) );
  NAND2_X1 U15203 ( .A1(n13115), .A2(n15198), .ZN(n12982) );
  INV_X1 U15204 ( .A(n12976), .ZN(n12977) );
  OAI22_X1 U15205 ( .A1(n15198), .A2(n12978), .B1(n12977), .B2(n15184), .ZN(
        n12979) );
  AOI21_X1 U15206 ( .B1(n12980), .B2(n14583), .A(n12979), .ZN(n12981) );
  OAI211_X1 U15207 ( .C1(n12983), .C2(n13113), .A(n12982), .B(n12981), .ZN(
        P3_U3210) );
  XOR2_X1 U15208 ( .A(n12984), .B(n12989), .Z(n12985) );
  OAI222_X1 U15209 ( .A1(n15195), .A2(n12987), .B1(n15193), .B2(n12986), .C1(
        n12985), .C2(n15191), .ZN(n13118) );
  INV_X1 U15210 ( .A(n13118), .ZN(n12994) );
  XOR2_X1 U15211 ( .A(n12988), .B(n12989), .Z(n13119) );
  AOI22_X1 U15212 ( .A1(n14582), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15178), 
        .B2(n12990), .ZN(n12991) );
  OAI21_X1 U15213 ( .B1(n7037), .B2(n13081), .A(n12991), .ZN(n12992) );
  AOI21_X1 U15214 ( .B1(n13119), .B2(n14611), .A(n12992), .ZN(n12993) );
  OAI21_X1 U15215 ( .B1(n12994), .B2(n14582), .A(n12993), .ZN(P3_U3211) );
  OR2_X1 U15216 ( .A1(n12995), .A2(n12996), .ZN(n13013) );
  NAND2_X1 U15217 ( .A1(n13013), .A2(n12997), .ZN(n12998) );
  XOR2_X1 U15218 ( .A(n12998), .B(n13001), .Z(n12999) );
  OAI222_X1 U15219 ( .A1(n15195), .A2(n13030), .B1(n15193), .B2(n7036), .C1(
        n15191), .C2(n12999), .ZN(n13122) );
  INV_X1 U15220 ( .A(n13122), .ZN(n13006) );
  XOR2_X1 U15221 ( .A(n13001), .B(n13000), .Z(n13123) );
  AOI22_X1 U15222 ( .A1(n14582), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15178), 
        .B2(n13002), .ZN(n13003) );
  OAI21_X1 U15223 ( .B1(n13187), .B2(n13081), .A(n13003), .ZN(n13004) );
  AOI21_X1 U15224 ( .B1(n13123), .B2(n14611), .A(n13004), .ZN(n13005) );
  OAI21_X1 U15225 ( .B1(n13006), .B2(n14582), .A(n13005), .ZN(P3_U3212) );
  OR2_X1 U15226 ( .A1(n12995), .A2(n13054), .ZN(n13008) );
  NAND2_X1 U15227 ( .A1(n13040), .A2(n13009), .ZN(n13011) );
  AND2_X1 U15228 ( .A1(n13011), .A2(n13010), .ZN(n13015) );
  AND2_X1 U15229 ( .A1(n13013), .A2(n13012), .ZN(n13014) );
  OAI211_X1 U15230 ( .C1(n13015), .C2(n12474), .A(n15149), .B(n13014), .ZN(
        n13018) );
  AOI22_X1 U15231 ( .A1(n6752), .A2(n15154), .B1(n15155), .B2(n13016), .ZN(
        n13017) );
  NAND2_X1 U15232 ( .A1(n13018), .A2(n13017), .ZN(n13126) );
  AOI21_X1 U15233 ( .B1(n15178), .B2(n13019), .A(n13126), .ZN(n13026) );
  AOI22_X1 U15234 ( .A1(n13020), .A2(n14583), .B1(P3_REG2_REG_20__SCAN_IN), 
        .B2(n14582), .ZN(n13025) );
  INV_X1 U15235 ( .A(n13021), .ZN(n13022) );
  AOI21_X1 U15236 ( .B1(n12474), .B2(n13023), .A(n13022), .ZN(n13127) );
  NAND2_X1 U15237 ( .A1(n13127), .A2(n14611), .ZN(n13024) );
  OAI211_X1 U15238 ( .C1(n13026), .C2(n14582), .A(n13025), .B(n13024), .ZN(
        P3_U3213) );
  NAND2_X1 U15239 ( .A1(n13040), .A2(n13048), .ZN(n13039) );
  NAND2_X1 U15240 ( .A1(n13039), .A2(n13027), .ZN(n13028) );
  XOR2_X1 U15241 ( .A(n13031), .B(n13028), .Z(n13029) );
  OAI222_X1 U15242 ( .A1(n15195), .A2(n13053), .B1(n15193), .B2(n13030), .C1(
        n15191), .C2(n13029), .ZN(n13130) );
  INV_X1 U15243 ( .A(n13130), .ZN(n13038) );
  OAI21_X1 U15244 ( .B1(n13033), .B2(n6800), .A(n13032), .ZN(n13131) );
  AOI22_X1 U15245 ( .A1(n14582), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15178), 
        .B2(n13034), .ZN(n13035) );
  OAI21_X1 U15246 ( .B1(n13193), .B2(n13081), .A(n13035), .ZN(n13036) );
  AOI21_X1 U15247 ( .B1(n13131), .B2(n14611), .A(n13036), .ZN(n13037) );
  OAI21_X1 U15248 ( .B1(n13038), .B2(n14582), .A(n13037), .ZN(P3_U3214) );
  OAI21_X1 U15249 ( .B1(n13040), .B2(n13048), .A(n13039), .ZN(n13044) );
  OAI22_X1 U15250 ( .A1(n13042), .A2(n15193), .B1(n13041), .B2(n15195), .ZN(
        n13043) );
  AOI21_X1 U15251 ( .B1(n13044), .B2(n15149), .A(n13043), .ZN(n13140) );
  INV_X1 U15252 ( .A(n13045), .ZN(n13046) );
  OAI22_X1 U15253 ( .A1(n15198), .A2(n12852), .B1(n13046), .B2(n15184), .ZN(
        n13047) );
  AOI21_X1 U15254 ( .B1(n13136), .B2(n14583), .A(n13047), .ZN(n13051) );
  NAND2_X1 U15255 ( .A1(n13049), .A2(n13048), .ZN(n13134) );
  NAND3_X1 U15256 ( .A1(n13135), .A2(n13134), .A3(n14611), .ZN(n13050) );
  OAI211_X1 U15257 ( .C1(n13140), .C2(n14582), .A(n13051), .B(n13050), .ZN(
        P3_U3215) );
  XNOR2_X1 U15258 ( .A(n12995), .B(n13054), .ZN(n13052) );
  OAI222_X1 U15259 ( .A1(n15193), .A2(n13053), .B1(n15195), .B2(n13076), .C1(
        n15191), .C2(n13052), .ZN(n13143) );
  INV_X1 U15260 ( .A(n13143), .ZN(n13060) );
  XNOR2_X1 U15261 ( .A(n13055), .B(n13054), .ZN(n13144) );
  AOI22_X1 U15262 ( .A1(n14582), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15178), 
        .B2(n13056), .ZN(n13057) );
  OAI21_X1 U15263 ( .B1(n13199), .B2(n13081), .A(n13057), .ZN(n13058) );
  AOI21_X1 U15264 ( .B1(n13144), .B2(n14611), .A(n13058), .ZN(n13059) );
  OAI21_X1 U15265 ( .B1(n13060), .B2(n14582), .A(n13059), .ZN(P3_U3216) );
  XNOR2_X1 U15266 ( .A(n13061), .B(n13066), .ZN(n13064) );
  AOI222_X1 U15267 ( .A1(n15149), .A2(n13064), .B1(n13063), .B2(n15155), .C1(
        n13062), .C2(n15154), .ZN(n13150) );
  OAI21_X1 U15268 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(n13148) );
  AOI22_X1 U15269 ( .A1(n14582), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15178), 
        .B2(n13068), .ZN(n13069) );
  OAI21_X1 U15270 ( .B1(n13070), .B2(n13081), .A(n13069), .ZN(n13071) );
  AOI21_X1 U15271 ( .B1(n13148), .B2(n14611), .A(n13071), .ZN(n13072) );
  OAI21_X1 U15272 ( .B1(n13150), .B2(n14582), .A(n13072), .ZN(P3_U3217) );
  XOR2_X1 U15273 ( .A(n13073), .B(n13077), .Z(n13074) );
  OAI222_X1 U15274 ( .A1(n15193), .A2(n13076), .B1(n15195), .B2(n13075), .C1(
        n13074), .C2(n15191), .ZN(n13151) );
  INV_X1 U15275 ( .A(n13151), .ZN(n13084) );
  XNOR2_X1 U15276 ( .A(n13078), .B(n13077), .ZN(n13152) );
  AOI22_X1 U15277 ( .A1(n14582), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15178), 
        .B2(n13079), .ZN(n13080) );
  OAI21_X1 U15278 ( .B1(n13204), .B2(n13081), .A(n13080), .ZN(n13082) );
  AOI21_X1 U15279 ( .B1(n13152), .B2(n14611), .A(n13082), .ZN(n13083) );
  OAI21_X1 U15280 ( .B1(n13084), .B2(n14582), .A(n13083), .ZN(P3_U3218) );
  INV_X1 U15281 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13085) );
  NOR2_X1 U15282 ( .A1(n15235), .A2(n13085), .ZN(n13086) );
  AOI21_X1 U15283 ( .B1(n14616), .B2(n15235), .A(n13086), .ZN(n13087) );
  OAI21_X1 U15284 ( .B1(n13167), .B2(n13163), .A(n13087), .ZN(P3_U3490) );
  MUX2_X1 U15285 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n13168), .S(n15235), .Z(
        P3_U3488) );
  OAI21_X1 U15286 ( .B1(n13112), .B2(n13092), .A(n13091), .ZN(n13169) );
  OAI21_X1 U15287 ( .B1(n13170), .B2(n13163), .A(n13093), .ZN(P3_U3487) );
  OAI22_X1 U15288 ( .A1(n13095), .A2(n13112), .B1(n13094), .B2(n15183), .ZN(
        n13096) );
  OR2_X1 U15289 ( .A1(n13097), .A2(n13096), .ZN(n13171) );
  MUX2_X1 U15290 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13171), .S(n15235), .Z(
        P3_U3486) );
  INV_X1 U15291 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13101) );
  INV_X1 U15292 ( .A(n13098), .ZN(n15217) );
  AOI21_X1 U15293 ( .B1(n15217), .B2(n13100), .A(n13099), .ZN(n13172) );
  MUX2_X1 U15294 ( .A(n13101), .B(n13172), .S(n15235), .Z(n13102) );
  OAI21_X1 U15295 ( .B1(n13175), .B2(n13163), .A(n13102), .ZN(P3_U3485) );
  NAND2_X1 U15296 ( .A1(n13103), .A2(n15210), .ZN(n13104) );
  OAI211_X1 U15297 ( .C1(n13112), .C2(n13106), .A(n13105), .B(n13104), .ZN(
        n13176) );
  MUX2_X1 U15298 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13176), .S(n15235), .Z(
        P3_U3484) );
  AOI22_X1 U15299 ( .A1(n13108), .A2(n15221), .B1(n15210), .B2(n13107), .ZN(
        n13109) );
  NAND2_X1 U15300 ( .A1(n13110), .A2(n13109), .ZN(n13177) );
  MUX2_X1 U15301 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13177), .S(n15235), .Z(
        P3_U3483) );
  INV_X1 U15302 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13116) );
  OAI22_X1 U15303 ( .A1(n13113), .A2(n13112), .B1(n13111), .B2(n15183), .ZN(
        n13114) );
  NOR2_X1 U15304 ( .A1(n13115), .A2(n13114), .ZN(n13178) );
  MUX2_X1 U15305 ( .A(n13116), .B(n13178), .S(n15235), .Z(n13117) );
  INV_X1 U15306 ( .A(n13117), .ZN(P3_U3482) );
  INV_X1 U15307 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13120) );
  AOI21_X1 U15308 ( .B1(n15221), .B2(n13119), .A(n13118), .ZN(n13181) );
  MUX2_X1 U15309 ( .A(n13120), .B(n13181), .S(n15235), .Z(n13121) );
  OAI21_X1 U15310 ( .B1(n7037), .B2(n13163), .A(n13121), .ZN(P3_U3481) );
  INV_X1 U15311 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13124) );
  AOI21_X1 U15312 ( .B1(n13123), .B2(n15221), .A(n13122), .ZN(n13184) );
  MUX2_X1 U15313 ( .A(n13124), .B(n13184), .S(n15235), .Z(n13125) );
  OAI21_X1 U15314 ( .B1(n13187), .B2(n13163), .A(n13125), .ZN(P3_U3480) );
  INV_X1 U15315 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13128) );
  AOI21_X1 U15316 ( .B1(n13127), .B2(n15221), .A(n13126), .ZN(n13188) );
  MUX2_X1 U15317 ( .A(n13128), .B(n13188), .S(n15235), .Z(n13129) );
  OAI21_X1 U15318 ( .B1(n13190), .B2(n13163), .A(n13129), .ZN(P3_U3479) );
  INV_X1 U15319 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13132) );
  AOI21_X1 U15320 ( .B1(n15221), .B2(n13131), .A(n13130), .ZN(n13191) );
  MUX2_X1 U15321 ( .A(n13132), .B(n13191), .S(n15235), .Z(n13133) );
  OAI21_X1 U15322 ( .B1(n13163), .B2(n13193), .A(n13133), .ZN(P3_U3478) );
  NAND3_X1 U15323 ( .A1(n13135), .A2(n13134), .A3(n15221), .ZN(n13138) );
  NAND2_X1 U15324 ( .A1(n13136), .A2(n15210), .ZN(n13137) );
  AND2_X1 U15325 ( .A1(n13138), .A2(n13137), .ZN(n13139) );
  AND2_X1 U15326 ( .A1(n13140), .A2(n13139), .ZN(n13194) );
  MUX2_X1 U15327 ( .A(n13141), .B(n13194), .S(n15235), .Z(n13142) );
  INV_X1 U15328 ( .A(n13142), .ZN(P3_U3477) );
  INV_X1 U15329 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13145) );
  AOI21_X1 U15330 ( .B1(n13144), .B2(n15221), .A(n13143), .ZN(n13196) );
  MUX2_X1 U15331 ( .A(n13145), .B(n13196), .S(n15235), .Z(n13146) );
  OAI21_X1 U15332 ( .B1(n13199), .B2(n13163), .A(n13146), .ZN(P3_U3476) );
  AOI22_X1 U15333 ( .A1(n13148), .A2(n15221), .B1(n15210), .B2(n13147), .ZN(
        n13149) );
  NAND2_X1 U15334 ( .A1(n13150), .A2(n13149), .ZN(n13200) );
  MUX2_X1 U15335 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13200), .S(n15235), .Z(
        P3_U3475) );
  INV_X1 U15336 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13153) );
  AOI21_X1 U15337 ( .B1(n13152), .B2(n15221), .A(n13151), .ZN(n13201) );
  MUX2_X1 U15338 ( .A(n13153), .B(n13201), .S(n15235), .Z(n13154) );
  OAI21_X1 U15339 ( .B1(n13204), .B2(n13163), .A(n13154), .ZN(P3_U3474) );
  AOI21_X1 U15340 ( .B1(n15221), .B2(n13156), .A(n13155), .ZN(n13205) );
  MUX2_X1 U15341 ( .A(n13157), .B(n13205), .S(n15235), .Z(n13158) );
  OAI21_X1 U15342 ( .B1(n13208), .B2(n13163), .A(n13158), .ZN(P3_U3473) );
  INV_X1 U15343 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13161) );
  AOI21_X1 U15344 ( .B1(n13160), .B2(n15221), .A(n13159), .ZN(n13209) );
  MUX2_X1 U15345 ( .A(n13161), .B(n13209), .S(n15235), .Z(n13162) );
  OAI21_X1 U15346 ( .B1(n13163), .B2(n13211), .A(n13162), .ZN(P3_U3472) );
  INV_X1 U15347 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13164) );
  NOR2_X1 U15348 ( .A1(n15225), .A2(n13164), .ZN(n13165) );
  AOI21_X1 U15349 ( .B1(n14616), .B2(n15225), .A(n13165), .ZN(n13166) );
  OAI21_X1 U15350 ( .B1(n13167), .B2(n13212), .A(n13166), .ZN(P3_U3458) );
  MUX2_X1 U15351 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n13168), .S(n15225), .Z(
        P3_U3456) );
  MUX2_X1 U15352 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13171), .S(n15225), .Z(
        P3_U3454) );
  INV_X1 U15353 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13173) );
  MUX2_X1 U15354 ( .A(n13173), .B(n13172), .S(n15225), .Z(n13174) );
  OAI21_X1 U15355 ( .B1(n13175), .B2(n13212), .A(n13174), .ZN(P3_U3453) );
  MUX2_X1 U15356 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13176), .S(n15225), .Z(
        P3_U3452) );
  MUX2_X1 U15357 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13177), .S(n15225), .Z(
        P3_U3451) );
  INV_X1 U15358 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13179) );
  MUX2_X1 U15359 ( .A(n13179), .B(n13178), .S(n15225), .Z(n13180) );
  INV_X1 U15360 ( .A(n13180), .ZN(P3_U3450) );
  INV_X1 U15361 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13182) );
  MUX2_X1 U15362 ( .A(n13182), .B(n13181), .S(n15225), .Z(n13183) );
  OAI21_X1 U15363 ( .B1(n7037), .B2(n13212), .A(n13183), .ZN(P3_U3449) );
  INV_X1 U15364 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13185) );
  MUX2_X1 U15365 ( .A(n13185), .B(n13184), .S(n15225), .Z(n13186) );
  OAI21_X1 U15366 ( .B1(n13187), .B2(n13212), .A(n13186), .ZN(P3_U3448) );
  INV_X1 U15367 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n15431) );
  MUX2_X1 U15368 ( .A(n15431), .B(n13188), .S(n15225), .Z(n13189) );
  OAI21_X1 U15369 ( .B1(n13190), .B2(n13212), .A(n13189), .ZN(P3_U3447) );
  INV_X1 U15370 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n15460) );
  MUX2_X1 U15371 ( .A(n15460), .B(n13191), .S(n15225), .Z(n13192) );
  OAI21_X1 U15372 ( .B1(n13212), .B2(n13193), .A(n13192), .ZN(P3_U3446) );
  INV_X1 U15373 ( .A(n13194), .ZN(n13195) );
  MUX2_X1 U15374 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13195), .S(n15225), .Z(
        P3_U3444) );
  INV_X1 U15375 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13197) );
  MUX2_X1 U15376 ( .A(n13197), .B(n13196), .S(n15225), .Z(n13198) );
  OAI21_X1 U15377 ( .B1(n13199), .B2(n13212), .A(n13198), .ZN(P3_U3441) );
  MUX2_X1 U15378 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13200), .S(n15225), .Z(
        P3_U3438) );
  INV_X1 U15379 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13202) );
  MUX2_X1 U15380 ( .A(n13202), .B(n13201), .S(n15225), .Z(n13203) );
  OAI21_X1 U15381 ( .B1(n13204), .B2(n13212), .A(n13203), .ZN(P3_U3435) );
  INV_X1 U15382 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13206) );
  MUX2_X1 U15383 ( .A(n13206), .B(n13205), .S(n15225), .Z(n13207) );
  OAI21_X1 U15384 ( .B1(n13208), .B2(n13212), .A(n13207), .ZN(P3_U3432) );
  INV_X1 U15385 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15433) );
  MUX2_X1 U15386 ( .A(n15433), .B(n13209), .S(n15225), .Z(n13210) );
  OAI21_X1 U15387 ( .B1(n13212), .B2(n13211), .A(n13210), .ZN(P3_U3429) );
  MUX2_X1 U15388 ( .A(n13214), .B(P3_D_REG_1__SCAN_IN), .S(n13213), .Z(
        P3_U3377) );
  MUX2_X1 U15389 ( .A(P3_D_REG_0__SCAN_IN), .B(n13216), .S(n13215), .Z(
        P3_U3376) );
  INV_X1 U15390 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13217) );
  NAND3_X1 U15391 ( .A1(n13217), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13219) );
  OAI22_X1 U15392 ( .A1(n7597), .A2(n13219), .B1(n13218), .B2(n13228), .ZN(
        n13220) );
  AOI21_X1 U15393 ( .B1(n13222), .B2(n13221), .A(n13220), .ZN(n13223) );
  INV_X1 U15394 ( .A(n13223), .ZN(P3_U3264) );
  INV_X1 U15395 ( .A(n13224), .ZN(n13226) );
  OAI222_X1 U15396 ( .A1(n13228), .A2(n15505), .B1(n13227), .B2(n13226), .C1(
        P3_U3151), .C2(n13225), .ZN(P3_U3266) );
  OAI22_X1 U15397 ( .A1(n14933), .A2(n13517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13232), .ZN(n13234) );
  OAI22_X1 U15398 ( .A1(n14932), .A2(n13519), .B1(n14947), .B2(n13551), .ZN(
        n13233) );
  AOI211_X1 U15399 ( .C1(n13717), .C2(n14943), .A(n13234), .B(n13233), .ZN(
        n13235) );
  XOR2_X1 U15400 ( .A(n13237), .B(n13236), .Z(n13242) );
  AOI22_X1 U15401 ( .A1(n13514), .A2(n13667), .B1(n13585), .B2(n13665), .ZN(
        n13615) );
  NOR2_X1 U15402 ( .A1(n13615), .A2(n13238), .ZN(n13240) );
  INV_X1 U15403 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n15367) );
  OAI22_X1 U15404 ( .A1(n13621), .A2(n14947), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15367), .ZN(n13239) );
  AOI211_X1 U15405 ( .C1(n7056), .C2(n14943), .A(n13240), .B(n13239), .ZN(
        n13241) );
  OAI21_X1 U15406 ( .B1(n13242), .B2(n14939), .A(n13241), .ZN(P2_U3188) );
  NAND2_X1 U15407 ( .A1(n6732), .A2(n13243), .ZN(n13244) );
  XNOR2_X1 U15408 ( .A(n13245), .B(n13244), .ZN(n13249) );
  OAI22_X1 U15409 ( .A1(n13513), .A2(n15039), .B1(n13477), .B2(n13595), .ZN(
        n13682) );
  AOI22_X1 U15410 ( .A1(n13682), .A2(n13285), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13246) );
  OAI21_X1 U15411 ( .B1(n13687), .B2(n14947), .A(n13246), .ZN(n13247) );
  AOI21_X1 U15412 ( .B1(n13757), .B2(n14943), .A(n13247), .ZN(n13248) );
  OAI21_X1 U15413 ( .B1(n13249), .B2(n14939), .A(n13248), .ZN(P2_U3191) );
  OAI22_X1 U15414 ( .A1(n13250), .A2(n15039), .B1(n13513), .B2(n13595), .ZN(
        n13648) );
  AOI22_X1 U15415 ( .A1(n13648), .A2(n13285), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13251) );
  OAI21_X1 U15416 ( .B1(n13652), .B2(n14947), .A(n13251), .ZN(n13256) );
  AOI211_X1 U15417 ( .C1(n13254), .C2(n13253), .A(n14939), .B(n13252), .ZN(
        n13255) );
  AOI211_X1 U15418 ( .C1(n13747), .C2(n14943), .A(n13256), .B(n13255), .ZN(
        n13257) );
  INV_X1 U15419 ( .A(n13257), .ZN(P2_U3195) );
  OAI21_X1 U15420 ( .B1(n13260), .B2(n13258), .A(n13259), .ZN(n13261) );
  NAND2_X1 U15421 ( .A1(n13261), .A2(n7445), .ZN(n13268) );
  AOI22_X1 U15422 ( .A1(n13294), .A2(n13320), .B1(n13262), .B2(n13318), .ZN(
        n13267) );
  INV_X1 U15423 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n15480) );
  NOR2_X1 U15424 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15480), .ZN(n13361) );
  NOR2_X1 U15425 ( .A1(n13297), .A2(n15084), .ZN(n13263) );
  AOI211_X1 U15426 ( .C1(n13265), .C2(n13264), .A(n13361), .B(n13263), .ZN(
        n13266) );
  NAND3_X1 U15427 ( .A1(n13268), .A2(n13267), .A3(n13266), .ZN(P2_U3199) );
  NOR2_X1 U15428 ( .A1(n13269), .A2(n6722), .ZN(n13270) );
  XNOR2_X1 U15429 ( .A(n13271), .B(n13270), .ZN(n13277) );
  INV_X1 U15430 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13272) );
  OAI22_X1 U15431 ( .A1(n13480), .A2(n14932), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13272), .ZN(n13275) );
  INV_X1 U15432 ( .A(n13674), .ZN(n13273) );
  OAI22_X1 U15433 ( .A1(n13507), .A2(n14933), .B1(n13273), .B2(n14947), .ZN(
        n13274) );
  AOI211_X1 U15434 ( .C1(n13752), .C2(n14943), .A(n13275), .B(n13274), .ZN(
        n13276) );
  OAI21_X1 U15435 ( .B1(n13277), .B2(n14939), .A(n13276), .ZN(P2_U3205) );
  OAI21_X1 U15436 ( .B1(n13280), .B2(n13279), .A(n13278), .ZN(n13281) );
  NAND2_X1 U15437 ( .A1(n13281), .A2(n7445), .ZN(n13287) );
  OAI22_X1 U15438 ( .A1(n13596), .A2(n15039), .B1(n13480), .B2(n13595), .ZN(
        n13632) );
  OAI22_X1 U15439 ( .A1(n13283), .A2(n14947), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13282), .ZN(n13284) );
  AOI21_X1 U15440 ( .B1(n13632), .B2(n13285), .A(n13284), .ZN(n13286) );
  OAI211_X1 U15441 ( .C1(n13741), .C2(n13297), .A(n13287), .B(n13286), .ZN(
        P2_U3207) );
  AOI211_X1 U15442 ( .C1(n13290), .C2(n13289), .A(n14939), .B(n13288), .ZN(
        n13291) );
  INV_X1 U15443 ( .A(n13291), .ZN(n13296) );
  AND2_X1 U15444 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13435) );
  OAI22_X1 U15445 ( .A1(n13507), .A2(n14932), .B1(n13292), .B2(n14947), .ZN(
        n13293) );
  AOI211_X1 U15446 ( .C1(n13294), .C2(n13308), .A(n13435), .B(n13293), .ZN(
        n13295) );
  OAI211_X1 U15447 ( .C1(n13478), .C2(n13297), .A(n13296), .B(n13295), .ZN(
        P2_U3210) );
  INV_X1 U15448 ( .A(n13299), .ZN(n13300) );
  AOI21_X1 U15449 ( .B1(n13301), .B2(n13298), .A(n13300), .ZN(n13306) );
  OAI22_X1 U15450 ( .A1(n14933), .A2(n13594), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13302), .ZN(n13304) );
  OAI22_X1 U15451 ( .A1(n14932), .A2(n13490), .B1(n14947), .B2(n13563), .ZN(
        n13303) );
  AOI211_X1 U15452 ( .C1(n13722), .C2(n14943), .A(n13304), .B(n13303), .ZN(
        n13305) );
  OAI21_X1 U15453 ( .B1(n13306), .B2(n14939), .A(n13305), .ZN(P2_U3212) );
  CLKBUF_X2 U15454 ( .A(P2_U3947), .Z(n14930) );
  MUX2_X1 U15455 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13307), .S(n14930), .Z(
        P2_U3562) );
  MUX2_X1 U15456 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13493), .S(n14930), .Z(
        P2_U3561) );
  MUX2_X1 U15457 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13528), .S(n14930), .Z(
        P2_U3560) );
  MUX2_X1 U15458 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13543), .S(n14930), .Z(
        P2_U3559) );
  MUX2_X1 U15459 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13571), .S(n14930), .Z(
        P2_U3558) );
  MUX2_X1 U15460 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13586), .S(n14930), .Z(
        P2_U3557) );
  MUX2_X1 U15461 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13570), .S(n14930), .Z(
        P2_U3556) );
  MUX2_X1 U15462 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13585), .S(n14930), .Z(
        P2_U3555) );
  MUX2_X1 U15463 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13483), .S(n14930), .Z(
        P2_U3554) );
  MUX2_X1 U15464 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13514), .S(n14930), .Z(
        P2_U3553) );
  MUX2_X1 U15465 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13666), .S(n14930), .Z(
        P2_U3552) );
  MUX2_X1 U15466 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13509), .S(n14930), .Z(
        P2_U3551) );
  MUX2_X1 U15467 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13668), .S(n14930), .Z(
        P2_U3550) );
  MUX2_X1 U15468 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13505), .S(n14930), .Z(
        P2_U3549) );
  MUX2_X1 U15469 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13308), .S(n14930), .Z(
        P2_U3548) );
  MUX2_X1 U15470 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13309), .S(n14930), .Z(
        P2_U3547) );
  MUX2_X1 U15471 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13310), .S(n14930), .Z(
        P2_U3546) );
  MUX2_X1 U15472 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13311), .S(n14930), .Z(
        P2_U3545) );
  MUX2_X1 U15473 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n7408), .S(n14930), .Z(
        P2_U3544) );
  MUX2_X1 U15474 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13312), .S(n14930), .Z(
        P2_U3543) );
  MUX2_X1 U15475 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13313), .S(n14930), .Z(
        P2_U3542) );
  MUX2_X1 U15476 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13314), .S(n14930), .Z(
        P2_U3541) );
  MUX2_X1 U15477 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13315), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15478 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13316), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15479 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13317), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15480 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13318), .S(n14930), .Z(
        P2_U3537) );
  MUX2_X1 U15481 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13319), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U15482 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13320), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15483 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13321), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15484 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13322), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U15485 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12147), .S(P2_U3947), .Z(
        P2_U3532) );
  MUX2_X1 U15486 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n12144), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI22_X1 U15487 ( .A1(n14996), .A2(n13325), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13323), .ZN(n13324) );
  AOI21_X1 U15488 ( .B1(n14949), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n13324), .ZN(
        n13335) );
  INV_X1 U15489 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13327) );
  MUX2_X1 U15490 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9493), .S(n13325), .Z(
        n13326) );
  OAI21_X1 U15491 ( .B1(n15047), .B2(n13327), .A(n13326), .ZN(n13328) );
  NAND3_X1 U15492 ( .A1(n15027), .A2(n13329), .A3(n13328), .ZN(n13334) );
  OAI211_X1 U15493 ( .C1(n13332), .C2(n13331), .A(n15002), .B(n13330), .ZN(
        n13333) );
  NAND3_X1 U15494 ( .A1(n13335), .A2(n13334), .A3(n13333), .ZN(P2_U3215) );
  NOR2_X1 U15495 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15314), .ZN(n13338) );
  NOR2_X1 U15496 ( .A1(n14996), .A2(n13336), .ZN(n13337) );
  AOI211_X1 U15497 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n14949), .A(n13338), .B(
        n13337), .ZN(n13346) );
  OAI211_X1 U15498 ( .C1(n13341), .C2(n13340), .A(n15002), .B(n13339), .ZN(
        n13345) );
  OAI211_X1 U15499 ( .C1(n13343), .C2(n13342), .A(n15027), .B(n13355), .ZN(
        n13344) );
  NAND3_X1 U15500 ( .A1(n13346), .A2(n13345), .A3(n13344), .ZN(P2_U3217) );
  NOR2_X1 U15501 ( .A1(n14996), .A2(n13352), .ZN(n13347) );
  AOI211_X1 U15502 ( .C1(n14949), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n13348), .B(
        n13347), .ZN(n13359) );
  OAI211_X1 U15503 ( .C1(n13351), .C2(n13350), .A(n15002), .B(n13349), .ZN(
        n13358) );
  MUX2_X1 U15504 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9821), .S(n13352), .Z(
        n13353) );
  NAND3_X1 U15505 ( .A1(n13355), .A2(n13354), .A3(n13353), .ZN(n13356) );
  NAND3_X1 U15506 ( .A1(n15027), .A2(n13368), .A3(n13356), .ZN(n13357) );
  NAND3_X1 U15507 ( .A1(n13359), .A2(n13358), .A3(n13357), .ZN(P2_U3218) );
  NOR2_X1 U15508 ( .A1(n14996), .A2(n13365), .ZN(n13360) );
  AOI211_X1 U15509 ( .C1(n14949), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n13361), .B(
        n13360), .ZN(n13373) );
  OAI211_X1 U15510 ( .C1(n13364), .C2(n13363), .A(n15002), .B(n13362), .ZN(
        n13372) );
  MUX2_X1 U15511 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9025), .S(n13365), .Z(
        n13366) );
  NAND3_X1 U15512 ( .A1(n13368), .A2(n13367), .A3(n13366), .ZN(n13369) );
  NAND3_X1 U15513 ( .A1(n15027), .A2(n13370), .A3(n13369), .ZN(n13371) );
  NAND3_X1 U15514 ( .A1(n13373), .A2(n13372), .A3(n13371), .ZN(P2_U3219) );
  NOR2_X1 U15515 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8561), .ZN(n13376) );
  NOR2_X1 U15516 ( .A1(n14996), .A2(n13374), .ZN(n13375) );
  AOI211_X1 U15517 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n14949), .A(n13376), .B(
        n13375), .ZN(n13386) );
  OAI211_X1 U15518 ( .C1(n13379), .C2(n13378), .A(n15002), .B(n13377), .ZN(
        n13385) );
  MUX2_X1 U15519 ( .A(n9539), .B(P2_REG2_REG_7__SCAN_IN), .S(n13380), .Z(
        n13381) );
  NAND3_X1 U15520 ( .A1(n14969), .A2(n13382), .A3(n13381), .ZN(n13383) );
  NAND3_X1 U15521 ( .A1(n15027), .A2(n13397), .A3(n13383), .ZN(n13384) );
  NAND3_X1 U15522 ( .A1(n13386), .A2(n13385), .A3(n13384), .ZN(P2_U3221) );
  INV_X1 U15523 ( .A(n13387), .ZN(n13390) );
  NOR2_X1 U15524 ( .A1(n14996), .A2(n13388), .ZN(n13389) );
  AOI211_X1 U15525 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n14949), .A(n13390), .B(
        n13389), .ZN(n13402) );
  OAI211_X1 U15526 ( .C1(n13393), .C2(n13392), .A(n13391), .B(n15002), .ZN(
        n13401) );
  MUX2_X1 U15527 ( .A(n9807), .B(P2_REG2_REG_8__SCAN_IN), .S(n13394), .Z(
        n13395) );
  NAND3_X1 U15528 ( .A1(n13397), .A2(n13396), .A3(n13395), .ZN(n13398) );
  NAND3_X1 U15529 ( .A1(n15027), .A2(n13399), .A3(n13398), .ZN(n13400) );
  NAND3_X1 U15530 ( .A1(n13402), .A2(n13401), .A3(n13400), .ZN(P2_U3222) );
  AOI21_X1 U15531 ( .B1(n13404), .B2(n13403), .A(n15018), .ZN(n13406) );
  NAND2_X1 U15532 ( .A1(n13406), .A2(n13405), .ZN(n13418) );
  NOR2_X1 U15533 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15436), .ZN(n13409) );
  NOR2_X1 U15534 ( .A1(n14996), .A2(n13407), .ZN(n13408) );
  AOI211_X1 U15535 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n14949), .A(n13409), 
        .B(n13408), .ZN(n13417) );
  INV_X1 U15536 ( .A(n13410), .ZN(n13415) );
  MUX2_X1 U15537 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n13412), .S(n13411), .Z(
        n13414) );
  OAI211_X1 U15538 ( .C1(n13415), .C2(n13414), .A(n15027), .B(n13413), .ZN(
        n13416) );
  NAND3_X1 U15539 ( .A1(n13418), .A2(n13417), .A3(n13416), .ZN(P2_U3224) );
  INV_X1 U15540 ( .A(n13419), .ZN(n13422) );
  INV_X1 U15541 ( .A(n13420), .ZN(n13421) );
  OAI211_X1 U15542 ( .C1(n13422), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15002), 
        .B(n13421), .ZN(n13431) );
  NOR2_X1 U15543 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13423), .ZN(n13426) );
  NOR2_X1 U15544 ( .A1(n14996), .A2(n13424), .ZN(n13425) );
  AOI211_X1 U15545 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14949), .A(n13426), 
        .B(n13425), .ZN(n13430) );
  OAI211_X1 U15546 ( .C1(n13428), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15027), 
        .B(n13427), .ZN(n13429) );
  NAND3_X1 U15547 ( .A1(n13431), .A2(n13430), .A3(n13429), .ZN(P2_U3229) );
  OAI21_X1 U15548 ( .B1(n13433), .B2(n11053), .A(n13432), .ZN(n13450) );
  XOR2_X1 U15549 ( .A(n13450), .B(n13445), .Z(n13434) );
  NOR2_X1 U15550 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13434), .ZN(n13453) );
  AOI21_X1 U15551 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13434), .A(n13453), 
        .ZN(n13444) );
  INV_X1 U15552 ( .A(n13435), .ZN(n13436) );
  OAI21_X1 U15553 ( .B1(n14996), .B2(n13445), .A(n13436), .ZN(n13442) );
  AOI21_X1 U15554 ( .B1(n13438), .B2(P2_REG1_REG_17__SCAN_IN), .A(n13437), 
        .ZN(n13446) );
  XNOR2_X1 U15555 ( .A(n13445), .B(n13446), .ZN(n13440) );
  INV_X1 U15556 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13439) );
  NOR2_X1 U15557 ( .A1(n13439), .A2(n13440), .ZN(n13448) );
  AOI211_X1 U15558 ( .C1(n13440), .C2(n13439), .A(n13448), .B(n15018), .ZN(
        n13441) );
  AOI211_X1 U15559 ( .C1(n14949), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13442), 
        .B(n13441), .ZN(n13443) );
  OAI21_X1 U15560 ( .B1(n13444), .B2(n14998), .A(n13443), .ZN(P2_U3232) );
  INV_X1 U15561 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n15349) );
  NOR2_X1 U15562 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  NOR2_X1 U15563 ( .A1(n13448), .A2(n13447), .ZN(n13449) );
  INV_X1 U15564 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15350) );
  XOR2_X1 U15565 ( .A(n13449), .B(n15350), .Z(n13458) );
  INV_X1 U15566 ( .A(n13458), .ZN(n13456) );
  NOR2_X1 U15567 ( .A1(n13451), .A2(n13450), .ZN(n13452) );
  NOR2_X1 U15568 ( .A1(n13453), .A2(n13452), .ZN(n13454) );
  XOR2_X1 U15569 ( .A(n13454), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13457) );
  OAI21_X1 U15570 ( .B1(n13457), .B2(n14998), .A(n14996), .ZN(n13455) );
  AOI21_X1 U15571 ( .B1(n13456), .B2(n15002), .A(n13455), .ZN(n13461) );
  AOI22_X1 U15572 ( .A1(n13458), .A2(n15002), .B1(n15027), .B2(n13457), .ZN(
        n13460) );
  MUX2_X1 U15573 ( .A(n13461), .B(n13460), .S(n13459), .Z(n13463) );
  NAND2_X1 U15574 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n13462)
         );
  OAI211_X1 U15575 ( .C1(n15349), .C2(n15032), .A(n13463), .B(n13462), .ZN(
        P2_U3233) );
  INV_X1 U15576 ( .A(n13722), .ZN(n13566) );
  OR2_X2 U15577 ( .A1(n13717), .A2(n13561), .ZN(n13548) );
  XNOR2_X1 U15578 ( .A(n13470), .B(n12364), .ZN(n13464) );
  NAND2_X1 U15579 ( .A1(n13464), .A2(n6577), .ZN(n13700) );
  OAI21_X1 U15580 ( .B1(n9010), .B2(n13465), .A(n13665), .ZN(n13494) );
  OR2_X1 U15581 ( .A1(n13466), .A2(n13494), .ZN(n13702) );
  NOR2_X1 U15582 ( .A1(n6578), .A2(n13702), .ZN(n13474) );
  INV_X1 U15583 ( .A(n12364), .ZN(n13701) );
  NOR2_X1 U15584 ( .A1(n13701), .A2(n13677), .ZN(n13467) );
  AOI211_X1 U15585 ( .C1(n6578), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13474), .B(
        n13467), .ZN(n13468) );
  OAI21_X1 U15586 ( .B1(n13700), .B2(n13639), .A(n13468), .ZN(P2_U3234) );
  INV_X1 U15587 ( .A(n13498), .ZN(n13472) );
  OAI211_X1 U15588 ( .C1(n13704), .C2(n13472), .A(n13471), .B(n6577), .ZN(
        n13703) );
  NOR2_X1 U15589 ( .A1(n13704), .A2(n13677), .ZN(n13473) );
  AOI211_X1 U15590 ( .C1(n6578), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13474), .B(
        n13473), .ZN(n13475) );
  OAI21_X1 U15591 ( .B1(n13639), .B2(n13703), .A(n13475), .ZN(P2_U3235) );
  NAND2_X1 U15592 ( .A1(n13663), .A2(n13664), .ZN(n13662) );
  NAND2_X1 U15593 ( .A1(n13655), .A2(n13666), .ZN(n13481) );
  NAND2_X1 U15594 ( .A1(n13631), .A2(n13636), .ZN(n13630) );
  NAND2_X1 U15595 ( .A1(n7056), .A2(n13596), .ZN(n13484) );
  INV_X1 U15596 ( .A(n13598), .ZN(n13593) );
  INV_X1 U15597 ( .A(n13487), .ZN(n13569) );
  NAND2_X1 U15598 ( .A1(n13717), .A2(n13490), .ZN(n13527) );
  INV_X1 U15599 ( .A(n13493), .ZN(n13495) );
  OAI22_X1 U15600 ( .A1(n13519), .A2(n13595), .B1(n13495), .B2(n13494), .ZN(
        n13496) );
  AOI21_X1 U15601 ( .B1(n13706), .B2(n13534), .A(n8705), .ZN(n13499) );
  OAI22_X1 U15602 ( .A1(n15045), .A2(n13501), .B1(n13500), .B2(n15037), .ZN(
        n13503) );
  NOR2_X1 U15603 ( .A1(n7041), .A2(n13677), .ZN(n13502) );
  AOI211_X1 U15604 ( .C1(n13694), .C2(n13705), .A(n13503), .B(n13502), .ZN(
        n13524) );
  NAND2_X1 U15605 ( .A1(n13510), .A2(n13513), .ZN(n13511) );
  OAI21_X1 U15606 ( .B1(n13510), .B2(n13513), .A(n13512), .ZN(n13656) );
  INV_X1 U15607 ( .A(n13625), .ZN(n13613) );
  NOR2_X1 U15608 ( .A1(n13722), .A2(n13586), .ZN(n13518) );
  INV_X1 U15609 ( .A(n13712), .ZN(n13536) );
  XNOR2_X1 U15610 ( .A(n13521), .B(n13492), .ZN(n13709) );
  INV_X1 U15611 ( .A(n13709), .ZN(n13522) );
  NAND2_X1 U15612 ( .A1(n13522), .A2(n13644), .ZN(n13523) );
  OAI211_X1 U15613 ( .C1(n13708), .C2(n6578), .A(n13524), .B(n13523), .ZN(
        P2_U3236) );
  NAND2_X1 U15614 ( .A1(n13525), .A2(n13683), .ZN(n13531) );
  AOI21_X1 U15615 ( .B1(n13542), .B2(n13527), .A(n13526), .ZN(n13530) );
  AOI22_X1 U15616 ( .A1(n13665), .A2(n13528), .B1(n13571), .B2(n13667), .ZN(
        n13529) );
  OAI21_X1 U15617 ( .B1(n13531), .B2(n13530), .A(n13529), .ZN(n13714) );
  NOR2_X1 U15618 ( .A1(n15037), .A2(n13532), .ZN(n13533) );
  OAI21_X1 U15619 ( .B1(n13714), .B2(n13533), .A(n15045), .ZN(n13539) );
  AOI211_X1 U15620 ( .C1(n13712), .C2(n13548), .A(n8705), .B(n7042), .ZN(
        n13711) );
  OAI22_X1 U15621 ( .A1(n13536), .A2(n13677), .B1(n15045), .B2(n13535), .ZN(
        n13537) );
  AOI21_X1 U15622 ( .B1(n13711), .B2(n13694), .A(n13537), .ZN(n13538) );
  OAI211_X1 U15623 ( .C1(n13540), .C2(n13710), .A(n13539), .B(n13538), .ZN(
        P2_U3237) );
  NAND2_X1 U15624 ( .A1(n13543), .A2(n13665), .ZN(n13545) );
  AOI21_X2 U15625 ( .B1(n13547), .B2(n13683), .A(n13546), .ZN(n13719) );
  INV_X1 U15626 ( .A(n13548), .ZN(n13549) );
  AOI211_X1 U15627 ( .C1(n13717), .C2(n13561), .A(n8705), .B(n13549), .ZN(
        n13716) );
  INV_X1 U15628 ( .A(n13717), .ZN(n13550) );
  NOR2_X1 U15629 ( .A1(n13550), .A2(n13677), .ZN(n13554) );
  OAI22_X1 U15630 ( .A1(n15045), .A2(n13552), .B1(n13551), .B2(n15037), .ZN(
        n13553) );
  AOI211_X1 U15631 ( .C1(n13716), .C2(n13694), .A(n13554), .B(n13553), .ZN(
        n13559) );
  XNOR2_X1 U15632 ( .A(n13556), .B(n13555), .ZN(n13720) );
  INV_X1 U15633 ( .A(n13720), .ZN(n13557) );
  NAND2_X1 U15634 ( .A1(n13557), .A2(n13644), .ZN(n13558) );
  OAI211_X1 U15635 ( .C1(n13719), .C2(n6578), .A(n13559), .B(n13558), .ZN(
        P2_U3238) );
  XNOR2_X1 U15636 ( .A(n13560), .B(n13569), .ZN(n13725) );
  INV_X1 U15637 ( .A(n13561), .ZN(n13562) );
  AOI211_X1 U15638 ( .C1(n13722), .C2(n7057), .A(n8705), .B(n13562), .ZN(
        n13721) );
  INV_X1 U15639 ( .A(n13563), .ZN(n13564) );
  AOI22_X1 U15640 ( .A1(n6578), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13564), 
        .B2(n13673), .ZN(n13565) );
  OAI21_X1 U15641 ( .B1(n13566), .B2(n13677), .A(n13565), .ZN(n13573) );
  NOR2_X1 U15642 ( .A1(n13724), .A2(n6578), .ZN(n13572) );
  AOI211_X1 U15643 ( .C1(n13721), .C2(n13694), .A(n13573), .B(n13572), .ZN(
        n13574) );
  OAI21_X1 U15644 ( .B1(n13697), .B2(n13725), .A(n13574), .ZN(P2_U3239) );
  XOR2_X1 U15645 ( .A(n13584), .B(n13575), .Z(n13730) );
  NAND2_X1 U15646 ( .A1(n13727), .A2(n13603), .ZN(n13576) );
  NAND2_X1 U15647 ( .A1(n13576), .A2(n6577), .ZN(n13577) );
  NOR2_X1 U15648 ( .A1(n13578), .A2(n13577), .ZN(n13726) );
  INV_X1 U15649 ( .A(n13579), .ZN(n13580) );
  AOI22_X1 U15650 ( .A1(n6578), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13580), 
        .B2(n13673), .ZN(n13581) );
  OAI21_X1 U15651 ( .B1(n7054), .B2(n13677), .A(n13581), .ZN(n13589) );
  OAI21_X1 U15652 ( .B1(n13584), .B2(n13583), .A(n13582), .ZN(n13587) );
  AOI222_X1 U15653 ( .A1(n13683), .A2(n13587), .B1(n13586), .B2(n13665), .C1(
        n13585), .C2(n13667), .ZN(n13729) );
  NOR2_X1 U15654 ( .A1(n13729), .A2(n6578), .ZN(n13588) );
  OAI21_X1 U15655 ( .B1(n13697), .B2(n13730), .A(n13590), .ZN(P2_U3240) );
  OAI21_X1 U15656 ( .B1(n13593), .B2(n13592), .A(n13591), .ZN(n13602) );
  OAI22_X1 U15657 ( .A1(n13596), .A2(n13595), .B1(n13594), .B2(n15039), .ZN(
        n13601) );
  OAI21_X1 U15658 ( .B1(n13599), .B2(n13598), .A(n13597), .ZN(n13735) );
  NOR2_X1 U15659 ( .A1(n13735), .A2(n9127), .ZN(n13600) );
  INV_X1 U15660 ( .A(n13603), .ZN(n13604) );
  AOI211_X1 U15661 ( .C1(n13732), .C2(n13618), .A(n8705), .B(n13604), .ZN(
        n13731) );
  INV_X1 U15662 ( .A(n13605), .ZN(n13606) );
  AOI22_X1 U15663 ( .A1(n13606), .A2(n13673), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n6578), .ZN(n13607) );
  OAI21_X1 U15664 ( .B1(n13608), .B2(n13677), .A(n13607), .ZN(n13611) );
  NOR2_X1 U15665 ( .A1(n13735), .A2(n13609), .ZN(n13610) );
  AOI211_X1 U15666 ( .C1(n13731), .C2(n13694), .A(n13611), .B(n13610), .ZN(
        n13612) );
  OAI21_X1 U15667 ( .B1(n13734), .B2(n6578), .A(n13612), .ZN(P2_U3241) );
  XNOR2_X1 U15668 ( .A(n13614), .B(n13613), .ZN(n13617) );
  INV_X1 U15669 ( .A(n13615), .ZN(n13616) );
  AOI21_X1 U15670 ( .B1(n13617), .B2(n13683), .A(n13616), .ZN(n13738) );
  INV_X1 U15671 ( .A(n13638), .ZN(n13620) );
  INV_X1 U15672 ( .A(n13618), .ZN(n13619) );
  AOI211_X1 U15673 ( .C1(n7056), .C2(n13620), .A(n8705), .B(n13619), .ZN(
        n13736) );
  INV_X1 U15674 ( .A(n13621), .ZN(n13622) );
  AOI22_X1 U15675 ( .A1(n13622), .A2(n13673), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n6578), .ZN(n13623) );
  OAI21_X1 U15676 ( .B1(n13624), .B2(n13677), .A(n13623), .ZN(n13628) );
  XNOR2_X1 U15677 ( .A(n13626), .B(n13625), .ZN(n13739) );
  NOR2_X1 U15678 ( .A1(n13739), .A2(n13697), .ZN(n13627) );
  AOI211_X1 U15679 ( .C1(n13736), .C2(n13694), .A(n13628), .B(n13627), .ZN(
        n13629) );
  OAI21_X1 U15680 ( .B1(n6578), .B2(n13738), .A(n13629), .ZN(P2_U3242) );
  OAI211_X1 U15681 ( .C1(n13631), .C2(n13636), .A(n13630), .B(n13683), .ZN(
        n13634) );
  INV_X1 U15682 ( .A(n13632), .ZN(n13633) );
  NAND2_X1 U15683 ( .A1(n13634), .A2(n13633), .ZN(n13742) );
  INV_X1 U15684 ( .A(n13742), .ZN(n13646) );
  AOI21_X1 U15685 ( .B1(n13636), .B2(n13635), .A(n6640), .ZN(n13744) );
  OAI21_X1 U15686 ( .B1(n13741), .B2(n13650), .A(n6577), .ZN(n13637) );
  OR2_X1 U15687 ( .A1(n13638), .A2(n13637), .ZN(n13740) );
  NOR2_X1 U15688 ( .A1(n13740), .A2(n13639), .ZN(n13643) );
  AOI22_X1 U15689 ( .A1(n13640), .A2(n13673), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n6578), .ZN(n13641) );
  OAI21_X1 U15690 ( .B1(n13741), .B2(n13677), .A(n13641), .ZN(n13642) );
  AOI211_X1 U15691 ( .C1(n13744), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13645) );
  OAI21_X1 U15692 ( .B1(n13646), .B2(n6578), .A(n13645), .ZN(P2_U3243) );
  XNOR2_X1 U15693 ( .A(n13647), .B(n13657), .ZN(n13649) );
  AOI21_X1 U15694 ( .B1(n13649), .B2(n13683), .A(n13648), .ZN(n13749) );
  INV_X1 U15695 ( .A(n13672), .ZN(n13651) );
  AOI211_X1 U15696 ( .C1(n13747), .C2(n13651), .A(n8705), .B(n13650), .ZN(
        n13746) );
  INV_X1 U15697 ( .A(n13652), .ZN(n13653) );
  AOI22_X1 U15698 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n6578), .B1(n13653), 
        .B2(n13673), .ZN(n13654) );
  OAI21_X1 U15699 ( .B1(n13655), .B2(n13677), .A(n13654), .ZN(n13659) );
  XOR2_X1 U15700 ( .A(n13657), .B(n13656), .Z(n13750) );
  NOR2_X1 U15701 ( .A1(n13750), .A2(n13697), .ZN(n13658) );
  AOI211_X1 U15702 ( .C1(n13746), .C2(n13694), .A(n13659), .B(n13658), .ZN(
        n13660) );
  OAI21_X1 U15703 ( .B1(n6578), .B2(n13749), .A(n13660), .ZN(P2_U3244) );
  XOR2_X1 U15704 ( .A(n13661), .B(n13664), .Z(n13755) );
  OAI21_X1 U15705 ( .B1(n13664), .B2(n13663), .A(n13662), .ZN(n13669) );
  AOI222_X1 U15706 ( .A1(n13683), .A2(n13669), .B1(n13668), .B2(n13667), .C1(
        n13666), .C2(n13665), .ZN(n13754) );
  INV_X1 U15707 ( .A(n13754), .ZN(n13679) );
  NAND2_X1 U15708 ( .A1(n13752), .A2(n13693), .ZN(n13670) );
  NAND2_X1 U15709 ( .A1(n13670), .A2(n6577), .ZN(n13671) );
  NOR2_X1 U15710 ( .A1(n13672), .A2(n13671), .ZN(n13751) );
  NAND2_X1 U15711 ( .A1(n13751), .A2(n13694), .ZN(n13676) );
  AOI22_X1 U15712 ( .A1(n6578), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13674), 
        .B2(n13673), .ZN(n13675) );
  OAI211_X1 U15713 ( .C1(n13510), .C2(n13677), .A(n13676), .B(n13675), .ZN(
        n13678) );
  AOI21_X1 U15714 ( .B1(n13679), .B2(n15045), .A(n13678), .ZN(n13680) );
  OAI21_X1 U15715 ( .B1(n13697), .B2(n13755), .A(n13680), .ZN(P2_U3245) );
  XOR2_X1 U15716 ( .A(n13685), .B(n13681), .Z(n13684) );
  AOI21_X1 U15717 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13759) );
  XOR2_X1 U15718 ( .A(n13686), .B(n13685), .Z(n13760) );
  INV_X1 U15719 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13688) );
  OAI22_X1 U15720 ( .A1(n15045), .A2(n13688), .B1(n13687), .B2(n15037), .ZN(
        n13689) );
  AOI21_X1 U15721 ( .B1(n13757), .B2(n13690), .A(n13689), .ZN(n13696) );
  AOI21_X1 U15722 ( .B1(n13691), .B2(n13757), .A(n8705), .ZN(n13692) );
  AND2_X1 U15723 ( .A1(n13693), .A2(n13692), .ZN(n13756) );
  NAND2_X1 U15724 ( .A1(n13756), .A2(n13694), .ZN(n13695) );
  OAI211_X1 U15725 ( .C1(n13760), .C2(n13697), .A(n13696), .B(n13695), .ZN(
        n13698) );
  INV_X1 U15726 ( .A(n13698), .ZN(n13699) );
  OAI21_X1 U15727 ( .B1(n13759), .B2(n6578), .A(n13699), .ZN(P2_U3246) );
  OAI211_X1 U15728 ( .C1(n13701), .C2(n15097), .A(n13700), .B(n13702), .ZN(
        n13782) );
  MUX2_X1 U15729 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13782), .S(n15141), .Z(
        P2_U3530) );
  OAI211_X1 U15730 ( .C1(n13704), .C2(n15097), .A(n13703), .B(n13702), .ZN(
        n13783) );
  MUX2_X1 U15731 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13783), .S(n15141), .Z(
        P2_U3529) );
  AOI21_X1 U15732 ( .B1(n15118), .B2(n13706), .A(n13705), .ZN(n13707) );
  OAI211_X1 U15733 ( .C1(n15078), .C2(n13709), .A(n13708), .B(n13707), .ZN(
        n13784) );
  MUX2_X1 U15734 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13784), .S(n15141), .Z(
        P2_U3528) );
  MUX2_X1 U15735 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13785), .S(n15141), .Z(
        P2_U3527) );
  AOI21_X1 U15736 ( .B1(n15118), .B2(n13717), .A(n13716), .ZN(n13718) );
  OAI211_X1 U15737 ( .C1(n15078), .C2(n13720), .A(n13719), .B(n13718), .ZN(
        n13786) );
  MUX2_X1 U15738 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13786), .S(n15141), .Z(
        P2_U3526) );
  AOI21_X1 U15739 ( .B1(n15118), .B2(n13722), .A(n13721), .ZN(n13723) );
  OAI211_X1 U15740 ( .C1(n15078), .C2(n13725), .A(n13724), .B(n13723), .ZN(
        n13787) );
  MUX2_X1 U15741 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13787), .S(n15141), .Z(
        P2_U3525) );
  AOI21_X1 U15742 ( .B1(n15118), .B2(n13727), .A(n13726), .ZN(n13728) );
  OAI211_X1 U15743 ( .C1(n15078), .C2(n13730), .A(n13729), .B(n13728), .ZN(
        n13788) );
  MUX2_X1 U15744 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13788), .S(n15141), .Z(
        P2_U3524) );
  AOI21_X1 U15745 ( .B1(n15118), .B2(n13732), .A(n13731), .ZN(n13733) );
  OAI211_X1 U15746 ( .C1(n12137), .C2(n13735), .A(n13734), .B(n13733), .ZN(
        n13789) );
  MUX2_X1 U15747 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13789), .S(n15141), .Z(
        P2_U3523) );
  AOI21_X1 U15748 ( .B1(n15118), .B2(n7056), .A(n13736), .ZN(n13737) );
  OAI211_X1 U15749 ( .C1(n15078), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        n13790) );
  MUX2_X1 U15750 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13790), .S(n15141), .Z(
        P2_U3522) );
  INV_X1 U15751 ( .A(n15078), .ZN(n15102) );
  OAI21_X1 U15752 ( .B1(n13741), .B2(n15097), .A(n13740), .ZN(n13743) );
  AOI211_X1 U15753 ( .C1(n13744), .C2(n15102), .A(n13743), .B(n13742), .ZN(
        n13745) );
  INV_X1 U15754 ( .A(n13745), .ZN(n13791) );
  MUX2_X1 U15755 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13791), .S(n15141), .Z(
        P2_U3521) );
  AOI21_X1 U15756 ( .B1(n15118), .B2(n13747), .A(n13746), .ZN(n13748) );
  OAI211_X1 U15757 ( .C1(n15078), .C2(n13750), .A(n13749), .B(n13748), .ZN(
        n13792) );
  MUX2_X1 U15758 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13792), .S(n15141), .Z(
        P2_U3520) );
  AOI21_X1 U15759 ( .B1(n15118), .B2(n13752), .A(n13751), .ZN(n13753) );
  OAI211_X1 U15760 ( .C1(n15078), .C2(n13755), .A(n13754), .B(n13753), .ZN(
        n13793) );
  MUX2_X1 U15761 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13793), .S(n15141), .Z(
        P2_U3519) );
  AOI21_X1 U15762 ( .B1(n15118), .B2(n13757), .A(n13756), .ZN(n13758) );
  OAI211_X1 U15763 ( .C1(n15078), .C2(n13760), .A(n13759), .B(n13758), .ZN(
        n13794) );
  MUX2_X1 U15764 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13794), .S(n15141), .Z(
        P2_U3518) );
  INV_X1 U15765 ( .A(n13761), .ZN(n13766) );
  AOI21_X1 U15766 ( .B1(n15118), .B2(n13763), .A(n13762), .ZN(n13764) );
  OAI211_X1 U15767 ( .C1(n15078), .C2(n13766), .A(n13765), .B(n13764), .ZN(
        n13795) );
  MUX2_X1 U15768 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13795), .S(n15141), .Z(
        P2_U3517) );
  AOI21_X1 U15769 ( .B1(n15118), .B2(n13768), .A(n13767), .ZN(n13769) );
  OAI211_X1 U15770 ( .C1(n13771), .C2(n15078), .A(n13770), .B(n13769), .ZN(
        n13796) );
  MUX2_X1 U15771 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13796), .S(n15141), .Z(
        P2_U3516) );
  AOI21_X1 U15772 ( .B1(n15118), .B2(n13773), .A(n13772), .ZN(n13774) );
  OAI211_X1 U15773 ( .C1(n13776), .C2(n15078), .A(n13775), .B(n13774), .ZN(
        n13797) );
  MUX2_X1 U15774 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13797), .S(n15141), .Z(
        P2_U3515) );
  AOI21_X1 U15775 ( .B1(n15118), .B2(n13778), .A(n13777), .ZN(n13779) );
  OAI211_X1 U15776 ( .C1(n13781), .C2(n15078), .A(n13780), .B(n13779), .ZN(
        n13798) );
  MUX2_X1 U15777 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13798), .S(n15141), .Z(
        P2_U3514) );
  MUX2_X1 U15778 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13782), .S(n15129), .Z(
        P2_U3498) );
  MUX2_X1 U15779 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13783), .S(n15129), .Z(
        P2_U3497) );
  MUX2_X1 U15780 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13784), .S(n15129), .Z(
        P2_U3496) );
  MUX2_X1 U15781 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13785), .S(n15129), .Z(
        P2_U3495) );
  MUX2_X1 U15782 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13786), .S(n15129), .Z(
        P2_U3494) );
  MUX2_X1 U15783 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13787), .S(n15129), .Z(
        P2_U3493) );
  MUX2_X1 U15784 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13788), .S(n15129), .Z(
        P2_U3492) );
  MUX2_X1 U15785 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13789), .S(n15129), .Z(
        P2_U3491) );
  MUX2_X1 U15786 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13790), .S(n15129), .Z(
        P2_U3490) );
  MUX2_X1 U15787 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13791), .S(n15129), .Z(
        P2_U3489) );
  MUX2_X1 U15788 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13792), .S(n15129), .Z(
        P2_U3488) );
  MUX2_X1 U15789 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13793), .S(n15129), .Z(
        P2_U3487) );
  MUX2_X1 U15790 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13794), .S(n15129), .Z(
        P2_U3486) );
  MUX2_X1 U15791 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13795), .S(n15129), .Z(
        P2_U3484) );
  MUX2_X1 U15792 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13796), .S(n15129), .Z(
        P2_U3481) );
  MUX2_X1 U15793 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13797), .S(n15129), .Z(
        P2_U3478) );
  MUX2_X1 U15794 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13798), .S(n15129), .Z(
        P2_U3475) );
  INV_X1 U15795 ( .A(n13799), .ZN(n14425) );
  NOR4_X1 U15796 ( .A1(n13801), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13800), .A4(
        P2_U3088), .ZN(n13802) );
  AOI21_X1 U15797 ( .B1(n13808), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13802), 
        .ZN(n13803) );
  OAI21_X1 U15798 ( .B1(n14425), .B2(n13818), .A(n13803), .ZN(P2_U3296) );
  OAI222_X1 U15799 ( .A1(n13818), .A2(n13806), .B1(P2_U3088), .B2(n13805), 
        .C1(n13804), .C2(n13820), .ZN(P2_U3298) );
  AOI21_X1 U15800 ( .B1(n13808), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13807), 
        .ZN(n13809) );
  OAI21_X1 U15801 ( .B1(n13810), .B2(n13818), .A(n13809), .ZN(P2_U3299) );
  INV_X1 U15802 ( .A(n13811), .ZN(n14427) );
  OAI222_X1 U15803 ( .A1(n13820), .A2(n13812), .B1(n13818), .B2(n14427), .C1(
        P2_U3088), .C2(n9010), .ZN(P2_U3300) );
  INV_X1 U15804 ( .A(n13813), .ZN(n14430) );
  OAI222_X1 U15805 ( .A1(P2_U3088), .A2(n13815), .B1(n13818), .B2(n14430), 
        .C1(n13814), .C2(n13820), .ZN(P2_U3301) );
  INV_X1 U15806 ( .A(n13816), .ZN(n14433) );
  OAI222_X1 U15807 ( .A1(n13820), .A2(n13819), .B1(n13818), .B2(n14433), .C1(
        P2_U3088), .C2(n13817), .ZN(P2_U3302) );
  MUX2_X1 U15808 ( .A(n13821), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U15809 ( .A(n13823), .B(n13822), .Z(n13829) );
  NAND2_X1 U15810 ( .A1(n14102), .A2(n13966), .ZN(n13825) );
  AOI22_X1 U15811 ( .A1(n14140), .A2(n13939), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13824) );
  OAI211_X1 U15812 ( .C1(n13963), .C2(n13826), .A(n13825), .B(n13824), .ZN(
        n13827) );
  AOI21_X1 U15813 ( .B1(n14337), .B2(n6564), .A(n13827), .ZN(n13828) );
  OAI21_X1 U15814 ( .B1(n13829), .B2(n13955), .A(n13828), .ZN(P1_U3214) );
  INV_X1 U15815 ( .A(n13831), .ZN(n13832) );
  AOI21_X1 U15816 ( .B1(n13833), .B2(n13830), .A(n13832), .ZN(n13840) );
  NAND2_X1 U15817 ( .A1(n13976), .A2(n14750), .ZN(n13835) );
  NAND2_X1 U15818 ( .A1(n13977), .A2(n14747), .ZN(n13834) );
  NAND2_X1 U15819 ( .A1(n13835), .A2(n13834), .ZN(n14654) );
  NAND2_X1 U15820 ( .A1(n14654), .A2(n13916), .ZN(n13836) );
  OAI211_X1 U15821 ( .C1(n13963), .C2(n14299), .A(n13837), .B(n13836), .ZN(
        n13838) );
  AOI21_X1 U15822 ( .B1(n11297), .B2(n6564), .A(n13838), .ZN(n13839) );
  OAI21_X1 U15823 ( .B1(n13840), .B2(n13955), .A(n13839), .ZN(P1_U3215) );
  XOR2_X1 U15824 ( .A(n13841), .B(n13842), .Z(n13847) );
  OAI22_X1 U15825 ( .A1(n13861), .A2(n13962), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15519), .ZN(n13843) );
  AOI21_X1 U15826 ( .B1(n14167), .B2(n13966), .A(n13843), .ZN(n13844) );
  OAI21_X1 U15827 ( .B1(n13963), .B2(n14171), .A(n13844), .ZN(n13845) );
  AOI21_X1 U15828 ( .B1(n14364), .B2(n6564), .A(n13845), .ZN(n13846) );
  OAI21_X1 U15829 ( .B1(n13847), .B2(n13955), .A(n13846), .ZN(P1_U3216) );
  OAI22_X1 U15830 ( .A1(n13860), .A2(n14189), .B1(n13903), .B2(n14191), .ZN(
        n14229) );
  NAND2_X1 U15831 ( .A1(n14229), .A2(n13916), .ZN(n13849) );
  OAI211_X1 U15832 ( .C1(n13963), .C2(n14221), .A(n13849), .B(n13848), .ZN(
        n13854) );
  AOI211_X1 U15833 ( .C1(n13852), .C2(n13851), .A(n13955), .B(n13850), .ZN(
        n13853) );
  AOI211_X1 U15834 ( .C1(n14388), .C2(n6564), .A(n13854), .B(n13853), .ZN(
        n13855) );
  INV_X1 U15835 ( .A(n13855), .ZN(P1_U3219) );
  OAI21_X1 U15836 ( .B1(n13858), .B2(n13857), .A(n13856), .ZN(n13859) );
  NAND2_X1 U15837 ( .A1(n13859), .A2(n13959), .ZN(n13867) );
  INV_X1 U15838 ( .A(n14211), .ZN(n13865) );
  OAI22_X1 U15839 ( .A1(n13861), .A2(n14189), .B1(n13860), .B2(n14191), .ZN(
        n14208) );
  INV_X1 U15840 ( .A(n14208), .ZN(n13863) );
  OAI22_X1 U15841 ( .A1(n13863), .A2(n13951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13862), .ZN(n13864) );
  AOI21_X1 U15842 ( .B1(n13865), .B2(n13949), .A(n13864), .ZN(n13866) );
  OAI211_X1 U15843 ( .C1(n7373), .C2(n13969), .A(n13867), .B(n13866), .ZN(
        P1_U3223) );
  AOI22_X1 U15844 ( .A1(n13868), .A2(n13916), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13869) );
  OAI21_X1 U15845 ( .B1(n13963), .B2(n13870), .A(n13869), .ZN(n13876) );
  INV_X1 U15846 ( .A(n13871), .ZN(n13872) );
  AOI211_X1 U15847 ( .C1(n13874), .C2(n13873), .A(n13955), .B(n13872), .ZN(
        n13875) );
  AOI211_X1 U15848 ( .C1(n13877), .C2(n6564), .A(n13876), .B(n13875), .ZN(
        n13878) );
  INV_X1 U15849 ( .A(n13878), .ZN(P1_U3224) );
  XOR2_X1 U15850 ( .A(n13880), .B(n13879), .Z(n13885) );
  NAND2_X1 U15851 ( .A1(n14140), .A2(n13966), .ZN(n13882) );
  AOI22_X1 U15852 ( .A1(n14167), .A2(n13939), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13881) );
  OAI211_X1 U15853 ( .C1(n13963), .C2(n14141), .A(n13882), .B(n13881), .ZN(
        n13883) );
  AOI21_X1 U15854 ( .B1(n14137), .B2(n6564), .A(n13883), .ZN(n13884) );
  OAI21_X1 U15855 ( .B1(n13885), .B2(n13955), .A(n13884), .ZN(P1_U3225) );
  OAI21_X1 U15856 ( .B1(n13888), .B2(n13887), .A(n13886), .ZN(n13889) );
  NAND2_X1 U15857 ( .A1(n13889), .A2(n13959), .ZN(n13896) );
  NAND2_X1 U15858 ( .A1(n14236), .A2(n14750), .ZN(n13891) );
  NAND2_X1 U15859 ( .A1(n13976), .A2(n14747), .ZN(n13890) );
  NAND2_X1 U15860 ( .A1(n13891), .A2(n13890), .ZN(n14263) );
  INV_X1 U15861 ( .A(n13892), .ZN(n13894) );
  NOR2_X1 U15862 ( .A1(n13963), .A2(n14268), .ZN(n13893) );
  AOI211_X1 U15863 ( .C1(n13916), .C2(n14263), .A(n13894), .B(n13893), .ZN(
        n13895) );
  OAI211_X1 U15864 ( .C1(n14647), .C2(n13969), .A(n13896), .B(n13895), .ZN(
        P1_U3226) );
  INV_X1 U15865 ( .A(n13897), .ZN(n13902) );
  AOI21_X1 U15866 ( .B1(n13899), .B2(n13901), .A(n13898), .ZN(n13900) );
  AOI21_X1 U15867 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13907) );
  NAND2_X1 U15868 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14076)
         );
  OAI22_X1 U15869 ( .A1(n13903), .A2(n14189), .B1(n6871), .B2(n14191), .ZN(
        n14252) );
  NAND2_X1 U15870 ( .A1(n14252), .A2(n13916), .ZN(n13904) );
  OAI211_X1 U15871 ( .C1(n13963), .C2(n14254), .A(n14076), .B(n13904), .ZN(
        n13905) );
  AOI21_X1 U15872 ( .B1(n14397), .B2(n6564), .A(n13905), .ZN(n13906) );
  OAI21_X1 U15873 ( .B1(n13907), .B2(n13955), .A(n13906), .ZN(P1_U3228) );
  XOR2_X1 U15874 ( .A(n13909), .B(n13908), .Z(n13915) );
  AND2_X1 U15875 ( .A1(n14183), .A2(n14747), .ZN(n13910) );
  AOI21_X1 U15876 ( .B1(n13972), .B2(n14750), .A(n13910), .ZN(n14150) );
  OAI22_X1 U15877 ( .A1(n14150), .A2(n13951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13911), .ZN(n13912) );
  AOI21_X1 U15878 ( .B1(n14156), .B2(n13949), .A(n13912), .ZN(n13914) );
  NAND2_X1 U15879 ( .A1(n14359), .A2(n6564), .ZN(n13913) );
  OAI211_X1 U15880 ( .C1(n13915), .C2(n13955), .A(n13914), .B(n13913), .ZN(
        P1_U3229) );
  AOI22_X1 U15881 ( .A1(n14380), .A2(n13916), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13917) );
  OAI21_X1 U15882 ( .B1(n13963), .B2(n13918), .A(n13917), .ZN(n13923) );
  AOI211_X1 U15883 ( .C1(n13921), .C2(n13920), .A(n13955), .B(n13919), .ZN(
        n13922) );
  AOI211_X1 U15884 ( .C1(n14381), .C2(n6564), .A(n13923), .B(n13922), .ZN(
        n13924) );
  INV_X1 U15885 ( .A(n13924), .ZN(P1_U3233) );
  OAI21_X1 U15886 ( .B1(n13927), .B2(n13926), .A(n13925), .ZN(n13928) );
  NAND2_X1 U15887 ( .A1(n13928), .A2(n13959), .ZN(n13933) );
  NOR2_X1 U15888 ( .A1(n13963), .A2(n14192), .ZN(n13931) );
  OAI22_X1 U15889 ( .A1(n14190), .A2(n13962), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13929), .ZN(n13930) );
  AOI211_X1 U15890 ( .C1(n13966), .C2(n14183), .A(n13931), .B(n13930), .ZN(
        n13932) );
  OAI211_X1 U15891 ( .C1(n13969), .C2(n14198), .A(n13933), .B(n13932), .ZN(
        P1_U3235) );
  OAI21_X1 U15892 ( .B1(n13936), .B2(n6777), .A(n13934), .ZN(n13937) );
  NAND2_X1 U15893 ( .A1(n13937), .A2(n13959), .ZN(n13945) );
  INV_X1 U15894 ( .A(n13938), .ZN(n14240) );
  AOI22_X1 U15895 ( .A1(n13939), .A2(n14236), .B1(P1_REG3_REG_18__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13940) );
  OAI21_X1 U15896 ( .B1(n13942), .B2(n13941), .A(n13940), .ZN(n13943) );
  AOI21_X1 U15897 ( .B1(n14240), .B2(n13949), .A(n13943), .ZN(n13944) );
  OAI211_X1 U15898 ( .C1(n14244), .C2(n13969), .A(n13945), .B(n13944), .ZN(
        P1_U3238) );
  XOR2_X1 U15899 ( .A(n13947), .B(n13946), .Z(n13956) );
  AND2_X1 U15900 ( .A1(n13972), .A2(n14747), .ZN(n13948) );
  AOI21_X1 U15901 ( .B1(n13971), .B2(n14750), .A(n13948), .ZN(n14343) );
  AOI22_X1 U15902 ( .A1(n14122), .A2(n13949), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13950) );
  OAI21_X1 U15903 ( .B1(n14343), .B2(n13951), .A(n13950), .ZN(n13952) );
  AOI21_X1 U15904 ( .B1(n14125), .B2(n6564), .A(n13952), .ZN(n13954) );
  OAI21_X1 U15905 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(P1_U3240) );
  OAI21_X1 U15906 ( .B1(n13958), .B2(n6730), .A(n13957), .ZN(n13960) );
  NAND2_X1 U15907 ( .A1(n13960), .A2(n13959), .ZN(n13968) );
  OAI22_X1 U15908 ( .A1(n13962), .A2(n13961), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15522), .ZN(n13965) );
  NOR2_X1 U15909 ( .A1(n13963), .A2(n14283), .ZN(n13964) );
  AOI211_X1 U15910 ( .C1(n13966), .C2(n14279), .A(n13965), .B(n13964), .ZN(
        n13967) );
  OAI211_X1 U15911 ( .C1(n6967), .C2(n13969), .A(n13968), .B(n13967), .ZN(
        P1_U3241) );
  MUX2_X1 U15912 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14084), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15913 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14104), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15914 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13970), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15915 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14102), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15916 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13971), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15917 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14140), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13972), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14167), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14183), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14168), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13973), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13974), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14237), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13975), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14236), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15927 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14279), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15928 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13976), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15929 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14278), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15930 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13977), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15931 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13978), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13979), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13980), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13981), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15935 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14749), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15936 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13982), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15937 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14748), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15938 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13983), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15939 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13984), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15940 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9650), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15941 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13985), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15942 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13986), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15943 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13987), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI22_X1 U15944 ( .A1(n14731), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14002) );
  MUX2_X1 U15945 ( .A(n14913), .B(P1_REG1_REG_2__SCAN_IN), .S(n13998), .Z(
        n13988) );
  NOR3_X1 U15946 ( .A1(n13990), .A2(n13989), .A3(n13988), .ZN(n13991) );
  NOR3_X1 U15947 ( .A1(n14721), .A2(n13992), .A3(n13991), .ZN(n14000) );
  MUX2_X1 U15948 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9079), .S(n13998), .Z(
        n13995) );
  NAND3_X1 U15949 ( .A1(n13995), .A2(n13994), .A3(n13993), .ZN(n13996) );
  NAND2_X1 U15950 ( .A1(n13996), .A2(n14014), .ZN(n13997) );
  OAI22_X1 U15951 ( .A1(n13998), .A2(n14725), .B1(n14723), .B2(n13997), .ZN(
        n13999) );
  NOR2_X1 U15952 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  NAND3_X1 U15953 ( .A1(n14003), .A2(n14002), .A3(n14001), .ZN(P1_U3245) );
  OAI22_X1 U15954 ( .A1(n14729), .A2(n15477), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14004), .ZN(n14005) );
  AOI21_X1 U15955 ( .B1(n14006), .B2(n14736), .A(n14005), .ZN(n14020) );
  NAND3_X1 U15956 ( .A1(n14009), .A2(n14008), .A3(n14007), .ZN(n14010) );
  NAND3_X1 U15957 ( .A1(n14738), .A2(n14011), .A3(n14010), .ZN(n14019) );
  MUX2_X1 U15958 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9323), .S(n14012), .Z(
        n14015) );
  NAND3_X1 U15959 ( .A1(n14015), .A2(n14014), .A3(n14013), .ZN(n14016) );
  NAND3_X1 U15960 ( .A1(n14733), .A2(n14017), .A3(n14016), .ZN(n14018) );
  NAND3_X1 U15961 ( .A1(n14020), .A2(n14019), .A3(n14018), .ZN(P1_U3246) );
  INV_X1 U15962 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14449) );
  NAND2_X1 U15963 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14021) );
  OAI21_X1 U15964 ( .B1(n14729), .B2(n14449), .A(n14021), .ZN(n14022) );
  AOI21_X1 U15965 ( .B1(n14027), .B2(n14736), .A(n14022), .ZN(n14035) );
  OAI21_X1 U15966 ( .B1(n14025), .B2(n14024), .A(n14023), .ZN(n14026) );
  NAND2_X1 U15967 ( .A1(n14738), .A2(n14026), .ZN(n14034) );
  MUX2_X1 U15968 ( .A(n9661), .B(P1_REG2_REG_5__SCAN_IN), .S(n14027), .Z(
        n14030) );
  NAND3_X1 U15969 ( .A1(n14030), .A2(n14029), .A3(n14028), .ZN(n14031) );
  NAND3_X1 U15970 ( .A1(n14733), .A2(n14032), .A3(n14031), .ZN(n14033) );
  NAND3_X1 U15971 ( .A1(n14035), .A2(n14034), .A3(n14033), .ZN(P1_U3248) );
  NOR2_X1 U15972 ( .A1(n14725), .A2(n14036), .ZN(n14037) );
  AOI211_X1 U15973 ( .C1(n14731), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14038), .B(
        n14037), .ZN(n14052) );
  OR3_X1 U15974 ( .A1(n14041), .A2(n14040), .A3(n14039), .ZN(n14042) );
  NAND3_X1 U15975 ( .A1(n14043), .A2(n14738), .A3(n14042), .ZN(n14051) );
  MUX2_X1 U15976 ( .A(n9698), .B(P1_REG2_REG_7__SCAN_IN), .S(n14044), .Z(
        n14045) );
  NAND3_X1 U15977 ( .A1(n14047), .A2(n14046), .A3(n14045), .ZN(n14048) );
  NAND3_X1 U15978 ( .A1(n14733), .A2(n14049), .A3(n14048), .ZN(n14050) );
  NAND3_X1 U15979 ( .A1(n14052), .A2(n14051), .A3(n14050), .ZN(P1_U3250) );
  INV_X1 U15980 ( .A(n14053), .ZN(n14058) );
  NOR3_X1 U15981 ( .A1(n14056), .A2(n14055), .A3(n14054), .ZN(n14057) );
  OAI21_X1 U15982 ( .B1(n14058), .B2(n14057), .A(n14738), .ZN(n14068) );
  INV_X1 U15983 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14460) );
  NAND2_X1 U15984 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14059) );
  OAI21_X1 U15985 ( .B1(n14729), .B2(n14460), .A(n14059), .ZN(n14060) );
  AOI21_X1 U15986 ( .B1(n14061), .B2(n14736), .A(n14060), .ZN(n14067) );
  MUX2_X1 U15987 ( .A(n10139), .B(P1_REG2_REG_9__SCAN_IN), .S(n14061), .Z(
        n14062) );
  NAND3_X1 U15988 ( .A1(n14064), .A2(n14063), .A3(n14062), .ZN(n14065) );
  NAND3_X1 U15989 ( .A1(n14733), .A2(n14707), .A3(n14065), .ZN(n14066) );
  NAND3_X1 U15990 ( .A1(n14068), .A2(n14067), .A3(n14066), .ZN(P1_U3252) );
  OAI211_X1 U15991 ( .C1(n14071), .C2(n14070), .A(n14733), .B(n14069), .ZN(
        n14079) );
  OAI211_X1 U15992 ( .C1(n14074), .C2(n14073), .A(n14072), .B(n14738), .ZN(
        n14075) );
  NAND2_X1 U15993 ( .A1(n14076), .A2(n14075), .ZN(n14077) );
  AOI21_X1 U15994 ( .B1(n14731), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14077), 
        .ZN(n14078) );
  OAI211_X1 U15995 ( .C1(n14725), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        P1_U3260) );
  NAND2_X1 U15996 ( .A1(n14319), .A2(n14100), .ZN(n14081) );
  XNOR2_X1 U15997 ( .A(n14081), .B(n14314), .ZN(n14316) );
  INV_X1 U15998 ( .A(P1_B_REG_SCAN_IN), .ZN(n14082) );
  NOR2_X1 U15999 ( .A1(n14426), .A2(n14082), .ZN(n14083) );
  NOR2_X1 U16000 ( .A1(n14189), .A2(n14083), .ZN(n14105) );
  AND2_X1 U16001 ( .A1(n14084), .A2(n14105), .ZN(n14313) );
  INV_X1 U16002 ( .A(n14313), .ZN(n14317) );
  NOR2_X1 U16003 ( .A1(n14317), .A2(n14286), .ZN(n14090) );
  AOI21_X1 U16004 ( .B1(n14797), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14090), 
        .ZN(n14086) );
  NAND2_X1 U16005 ( .A1(n14314), .A2(n14303), .ZN(n14085) );
  OAI211_X1 U16006 ( .C1(n14316), .C2(n14087), .A(n14086), .B(n14085), .ZN(
        P1_U3263) );
  XNOR2_X1 U16007 ( .A(n14100), .B(n14091), .ZN(n14088) );
  NAND2_X1 U16008 ( .A1(n14088), .A2(n14790), .ZN(n14318) );
  AND2_X1 U16009 ( .A1(n14797), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14089) );
  NOR2_X1 U16010 ( .A1(n14090), .A2(n14089), .ZN(n14093) );
  NAND2_X1 U16011 ( .A1(n14091), .A2(n14303), .ZN(n14092) );
  OAI211_X1 U16012 ( .C1(n14318), .C2(n14273), .A(n14093), .B(n14092), .ZN(
        P1_U3264) );
  NAND2_X1 U16013 ( .A1(n14098), .A2(n14102), .ZN(n14096) );
  AOI211_X1 U16014 ( .C1(n14113), .C2(n14101), .A(n14837), .B(n14100), .ZN(
        n14324) );
  INV_X1 U16015 ( .A(n14324), .ZN(n14115) );
  NAND2_X1 U16016 ( .A1(n14102), .A2(n14747), .ZN(n14320) );
  NOR2_X1 U16017 ( .A1(n14320), .A2(n14286), .ZN(n14112) );
  NAND2_X1 U16018 ( .A1(n14284), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14109) );
  INV_X1 U16019 ( .A(n14103), .ZN(n14107) );
  NAND2_X1 U16020 ( .A1(n14105), .A2(n14104), .ZN(n14321) );
  INV_X1 U16021 ( .A(n14321), .ZN(n14106) );
  AOI22_X1 U16022 ( .A1(n14797), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n14107), 
        .B2(n14106), .ZN(n14108) );
  OAI21_X1 U16023 ( .B1(n14110), .B2(n14109), .A(n14108), .ZN(n14111) );
  AOI211_X1 U16024 ( .C1(n14113), .C2(n14303), .A(n14112), .B(n14111), .ZN(
        n14114) );
  OAI21_X1 U16025 ( .B1(n14115), .B2(n14273), .A(n14114), .ZN(n14116) );
  AOI21_X1 U16026 ( .B1(n14325), .B2(n14136), .A(n14116), .ZN(n14117) );
  OAI21_X1 U16027 ( .B1(n14328), .B2(n14292), .A(n14117), .ZN(P1_U3356) );
  XNOR2_X1 U16028 ( .A(n14119), .B(n14118), .ZN(n14349) );
  AOI21_X1 U16029 ( .B1(n6700), .B2(n14120), .A(n6610), .ZN(n14347) );
  OAI211_X1 U16030 ( .C1(n14345), .C2(n14139), .A(n14790), .B(n14121), .ZN(
        n14344) );
  AOI22_X1 U16031 ( .A1(n14122), .A2(n14284), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n14797), .ZN(n14123) );
  OAI21_X1 U16032 ( .B1(n14343), .B2(n14286), .A(n14123), .ZN(n14124) );
  AOI21_X1 U16033 ( .B1(n14125), .B2(n14303), .A(n14124), .ZN(n14126) );
  OAI21_X1 U16034 ( .B1(n14344), .B2(n14273), .A(n14126), .ZN(n14127) );
  AOI21_X1 U16035 ( .B1(n14347), .B2(n14306), .A(n14127), .ZN(n14128) );
  OAI21_X1 U16036 ( .B1(n14349), .B2(n14129), .A(n14128), .ZN(P1_U3267) );
  AOI21_X1 U16037 ( .B1(n14134), .B2(n14131), .A(n14130), .ZN(n14132) );
  INV_X1 U16038 ( .A(n14132), .ZN(n14357) );
  OAI21_X1 U16039 ( .B1(n14135), .B2(n14134), .A(n14133), .ZN(n14355) );
  NAND2_X1 U16040 ( .A1(n14355), .A2(n14136), .ZN(n14147) );
  AND2_X1 U16041 ( .A1(n14137), .A2(n14154), .ZN(n14138) );
  NOR2_X1 U16042 ( .A1(n14139), .A2(n14138), .ZN(n14350) );
  AOI22_X1 U16043 ( .A1(n14140), .A2(n14750), .B1(n14747), .B2(n14167), .ZN(
        n14351) );
  OAI21_X1 U16044 ( .B1(n14141), .B2(n14783), .A(n14351), .ZN(n14142) );
  MUX2_X1 U16045 ( .A(P1_REG2_REG_25__SCAN_IN), .B(n14142), .S(n14301), .Z(
        n14144) );
  NOR2_X1 U16046 ( .A1(n14353), .A2(n14786), .ZN(n14143) );
  AOI211_X1 U16047 ( .C1(n14350), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        n14146) );
  OAI211_X1 U16048 ( .C1(n14357), .C2(n14292), .A(n14147), .B(n14146), .ZN(
        P1_U3268) );
  AOI211_X1 U16049 ( .C1(n14160), .C2(n14149), .A(n14863), .B(n14148), .ZN(
        n14152) );
  INV_X1 U16050 ( .A(n14150), .ZN(n14151) );
  NOR2_X1 U16051 ( .A1(n14152), .A2(n14151), .ZN(n14361) );
  INV_X1 U16052 ( .A(n14154), .ZN(n14155) );
  AOI211_X1 U16053 ( .C1(n14359), .C2(n14170), .A(n14837), .B(n14155), .ZN(
        n14358) );
  AOI22_X1 U16054 ( .A1(n14156), .A2(n14284), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n14286), .ZN(n14157) );
  OAI21_X1 U16055 ( .B1(n14158), .B2(n14786), .A(n14157), .ZN(n14164) );
  OAI21_X1 U16056 ( .B1(n14161), .B2(n14160), .A(n14159), .ZN(n14162) );
  INV_X1 U16057 ( .A(n14162), .ZN(n14362) );
  NOR2_X1 U16058 ( .A1(n14362), .A2(n14292), .ZN(n14163) );
  AOI211_X1 U16059 ( .C1(n14358), .C2(n14793), .A(n14164), .B(n14163), .ZN(
        n14165) );
  OAI21_X1 U16060 ( .B1(n14361), .B2(n14797), .A(n14165), .ZN(P1_U3269) );
  XNOR2_X1 U16061 ( .A(n6694), .B(n14166), .ZN(n14169) );
  AOI222_X1 U16062 ( .A1(n14902), .A2(n14169), .B1(n14168), .B2(n14747), .C1(
        n14167), .C2(n14750), .ZN(n14366) );
  AOI211_X1 U16063 ( .C1(n14364), .C2(n14194), .A(n14837), .B(n14153), .ZN(
        n14363) );
  INV_X1 U16064 ( .A(n14171), .ZN(n14172) );
  AOI22_X1 U16065 ( .A1(n14172), .A2(n14284), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n14286), .ZN(n14173) );
  OAI21_X1 U16066 ( .B1(n14174), .B2(n14786), .A(n14173), .ZN(n14180) );
  AND2_X1 U16067 ( .A1(n14176), .A2(n14175), .ZN(n14177) );
  OR2_X1 U16068 ( .A1(n14178), .A2(n14177), .ZN(n14367) );
  NOR2_X1 U16069 ( .A1(n14367), .A2(n14292), .ZN(n14179) );
  AOI211_X1 U16070 ( .C1(n14363), .C2(n14793), .A(n14180), .B(n14179), .ZN(
        n14181) );
  OAI21_X1 U16071 ( .B1(n14366), .B2(n14797), .A(n14181), .ZN(P1_U3270) );
  XOR2_X1 U16072 ( .A(n14182), .B(n14186), .Z(n14372) );
  INV_X1 U16073 ( .A(n14183), .ZN(n14188) );
  AOI21_X1 U16074 ( .B1(n14186), .B2(n14185), .A(n14184), .ZN(n14187) );
  OAI222_X1 U16075 ( .A1(n14191), .A2(n14190), .B1(n14189), .B2(n14188), .C1(
        n14863), .C2(n14187), .ZN(n14368) );
  NOR2_X1 U16076 ( .A1(n14192), .A2(n14783), .ZN(n14193) );
  OAI21_X1 U16077 ( .B1(n14368), .B2(n14193), .A(n14301), .ZN(n14201) );
  INV_X1 U16078 ( .A(n14213), .ZN(n14196) );
  INV_X1 U16079 ( .A(n14194), .ZN(n14195) );
  AOI211_X1 U16080 ( .C1(n14370), .C2(n14196), .A(n14837), .B(n14195), .ZN(
        n14369) );
  INV_X1 U16081 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14197) );
  OAI22_X1 U16082 ( .A1(n14198), .A2(n14786), .B1(n14197), .B2(n14301), .ZN(
        n14199) );
  AOI21_X1 U16083 ( .B1(n14369), .B2(n14793), .A(n14199), .ZN(n14200) );
  OAI211_X1 U16084 ( .C1(n14372), .C2(n14292), .A(n14201), .B(n14200), .ZN(
        P1_U3271) );
  NAND2_X1 U16085 ( .A1(n14202), .A2(n14205), .ZN(n14203) );
  NOR3_X1 U16086 ( .A1(n11839), .A2(n14206), .A3(n14205), .ZN(n14207) );
  NOR2_X1 U16087 ( .A1(n14207), .A2(n14863), .ZN(n14210) );
  AOI21_X1 U16088 ( .B1(n14210), .B2(n14209), .A(n14208), .ZN(n14376) );
  OAI21_X1 U16089 ( .B1(n14211), .B2(n14783), .A(n14376), .ZN(n14212) );
  NAND2_X1 U16090 ( .A1(n14212), .A2(n14301), .ZN(n14218) );
  AOI211_X1 U16091 ( .C1(n14374), .C2(n14214), .A(n14837), .B(n14213), .ZN(
        n14373) );
  INV_X1 U16092 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14215) );
  OAI22_X1 U16093 ( .A1(n7373), .A2(n14786), .B1(n14301), .B2(n14215), .ZN(
        n14216) );
  AOI21_X1 U16094 ( .B1(n14373), .B2(n14793), .A(n14216), .ZN(n14217) );
  OAI211_X1 U16095 ( .C1(n14377), .C2(n14292), .A(n14218), .B(n14217), .ZN(
        P1_U3272) );
  XNOR2_X1 U16096 ( .A(n14219), .B(n14227), .ZN(n14391) );
  AOI211_X1 U16097 ( .C1(n14388), .C2(n14242), .A(n14837), .B(n11812), .ZN(
        n14387) );
  INV_X1 U16098 ( .A(n14388), .ZN(n14224) );
  INV_X1 U16099 ( .A(n14221), .ZN(n14222) );
  AOI22_X1 U16100 ( .A1(n14286), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14222), 
        .B2(n14284), .ZN(n14223) );
  OAI21_X1 U16101 ( .B1(n14224), .B2(n14786), .A(n14223), .ZN(n14232) );
  AND2_X1 U16102 ( .A1(n14234), .A2(n14225), .ZN(n14228) );
  OAI21_X1 U16103 ( .B1(n14228), .B2(n14227), .A(n14226), .ZN(n14230) );
  AOI21_X1 U16104 ( .B1(n14230), .B2(n14902), .A(n14229), .ZN(n14390) );
  NOR2_X1 U16105 ( .A1(n14390), .A2(n14286), .ZN(n14231) );
  AOI211_X1 U16106 ( .C1(n14387), .C2(n14793), .A(n14232), .B(n14231), .ZN(
        n14233) );
  OAI21_X1 U16107 ( .B1(n14391), .B2(n14292), .A(n14233), .ZN(P1_U3274) );
  OAI211_X1 U16108 ( .C1(n14235), .C2(n14245), .A(n14234), .B(n14902), .ZN(
        n14239) );
  AOI22_X1 U16109 ( .A1(n14237), .A2(n14750), .B1(n14747), .B2(n14236), .ZN(
        n14238) );
  NAND2_X1 U16110 ( .A1(n14239), .A2(n14238), .ZN(n14392) );
  AOI21_X1 U16111 ( .B1(n14240), .B2(n14284), .A(n14392), .ZN(n14250) );
  OR2_X1 U16112 ( .A1(n6720), .A2(n14244), .ZN(n14241) );
  AND3_X1 U16113 ( .A1(n14242), .A2(n14790), .A3(n14241), .ZN(n14393) );
  OAI22_X1 U16114 ( .A1(n14244), .A2(n14786), .B1(n14243), .B2(n14301), .ZN(
        n14248) );
  XOR2_X1 U16115 ( .A(n14246), .B(n14245), .Z(n14395) );
  NOR2_X1 U16116 ( .A1(n14395), .A2(n14292), .ZN(n14247) );
  AOI211_X1 U16117 ( .C1(n14393), .C2(n14793), .A(n14248), .B(n14247), .ZN(
        n14249) );
  OAI21_X1 U16118 ( .B1(n14797), .B2(n14250), .A(n14249), .ZN(P1_U3275) );
  XNOR2_X1 U16119 ( .A(n14251), .B(n14257), .ZN(n14253) );
  AOI21_X1 U16120 ( .B1(n14253), .B2(n14902), .A(n14252), .ZN(n14399) );
  AOI211_X1 U16121 ( .C1(n14397), .C2(n14267), .A(n14837), .B(n6720), .ZN(
        n14396) );
  INV_X1 U16122 ( .A(n14254), .ZN(n14255) );
  AOI22_X1 U16123 ( .A1(n14286), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14255), 
        .B2(n14284), .ZN(n14256) );
  OAI21_X1 U16124 ( .B1(n7062), .B2(n14786), .A(n14256), .ZN(n14260) );
  XNOR2_X1 U16125 ( .A(n14258), .B(n14257), .ZN(n14400) );
  NOR2_X1 U16126 ( .A1(n14400), .A2(n14292), .ZN(n14259) );
  AOI211_X1 U16127 ( .C1(n14396), .C2(n14793), .A(n14260), .B(n14259), .ZN(
        n14261) );
  OAI21_X1 U16128 ( .B1(n14797), .B2(n14399), .A(n14261), .ZN(P1_U3276) );
  XNOR2_X1 U16129 ( .A(n14262), .B(n14266), .ZN(n14264) );
  AOI21_X1 U16130 ( .B1(n14264), .B2(n14902), .A(n14263), .ZN(n14648) );
  XNOR2_X1 U16131 ( .A(n14265), .B(n14266), .ZN(n14651) );
  OAI211_X1 U16132 ( .C1(n6719), .C2(n14647), .A(n14790), .B(n14267), .ZN(
        n14646) );
  OAI22_X1 U16133 ( .A1(n14301), .A2(n14269), .B1(n14268), .B2(n14783), .ZN(
        n14270) );
  AOI21_X1 U16134 ( .B1(n14271), .B2(n14303), .A(n14270), .ZN(n14272) );
  OAI21_X1 U16135 ( .B1(n14646), .B2(n14273), .A(n14272), .ZN(n14274) );
  AOI21_X1 U16136 ( .B1(n14651), .B2(n14306), .A(n14274), .ZN(n14275) );
  OAI21_X1 U16137 ( .B1(n14648), .B2(n14797), .A(n14275), .ZN(P1_U3277) );
  OAI211_X1 U16138 ( .C1(n14277), .C2(n14291), .A(n14276), .B(n14902), .ZN(
        n14281) );
  AOI22_X1 U16139 ( .A1(n14750), .A2(n14279), .B1(n14278), .B2(n14747), .ZN(
        n14280) );
  AND2_X1 U16140 ( .A1(n14281), .A2(n14280), .ZN(n14404) );
  INV_X1 U16141 ( .A(n14282), .ZN(n14307) );
  AOI211_X1 U16142 ( .C1(n14402), .C2(n14307), .A(n14837), .B(n6719), .ZN(
        n14401) );
  INV_X1 U16143 ( .A(n14283), .ZN(n14285) );
  AOI22_X1 U16144 ( .A1(n14286), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14285), 
        .B2(n14284), .ZN(n14287) );
  OAI21_X1 U16145 ( .B1(n6967), .B2(n14786), .A(n14287), .ZN(n14294) );
  INV_X1 U16146 ( .A(n14288), .ZN(n14289) );
  AOI21_X1 U16147 ( .B1(n14291), .B2(n14290), .A(n14289), .ZN(n14405) );
  NOR2_X1 U16148 ( .A1(n14405), .A2(n14292), .ZN(n14293) );
  AOI211_X1 U16149 ( .C1(n14401), .C2(n14793), .A(n14294), .B(n14293), .ZN(
        n14295) );
  OAI21_X1 U16150 ( .B1(n14797), .B2(n14404), .A(n14295), .ZN(P1_U3278) );
  OAI211_X1 U16151 ( .C1(n14297), .C2(n14305), .A(n14902), .B(n14296), .ZN(
        n14657) );
  INV_X1 U16152 ( .A(n14657), .ZN(n14298) );
  OAI21_X1 U16153 ( .B1(n14298), .B2(n14654), .A(n14301), .ZN(n14312) );
  OAI22_X1 U16154 ( .A1(n14301), .A2(n14300), .B1(n14299), .B2(n14783), .ZN(
        n14302) );
  AOI21_X1 U16155 ( .B1(n11297), .B2(n14303), .A(n14302), .ZN(n14311) );
  NAND2_X1 U16156 ( .A1(n14304), .A2(n14305), .ZN(n14655) );
  NAND3_X1 U16157 ( .A1(n6615), .A2(n14655), .A3(n14306), .ZN(n14310) );
  AOI211_X1 U16158 ( .C1(n11297), .C2(n14308), .A(n14837), .B(n14282), .ZN(
        n14653) );
  NAND2_X1 U16159 ( .A1(n14653), .A2(n14793), .ZN(n14309) );
  NAND4_X1 U16160 ( .A1(n14312), .A2(n14311), .A3(n14310), .A4(n14309), .ZN(
        P1_U3279) );
  AOI21_X1 U16161 ( .B1(n14314), .B2(n14876), .A(n14313), .ZN(n14315) );
  OAI21_X1 U16162 ( .B1(n14316), .B2(n14837), .A(n14315), .ZN(n14406) );
  MUX2_X1 U16163 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14406), .S(n14929), .Z(
        P1_U3559) );
  OAI211_X1 U16164 ( .C1(n14319), .C2(n14899), .A(n14318), .B(n14317), .ZN(
        n14407) );
  MUX2_X1 U16165 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14407), .S(n14929), .Z(
        P1_U3558) );
  OAI211_X1 U16166 ( .C1(n14322), .C2(n14899), .A(n14321), .B(n14320), .ZN(
        n14323) );
  NAND2_X1 U16167 ( .A1(n14329), .A2(n14906), .ZN(n14334) );
  AOI22_X1 U16168 ( .A1(n14331), .A2(n14790), .B1(n14876), .B2(n14330), .ZN(
        n14332) );
  OAI211_X1 U16169 ( .C1(n14335), .C2(n14334), .A(n14333), .B(n14332), .ZN(
        n14408) );
  MUX2_X1 U16170 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14408), .S(n14929), .Z(
        P1_U3556) );
  AOI21_X1 U16171 ( .B1(n14876), .B2(n14337), .A(n14336), .ZN(n14338) );
  MUX2_X1 U16172 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14409), .S(n14929), .Z(
        P1_U3555) );
  OAI211_X1 U16173 ( .C1(n14345), .C2(n14899), .A(n14344), .B(n14343), .ZN(
        n14346) );
  AOI21_X1 U16174 ( .B1(n14347), .B2(n14906), .A(n14346), .ZN(n14348) );
  OAI21_X1 U16175 ( .B1(n14349), .B2(n14863), .A(n14348), .ZN(n14410) );
  MUX2_X1 U16176 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14410), .S(n14929), .Z(
        P1_U3554) );
  NAND2_X1 U16177 ( .A1(n14350), .A2(n14790), .ZN(n14352) );
  OAI211_X1 U16178 ( .C1(n14353), .C2(n14899), .A(n14352), .B(n14351), .ZN(
        n14354) );
  AOI21_X1 U16179 ( .B1(n14355), .B2(n14902), .A(n14354), .ZN(n14356) );
  OAI21_X1 U16180 ( .B1(n14828), .B2(n14357), .A(n14356), .ZN(n14411) );
  MUX2_X1 U16181 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14411), .S(n14929), .Z(
        P1_U3553) );
  AOI21_X1 U16182 ( .B1(n14876), .B2(n14359), .A(n14358), .ZN(n14360) );
  OAI211_X1 U16183 ( .C1(n14828), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14412) );
  MUX2_X1 U16184 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14412), .S(n14929), .Z(
        P1_U3552) );
  AOI21_X1 U16185 ( .B1(n14876), .B2(n14364), .A(n14363), .ZN(n14365) );
  OAI211_X1 U16186 ( .C1(n14828), .C2(n14367), .A(n14366), .B(n14365), .ZN(
        n14413) );
  MUX2_X1 U16187 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14413), .S(n14929), .Z(
        P1_U3551) );
  AOI211_X1 U16188 ( .C1(n14876), .C2(n14370), .A(n14369), .B(n14368), .ZN(
        n14371) );
  OAI21_X1 U16189 ( .B1(n14828), .B2(n14372), .A(n14371), .ZN(n14414) );
  MUX2_X1 U16190 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14414), .S(n14929), .Z(
        P1_U3550) );
  AOI21_X1 U16191 ( .B1(n14876), .B2(n14374), .A(n14373), .ZN(n14375) );
  OAI211_X1 U16192 ( .C1(n14828), .C2(n14377), .A(n14376), .B(n14375), .ZN(
        n14415) );
  MUX2_X1 U16193 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14415), .S(n14929), .Z(
        P1_U3549) );
  NAND2_X1 U16194 ( .A1(n14378), .A2(n14902), .ZN(n14386) );
  AOI211_X1 U16195 ( .C1(n14876), .C2(n14381), .A(n14380), .B(n14379), .ZN(
        n14385) );
  NAND3_X1 U16196 ( .A1(n14383), .A2(n14906), .A3(n14382), .ZN(n14384) );
  OAI211_X1 U16197 ( .C1(n11839), .C2(n14386), .A(n14385), .B(n14384), .ZN(
        n14416) );
  MUX2_X1 U16198 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14416), .S(n14929), .Z(
        P1_U3548) );
  AOI21_X1 U16199 ( .B1(n14876), .B2(n14388), .A(n14387), .ZN(n14389) );
  OAI211_X1 U16200 ( .C1(n14828), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        n14417) );
  MUX2_X1 U16201 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14417), .S(n14929), .Z(
        P1_U3547) );
  AOI211_X1 U16202 ( .C1(n14876), .C2(n11350), .A(n14393), .B(n14392), .ZN(
        n14394) );
  OAI21_X1 U16203 ( .B1(n14828), .B2(n14395), .A(n14394), .ZN(n14418) );
  MUX2_X1 U16204 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14418), .S(n14929), .Z(
        P1_U3546) );
  AOI21_X1 U16205 ( .B1(n14876), .B2(n14397), .A(n14396), .ZN(n14398) );
  OAI211_X1 U16206 ( .C1(n14828), .C2(n14400), .A(n14399), .B(n14398), .ZN(
        n14419) );
  MUX2_X1 U16207 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14419), .S(n14929), .Z(
        P1_U3545) );
  AOI21_X1 U16208 ( .B1(n14876), .B2(n14402), .A(n14401), .ZN(n14403) );
  OAI211_X1 U16209 ( .C1(n14405), .C2(n14828), .A(n14404), .B(n14403), .ZN(
        n14420) );
  MUX2_X1 U16210 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14420), .S(n14929), .Z(
        P1_U3543) );
  MUX2_X1 U16211 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14406), .S(n14909), .Z(
        P1_U3527) );
  MUX2_X1 U16212 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14407), .S(n14909), .Z(
        P1_U3526) );
  MUX2_X1 U16213 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14408), .S(n14909), .Z(
        P1_U3524) );
  MUX2_X1 U16214 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14409), .S(n14909), .Z(
        P1_U3523) );
  MUX2_X1 U16215 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14410), .S(n14909), .Z(
        P1_U3522) );
  MUX2_X1 U16216 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14411), .S(n14909), .Z(
        P1_U3521) );
  MUX2_X1 U16217 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14412), .S(n14909), .Z(
        P1_U3520) );
  MUX2_X1 U16218 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14413), .S(n14909), .Z(
        P1_U3519) );
  MUX2_X1 U16219 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14414), .S(n14909), .Z(
        P1_U3518) );
  MUX2_X1 U16220 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14415), .S(n14909), .Z(
        P1_U3517) );
  MUX2_X1 U16221 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14416), .S(n14909), .Z(
        P1_U3516) );
  MUX2_X1 U16222 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14417), .S(n14909), .Z(
        P1_U3515) );
  MUX2_X1 U16223 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14418), .S(n14909), .Z(
        P1_U3513) );
  MUX2_X1 U16224 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14419), .S(n14909), .Z(
        P1_U3510) );
  MUX2_X1 U16225 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14420), .S(n14909), .Z(
        P1_U3504) );
  NOR4_X1 U16226 ( .A1(n14421), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8966), .A4(
        P1_U3086), .ZN(n14422) );
  AOI21_X1 U16227 ( .B1(n14423), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14422), 
        .ZN(n14424) );
  OAI21_X1 U16228 ( .B1(n14425), .B2(n14434), .A(n14424), .ZN(P1_U3324) );
  OAI222_X1 U16229 ( .A1(n14436), .A2(n14429), .B1(n14428), .B2(n14427), .C1(
        P1_U3086), .C2(n14426), .ZN(P1_U3328) );
  OAI222_X1 U16230 ( .A1(n14431), .A2(P1_U3086), .B1(n14434), .B2(n14430), 
        .C1(n15333), .C2(n14436), .ZN(P1_U3329) );
  OAI222_X1 U16231 ( .A1(n14436), .A2(n14435), .B1(n14434), .B2(n14433), .C1(
        n14432), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U16232 ( .A(n14437), .B(n10306), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16233 ( .A(n14438), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16234 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15313) );
  INV_X1 U16235 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15453) );
  NOR2_X1 U16236 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15303), .ZN(n14471) );
  INV_X1 U16237 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14730) );
  NOR2_X1 U16238 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14730), .ZN(n14470) );
  INV_X1 U16239 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14439) );
  NOR2_X1 U16240 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14439), .ZN(n14468) );
  INV_X1 U16241 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14477) );
  INV_X1 U16242 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14466) );
  XNOR2_X1 U16243 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14466), .ZN(n14524) );
  INV_X1 U16244 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14464) );
  XOR2_X1 U16245 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Z(
        n14517) );
  XOR2_X1 U16246 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14458), .Z(n14484) );
  XNOR2_X1 U16247 ( .A(n6905), .B(n14442), .ZN(n14489) );
  NAND2_X1 U16248 ( .A1(n14492), .A2(n14491), .ZN(n14440) );
  NAND2_X1 U16249 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14443), .ZN(n14445) );
  NAND2_X1 U16250 ( .A1(n14498), .A2(n15477), .ZN(n14444) );
  NAND2_X1 U16251 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14446), .ZN(n14447) );
  NAND2_X1 U16252 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14448), .ZN(n14451) );
  NAND2_X1 U16253 ( .A1(n14502), .A2(n14449), .ZN(n14450) );
  NAND2_X1 U16254 ( .A1(n14454), .A2(n14453), .ZN(n14456) );
  XOR2_X1 U16255 ( .A(n14454), .B(n14453), .Z(n14511) );
  NAND2_X1 U16256 ( .A1(n14511), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14455) );
  NAND2_X1 U16257 ( .A1(n14456), .A2(n14455), .ZN(n14485) );
  NAND2_X1 U16258 ( .A1(n14484), .A2(n14485), .ZN(n14457) );
  NAND2_X1 U16259 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14482), .ZN(n14462) );
  NOR2_X1 U16260 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14482), .ZN(n14461) );
  XNOR2_X1 U16261 ( .A(n15383), .B(n14464), .ZN(n14480) );
  NAND2_X1 U16262 ( .A1(n14481), .A2(n14480), .ZN(n14463) );
  AND2_X1 U16263 ( .A1(n14477), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14467) );
  OAI22_X1 U16264 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15504), .B1(n14468), 
        .B2(n14528), .ZN(n14533) );
  OAI22_X1 U16265 ( .A1(n14470), .A2(n14533), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14469), .ZN(n14475) );
  OAI22_X1 U16266 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15453), .B1(n14471), 
        .B2(n14475), .ZN(n14472) );
  NOR2_X1 U16267 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14472), .ZN(n14474) );
  XOR2_X1 U16268 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14472), .Z(n14537) );
  AND2_X1 U16269 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14537), .ZN(n14473) );
  NOR2_X1 U16270 ( .A1(n14474), .A2(n14473), .ZN(n14575) );
  INV_X1 U16271 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14577) );
  XNOR2_X1 U16272 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n14577), .ZN(n14574) );
  XNOR2_X1 U16273 ( .A(n14575), .B(n14574), .ZN(n14572) );
  INV_X1 U16274 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14540) );
  INV_X1 U16275 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15320) );
  XOR2_X1 U16276 ( .A(n15453), .B(P3_ADDR_REG_16__SCAN_IN), .Z(n14476) );
  XNOR2_X1 U16277 ( .A(n14476), .B(n14475), .ZN(n14697) );
  INV_X1 U16278 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15017) );
  XNOR2_X1 U16279 ( .A(n14477), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14478) );
  XNOR2_X1 U16280 ( .A(n14479), .B(n14478), .ZN(n14687) );
  XOR2_X1 U16281 ( .A(n14481), .B(n14480), .Z(n14682) );
  INV_X1 U16282 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15434) );
  XOR2_X1 U16283 ( .A(n15434), .B(P3_ADDR_REG_10__SCAN_IN), .Z(n14483) );
  XOR2_X1 U16284 ( .A(n14483), .B(n14482), .Z(n14553) );
  XOR2_X1 U16285 ( .A(n14485), .B(n14484), .Z(n14515) );
  NAND2_X1 U16286 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14488), .ZN(n14501) );
  INV_X1 U16287 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15365) );
  XNOR2_X1 U16288 ( .A(n14490), .B(n14489), .ZN(n14544) );
  XNOR2_X1 U16289 ( .A(n14492), .B(n14491), .ZN(n14494) );
  NAND2_X1 U16290 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14494), .ZN(n14496) );
  AOI21_X1 U16291 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14493), .A(n14492), .ZN(
        n15545) );
  NOR2_X1 U16292 ( .A1(n15545), .A2(n9049), .ZN(n15554) );
  XOR2_X1 U16293 ( .A(n14494), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15553) );
  NAND2_X1 U16294 ( .A1(n15554), .A2(n15553), .ZN(n14495) );
  NAND2_X1 U16295 ( .A1(n14496), .A2(n14495), .ZN(n14545) );
  NAND2_X1 U16296 ( .A1(n14544), .A2(n14545), .ZN(n14497) );
  NOR2_X1 U16297 ( .A1(n14544), .A2(n14545), .ZN(n14543) );
  AOI21_X1 U16298 ( .B1(n15365), .B2(n14497), .A(n14543), .ZN(n15549) );
  XOR2_X1 U16299 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14498), .Z(n15550) );
  NOR2_X1 U16300 ( .A1(n15549), .A2(n15550), .ZN(n14499) );
  INV_X1 U16301 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U16302 ( .A1(n15549), .A2(n15550), .ZN(n15548) );
  OAI21_X1 U16303 ( .B1(n14499), .B2(n15551), .A(n15548), .ZN(n15542) );
  NAND2_X1 U16304 ( .A1(n15543), .A2(n15542), .ZN(n14500) );
  NAND2_X1 U16305 ( .A1(n14501), .A2(n14500), .ZN(n14504) );
  XOR2_X1 U16306 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14502), .Z(n14503) );
  NAND2_X1 U16307 ( .A1(n14505), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14510) );
  INV_X1 U16308 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14974) );
  XOR2_X1 U16309 ( .A(n14506), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14508) );
  XNOR2_X1 U16310 ( .A(n14508), .B(n14507), .ZN(n14547) );
  NAND2_X1 U16311 ( .A1(n14548), .A2(n14547), .ZN(n14509) );
  XOR2_X1 U16312 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14511), .Z(n15547) );
  NAND2_X1 U16313 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14512), .ZN(n14513) );
  XNOR2_X1 U16314 ( .A(n14517), .B(n14516), .ZN(n14519) );
  NAND2_X1 U16315 ( .A1(n14518), .A2(n14519), .ZN(n14520) );
  NOR2_X1 U16316 ( .A1(n14553), .A2(n14552), .ZN(n14521) );
  INV_X1 U16317 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U16318 ( .A1(n14553), .A2(n14552), .ZN(n14551) );
  NOR2_X1 U16319 ( .A1(n14682), .A2(n14683), .ZN(n14522) );
  INV_X1 U16320 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14989) );
  NAND2_X1 U16321 ( .A1(n14682), .A2(n14683), .ZN(n14681) );
  OAI21_X1 U16322 ( .B1(n14522), .B2(n14989), .A(n14681), .ZN(n14526) );
  XNOR2_X1 U16323 ( .A(n14524), .B(n14523), .ZN(n14525) );
  NOR2_X1 U16324 ( .A1(n14526), .A2(n14525), .ZN(n14527) );
  XNOR2_X1 U16325 ( .A(n14526), .B(n14525), .ZN(n14685) );
  XOR2_X1 U16326 ( .A(n15504), .B(P3_ADDR_REG_14__SCAN_IN), .Z(n14529) );
  XNOR2_X1 U16327 ( .A(n14529), .B(n14528), .ZN(n14691) );
  AND2_X1 U16328 ( .A1(n14690), .A2(n14691), .ZN(n14531) );
  OAI21_X1 U16329 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n14531), .A(n14530), 
        .ZN(n14534) );
  XNOR2_X1 U16330 ( .A(n14730), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n14532) );
  XOR2_X1 U16331 ( .A(n14533), .B(n14532), .Z(n14535) );
  NAND2_X1 U16332 ( .A1(n14697), .A2(n14698), .ZN(n14536) );
  XOR2_X1 U16333 ( .A(n14538), .B(n14537), .Z(n14568) );
  NAND2_X1 U16334 ( .A1(n14569), .A2(n14568), .ZN(n14539) );
  NOR2_X1 U16335 ( .A1(n14569), .A2(n14568), .ZN(n14567) );
  XOR2_X1 U16336 ( .A(n15313), .B(n14571), .Z(SUB_1596_U62) );
  AOI21_X1 U16337 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14541) );
  OAI21_X1 U16338 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14541), 
        .ZN(U28) );
  AOI21_X1 U16339 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14542) );
  OAI21_X1 U16340 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14542), 
        .ZN(U29) );
  AOI21_X1 U16341 ( .B1(n14545), .B2(n14544), .A(n14543), .ZN(n14546) );
  XOR2_X1 U16342 ( .A(n14546), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16343 ( .A(n14548), .B(n14547), .Z(SUB_1596_U57) );
  XNOR2_X1 U16344 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14549), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16345 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14550), .Z(SUB_1596_U54) );
  OAI21_X1 U16346 ( .B1(n14553), .B2(n14552), .A(n14551), .ZN(n14555) );
  XOR2_X1 U16347 ( .A(n14555), .B(n14554), .Z(SUB_1596_U70) );
  INV_X1 U16348 ( .A(n14557), .ZN(n14563) );
  NOR2_X1 U16349 ( .A1(n14557), .A2(n14879), .ZN(n14562) );
  OAI211_X1 U16350 ( .C1(n14560), .C2(n14899), .A(n14559), .B(n14558), .ZN(
        n14561) );
  AOI211_X1 U16351 ( .C1(n14563), .C2(n14882), .A(n14562), .B(n14561), .ZN(
        n14566) );
  INV_X1 U16352 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16353 ( .A1(n14909), .A2(n14566), .B1(n14564), .B2(n14908), .ZN(
        P1_U3495) );
  AOI22_X1 U16354 ( .A1(n14929), .A2(n14566), .B1(n14565), .B2(n14926), .ZN(
        P1_U3540) );
  AOI21_X1 U16355 ( .B1(n14569), .B2(n14568), .A(n14567), .ZN(n14570) );
  XOR2_X1 U16356 ( .A(n14570), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16357 ( .A1(n14575), .A2(n14574), .ZN(n14576) );
  AOI21_X1 U16358 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14577), .A(n14576), 
        .ZN(n14581) );
  XNOR2_X1 U16359 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14579) );
  XNOR2_X1 U16360 ( .A(n14579), .B(n14578), .ZN(n14580) );
  AOI22_X1 U16361 ( .A1(n14617), .A2(n14583), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14582), .ZN(n14585) );
  NAND2_X1 U16362 ( .A1(n14585), .A2(n14584), .ZN(P3_U3203) );
  NAND2_X1 U16363 ( .A1(n15150), .A2(n14586), .ZN(n14600) );
  NAND2_X1 U16364 ( .A1(n14600), .A2(n14587), .ZN(n14589) );
  NAND2_X1 U16365 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  XNOR2_X1 U16366 ( .A(n14590), .B(n14594), .ZN(n14592) );
  AOI222_X1 U16367 ( .A1(n15149), .A2(n14592), .B1(n14591), .B2(n15155), .C1(
        n15156), .C2(n15154), .ZN(n14619) );
  AOI22_X1 U16368 ( .A1(n14582), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15178), 
        .B2(n14593), .ZN(n14599) );
  XNOR2_X1 U16369 ( .A(n14595), .B(n14594), .ZN(n14622) );
  INV_X1 U16370 ( .A(n14596), .ZN(n15161) );
  NOR2_X1 U16371 ( .A1(n14597), .A2(n15183), .ZN(n14621) );
  AOI22_X1 U16372 ( .A1(n14622), .A2(n14611), .B1(n15161), .B2(n14621), .ZN(
        n14598) );
  OAI211_X1 U16373 ( .C1(n14582), .C2(n14619), .A(n14599), .B(n14598), .ZN(
        P3_U3221) );
  XOR2_X1 U16374 ( .A(n14608), .B(n14600), .Z(n14601) );
  OAI222_X1 U16375 ( .A1(n15193), .A2(n14603), .B1(n15195), .B2(n14602), .C1(
        n14601), .C2(n15191), .ZN(n14624) );
  INV_X1 U16376 ( .A(n14604), .ZN(n14605) );
  OAI22_X1 U16377 ( .A1(n15198), .A2(n14606), .B1(n15184), .B2(n14605), .ZN(
        n14614) );
  OAI21_X1 U16378 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14626) );
  NOR2_X1 U16379 ( .A1(n14610), .A2(n15183), .ZN(n14625) );
  AOI22_X1 U16380 ( .A1(n14626), .A2(n14611), .B1(n15161), .B2(n14625), .ZN(
        n14612) );
  INV_X1 U16381 ( .A(n14612), .ZN(n14613) );
  AOI211_X1 U16382 ( .C1(n15198), .C2(n14624), .A(n14614), .B(n14613), .ZN(
        n14615) );
  INV_X1 U16383 ( .A(n14615), .ZN(P3_U3222) );
  AOI21_X1 U16384 ( .B1(n14617), .B2(n15210), .A(n14616), .ZN(n14629) );
  AOI22_X1 U16385 ( .A1(n15235), .A2(n14629), .B1(n14618), .B2(n15233), .ZN(
        P3_U3489) );
  INV_X1 U16386 ( .A(n14619), .ZN(n14620) );
  AOI211_X1 U16387 ( .C1(n14622), .C2(n15221), .A(n14621), .B(n14620), .ZN(
        n14631) );
  AOI22_X1 U16388 ( .A1(n15235), .A2(n14631), .B1(n14623), .B2(n15233), .ZN(
        P3_U3471) );
  AOI211_X1 U16389 ( .C1(n15221), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        n14632) );
  INV_X1 U16390 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U16391 ( .A1(n15235), .A2(n14632), .B1(n14627), .B2(n15233), .ZN(
        P3_U3470) );
  INV_X1 U16392 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U16393 ( .A1(n15225), .A2(n14629), .B1(n14628), .B2(n15223), .ZN(
        P3_U3457) );
  INV_X1 U16394 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14630) );
  AOI22_X1 U16395 ( .A1(n15225), .A2(n14631), .B1(n14630), .B2(n15223), .ZN(
        P3_U3426) );
  INV_X1 U16396 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U16397 ( .A1(n15225), .A2(n14632), .B1(n15449), .B2(n15223), .ZN(
        P3_U3423) );
  OAI21_X1 U16398 ( .B1(n14634), .B2(n15097), .A(n14633), .ZN(n14635) );
  AOI211_X1 U16399 ( .C1(n14637), .C2(n15102), .A(n14636), .B(n14635), .ZN(
        n14644) );
  AOI22_X1 U16400 ( .A1(n15141), .A2(n14644), .B1(n9438), .B2(n15139), .ZN(
        P2_U3512) );
  INV_X1 U16401 ( .A(n14638), .ZN(n14643) );
  OAI21_X1 U16402 ( .B1(n14640), .B2(n15097), .A(n14639), .ZN(n14642) );
  AOI211_X1 U16403 ( .C1(n15088), .C2(n14643), .A(n14642), .B(n14641), .ZN(
        n14645) );
  AOI22_X1 U16404 ( .A1(n15141), .A2(n14645), .B1(n8662), .B2(n15139), .ZN(
        P2_U3511) );
  AOI22_X1 U16405 ( .A1(n15129), .A2(n14644), .B1(n8683), .B2(n15127), .ZN(
        P2_U3469) );
  INV_X1 U16406 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U16407 ( .A1(n15129), .A2(n14645), .B1(n15421), .B2(n15127), .ZN(
        P2_U3466) );
  OAI21_X1 U16408 ( .B1(n14647), .B2(n14899), .A(n14646), .ZN(n14650) );
  INV_X1 U16409 ( .A(n14648), .ZN(n14649) );
  AOI211_X1 U16410 ( .C1(n14651), .C2(n14906), .A(n14650), .B(n14649), .ZN(
        n14674) );
  AOI22_X1 U16411 ( .A1(n14929), .A2(n14674), .B1(n14652), .B2(n14926), .ZN(
        P1_U3544) );
  AOI211_X1 U16412 ( .C1(n14876), .C2(n11297), .A(n14654), .B(n14653), .ZN(
        n14658) );
  NAND3_X1 U16413 ( .A1(n6615), .A2(n14655), .A3(n14906), .ZN(n14656) );
  AOI22_X1 U16414 ( .A1(n14929), .A2(n14676), .B1(n15332), .B2(n14926), .ZN(
        P1_U3542) );
  AOI21_X1 U16415 ( .B1(n14660), .B2(n14876), .A(n14659), .ZN(n14662) );
  OAI211_X1 U16416 ( .C1(n14663), .C2(n14863), .A(n14662), .B(n14661), .ZN(
        n14664) );
  AOI21_X1 U16417 ( .B1(n14665), .B2(n14906), .A(n14664), .ZN(n14678) );
  AOI22_X1 U16418 ( .A1(n14929), .A2(n14678), .B1(n10579), .B2(n14926), .ZN(
        P1_U3541) );
  AND2_X1 U16419 ( .A1(n14666), .A2(n14906), .ZN(n14671) );
  INV_X1 U16420 ( .A(n14667), .ZN(n14668) );
  OAI22_X1 U16421 ( .A1(n14669), .A2(n14837), .B1(n14668), .B2(n14899), .ZN(
        n14670) );
  NOR3_X1 U16422 ( .A1(n14672), .A2(n14671), .A3(n14670), .ZN(n14680) );
  AOI22_X1 U16423 ( .A1(n14929), .A2(n14680), .B1(n14673), .B2(n14926), .ZN(
        P1_U3539) );
  INV_X1 U16424 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U16425 ( .A1(n14909), .A2(n14674), .B1(n15490), .B2(n14908), .ZN(
        P1_U3507) );
  INV_X1 U16426 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14675) );
  AOI22_X1 U16427 ( .A1(n14909), .A2(n14676), .B1(n14675), .B2(n14908), .ZN(
        P1_U3501) );
  INV_X1 U16428 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14677) );
  AOI22_X1 U16429 ( .A1(n14909), .A2(n14678), .B1(n14677), .B2(n14908), .ZN(
        P1_U3498) );
  INV_X1 U16430 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14679) );
  AOI22_X1 U16431 ( .A1(n14909), .A2(n14680), .B1(n14679), .B2(n14908), .ZN(
        P1_U3492) );
  OAI21_X1 U16432 ( .B1(n14683), .B2(n14682), .A(n14681), .ZN(n14684) );
  XOR2_X1 U16433 ( .A(n14684), .B(n14989), .Z(SUB_1596_U69) );
  INV_X1 U16434 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15005) );
  XOR2_X1 U16435 ( .A(n15005), .B(n14685), .Z(SUB_1596_U68) );
  AOI21_X1 U16436 ( .B1(n6721), .B2(n14687), .A(n14686), .ZN(n14688) );
  XOR2_X1 U16437 ( .A(n14688), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16438 ( .B1(n14691), .B2(n14690), .A(n14689), .ZN(n14692) );
  XOR2_X1 U16439 ( .A(n14692), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16440 ( .A1(n14694), .A2(n14693), .ZN(n14695) );
  XOR2_X1 U16441 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14695), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16442 ( .B1(n14698), .B2(n14697), .A(n14696), .ZN(n14699) );
  XOR2_X1 U16443 ( .A(n14699), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  INV_X1 U16444 ( .A(n14700), .ZN(n14703) );
  MUX2_X1 U16445 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14927), .S(n14704), .Z(
        n14702) );
  OAI211_X1 U16446 ( .C1(n14703), .C2(n14702), .A(n14738), .B(n14701), .ZN(
        n14711) );
  MUX2_X1 U16447 ( .A(n10156), .B(P1_REG2_REG_10__SCAN_IN), .S(n14704), .Z(
        n14705) );
  NAND3_X1 U16448 ( .A1(n14707), .A2(n14706), .A3(n14705), .ZN(n14708) );
  NAND3_X1 U16449 ( .A1(n14733), .A2(n14709), .A3(n14708), .ZN(n14710) );
  OAI211_X1 U16450 ( .C1(n14725), .C2(n14712), .A(n14711), .B(n14710), .ZN(
        n14713) );
  AOI211_X1 U16451 ( .C1(P1_ADDR_REG_10__SCAN_IN), .C2(n14731), .A(n14714), 
        .B(n14713), .ZN(n14715) );
  INV_X1 U16452 ( .A(n14715), .ZN(P1_U3253) );
  AOI21_X1 U16453 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14717), .A(n14716), 
        .ZN(n14722) );
  AOI21_X1 U16454 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14719), .A(n14718), 
        .ZN(n14720) );
  OAI222_X1 U16455 ( .A1(n14725), .A2(n14724), .B1(n14723), .B2(n14722), .C1(
        n14721), .C2(n14720), .ZN(n14726) );
  INV_X1 U16456 ( .A(n14726), .ZN(n14728) );
  NAND2_X1 U16457 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14727)
         );
  OAI211_X1 U16458 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        P1_U3258) );
  AOI22_X1 U16459 ( .A1(n14731), .A2(P1_ADDR_REG_18__SCAN_IN), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(P1_U3086), .ZN(n14743) );
  OAI211_X1 U16460 ( .C1(n14734), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14733), 
        .B(n14732), .ZN(n14742) );
  NAND2_X1 U16461 ( .A1(n14736), .A2(n14735), .ZN(n14741) );
  OAI211_X1 U16462 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14739), .A(n14738), 
        .B(n14737), .ZN(n14740) );
  NAND4_X1 U16463 ( .A1(n14743), .A2(n14742), .A3(n14741), .A4(n14740), .ZN(
        P1_U3261) );
  XNOR2_X1 U16464 ( .A(n14744), .B(n14746), .ZN(n14888) );
  XNOR2_X1 U16465 ( .A(n14745), .B(n14746), .ZN(n14752) );
  AOI22_X1 U16466 ( .A1(n14750), .A2(n14749), .B1(n14748), .B2(n14747), .ZN(
        n14751) );
  OAI21_X1 U16467 ( .B1(n14752), .B2(n14863), .A(n14751), .ZN(n14753) );
  AOI21_X1 U16468 ( .B1(n14882), .B2(n14888), .A(n14753), .ZN(n14885) );
  NOR2_X1 U16469 ( .A1(n14783), .A2(n14754), .ZN(n14755) );
  AOI21_X1 U16470 ( .B1(n14797), .B2(P1_REG2_REG_7__SCAN_IN), .A(n14755), .ZN(
        n14756) );
  OAI21_X1 U16471 ( .B1(n14786), .B2(n7065), .A(n14756), .ZN(n14757) );
  INV_X1 U16472 ( .A(n14757), .ZN(n14761) );
  OAI211_X1 U16473 ( .C1(n6731), .C2(n7065), .A(n14790), .B(n14758), .ZN(
        n14884) );
  INV_X1 U16474 ( .A(n14884), .ZN(n14759) );
  AOI22_X1 U16475 ( .A1(n14888), .A2(n14794), .B1(n14793), .B2(n14759), .ZN(
        n14760) );
  OAI211_X1 U16476 ( .C1(n14797), .C2(n14885), .A(n14761), .B(n14760), .ZN(
        P1_U3286) );
  XNOR2_X1 U16477 ( .A(n14762), .B(n14764), .ZN(n14872) );
  XNOR2_X1 U16478 ( .A(n14763), .B(n14764), .ZN(n14765) );
  NOR2_X1 U16479 ( .A1(n14765), .A2(n14863), .ZN(n14766) );
  AOI211_X1 U16480 ( .C1(n14882), .C2(n14872), .A(n14767), .B(n14766), .ZN(
        n14869) );
  NOR2_X1 U16481 ( .A1(n14783), .A2(n14768), .ZN(n14769) );
  AOI21_X1 U16482 ( .B1(n14797), .B2(P1_REG2_REG_5__SCAN_IN), .A(n14769), .ZN(
        n14770) );
  OAI21_X1 U16483 ( .B1(n14786), .B2(n14868), .A(n14770), .ZN(n14771) );
  INV_X1 U16484 ( .A(n14771), .ZN(n14776) );
  OAI211_X1 U16485 ( .C1(n14868), .C2(n14773), .A(n14772), .B(n14790), .ZN(
        n14867) );
  INV_X1 U16486 ( .A(n14867), .ZN(n14774) );
  AOI22_X1 U16487 ( .A1(n14872), .A2(n14794), .B1(n14793), .B2(n14774), .ZN(
        n14775) );
  OAI211_X1 U16488 ( .C1(n14797), .C2(n14869), .A(n14776), .B(n14775), .ZN(
        P1_U3288) );
  XNOR2_X1 U16489 ( .A(n14778), .B(n14777), .ZN(n14856) );
  XNOR2_X1 U16490 ( .A(n14779), .B(n14778), .ZN(n14780) );
  NOR2_X1 U16491 ( .A1(n14780), .A2(n14863), .ZN(n14781) );
  AOI211_X1 U16492 ( .C1(n14882), .C2(n14856), .A(n14782), .B(n14781), .ZN(
        n14853) );
  NOR2_X1 U16493 ( .A1(n14783), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n14784) );
  AOI21_X1 U16494 ( .B1(n14797), .B2(P1_REG2_REG_3__SCAN_IN), .A(n14784), .ZN(
        n14785) );
  OAI21_X1 U16495 ( .B1(n14786), .B2(n14852), .A(n14785), .ZN(n14787) );
  INV_X1 U16496 ( .A(n14787), .ZN(n14796) );
  INV_X1 U16497 ( .A(n14788), .ZN(n14791) );
  OAI211_X1 U16498 ( .C1(n14791), .C2(n14852), .A(n14790), .B(n14789), .ZN(
        n14851) );
  INV_X1 U16499 ( .A(n14851), .ZN(n14792) );
  AOI22_X1 U16500 ( .A1(n14856), .A2(n14794), .B1(n14793), .B2(n14792), .ZN(
        n14795) );
  OAI211_X1 U16501 ( .C1(n14797), .C2(n14853), .A(n14796), .B(n14795), .ZN(
        P1_U3290) );
  INV_X1 U16502 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14798) );
  NOR2_X1 U16503 ( .A1(n14825), .A2(n14798), .ZN(P1_U3294) );
  INV_X1 U16504 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14799) );
  NOR2_X1 U16505 ( .A1(n14825), .A2(n14799), .ZN(P1_U3295) );
  INV_X1 U16506 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14800) );
  NOR2_X1 U16507 ( .A1(n14825), .A2(n14800), .ZN(P1_U3296) );
  INV_X1 U16508 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14801) );
  NOR2_X1 U16509 ( .A1(n14810), .A2(n14801), .ZN(P1_U3297) );
  INV_X1 U16510 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14802) );
  NOR2_X1 U16511 ( .A1(n14810), .A2(n14802), .ZN(P1_U3298) );
  INV_X1 U16512 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14803) );
  NOR2_X1 U16513 ( .A1(n14810), .A2(n14803), .ZN(P1_U3299) );
  INV_X1 U16514 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14804) );
  NOR2_X1 U16515 ( .A1(n14810), .A2(n14804), .ZN(P1_U3300) );
  INV_X1 U16516 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14805) );
  NOR2_X1 U16517 ( .A1(n14810), .A2(n14805), .ZN(P1_U3301) );
  INV_X1 U16518 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14806) );
  NOR2_X1 U16519 ( .A1(n14810), .A2(n14806), .ZN(P1_U3302) );
  NOR2_X1 U16520 ( .A1(n14810), .A2(n15423), .ZN(P1_U3303) );
  INV_X1 U16521 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14807) );
  NOR2_X1 U16522 ( .A1(n14810), .A2(n14807), .ZN(P1_U3304) );
  NOR2_X1 U16523 ( .A1(n14810), .A2(n15402), .ZN(P1_U3305) );
  INV_X1 U16524 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14808) );
  NOR2_X1 U16525 ( .A1(n14810), .A2(n14808), .ZN(P1_U3306) );
  INV_X1 U16526 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14809) );
  NOR2_X1 U16527 ( .A1(n14810), .A2(n14809), .ZN(P1_U3307) );
  NOR2_X1 U16528 ( .A1(n14810), .A2(n15305), .ZN(P1_U3308) );
  NOR2_X1 U16529 ( .A1(n14825), .A2(n15521), .ZN(P1_U3309) );
  INV_X1 U16530 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14811) );
  NOR2_X1 U16531 ( .A1(n14825), .A2(n14811), .ZN(P1_U3310) );
  INV_X1 U16532 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14812) );
  NOR2_X1 U16533 ( .A1(n14825), .A2(n14812), .ZN(P1_U3311) );
  INV_X1 U16534 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14813) );
  NOR2_X1 U16535 ( .A1(n14825), .A2(n14813), .ZN(P1_U3312) );
  INV_X1 U16536 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14814) );
  NOR2_X1 U16537 ( .A1(n14825), .A2(n14814), .ZN(P1_U3313) );
  INV_X1 U16538 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U16539 ( .A1(n14825), .A2(n14815), .ZN(P1_U3314) );
  INV_X1 U16540 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14816) );
  NOR2_X1 U16541 ( .A1(n14825), .A2(n14816), .ZN(P1_U3315) );
  INV_X1 U16542 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14817) );
  NOR2_X1 U16543 ( .A1(n14825), .A2(n14817), .ZN(P1_U3316) );
  INV_X1 U16544 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14818) );
  NOR2_X1 U16545 ( .A1(n14825), .A2(n14818), .ZN(P1_U3317) );
  INV_X1 U16546 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14819) );
  NOR2_X1 U16547 ( .A1(n14825), .A2(n14819), .ZN(P1_U3318) );
  INV_X1 U16548 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14820) );
  NOR2_X1 U16549 ( .A1(n14825), .A2(n14820), .ZN(P1_U3319) );
  INV_X1 U16550 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14821) );
  NOR2_X1 U16551 ( .A1(n14825), .A2(n14821), .ZN(P1_U3320) );
  INV_X1 U16552 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14822) );
  NOR2_X1 U16553 ( .A1(n14825), .A2(n14822), .ZN(P1_U3321) );
  INV_X1 U16554 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14823) );
  NOR2_X1 U16555 ( .A1(n14825), .A2(n14823), .ZN(P1_U3322) );
  INV_X1 U16556 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14824) );
  NOR2_X1 U16557 ( .A1(n14825), .A2(n14824), .ZN(P1_U3323) );
  INV_X1 U16558 ( .A(n14826), .ZN(n14830) );
  AOI21_X1 U16559 ( .B1(n14828), .B2(n14863), .A(n14827), .ZN(n14829) );
  AOI211_X1 U16560 ( .C1(n14832), .C2(n14831), .A(n14830), .B(n14829), .ZN(
        n14910) );
  AOI22_X1 U16561 ( .A1(n14909), .A2(n14910), .B1(n9239), .B2(n14908), .ZN(
        P1_U3459) );
  INV_X1 U16562 ( .A(n14833), .ZN(n14842) );
  NAND2_X1 U16563 ( .A1(n14876), .A2(n14834), .ZN(n14835) );
  OAI211_X1 U16564 ( .C1(n14838), .C2(n14837), .A(n14836), .B(n14835), .ZN(
        n14841) );
  INV_X1 U16565 ( .A(n14839), .ZN(n14840) );
  AOI211_X1 U16566 ( .C1(n14842), .C2(n14906), .A(n14841), .B(n14840), .ZN(
        n14912) );
  INV_X1 U16567 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14843) );
  AOI22_X1 U16568 ( .A1(n14909), .A2(n14912), .B1(n14843), .B2(n14908), .ZN(
        P1_U3462) );
  INV_X1 U16569 ( .A(n14844), .ZN(n14850) );
  NOR2_X1 U16570 ( .A1(n14844), .A2(n14879), .ZN(n14849) );
  OAI211_X1 U16571 ( .C1(n14847), .C2(n14899), .A(n14846), .B(n14845), .ZN(
        n14848) );
  AOI211_X1 U16572 ( .C1(n14850), .C2(n14882), .A(n14849), .B(n14848), .ZN(
        n14914) );
  AOI22_X1 U16573 ( .A1(n14909), .A2(n14914), .B1(n9306), .B2(n14908), .ZN(
        P1_U3465) );
  INV_X1 U16574 ( .A(n14879), .ZN(n14889) );
  OAI21_X1 U16575 ( .B1(n14852), .B2(n14899), .A(n14851), .ZN(n14855) );
  INV_X1 U16576 ( .A(n14853), .ZN(n14854) );
  AOI211_X1 U16577 ( .C1(n14889), .C2(n14856), .A(n14855), .B(n14854), .ZN(
        n14916) );
  INV_X1 U16578 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U16579 ( .A1(n14909), .A2(n14916), .B1(n14857), .B2(n14908), .ZN(
        P1_U3468) );
  AOI211_X1 U16580 ( .C1(n14876), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14861) );
  OAI21_X1 U16581 ( .B1(n14863), .B2(n14862), .A(n14861), .ZN(n14864) );
  AOI21_X1 U16582 ( .B1(n14865), .B2(n14906), .A(n14864), .ZN(n14918) );
  INV_X1 U16583 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U16584 ( .A1(n14909), .A2(n14918), .B1(n14866), .B2(n14908), .ZN(
        P1_U3471) );
  OAI21_X1 U16585 ( .B1(n14868), .B2(n14899), .A(n14867), .ZN(n14871) );
  INV_X1 U16586 ( .A(n14869), .ZN(n14870) );
  AOI211_X1 U16587 ( .C1(n14889), .C2(n14872), .A(n14871), .B(n14870), .ZN(
        n14920) );
  INV_X1 U16588 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U16589 ( .A1(n14909), .A2(n14920), .B1(n15355), .B2(n14908), .ZN(
        P1_U3474) );
  INV_X1 U16590 ( .A(n14878), .ZN(n14881) );
  AOI211_X1 U16591 ( .C1(n14876), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        n14877) );
  OAI21_X1 U16592 ( .B1(n14879), .B2(n14878), .A(n14877), .ZN(n14880) );
  AOI21_X1 U16593 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14922) );
  INV_X1 U16594 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U16595 ( .A1(n14909), .A2(n14922), .B1(n14883), .B2(n14908), .ZN(
        P1_U3477) );
  OAI21_X1 U16596 ( .B1(n7065), .B2(n14899), .A(n14884), .ZN(n14887) );
  INV_X1 U16597 ( .A(n14885), .ZN(n14886) );
  AOI211_X1 U16598 ( .C1(n14889), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n14924) );
  INV_X1 U16599 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14890) );
  AOI22_X1 U16600 ( .A1(n14909), .A2(n14924), .B1(n14890), .B2(n14908), .ZN(
        P1_U3480) );
  OAI211_X1 U16601 ( .C1(n7064), .C2(n14899), .A(n14893), .B(n14892), .ZN(
        n14894) );
  AOI21_X1 U16602 ( .B1(n14895), .B2(n14906), .A(n14894), .ZN(n14925) );
  INV_X1 U16603 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14896) );
  AOI22_X1 U16604 ( .A1(n14909), .A2(n14925), .B1(n14896), .B2(n14908), .ZN(
        P1_U3483) );
  OAI211_X1 U16605 ( .C1(n14900), .C2(n14899), .A(n14898), .B(n14897), .ZN(
        n14905) );
  AND3_X1 U16606 ( .A1(n14903), .A2(n14902), .A3(n14901), .ZN(n14904) );
  AOI211_X1 U16607 ( .C1(n14907), .C2(n14906), .A(n14905), .B(n14904), .ZN(
        n14928) );
  INV_X1 U16608 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U16609 ( .A1(n14909), .A2(n14928), .B1(n15390), .B2(n14908), .ZN(
        P1_U3489) );
  AOI22_X1 U16610 ( .A1(n14929), .A2(n14910), .B1(n9237), .B2(n14926), .ZN(
        P1_U3528) );
  AOI22_X1 U16611 ( .A1(n14929), .A2(n14912), .B1(n14911), .B2(n14926), .ZN(
        P1_U3529) );
  AOI22_X1 U16612 ( .A1(n14929), .A2(n14914), .B1(n14913), .B2(n14926), .ZN(
        P1_U3530) );
  AOI22_X1 U16613 ( .A1(n14929), .A2(n14916), .B1(n14915), .B2(n14926), .ZN(
        P1_U3531) );
  AOI22_X1 U16614 ( .A1(n14929), .A2(n14918), .B1(n14917), .B2(n14926), .ZN(
        P1_U3532) );
  AOI22_X1 U16615 ( .A1(n14929), .A2(n14920), .B1(n14919), .B2(n14926), .ZN(
        P1_U3533) );
  AOI22_X1 U16616 ( .A1(n14929), .A2(n14922), .B1(n14921), .B2(n14926), .ZN(
        P1_U3534) );
  AOI22_X1 U16617 ( .A1(n14929), .A2(n14924), .B1(n14923), .B2(n14926), .ZN(
        P1_U3535) );
  AOI22_X1 U16618 ( .A1(n14929), .A2(n14925), .B1(n10126), .B2(n14926), .ZN(
        P1_U3536) );
  AOI22_X1 U16619 ( .A1(n14929), .A2(n14928), .B1(n14927), .B2(n14926), .ZN(
        P1_U3538) );
  NOR2_X1 U16620 ( .A1(n14949), .A2(n14930), .ZN(P2_U3087) );
  OAI22_X1 U16621 ( .A1(n14934), .A2(n14933), .B1(n14932), .B2(n14931), .ZN(
        n14942) );
  NAND2_X1 U16622 ( .A1(n14937), .A2(n14938), .ZN(n14940) );
  AOI21_X1 U16623 ( .B1(n14936), .B2(n14940), .A(n14939), .ZN(n14941) );
  AOI211_X1 U16624 ( .C1(n14944), .C2(n14943), .A(n14942), .B(n14941), .ZN(
        n14945) );
  NAND2_X1 U16625 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15003)
         );
  OAI211_X1 U16626 ( .C1(n14947), .C2(n14946), .A(n14945), .B(n15003), .ZN(
        P2_U3196) );
  AOI22_X1 U16627 ( .A1(n14949), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14961) );
  OAI211_X1 U16628 ( .C1(n14952), .C2(n14951), .A(n15002), .B(n14950), .ZN(
        n14953) );
  OAI21_X1 U16629 ( .B1(n14996), .B2(n14954), .A(n14953), .ZN(n14955) );
  INV_X1 U16630 ( .A(n14955), .ZN(n14960) );
  XOR2_X1 U16631 ( .A(n14957), .B(n14956), .Z(n14958) );
  NAND2_X1 U16632 ( .A1(n15027), .A2(n14958), .ZN(n14959) );
  NAND3_X1 U16633 ( .A1(n14961), .A2(n14960), .A3(n14959), .ZN(P2_U3216) );
  OAI211_X1 U16634 ( .C1(n14964), .C2(n14963), .A(n15002), .B(n14962), .ZN(
        n14966) );
  OAI211_X1 U16635 ( .C1(n14996), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n14968) );
  INV_X1 U16636 ( .A(n14968), .ZN(n14973) );
  OAI211_X1 U16637 ( .C1(n14971), .C2(n14970), .A(n15027), .B(n14969), .ZN(
        n14972) );
  OAI211_X1 U16638 ( .C1(n15032), .C2(n14974), .A(n14973), .B(n14972), .ZN(
        P2_U3220) );
  OAI21_X1 U16639 ( .B1(n14976), .B2(n14975), .A(n15002), .ZN(n14984) );
  NOR2_X1 U16640 ( .A1(n14978), .A2(n14977), .ZN(n14979) );
  OAI21_X1 U16641 ( .B1(n14980), .B2(n14979), .A(n15027), .ZN(n14983) );
  NAND2_X1 U16642 ( .A1(n15025), .A2(n14981), .ZN(n14982) );
  OAI211_X1 U16643 ( .C1(n14985), .C2(n14984), .A(n14983), .B(n14982), .ZN(
        n14986) );
  INV_X1 U16644 ( .A(n14986), .ZN(n14988) );
  OAI211_X1 U16645 ( .C1(n14989), .C2(n15032), .A(n14988), .B(n14987), .ZN(
        P2_U3225) );
  OAI21_X1 U16646 ( .B1(n14992), .B2(n14991), .A(n14990), .ZN(n15001) );
  AOI21_X1 U16647 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14999) );
  OAI22_X1 U16648 ( .A1(n14999), .A2(n14998), .B1(n14997), .B2(n14996), .ZN(
        n15000) );
  AOI21_X1 U16649 ( .B1(n15002), .B2(n15001), .A(n15000), .ZN(n15004) );
  OAI211_X1 U16650 ( .C1(n15005), .C2(n15032), .A(n15004), .B(n15003), .ZN(
        P2_U3226) );
  NOR2_X1 U16651 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8680), .ZN(n15010) );
  AOI211_X1 U16652 ( .C1(n15008), .C2(n15007), .A(n15006), .B(n15018), .ZN(
        n15009) );
  AOI211_X1 U16653 ( .C1(n15025), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        n15016) );
  OAI211_X1 U16654 ( .C1(n15014), .C2(n15013), .A(n15027), .B(n15012), .ZN(
        n15015) );
  OAI211_X1 U16655 ( .C1(n15032), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        P2_U3227) );
  NOR2_X1 U16656 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15518), .ZN(n15023) );
  AOI211_X1 U16657 ( .C1(n15021), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15022) );
  AOI211_X1 U16658 ( .C1(n15025), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15031) );
  OAI211_X1 U16659 ( .C1(n15029), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        n15030) );
  OAI211_X1 U16660 ( .C1(n15032), .C2(n15320), .A(n15031), .B(n15030), .ZN(
        P2_U3230) );
  INV_X1 U16661 ( .A(n15042), .ZN(n15059) );
  INV_X1 U16662 ( .A(n15033), .ZN(n15034) );
  AND2_X1 U16663 ( .A1(n15035), .A2(n15034), .ZN(n15058) );
  NAND2_X1 U16664 ( .A1(n15058), .A2(n12351), .ZN(n15036) );
  OAI21_X1 U16665 ( .B1(n15038), .B2(n15037), .A(n15036), .ZN(n15043) );
  NOR2_X1 U16666 ( .A1(n15126), .A2(n13683), .ZN(n15041) );
  OAI22_X1 U16667 ( .A1(n15042), .A2(n15041), .B1(n15040), .B2(n15039), .ZN(
        n15057) );
  AOI211_X1 U16668 ( .C1(n15059), .C2(n15044), .A(n15043), .B(n15057), .ZN(
        n15046) );
  AOI22_X1 U16669 ( .A1(n6578), .A2(n15047), .B1(n15046), .B2(n15045), .ZN(
        P2_U3265) );
  INV_X1 U16670 ( .A(n15049), .ZN(n15050) );
  AND2_X1 U16671 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15050), .ZN(P2_U3266) );
  AND2_X1 U16672 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15050), .ZN(P2_U3267) );
  AND2_X1 U16673 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15050), .ZN(P2_U3268) );
  AND2_X1 U16674 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15050), .ZN(P2_U3269) );
  AND2_X1 U16675 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15050), .ZN(P2_U3270) );
  AND2_X1 U16676 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15050), .ZN(P2_U3271) );
  AND2_X1 U16677 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15050), .ZN(P2_U3272) );
  AND2_X1 U16678 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15050), .ZN(P2_U3273) );
  AND2_X1 U16679 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15050), .ZN(P2_U3274) );
  AND2_X1 U16680 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15050), .ZN(P2_U3275) );
  AND2_X1 U16681 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15050), .ZN(P2_U3276) );
  INV_X1 U16682 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15459) );
  NOR2_X1 U16683 ( .A1(n15049), .A2(n15459), .ZN(P2_U3277) );
  AND2_X1 U16684 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15050), .ZN(P2_U3278) );
  AND2_X1 U16685 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15050), .ZN(P2_U3279) );
  AND2_X1 U16686 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15050), .ZN(P2_U3280) );
  INV_X1 U16687 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U16688 ( .A1(n15049), .A2(n15335), .ZN(P2_U3281) );
  AND2_X1 U16689 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15050), .ZN(P2_U3282) );
  AND2_X1 U16690 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15050), .ZN(P2_U3283) );
  AND2_X1 U16691 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15050), .ZN(P2_U3284) );
  AND2_X1 U16692 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15050), .ZN(P2_U3285) );
  AND2_X1 U16693 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15050), .ZN(P2_U3286) );
  AND2_X1 U16694 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15050), .ZN(P2_U3287) );
  AND2_X1 U16695 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15050), .ZN(P2_U3288) );
  AND2_X1 U16696 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15050), .ZN(P2_U3289) );
  INV_X1 U16697 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15437) );
  NOR2_X1 U16698 ( .A1(n15049), .A2(n15437), .ZN(P2_U3290) );
  AND2_X1 U16699 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15050), .ZN(P2_U3291) );
  AND2_X1 U16700 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15050), .ZN(P2_U3292) );
  AND2_X1 U16701 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15050), .ZN(P2_U3293) );
  AND2_X1 U16702 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15050), .ZN(P2_U3294) );
  AND2_X1 U16703 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15050), .ZN(P2_U3295) );
  AOI22_X1 U16704 ( .A1(n15056), .A2(n15053), .B1(n15052), .B2(n15051), .ZN(
        P2_U3416) );
  OAI21_X1 U16705 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(P2_U3417) );
  AOI211_X1 U16706 ( .C1(n15059), .C2(n15088), .A(n15058), .B(n15057), .ZN(
        n15130) );
  AOI22_X1 U16707 ( .A1(n15129), .A2(n15130), .B1(n8437), .B2(n15127), .ZN(
        P2_U3430) );
  AOI22_X1 U16708 ( .A1(n15129), .A2(n15060), .B1(n8427), .B2(n15127), .ZN(
        P2_U3433) );
  INV_X1 U16709 ( .A(n15065), .ZN(n15067) );
  AOI21_X1 U16710 ( .B1(n15118), .B2(n15062), .A(n15061), .ZN(n15063) );
  OAI211_X1 U16711 ( .C1(n15065), .C2(n12137), .A(n15064), .B(n15063), .ZN(
        n15066) );
  AOI21_X1 U16712 ( .B1(n15126), .B2(n15067), .A(n15066), .ZN(n15131) );
  AOI22_X1 U16713 ( .A1(n15129), .A2(n15131), .B1(n8450), .B2(n15127), .ZN(
        P2_U3436) );
  INV_X1 U16714 ( .A(n15072), .ZN(n15074) );
  AOI211_X1 U16715 ( .C1(n15118), .C2(n15070), .A(n15069), .B(n15068), .ZN(
        n15071) );
  OAI21_X1 U16716 ( .B1(n15072), .B2(n12137), .A(n15071), .ZN(n15073) );
  AOI21_X1 U16717 ( .B1(n15126), .B2(n15074), .A(n15073), .ZN(n15132) );
  AOI22_X1 U16718 ( .A1(n15129), .A2(n15132), .B1(n8487), .B2(n15127), .ZN(
        P2_U3439) );
  AND2_X1 U16719 ( .A1(n15075), .A2(n15118), .ZN(n15076) );
  NOR2_X1 U16720 ( .A1(n15077), .A2(n15076), .ZN(n15081) );
  OR2_X1 U16721 ( .A1(n15079), .A2(n15078), .ZN(n15080) );
  AND3_X1 U16722 ( .A1(n15082), .A2(n15081), .A3(n15080), .ZN(n15133) );
  AOI22_X1 U16723 ( .A1(n15129), .A2(n15133), .B1(n8501), .B2(n15127), .ZN(
        P2_U3442) );
  OAI21_X1 U16724 ( .B1(n15084), .B2(n15097), .A(n15083), .ZN(n15086) );
  AOI211_X1 U16725 ( .C1(n15088), .C2(n15087), .A(n15086), .B(n15085), .ZN(
        n15134) );
  AOI22_X1 U16726 ( .A1(n15129), .A2(n15134), .B1(n8515), .B2(n15127), .ZN(
        P2_U3445) );
  AOI21_X1 U16727 ( .B1(n15118), .B2(n15090), .A(n15089), .ZN(n15091) );
  OAI211_X1 U16728 ( .C1(n15093), .C2(n12137), .A(n15092), .B(n15091), .ZN(
        n15094) );
  INV_X1 U16729 ( .A(n15094), .ZN(n15135) );
  INV_X1 U16730 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15095) );
  AOI22_X1 U16731 ( .A1(n15129), .A2(n15135), .B1(n15095), .B2(n15127), .ZN(
        P2_U3448) );
  OAI21_X1 U16732 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15100) );
  AOI211_X1 U16733 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15136) );
  INV_X1 U16734 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U16735 ( .A1(n15129), .A2(n15136), .B1(n15481), .B2(n15127), .ZN(
        P2_U3451) );
  NAND2_X1 U16736 ( .A1(n15103), .A2(n15118), .ZN(n15104) );
  OAI211_X1 U16737 ( .C1(n15106), .C2(n12137), .A(n15105), .B(n15104), .ZN(
        n15107) );
  AOI211_X1 U16738 ( .C1(n15126), .C2(n15109), .A(n15108), .B(n15107), .ZN(
        n15137) );
  INV_X1 U16739 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15110) );
  AOI22_X1 U16740 ( .A1(n15129), .A2(n15137), .B1(n15110), .B2(n15127), .ZN(
        P2_U3454) );
  NAND2_X1 U16741 ( .A1(n15111), .A2(n15118), .ZN(n15112) );
  OAI211_X1 U16742 ( .C1(n15114), .C2(n12137), .A(n15113), .B(n15112), .ZN(
        n15117) );
  NOR2_X1 U16743 ( .A1(n15114), .A2(n9127), .ZN(n15116) );
  NOR3_X1 U16744 ( .A1(n15117), .A2(n15116), .A3(n15115), .ZN(n15138) );
  AOI22_X1 U16745 ( .A1(n15129), .A2(n15138), .B1(n8606), .B2(n15127), .ZN(
        P2_U3457) );
  NAND2_X1 U16746 ( .A1(n15119), .A2(n15118), .ZN(n15120) );
  OAI211_X1 U16747 ( .C1(n15122), .C2(n12137), .A(n15121), .B(n15120), .ZN(
        n15123) );
  AOI211_X1 U16748 ( .C1(n15126), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15140) );
  INV_X1 U16749 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16750 ( .A1(n15129), .A2(n15140), .B1(n15128), .B2(n15127), .ZN(
        P2_U3460) );
  AOI22_X1 U16751 ( .A1(n15141), .A2(n15130), .B1(n9045), .B2(n15139), .ZN(
        P2_U3499) );
  AOI22_X1 U16752 ( .A1(n15141), .A2(n15131), .B1(n8993), .B2(n15139), .ZN(
        P2_U3501) );
  AOI22_X1 U16753 ( .A1(n15141), .A2(n15132), .B1(n8995), .B2(n15139), .ZN(
        P2_U3502) );
  AOI22_X1 U16754 ( .A1(n15141), .A2(n15133), .B1(n8997), .B2(n15139), .ZN(
        P2_U3503) );
  AOI22_X1 U16755 ( .A1(n15141), .A2(n15134), .B1(n8514), .B2(n15139), .ZN(
        P2_U3504) );
  AOI22_X1 U16756 ( .A1(n15141), .A2(n15135), .B1(n8545), .B2(n15139), .ZN(
        P2_U3505) );
  AOI22_X1 U16757 ( .A1(n15141), .A2(n15136), .B1(n8560), .B2(n15139), .ZN(
        P2_U3506) );
  AOI22_X1 U16758 ( .A1(n15141), .A2(n15137), .B1(n8579), .B2(n15139), .ZN(
        P2_U3507) );
  AOI22_X1 U16759 ( .A1(n15141), .A2(n15138), .B1(n9431), .B2(n15139), .ZN(
        P2_U3508) );
  AOI22_X1 U16760 ( .A1(n15141), .A2(n15140), .B1(n9435), .B2(n15139), .ZN(
        P2_U3509) );
  NOR2_X1 U16761 ( .A1(P3_U3897), .A2(n15142), .ZN(P3_U3150) );
  NAND2_X1 U16762 ( .A1(n15144), .A2(n15143), .ZN(n15146) );
  AND2_X1 U16763 ( .A1(n15146), .A2(n15145), .ZN(n15148) );
  XNOR2_X1 U16764 ( .A(n15148), .B(n15147), .ZN(n15222) );
  OAI211_X1 U16765 ( .C1(n15152), .C2(n15151), .A(n15150), .B(n15149), .ZN(
        n15158) );
  AOI22_X1 U16766 ( .A1(n15156), .A2(n15155), .B1(n15154), .B2(n15153), .ZN(
        n15157) );
  NAND2_X1 U16767 ( .A1(n15158), .A2(n15157), .ZN(n15219) );
  AOI21_X1 U16768 ( .B1(n15222), .B2(n15197), .A(n15219), .ZN(n15163) );
  AND2_X1 U16769 ( .A1(n15159), .A2(n15210), .ZN(n15220) );
  AOI22_X1 U16770 ( .A1(n15161), .A2(n15220), .B1(n15178), .B2(n15160), .ZN(
        n15162) );
  OAI221_X1 U16771 ( .B1(n14582), .B2(n15163), .C1(n15198), .C2(n10547), .A(
        n15162), .ZN(P3_U3223) );
  XNOR2_X1 U16772 ( .A(n15166), .B(n15164), .ZN(n15172) );
  OAI21_X1 U16773 ( .B1(n15167), .B2(n15166), .A(n15165), .ZN(n15207) );
  AOI21_X1 U16774 ( .B1(n15207), .B2(n15170), .A(n15169), .ZN(n15171) );
  OAI21_X1 U16775 ( .B1(n15191), .B2(n15172), .A(n15171), .ZN(n15205) );
  INV_X1 U16776 ( .A(n15207), .ZN(n15176) );
  NOR2_X1 U16777 ( .A1(n15173), .A2(n15183), .ZN(n15206) );
  INV_X1 U16778 ( .A(n15206), .ZN(n15174) );
  OAI22_X1 U16779 ( .A1(n15176), .A2(n15175), .B1(n15186), .B2(n15174), .ZN(
        n15177) );
  AOI211_X1 U16780 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15178), .A(n15205), .B(
        n15177), .ZN(n15179) );
  AOI22_X1 U16781 ( .A1(n14582), .A2(n15180), .B1(n15179), .B2(n15198), .ZN(
        P3_U3231) );
  XNOR2_X1 U16782 ( .A(n15182), .B(n15181), .ZN(n15203) );
  NOR2_X1 U16783 ( .A1(n10201), .A2(n15183), .ZN(n15202) );
  INV_X1 U16784 ( .A(n15202), .ZN(n15187) );
  OAI22_X1 U16785 ( .A1(n15187), .A2(n15186), .B1(n15185), .B2(n15184), .ZN(
        n15196) );
  XNOR2_X1 U16786 ( .A(n15189), .B(n15188), .ZN(n15190) );
  OAI222_X1 U16787 ( .A1(n15195), .A2(n15194), .B1(n15193), .B2(n15192), .C1(
        n15191), .C2(n15190), .ZN(n15201) );
  AOI211_X1 U16788 ( .C1(n15197), .C2(n15203), .A(n15196), .B(n15201), .ZN(
        n15199) );
  AOI22_X1 U16789 ( .A1(n14582), .A2(n15200), .B1(n15199), .B2(n15198), .ZN(
        P3_U3232) );
  AOI211_X1 U16790 ( .C1(n15221), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15226) );
  INV_X1 U16791 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15204) );
  AOI22_X1 U16792 ( .A1(n15225), .A2(n15226), .B1(n15204), .B2(n15223), .ZN(
        P3_U3393) );
  AOI211_X1 U16793 ( .C1(n15217), .C2(n15207), .A(n15206), .B(n15205), .ZN(
        n15227) );
  INV_X1 U16794 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15208) );
  AOI22_X1 U16795 ( .A1(n15225), .A2(n15227), .B1(n15208), .B2(n15223), .ZN(
        P3_U3396) );
  AOI22_X1 U16796 ( .A1(n15211), .A2(n15221), .B1(n15210), .B2(n15209), .ZN(
        n15212) );
  AND2_X1 U16797 ( .A1(n15213), .A2(n15212), .ZN(n15228) );
  INV_X1 U16798 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U16799 ( .A1(n15225), .A2(n15228), .B1(n15508), .B2(n15223), .ZN(
        P3_U3411) );
  INV_X1 U16800 ( .A(n15214), .ZN(n15216) );
  AOI211_X1 U16801 ( .C1(n15218), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15232) );
  INV_X1 U16802 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U16803 ( .A1(n15225), .A2(n15232), .B1(n15451), .B2(n15223), .ZN(
        P3_U3414) );
  AOI211_X1 U16804 ( .C1(n15222), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        n15234) );
  INV_X1 U16805 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15224) );
  AOI22_X1 U16806 ( .A1(n15225), .A2(n15234), .B1(n15224), .B2(n15223), .ZN(
        P3_U3420) );
  AOI22_X1 U16807 ( .A1(n15235), .A2(n15226), .B1(n9561), .B2(n15233), .ZN(
        P3_U3460) );
  AOI22_X1 U16808 ( .A1(n15235), .A2(n15227), .B1(n9557), .B2(n15233), .ZN(
        P3_U3461) );
  INV_X1 U16809 ( .A(n15228), .ZN(n15229) );
  OAI22_X1 U16810 ( .A1(n15233), .A2(n15229), .B1(P3_REG1_REG_7__SCAN_IN), 
        .B2(n15235), .ZN(n15230) );
  INV_X1 U16811 ( .A(n15230), .ZN(P3_U3466) );
  AOI22_X1 U16812 ( .A1(n15235), .A2(n15232), .B1(n15231), .B2(n15233), .ZN(
        P3_U3467) );
  AOI22_X1 U16813 ( .A1(n15235), .A2(n15234), .B1(n10558), .B2(n15233), .ZN(
        P3_U3469) );
  NAND2_X1 U16814 ( .A1(n15236), .A2(P3_D_REG_19__SCAN_IN), .ZN(n15541) );
  NAND2_X1 U16815 ( .A1(keyinput97), .A2(keyinput79), .ZN(n15237) );
  NOR3_X1 U16816 ( .A1(keyinput124), .A2(keyinput2), .A3(n15237), .ZN(n15238)
         );
  NAND3_X1 U16817 ( .A1(keyinput104), .A2(keyinput49), .A3(n15238), .ZN(n15251) );
  NOR2_X1 U16818 ( .A1(keyinput76), .A2(keyinput26), .ZN(n15239) );
  NAND3_X1 U16819 ( .A1(keyinput89), .A2(keyinput61), .A3(n15239), .ZN(n15240)
         );
  NOR3_X1 U16820 ( .A1(keyinput29), .A2(keyinput13), .A3(n15240), .ZN(n15249)
         );
  NOR2_X1 U16821 ( .A1(keyinput64), .A2(keyinput125), .ZN(n15241) );
  NAND3_X1 U16822 ( .A1(keyinput62), .A2(keyinput96), .A3(n15241), .ZN(n15247)
         );
  OR4_X1 U16823 ( .A1(keyinput65), .A2(keyinput3), .A3(keyinput50), .A4(
        keyinput116), .ZN(n15246) );
  INV_X1 U16824 ( .A(keyinput55), .ZN(n15242) );
  NAND4_X1 U16825 ( .A1(keyinput100), .A2(keyinput63), .A3(keyinput71), .A4(
        n15242), .ZN(n15245) );
  NOR2_X1 U16826 ( .A1(keyinput66), .A2(keyinput110), .ZN(n15243) );
  NAND3_X1 U16827 ( .A1(keyinput75), .A2(keyinput9), .A3(n15243), .ZN(n15244)
         );
  NOR4_X1 U16828 ( .A1(n15247), .A2(n15246), .A3(n15245), .A4(n15244), .ZN(
        n15248) );
  NAND4_X1 U16829 ( .A1(keyinput67), .A2(keyinput85), .A3(n15249), .A4(n15248), 
        .ZN(n15250) );
  NOR4_X1 U16830 ( .A1(keyinput102), .A2(keyinput44), .A3(n15251), .A4(n15250), 
        .ZN(n15301) );
  NOR2_X1 U16831 ( .A1(keyinput68), .A2(keyinput58), .ZN(n15252) );
  NAND3_X1 U16832 ( .A1(keyinput113), .A2(keyinput70), .A3(n15252), .ZN(n15299) );
  NAND4_X1 U16833 ( .A1(keyinput11), .A2(keyinput87), .A3(keyinput92), .A4(
        keyinput99), .ZN(n15298) );
  NOR2_X1 U16834 ( .A1(keyinput6), .A2(keyinput42), .ZN(n15253) );
  NAND3_X1 U16835 ( .A1(keyinput54), .A2(keyinput82), .A3(n15253), .ZN(n15254)
         );
  NOR3_X1 U16836 ( .A1(keyinput90), .A2(keyinput7), .A3(n15254), .ZN(n15264)
         );
  INV_X1 U16837 ( .A(keyinput17), .ZN(n15255) );
  NAND4_X1 U16838 ( .A1(keyinput16), .A2(keyinput98), .A3(keyinput8), .A4(
        n15255), .ZN(n15262) );
  NOR2_X1 U16839 ( .A1(keyinput28), .A2(keyinput80), .ZN(n15256) );
  NAND3_X1 U16840 ( .A1(keyinput1), .A2(keyinput41), .A3(n15256), .ZN(n15261)
         );
  NOR2_X1 U16841 ( .A1(keyinput83), .A2(keyinput45), .ZN(n15257) );
  NAND3_X1 U16842 ( .A1(keyinput22), .A2(keyinput73), .A3(n15257), .ZN(n15260)
         );
  NOR2_X1 U16843 ( .A1(keyinput10), .A2(keyinput23), .ZN(n15258) );
  NAND3_X1 U16844 ( .A1(keyinput111), .A2(keyinput4), .A3(n15258), .ZN(n15259)
         );
  NOR4_X1 U16845 ( .A1(n15262), .A2(n15261), .A3(n15260), .A4(n15259), .ZN(
        n15263) );
  NAND4_X1 U16846 ( .A1(keyinput43), .A2(keyinput53), .A3(n15264), .A4(n15263), 
        .ZN(n15297) );
  NAND2_X1 U16847 ( .A1(keyinput95), .A2(keyinput57), .ZN(n15265) );
  NOR3_X1 U16848 ( .A1(keyinput81), .A2(keyinput0), .A3(n15265), .ZN(n15295)
         );
  NOR4_X1 U16849 ( .A1(keyinput27), .A2(keyinput74), .A3(keyinput101), .A4(
        keyinput115), .ZN(n15294) );
  NAND2_X1 U16850 ( .A1(keyinput14), .A2(keyinput126), .ZN(n15266) );
  NOR3_X1 U16851 ( .A1(keyinput25), .A2(keyinput36), .A3(n15266), .ZN(n15267)
         );
  NAND3_X1 U16852 ( .A1(keyinput109), .A2(keyinput47), .A3(n15267), .ZN(n15275) );
  INV_X1 U16853 ( .A(keyinput34), .ZN(n15268) );
  NAND4_X1 U16854 ( .A1(keyinput31), .A2(keyinput37), .A3(keyinput105), .A4(
        n15268), .ZN(n15269) );
  NOR4_X1 U16855 ( .A1(keyinput120), .A2(keyinput84), .A3(keyinput78), .A4(
        n15269), .ZN(n15273) );
  NOR2_X1 U16856 ( .A1(keyinput123), .A2(keyinput69), .ZN(n15270) );
  NAND3_X1 U16857 ( .A1(keyinput112), .A2(keyinput20), .A3(n15270), .ZN(n15271) );
  NOR3_X1 U16858 ( .A1(keyinput77), .A2(keyinput117), .A3(n15271), .ZN(n15272)
         );
  NAND4_X1 U16859 ( .A1(n15273), .A2(keyinput15), .A3(keyinput91), .A4(n15272), 
        .ZN(n15274) );
  NOR4_X1 U16860 ( .A1(keyinput32), .A2(keyinput5), .A3(n15275), .A4(n15274), 
        .ZN(n15293) );
  INV_X1 U16861 ( .A(keyinput121), .ZN(n15276) );
  NOR4_X1 U16862 ( .A1(keyinput118), .A2(keyinput48), .A3(keyinput122), .A4(
        n15276), .ZN(n15277) );
  NAND3_X1 U16863 ( .A1(keyinput114), .A2(keyinput39), .A3(n15277), .ZN(n15291) );
  INV_X1 U16864 ( .A(keyinput21), .ZN(n15278) );
  NOR4_X1 U16865 ( .A1(keyinput40), .A2(keyinput106), .A3(keyinput88), .A4(
        n15278), .ZN(n15289) );
  NAND2_X1 U16866 ( .A1(keyinput59), .A2(keyinput51), .ZN(n15279) );
  NOR3_X1 U16867 ( .A1(keyinput72), .A2(keyinput19), .A3(n15279), .ZN(n15288)
         );
  NOR2_X1 U16868 ( .A1(keyinput108), .A2(keyinput119), .ZN(n15280) );
  NAND3_X1 U16869 ( .A1(keyinput38), .A2(keyinput103), .A3(n15280), .ZN(n15286) );
  INV_X1 U16870 ( .A(keyinput33), .ZN(n15281) );
  NAND4_X1 U16871 ( .A1(keyinput30), .A2(keyinput24), .A3(keyinput52), .A4(
        n15281), .ZN(n15285) );
  NOR2_X1 U16872 ( .A1(keyinput93), .A2(keyinput56), .ZN(n15282) );
  NAND3_X1 U16873 ( .A1(keyinput60), .A2(keyinput46), .A3(n15282), .ZN(n15284)
         );
  NAND4_X1 U16874 ( .A1(keyinput107), .A2(keyinput86), .A3(keyinput18), .A4(
        keyinput12), .ZN(n15283) );
  NOR4_X1 U16875 ( .A1(n15286), .A2(n15285), .A3(n15284), .A4(n15283), .ZN(
        n15287) );
  NAND3_X1 U16876 ( .A1(n15289), .A2(n15288), .A3(n15287), .ZN(n15290) );
  NOR4_X1 U16877 ( .A1(keyinput35), .A2(keyinput94), .A3(n15291), .A4(n15290), 
        .ZN(n15292) );
  NAND4_X1 U16878 ( .A1(n15295), .A2(n15294), .A3(n15293), .A4(n15292), .ZN(
        n15296) );
  NOR4_X1 U16879 ( .A1(n15299), .A2(n15298), .A3(n15297), .A4(n15296), .ZN(
        n15300) );
  AOI21_X1 U16880 ( .B1(n15301), .B2(n15300), .A(keyinput127), .ZN(n15539) );
  INV_X1 U16881 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U16882 ( .A1(n15304), .A2(keyinput3), .B1(n15303), .B2(keyinput64), 
        .ZN(n15302) );
  OAI221_X1 U16883 ( .B1(n15304), .B2(keyinput3), .C1(n15303), .C2(keyinput64), 
        .A(n15302), .ZN(n15311) );
  XNOR2_X1 U16884 ( .A(n15305), .B(keyinput50), .ZN(n15310) );
  XNOR2_X1 U16885 ( .A(n15306), .B(keyinput62), .ZN(n15309) );
  XNOR2_X1 U16886 ( .A(n15307), .B(keyinput96), .ZN(n15308) );
  OR4_X1 U16887 ( .A1(n15311), .A2(n15310), .A3(n15309), .A4(n15308), .ZN(
        n15318) );
  AOI22_X1 U16888 ( .A1(n15314), .A2(keyinput116), .B1(keyinput67), .B2(n15313), .ZN(n15312) );
  OAI221_X1 U16889 ( .B1(n15314), .B2(keyinput116), .C1(n15313), .C2(
        keyinput67), .A(n15312), .ZN(n15317) );
  XNOR2_X1 U16890 ( .A(n15315), .B(keyinput125), .ZN(n15316) );
  NOR3_X1 U16891 ( .A1(n15318), .A2(n15317), .A3(n15316), .ZN(n15363) );
  AOI22_X1 U16892 ( .A1(n15320), .A2(keyinput26), .B1(n6905), .B2(keyinput76), 
        .ZN(n15319) );
  OAI221_X1 U16893 ( .B1(n15320), .B2(keyinput26), .C1(n6905), .C2(keyinput76), 
        .A(n15319), .ZN(n15330) );
  AOI22_X1 U16894 ( .A1(n15323), .A2(keyinput61), .B1(keyinput29), .B2(n15322), 
        .ZN(n15321) );
  OAI221_X1 U16895 ( .B1(n15323), .B2(keyinput61), .C1(n15322), .C2(keyinput29), .A(n15321), .ZN(n15329) );
  XNOR2_X1 U16896 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput89), .ZN(n15327) );
  XNOR2_X1 U16897 ( .A(P3_REG1_REG_30__SCAN_IN), .B(keyinput85), .ZN(n15326)
         );
  XNOR2_X1 U16898 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput124), .ZN(n15325) );
  XNOR2_X1 U16899 ( .A(SI_3_), .B(keyinput13), .ZN(n15324) );
  NAND4_X1 U16900 ( .A1(n15327), .A2(n15326), .A3(n15325), .A4(n15324), .ZN(
        n15328) );
  NOR3_X1 U16901 ( .A1(n15330), .A2(n15329), .A3(n15328), .ZN(n15362) );
  AOI22_X1 U16902 ( .A1(n15333), .A2(keyinput2), .B1(keyinput66), .B2(n15332), 
        .ZN(n15331) );
  OAI221_X1 U16903 ( .B1(n15333), .B2(keyinput2), .C1(n15332), .C2(keyinput66), 
        .A(n15331), .ZN(n15345) );
  INV_X1 U16904 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15336) );
  AOI22_X1 U16905 ( .A1(n15336), .A2(keyinput49), .B1(keyinput102), .B2(n15335), .ZN(n15334) );
  OAI221_X1 U16906 ( .B1(n15336), .B2(keyinput49), .C1(n15335), .C2(
        keyinput102), .A(n15334), .ZN(n15344) );
  AOI22_X1 U16907 ( .A1(n15339), .A2(keyinput79), .B1(n15338), .B2(keyinput104), .ZN(n15337) );
  OAI221_X1 U16908 ( .B1(n15339), .B2(keyinput79), .C1(n15338), .C2(
        keyinput104), .A(n15337), .ZN(n15343) );
  XNOR2_X1 U16909 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput97), .ZN(n15341)
         );
  XNOR2_X1 U16910 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput44), .ZN(n15340) );
  NAND2_X1 U16911 ( .A1(n15341), .A2(n15340), .ZN(n15342) );
  NOR4_X1 U16912 ( .A1(n15345), .A2(n15344), .A3(n15343), .A4(n15342), .ZN(
        n15361) );
  AOI22_X1 U16913 ( .A1(n11344), .A2(keyinput75), .B1(n15347), .B2(keyinput110), .ZN(n15346) );
  OAI221_X1 U16914 ( .B1(n11344), .B2(keyinput75), .C1(n15347), .C2(
        keyinput110), .A(n15346), .ZN(n15359) );
  AOI22_X1 U16915 ( .A1(n15350), .A2(keyinput9), .B1(n15349), .B2(keyinput63), 
        .ZN(n15348) );
  OAI221_X1 U16916 ( .B1(n15350), .B2(keyinput9), .C1(n15349), .C2(keyinput63), 
        .A(n15348), .ZN(n15358) );
  INV_X1 U16917 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U16918 ( .A1(n15353), .A2(keyinput100), .B1(n15352), .B2(keyinput55), .ZN(n15351) );
  OAI221_X1 U16919 ( .B1(n15353), .B2(keyinput100), .C1(n15352), .C2(
        keyinput55), .A(n15351), .ZN(n15357) );
  AOI22_X1 U16920 ( .A1(n8234), .A2(keyinput71), .B1(keyinput24), .B2(n15355), 
        .ZN(n15354) );
  OAI221_X1 U16921 ( .B1(n8234), .B2(keyinput71), .C1(n15355), .C2(keyinput24), 
        .A(n15354), .ZN(n15356) );
  NOR4_X1 U16922 ( .A1(n15359), .A2(n15358), .A3(n15357), .A4(n15356), .ZN(
        n15360) );
  NAND4_X1 U16923 ( .A1(n15363), .A2(n15362), .A3(n15361), .A4(n15360), .ZN(
        n15537) );
  AOI22_X1 U16924 ( .A1(n15365), .A2(keyinput33), .B1(n9079), .B2(keyinput38), 
        .ZN(n15364) );
  OAI221_X1 U16925 ( .B1(n15365), .B2(keyinput33), .C1(n9079), .C2(keyinput38), 
        .A(n15364), .ZN(n15375) );
  INV_X1 U16926 ( .A(SI_26_), .ZN(n15368) );
  AOI22_X1 U16927 ( .A1(n15368), .A2(keyinput119), .B1(keyinput108), .B2(
        n15367), .ZN(n15366) );
  OAI221_X1 U16928 ( .B1(n15368), .B2(keyinput119), .C1(n15367), .C2(
        keyinput108), .A(n15366), .ZN(n15374) );
  XNOR2_X1 U16929 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput52), .ZN(n15372) );
  XNOR2_X1 U16930 ( .A(P3_IR_REG_4__SCAN_IN), .B(keyinput30), .ZN(n15371) );
  XNOR2_X1 U16931 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput35), .ZN(n15370) );
  XNOR2_X1 U16932 ( .A(P1_REG1_REG_31__SCAN_IN), .B(keyinput103), .ZN(n15369)
         );
  NAND4_X1 U16933 ( .A1(n15372), .A2(n15371), .A3(n15370), .A4(n15369), .ZN(
        n15373) );
  NOR3_X1 U16934 ( .A1(n15375), .A2(n15374), .A3(n15373), .ZN(n15416) );
  AOI22_X1 U16935 ( .A1(n15377), .A2(keyinput48), .B1(keyinput114), .B2(n9239), 
        .ZN(n15376) );
  OAI221_X1 U16936 ( .B1(n15377), .B2(keyinput48), .C1(n9239), .C2(keyinput114), .A(n15376), .ZN(n15387) );
  AOI22_X1 U16937 ( .A1(n10014), .A2(keyinput121), .B1(n15379), .B2(
        keyinput107), .ZN(n15378) );
  OAI221_X1 U16938 ( .B1(n10014), .B2(keyinput121), .C1(n15379), .C2(
        keyinput107), .A(n15378), .ZN(n15386) );
  XNOR2_X1 U16939 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput118), .ZN(n15382) );
  XNOR2_X1 U16940 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput39), .ZN(n15381) );
  XNOR2_X1 U16941 ( .A(keyinput122), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n15380)
         );
  NAND3_X1 U16942 ( .A1(n15382), .A2(n15381), .A3(n15380), .ZN(n15385) );
  XNOR2_X1 U16943 ( .A(n15383), .B(keyinput94), .ZN(n15384) );
  NOR4_X1 U16944 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15415) );
  AOI22_X1 U16945 ( .A1(n7630), .A2(keyinput56), .B1(keyinput18), .B2(n15389), 
        .ZN(n15388) );
  OAI221_X1 U16946 ( .B1(n7630), .B2(keyinput56), .C1(n15389), .C2(keyinput18), 
        .A(n15388), .ZN(n15398) );
  XNOR2_X1 U16947 ( .A(keyinput86), .B(n15390), .ZN(n15397) );
  XNOR2_X1 U16948 ( .A(keyinput46), .B(n11457), .ZN(n15396) );
  XNOR2_X1 U16949 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput93), .ZN(n15394) );
  XNOR2_X1 U16950 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput60), .ZN(n15393) );
  XNOR2_X1 U16951 ( .A(P3_REG0_REG_25__SCAN_IN), .B(keyinput51), .ZN(n15392)
         );
  XNOR2_X1 U16952 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput12), .ZN(n15391) );
  NAND4_X1 U16953 ( .A1(n15394), .A2(n15393), .A3(n15392), .A4(n15391), .ZN(
        n15395) );
  NOR4_X1 U16954 ( .A1(n15398), .A2(n15397), .A3(n15396), .A4(n15395), .ZN(
        n15414) );
  AOI22_X1 U16955 ( .A1(n15400), .A2(keyinput59), .B1(keyinput40), .B2(n8501), 
        .ZN(n15399) );
  OAI221_X1 U16956 ( .B1(n15400), .B2(keyinput59), .C1(n8501), .C2(keyinput40), 
        .A(n15399), .ZN(n15412) );
  INV_X1 U16957 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U16958 ( .A1(n15403), .A2(keyinput19), .B1(keyinput72), .B2(n15402), 
        .ZN(n15401) );
  OAI221_X1 U16959 ( .B1(n15403), .B2(keyinput19), .C1(n15402), .C2(keyinput72), .A(n15401), .ZN(n15411) );
  AOI22_X1 U16960 ( .A1(n15406), .A2(keyinput106), .B1(keyinput21), .B2(n15405), .ZN(n15404) );
  OAI221_X1 U16961 ( .B1(n15406), .B2(keyinput106), .C1(n15405), .C2(
        keyinput21), .A(n15404), .ZN(n15410) );
  XNOR2_X1 U16962 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput88), .ZN(n15408) );
  XNOR2_X1 U16963 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput120), .ZN(n15407)
         );
  NAND2_X1 U16964 ( .A1(n15408), .A2(n15407), .ZN(n15409) );
  NOR4_X1 U16965 ( .A1(n15412), .A2(n15411), .A3(n15410), .A4(n15409), .ZN(
        n15413) );
  NAND4_X1 U16966 ( .A1(n15416), .A2(n15415), .A3(n15414), .A4(n15413), .ZN(
        n15536) );
  INV_X1 U16967 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U16968 ( .A1(n15419), .A2(keyinput70), .B1(keyinput92), .B2(n15418), 
        .ZN(n15417) );
  OAI221_X1 U16969 ( .B1(n15419), .B2(keyinput70), .C1(n15418), .C2(keyinput92), .A(n15417), .ZN(n15429) );
  AOI22_X1 U16970 ( .A1(n15421), .A2(keyinput113), .B1(keyinput58), .B2(n9807), 
        .ZN(n15420) );
  OAI221_X1 U16971 ( .B1(n15421), .B2(keyinput113), .C1(n9807), .C2(keyinput58), .A(n15420), .ZN(n15428) );
  AOI22_X1 U16972 ( .A1(n14269), .A2(keyinput99), .B1(n15423), .B2(keyinput1), 
        .ZN(n15422) );
  OAI221_X1 U16973 ( .B1(n14269), .B2(keyinput99), .C1(n15423), .C2(keyinput1), 
        .A(n15422), .ZN(n15427) );
  XNOR2_X1 U16974 ( .A(P3_D_REG_1__SCAN_IN), .B(keyinput68), .ZN(n15425) );
  NAND2_X1 U16975 ( .A1(n15425), .A2(n15424), .ZN(n15426) );
  NOR4_X1 U16976 ( .A1(n15429), .A2(n15428), .A3(n15427), .A4(n15426), .ZN(
        n15475) );
  AOI22_X1 U16977 ( .A1(n11315), .A2(keyinput53), .B1(n15431), .B2(keyinput6), 
        .ZN(n15430) );
  OAI221_X1 U16978 ( .B1(n11315), .B2(keyinput53), .C1(n15431), .C2(keyinput6), 
        .A(n15430), .ZN(n15443) );
  AOI22_X1 U16979 ( .A1(n15434), .A2(keyinput82), .B1(n15433), .B2(keyinput11), 
        .ZN(n15432) );
  OAI221_X1 U16980 ( .B1(n15434), .B2(keyinput82), .C1(n15433), .C2(keyinput11), .A(n15432), .ZN(n15442) );
  AOI22_X1 U16981 ( .A1(n15437), .A2(keyinput42), .B1(keyinput90), .B2(n15436), 
        .ZN(n15435) );
  OAI221_X1 U16982 ( .B1(n15437), .B2(keyinput42), .C1(n15436), .C2(keyinput90), .A(n15435), .ZN(n15441) );
  XOR2_X1 U16983 ( .A(n9731), .B(keyinput43), .Z(n15439) );
  XNOR2_X1 U16984 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput7), .ZN(n15438) );
  NAND2_X1 U16985 ( .A1(n15439), .A2(n15438), .ZN(n15440) );
  NOR4_X1 U16986 ( .A1(n15443), .A2(n15442), .A3(n15441), .A4(n15440), .ZN(
        n15474) );
  AOI22_X1 U16987 ( .A1(n15446), .A2(keyinput23), .B1(n15445), .B2(keyinput22), 
        .ZN(n15444) );
  OAI221_X1 U16988 ( .B1(n15446), .B2(keyinput23), .C1(n15445), .C2(keyinput22), .A(n15444), .ZN(n15457) );
  AOI22_X1 U16989 ( .A1(n15449), .A2(keyinput111), .B1(keyinput4), .B2(n15448), 
        .ZN(n15447) );
  OAI221_X1 U16990 ( .B1(n15449), .B2(keyinput111), .C1(n15448), .C2(keyinput4), .A(n15447), .ZN(n15456) );
  AOI22_X1 U16991 ( .A1(n8814), .A2(keyinput73), .B1(n15451), .B2(keyinput65), 
        .ZN(n15450) );
  OAI221_X1 U16992 ( .B1(n8814), .B2(keyinput73), .C1(n15451), .C2(keyinput65), 
        .A(n15450), .ZN(n15455) );
  AOI22_X1 U16993 ( .A1(n8641), .A2(keyinput45), .B1(keyinput83), .B2(n15453), 
        .ZN(n15452) );
  OAI221_X1 U16994 ( .B1(n8641), .B2(keyinput45), .C1(n15453), .C2(keyinput83), 
        .A(n15452), .ZN(n15454) );
  NOR4_X1 U16995 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15473) );
  AOI22_X1 U16996 ( .A1(n15460), .A2(keyinput80), .B1(keyinput28), .B2(n15459), 
        .ZN(n15458) );
  OAI221_X1 U16997 ( .B1(n15460), .B2(keyinput80), .C1(n15459), .C2(keyinput28), .A(n15458), .ZN(n15471) );
  AOI22_X1 U16998 ( .A1(n15462), .A2(keyinput8), .B1(keyinput10), .B2(n9248), 
        .ZN(n15461) );
  OAI221_X1 U16999 ( .B1(n15462), .B2(keyinput8), .C1(n9248), .C2(keyinput10), 
        .A(n15461), .ZN(n15470) );
  AOI22_X1 U17000 ( .A1(n15465), .A2(keyinput16), .B1(n15464), .B2(keyinput98), 
        .ZN(n15463) );
  OAI221_X1 U17001 ( .B1(n15465), .B2(keyinput16), .C1(n15464), .C2(keyinput98), .A(n15463), .ZN(n15469) );
  XNOR2_X1 U17002 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput41), .ZN(n15467)
         );
  XNOR2_X1 U17003 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput17), .ZN(n15466) );
  NAND2_X1 U17004 ( .A1(n15467), .A2(n15466), .ZN(n15468) );
  NOR4_X1 U17005 ( .A1(n15471), .A2(n15470), .A3(n15469), .A4(n15468), .ZN(
        n15472) );
  NAND4_X1 U17006 ( .A1(n15475), .A2(n15474), .A3(n15473), .A4(n15472), .ZN(
        n15535) );
  AOI22_X1 U17007 ( .A1(n15477), .A2(keyinput74), .B1(n10125), .B2(keyinput101), .ZN(n15476) );
  OAI221_X1 U17008 ( .B1(n15477), .B2(keyinput74), .C1(n10125), .C2(
        keyinput101), .A(n15476), .ZN(n15488) );
  AOI22_X1 U17009 ( .A1(n15480), .A2(keyinput115), .B1(keyinput57), .B2(n15479), .ZN(n15478) );
  OAI221_X1 U17010 ( .B1(n15480), .B2(keyinput115), .C1(n15479), .C2(
        keyinput57), .A(n15478), .ZN(n15487) );
  XOR2_X1 U17011 ( .A(n15481), .B(keyinput0), .Z(n15485) );
  XNOR2_X1 U17012 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput25), .ZN(n15484) );
  XNOR2_X1 U17013 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput81), .ZN(n15483) );
  XNOR2_X1 U17014 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput95), .ZN(n15482)
         );
  NAND4_X1 U17015 ( .A1(n15485), .A2(n15484), .A3(n15483), .A4(n15482), .ZN(
        n15486) );
  NOR3_X1 U17016 ( .A1(n15488), .A2(n15487), .A3(n15486), .ZN(n15533) );
  AOI22_X1 U17017 ( .A1(n9972), .A2(keyinput34), .B1(keyinput84), .B2(n15490), 
        .ZN(n15489) );
  OAI221_X1 U17018 ( .B1(n9972), .B2(keyinput34), .C1(n15490), .C2(keyinput84), 
        .A(n15489), .ZN(n15500) );
  AOI22_X1 U17019 ( .A1(n15492), .A2(keyinput78), .B1(keyinput27), .B2(n12516), 
        .ZN(n15491) );
  OAI221_X1 U17020 ( .B1(n15492), .B2(keyinput78), .C1(n12516), .C2(keyinput27), .A(n15491), .ZN(n15499) );
  AOI22_X1 U17021 ( .A1(n15495), .A2(keyinput37), .B1(keyinput31), .B2(n15494), 
        .ZN(n15493) );
  OAI221_X1 U17022 ( .B1(n15495), .B2(keyinput37), .C1(n15494), .C2(keyinput31), .A(n15493), .ZN(n15498) );
  XNOR2_X1 U17023 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput105), .ZN(n15496) );
  OAI21_X1 U17024 ( .B1(keyinput127), .B2(n12124), .A(n15496), .ZN(n15497) );
  NOR4_X1 U17025 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15532) );
  INV_X1 U17026 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U17027 ( .A1(n15502), .A2(keyinput117), .B1(keyinput54), .B2(n14215), .ZN(n15501) );
  OAI221_X1 U17028 ( .B1(n15502), .B2(keyinput117), .C1(n14215), .C2(
        keyinput54), .A(n15501), .ZN(n15514) );
  AOI22_X1 U17029 ( .A1(n15505), .A2(keyinput112), .B1(keyinput69), .B2(n15504), .ZN(n15503) );
  OAI221_X1 U17030 ( .B1(n15505), .B2(keyinput112), .C1(n15504), .C2(
        keyinput69), .A(n15503), .ZN(n15513) );
  AOI22_X1 U17031 ( .A1(n15508), .A2(keyinput20), .B1(n15507), .B2(keyinput15), 
        .ZN(n15506) );
  OAI221_X1 U17032 ( .B1(n15508), .B2(keyinput20), .C1(n15507), .C2(keyinput15), .A(n15506), .ZN(n15512) );
  XNOR2_X1 U17033 ( .A(P2_REG1_REG_26__SCAN_IN), .B(keyinput91), .ZN(n15510)
         );
  XNOR2_X1 U17034 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput77), .ZN(n15509) );
  NAND2_X1 U17035 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  NOR4_X1 U17036 ( .A1(n15514), .A2(n15513), .A3(n15512), .A4(n15511), .ZN(
        n15531) );
  AOI22_X1 U17037 ( .A1(n7160), .A2(keyinput5), .B1(keyinput36), .B2(n15516), 
        .ZN(n15515) );
  OAI221_X1 U17038 ( .B1(n7160), .B2(keyinput5), .C1(n15516), .C2(keyinput36), 
        .A(n15515), .ZN(n15529) );
  AOI22_X1 U17039 ( .A1(n15519), .A2(keyinput126), .B1(keyinput32), .B2(n15518), .ZN(n15517) );
  OAI221_X1 U17040 ( .B1(n15519), .B2(keyinput126), .C1(n15518), .C2(
        keyinput32), .A(n15517), .ZN(n15528) );
  AOI22_X1 U17041 ( .A1(n15522), .A2(keyinput47), .B1(n15521), .B2(keyinput123), .ZN(n15520) );
  OAI221_X1 U17042 ( .B1(n15522), .B2(keyinput47), .C1(n15521), .C2(
        keyinput123), .A(n15520), .ZN(n15527) );
  AOI22_X1 U17043 ( .A1(n15525), .A2(keyinput14), .B1(n15524), .B2(keyinput109), .ZN(n15523) );
  OAI221_X1 U17044 ( .B1(n15525), .B2(keyinput14), .C1(n15524), .C2(
        keyinput109), .A(n15523), .ZN(n15526) );
  NOR4_X1 U17045 ( .A1(n15529), .A2(n15528), .A3(n15527), .A4(n15526), .ZN(
        n15530) );
  NAND4_X1 U17046 ( .A1(n15533), .A2(n15532), .A3(n15531), .A4(n15530), .ZN(
        n15534) );
  NOR4_X1 U17047 ( .A1(n15537), .A2(n15536), .A3(n15535), .A4(n15534), .ZN(
        n15538) );
  OAI21_X1 U17048 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(n15539), .A(n15538), 
        .ZN(n15540) );
  XOR2_X1 U17049 ( .A(n15541), .B(n15540), .Z(P3_U3246) );
  XOR2_X1 U17050 ( .A(n15543), .B(n15542), .Z(SUB_1596_U59) );
  XNOR2_X1 U17051 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15544), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17052 ( .B1(n15545), .B2(n9049), .A(n15554), .ZN(SUB_1596_U53) );
  XOR2_X1 U17053 ( .A(n15547), .B(n15546), .Z(SUB_1596_U56) );
  OAI21_X1 U17054 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15552) );
  XOR2_X1 U17055 ( .A(n15552), .B(n15551), .Z(SUB_1596_U60) );
  XOR2_X1 U17056 ( .A(n15554), .B(n15553), .Z(SUB_1596_U5) );
  OR2_X1 U7400 ( .A1(n8397), .A2(n13800), .ZN(n8398) );
  NAND2_X1 U7420 ( .A1(n13801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8396) );
  BUF_X2 U7321 ( .A(n10100), .Z(n11757) );
  INV_X2 U7327 ( .A(n9552), .ZN(n8005) );
  CLKBUF_X1 U7334 ( .A(n12322), .Z(n6568) );
  CLKBUF_X1 U7358 ( .A(n8724), .Z(n6586) );
  INV_X1 U7378 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13800) );
  CLKBUF_X1 U7379 ( .A(n13935), .Z(n6777) );
  CLKBUF_X1 U7390 ( .A(n12640), .Z(n6813) );
  CLKBUF_X1 U7391 ( .A(n9358), .Z(n14837) );
  CLKBUF_X1 U7414 ( .A(n12882), .Z(n6589) );
  AOI211_X1 U7438 ( .C1(n13726), .C2(n13694), .A(n13589), .B(n13588), .ZN(
        n13590) );
  CLKBUF_X1 U8127 ( .A(n11642), .Z(n12322) );
endmodule

