

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068;

  INV_X1 U3547 ( .A(n6309), .ZN(n6326) );
  CLKBUF_X2 U3548 ( .A(n5363), .Z(n3104) );
  INV_X1 U3549 ( .A(n6305), .ZN(n6334) );
  NAND2_X1 U3550 ( .A1(n6463), .A2(n6069), .ZN(n5903) );
  BUF_X1 U3551 ( .A(n3431), .Z(n3977) );
  INV_X1 U3553 ( .A(n4391), .ZN(n5280) );
  CLKBUF_X1 U3554 ( .A(n3493), .Z(n4680) );
  CLKBUF_X2 U3555 ( .A(n3483), .Z(n3971) );
  BUF_X1 U3556 ( .A(n3497), .Z(n4688) );
  INV_X2 U3557 ( .A(n4703), .ZN(n3519) );
  AND2_X1 U3558 ( .A1(n4538), .A2(n4717), .ZN(n3483) );
  AND2_X1 U3559 ( .A1(n3218), .A2(n4537), .ZN(n3543) );
  BUF_X1 U3560 ( .A(n3541), .Z(n3530) );
  CLKBUF_X2 U3561 ( .A(n3462), .Z(n3991) );
  AND2_X1 U3563 ( .A1(n3271), .A2(n4537), .ZN(n3531) );
  AND3_X1 U3564 ( .A1(n4579), .A2(STATE2_REG_0__SCAN_IN), .A3(n3554), .ZN(
        n4078) );
  NAND2_X1 U3565 ( .A1(n3628), .A2(n3627), .ZN(n4123) );
  AOI21_X1 U3566 ( .B1(n4522), .B2(n5282), .A(n3592), .ZN(n3687) );
  INV_X1 U3567 ( .A(n4064), .ZN(n4353) );
  NAND2_X1 U3568 ( .A1(n5439), .A2(n6752), .ZN(n5272) );
  CLKBUF_X2 U3569 ( .A(n4327), .Z(n3099) );
  NAND2_X1 U3572 ( .A1(n3497), .A2(n3453), .ZN(n4239) );
  INV_X2 U3573 ( .A(n3224), .ZN(n5865) );
  INV_X1 U3574 ( .A(n6319), .ZN(n6294) );
  NAND2_X1 U3575 ( .A1(n4175), .A2(n4174), .ZN(n6100) );
  AND2_X2 U3576 ( .A1(n5346), .A2(n5348), .ZN(n5336) );
  AND2_X1 U3577 ( .A1(n4260), .A2(n6401), .ZN(n4649) );
  NAND2_X1 U3578 ( .A1(n4497), .A2(n4496), .ZN(n6756) );
  AOI211_X1 U3579 ( .C1(n5924), .C2(n6305), .A(n5309), .B(n5308), .ZN(n5310)
         );
  OR2_X1 U3580 ( .A1(n4595), .A2(n4869), .ZN(n6226) );
  NOR2_X4 U3582 ( .A1(n5361), .A2(n5362), .ZN(n5346) );
  OAI22_X2 U3583 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5744), .B1(n5753), .B2(n5736), .ZN(n5737) );
  XNOR2_X2 U3584 ( .A(n3595), .B(n3593), .ZN(n3686) );
  NAND2_X1 U3585 ( .A1(n4304), .A2(n4307), .ZN(n4327) );
  OR2_X1 U3586 ( .A1(n6031), .A2(n6028), .ZN(n6021) );
  NAND2_X1 U3587 ( .A1(n3719), .A2(n3674), .ZN(n4304) );
  OAI211_X1 U3588 ( .C1(n3144), .C2(n3553), .A(n3143), .B(n4306), .ZN(n3595)
         );
  NAND2_X1 U3589 ( .A1(n4502), .A2(n3502), .ZN(n4736) );
  BUF_X2 U3590 ( .A(n3372), .Z(n3905) );
  CLKBUF_X2 U3591 ( .A(n3476), .Z(n3818) );
  AOI21_X1 U3592 ( .B1(n5326), .B2(n5325), .A(n4336), .ZN(n5705) );
  XNOR2_X1 U3593 ( .A(n4355), .B(n4354), .ZN(n5291) );
  OAI21_X1 U3594 ( .B1(n4336), .B2(n4337), .A(n4069), .ZN(n5312) );
  AOI21_X1 U3595 ( .B1(n4070), .B2(n4069), .A(n4355), .ZN(n5694) );
  NAND2_X1 U3596 ( .A1(n3183), .A2(n3107), .ZN(n3197) );
  XNOR2_X1 U3597 ( .A(n5299), .B(n5298), .ZN(n5924) );
  NAND2_X2 U3598 ( .A1(n3852), .A2(n3172), .ZN(n5485) );
  AND2_X1 U3599 ( .A1(n4227), .A2(n5293), .ZN(n4228) );
  OR2_X1 U3600 ( .A1(n3838), .A2(n3837), .ZN(n3852) );
  AND3_X1 U3601 ( .A1(n3742), .A2(n4612), .A3(n4755), .ZN(n3169) );
  INV_X2 U3602 ( .A(n5070), .ZN(n5680) );
  XNOR2_X1 U3603 ( .A(n4304), .B(n3745), .ZN(n4298) );
  OR2_X1 U3604 ( .A1(n4893), .A2(n3904), .ZN(n3741) );
  AND3_X1 U3605 ( .A1(n3729), .A2(n3198), .A3(n3170), .ZN(n3719) );
  XNOR2_X1 U3606 ( .A(n3731), .B(n3712), .ZN(n4276) );
  NAND2_X1 U3607 ( .A1(n3729), .A2(n4770), .ZN(n3731) );
  AND2_X1 U3608 ( .A1(n4608), .A2(n4609), .ZN(n3709) );
  AND2_X1 U3609 ( .A1(n4770), .A2(n3651), .ZN(n3198) );
  NAND2_X1 U3610 ( .A1(n3213), .A2(n3212), .ZN(n5514) );
  XNOR2_X1 U3611 ( .A(n3684), .B(n4622), .ZN(n4661) );
  INV_X1 U3612 ( .A(n6100), .ZN(n3213) );
  CLKBUF_X1 U3613 ( .A(n4664), .Z(n6141) );
  NAND2_X1 U3614 ( .A1(n3683), .A2(n4622), .ZN(n3730) );
  NAND2_X1 U3615 ( .A1(n3618), .A2(n3617), .ZN(n4622) );
  NAND2_X1 U3616 ( .A1(n3697), .A2(n3696), .ZN(n5163) );
  NAND2_X1 U3617 ( .A1(n3621), .A2(n3620), .ZN(n4516) );
  INV_X1 U3618 ( .A(n5625), .ZN(n4175) );
  CLKBUF_X1 U3619 ( .A(n4522), .Z(n5582) );
  NAND2_X1 U3620 ( .A1(n3123), .A2(n3234), .ZN(n3236) );
  OR2_X1 U3621 ( .A1(n3603), .A2(n3263), .ZN(n3234) );
  NOR2_X1 U3622 ( .A1(n3214), .A2(n5512), .ZN(n3212) );
  INV_X1 U3623 ( .A(n3622), .ZN(n3603) );
  AND3_X1 U3624 ( .A1(n3517), .A2(n4505), .A3(n3253), .ZN(n3523) );
  AND3_X1 U3625 ( .A1(n3575), .A2(n3574), .A3(n3573), .ZN(n3593) );
  NAND2_X1 U3626 ( .A1(n3419), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3898)
         );
  AND2_X1 U3627 ( .A1(n3580), .A2(n3258), .ZN(n4502) );
  AND2_X1 U3628 ( .A1(n3694), .A2(n5282), .ZN(n3145) );
  INV_X1 U3629 ( .A(n4078), .ZN(n4109) );
  OR2_X1 U3630 ( .A1(n4533), .A2(n4617), .ZN(n4580) );
  AND2_X1 U3631 ( .A1(n3578), .A2(n3577), .ZN(n4578) );
  AND2_X1 U3632 ( .A1(n4133), .A2(n3540), .ZN(n3559) );
  NOR2_X1 U3633 ( .A1(n3508), .A2(n4524), .ZN(n4238) );
  NAND2_X1 U3634 ( .A1(n5424), .A2(n4221), .ZN(n5297) );
  NAND2_X1 U3635 ( .A1(n3548), .A2(n3109), .ZN(n4253) );
  NAND2_X1 U3637 ( .A1(n4128), .A2(n3259), .ZN(n3492) );
  NAND2_X1 U3638 ( .A1(n4075), .A2(n3493), .ZN(n4128) );
  INV_X2 U3639 ( .A(n5439), .ZN(n5424) );
  INV_X1 U3640 ( .A(n3453), .ZN(n3494) );
  NAND2_X2 U3641 ( .A1(n4130), .A2(n3554), .ZN(n4221) );
  NOR2_X2 U3642 ( .A1(n4680), .A2(n6632), .ZN(n3878) );
  OR2_X1 U3643 ( .A1(n3571), .A2(n3570), .ZN(n4245) );
  NAND4_X1 U3644 ( .A1(n3538), .A2(n3190), .A3(n3108), .A4(n3539), .ZN(n4308)
         );
  CLKBUF_X2 U3645 ( .A(n3453), .Z(n4697) );
  INV_X2 U3646 ( .A(n4134), .ZN(n3502) );
  AOI21_X1 U3647 ( .B1(n3353), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n3191), 
        .ZN(n3190) );
  AND2_X2 U3648 ( .A1(n4668), .A2(n4134), .ZN(n5439) );
  AND3_X1 U3649 ( .A1(n3392), .A2(n3391), .A3(n3390), .ZN(n3403) );
  OR2_X2 U3650 ( .A1(n3452), .A2(n3451), .ZN(n4668) );
  NAND2_X2 U3651 ( .A1(n3414), .A2(n3413), .ZN(n4693) );
  AND4_X2 U3652 ( .A1(n3442), .A2(n3117), .A3(n3441), .A4(n3440), .ZN(n4703)
         );
  AND4_X1 U3653 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3472)
         );
  AND4_X1 U3654 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3473)
         );
  AND4_X1 U3655 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3413)
         );
  AND4_X1 U3656 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3404)
         );
  AND4_X1 U3657 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(n3440)
         );
  AND4_X1 U3658 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3414)
         );
  AND4_X1 U3659 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3370)
         );
  AND4_X1 U3660 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3402)
         );
  AND4_X1 U3661 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3371)
         );
  AND4_X1 U3662 ( .A1(n3435), .A2(n3434), .A3(n3433), .A4(n3432), .ZN(n3441)
         );
  AND4_X1 U3663 ( .A1(n3457), .A2(n3456), .A3(n3455), .A4(n3454), .ZN(n3474)
         );
  AND4_X1 U3664 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(n3489)
         );
  AND4_X1 U3665 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  BUF_X2 U3666 ( .A(n3564), .Z(n3990) );
  CLKBUF_X1 U3667 ( .A(n3840), .Z(n3989) );
  BUF_X2 U3668 ( .A(n3565), .Z(n3998) );
  BUF_X2 U3669 ( .A(n3482), .Z(n3956) );
  INV_X2 U3670 ( .A(n4460), .ZN(n3100) );
  AND2_X2 U3671 ( .A1(n3271), .A2(n4538), .ZN(n3431) );
  INV_X1 U3672 ( .A(n3477), .ZN(n4725) );
  AND2_X2 U3673 ( .A1(n3272), .A2(n4717), .ZN(n3565) );
  AND2_X2 U3674 ( .A1(n4537), .A2(n4717), .ZN(n3477) );
  INV_X2 U3675 ( .A(n4019), .ZN(n3101) );
  INV_X1 U3676 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5262) );
  AND2_X2 U3677 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4717) );
  NOR2_X2 U3678 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4718) );
  AND2_X2 U3679 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4537) );
  INV_X4 U3680 ( .A(n4633), .ZN(n3554) );
  NAND2_X1 U3681 ( .A1(n4664), .A2(n5282), .ZN(n3640) );
  XNOR2_X1 U3682 ( .A(n4516), .B(n5075), .ZN(n4664) );
  OAI21_X2 U3683 ( .B1(n5814), .B2(n5813), .A(n5811), .ZN(n5802) );
  NAND2_X2 U3684 ( .A1(n5485), .A2(n3111), .ZN(n5411) );
  NOR2_X2 U3685 ( .A1(n3765), .A2(n6809), .ZN(n3807) );
  AOI211_X2 U3686 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6319), .A(n5463), .B(n5462), 
        .ZN(n5464) );
  AOI211_X2 U3687 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n6330), .A(n6329), 
        .B(n6328), .ZN(n6331) );
  XNOR2_X2 U3688 ( .A(n3138), .B(n5307), .ZN(n4398) );
  OAI21_X1 U3689 ( .B1(n5346), .B2(n5348), .A(n5347), .ZN(n5722) );
  XNOR2_X1 U3690 ( .A(n3686), .B(n3687), .ZN(n4625) );
  BUF_X4 U3692 ( .A(n5363), .Z(n3105) );
  NAND3_X2 U3693 ( .A1(n4398), .A2(STATE2_REG_1__SCAN_IN), .A3(n6278), .ZN(
        n5363) );
  NAND2_X1 U3694 ( .A1(n3107), .A2(n3120), .ZN(n3186) );
  OAI21_X1 U3695 ( .B1(n3719), .B2(n3674), .A(n4304), .ZN(n4288) );
  INV_X1 U3696 ( .A(n4308), .ZN(n3540) );
  AND2_X1 U3697 ( .A1(n4133), .A2(n4308), .ZN(n3558) );
  INV_X1 U3698 ( .A(n4668), .ZN(n4130) );
  NOR2_X1 U3699 ( .A1(n4852), .A2(n5282), .ZN(n4066) );
  NAND2_X1 U3700 ( .A1(n4413), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4064) );
  AND2_X1 U3701 ( .A1(n3207), .A2(n5409), .ZN(n3206) );
  NAND2_X1 U3702 ( .A1(n3224), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U3703 ( .A1(n3197), .A2(n3119), .ZN(n3194) );
  AND2_X1 U3704 ( .A1(n3228), .A2(n4319), .ZN(n3227) );
  NAND2_X1 U3705 ( .A1(n3219), .A2(n5246), .ZN(n3173) );
  AND2_X1 U3706 ( .A1(n5247), .A2(n5875), .ZN(n3219) );
  OAI211_X1 U3707 ( .C1(n4109), .C2(n3557), .A(n3556), .B(n3555), .ZN(n3694)
         );
  INV_X1 U3708 ( .A(n4200), .ZN(n5441) );
  NAND2_X1 U3709 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4048)
         );
  AND2_X1 U3710 ( .A1(n3210), .A2(n3209), .ZN(n3208) );
  INV_X1 U3711 ( .A(n5322), .ZN(n3209) );
  INV_X1 U3712 ( .A(n3185), .ZN(n3184) );
  OAI21_X1 U3713 ( .B1(n3187), .B2(n3186), .A(n4330), .ZN(n3185) );
  OR2_X1 U3714 ( .A1(n4595), .A2(n4570), .ZN(n4571) );
  NAND2_X2 U3715 ( .A1(n4125), .A2(n4124), .ZN(n4876) );
  NAND2_X1 U3716 ( .A1(n4363), .A2(n4123), .ZN(n4124) );
  NAND2_X1 U3717 ( .A1(n4122), .A2(n4121), .ZN(n4125) );
  NAND2_X1 U3718 ( .A1(n3537), .A2(n3192), .ZN(n3191) );
  NAND2_X1 U3719 ( .A1(n3976), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3192) );
  AND2_X2 U3720 ( .A1(n5262), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3272)
         );
  AND2_X1 U3721 ( .A1(n4102), .A2(n4101), .ZN(n4108) );
  INV_X1 U3722 ( .A(n3721), .ZN(n3170) );
  OR2_X1 U3723 ( .A1(n3231), .A2(n5855), .ZN(n3148) );
  INV_X1 U3724 ( .A(n4315), .ZN(n3231) );
  OR2_X1 U3725 ( .A1(n3671), .A2(n3670), .ZN(n4292) );
  AOI21_X1 U3726 ( .B1(n5129), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4108), 
        .ZN(n4119) );
  NAND2_X1 U3727 ( .A1(n4697), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U3728 ( .A1(n3238), .A2(n5374), .ZN(n3237) );
  INV_X1 U3729 ( .A(n3239), .ZN(n3238) );
  OR2_X1 U3730 ( .A1(n3240), .A2(n5386), .ZN(n3239) );
  INV_X1 U3731 ( .A(n4066), .ZN(n4036) );
  NAND2_X1 U3732 ( .A1(n3256), .A2(n5471), .ZN(n3247) );
  INV_X1 U3733 ( .A(n5485), .ZN(n3248) );
  AND2_X1 U3734 ( .A1(n3836), .A2(n3835), .ZN(n3837) );
  AND2_X1 U3735 ( .A1(n4995), .A2(n4643), .ZN(n3742) );
  NAND2_X1 U3736 ( .A1(n3685), .A2(n3899), .ZN(n3708) );
  NAND2_X1 U3737 ( .A1(n3257), .A2(n3178), .ZN(n3177) );
  NAND2_X1 U3738 ( .A1(n3215), .A2(n5615), .ZN(n3214) );
  INV_X1 U3739 ( .A(n3216), .ZN(n3215) );
  INV_X1 U3740 ( .A(n3148), .ZN(n3230) );
  AOI21_X1 U3741 ( .B1(n3221), .B2(n5875), .A(n3124), .ZN(n3220) );
  INV_X1 U3742 ( .A(n4303), .ZN(n3221) );
  AND2_X1 U3743 ( .A1(n6752), .A2(n5424), .ZN(n4152) );
  OAI21_X1 U3744 ( .B1(n4276), .B2(n4305), .A(n4275), .ZN(n4278) );
  NAND2_X1 U3745 ( .A1(n4152), .A2(n3205), .ZN(n3204) );
  AOI21_X1 U3746 ( .B1(n5281), .B2(n4628), .A(n5267), .ZN(n4630) );
  INV_X1 U3747 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U3748 ( .A1(n3502), .A2(n3554), .ZN(n4391) );
  NOR2_X1 U3749 ( .A1(n4059), .A2(n4344), .ZN(n3139) );
  AND2_X1 U3750 ( .A1(n5336), .A2(n3249), .ZN(n4355) );
  AND2_X1 U3751 ( .A1(n3110), .A2(n3250), .ZN(n3249) );
  INV_X1 U3752 ( .A(n4070), .ZN(n3250) );
  NOR2_X1 U3753 ( .A1(n4048), .A2(n3140), .ZN(n4055) );
  NAND2_X1 U3754 ( .A1(n4055), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4059)
         );
  MUX2_X1 U3755 ( .A(n4049), .B(n5708), .S(n3101), .Z(n5337) );
  NAND2_X1 U3756 ( .A1(n5336), .A2(n5337), .ZN(n5325) );
  INV_X1 U3757 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3881) );
  AND4_X1 U3758 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n5499)
         );
  OR2_X1 U3759 ( .A1(n5515), .A2(n5499), .ZN(n5501) );
  INV_X1 U3760 ( .A(n3896), .ZN(n3419) );
  NAND2_X1 U3761 ( .A1(n3839), .A2(n5614), .ZN(n3172) );
  NAND2_X1 U3762 ( .A1(n3746), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3792)
         );
  NOR2_X1 U3763 ( .A1(n4334), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U3764 ( .A1(n3176), .A2(n3174), .ZN(n5688) );
  NOR2_X1 U3765 ( .A1(n3177), .A2(n3175), .ZN(n3174) );
  INV_X1 U3766 ( .A(n4334), .ZN(n3195) );
  NAND2_X1 U3767 ( .A1(n3176), .A2(n3257), .ZN(n5696) );
  NAND2_X1 U3768 ( .A1(n3182), .A2(n3180), .ZN(n5726) );
  AOI21_X1 U3769 ( .B1(n3184), .B2(n3186), .A(n3181), .ZN(n3180) );
  INV_X1 U3770 ( .A(n5727), .ZN(n3181) );
  INV_X1 U3771 ( .A(n5734), .ZN(n3152) );
  AND2_X1 U3772 ( .A1(n3153), .A2(n3150), .ZN(n3149) );
  NAND2_X1 U3773 ( .A1(n3151), .A2(n5734), .ZN(n3150) );
  NOR2_X1 U3774 ( .A1(n4203), .A2(n5442), .ZN(n3207) );
  NAND2_X1 U3775 ( .A1(n3194), .A2(n3223), .ZN(n5770) );
  NOR2_X1 U3776 ( .A1(n6100), .A2(n3216), .ZN(n5616) );
  OR2_X1 U3777 ( .A1(n3201), .A2(n3200), .ZN(n3199) );
  INV_X1 U3778 ( .A(n5626), .ZN(n3200) );
  AND2_X1 U3779 ( .A1(n4173), .A2(n4172), .ZN(n5543) );
  AOI21_X1 U3780 ( .B1(n5229), .B2(n3157), .A(n3121), .ZN(n3156) );
  INV_X1 U3781 ( .A(n4502), .ZN(n4880) );
  NAND2_X1 U3782 ( .A1(n3693), .A2(n3553), .ZN(n3697) );
  NAND2_X1 U3783 ( .A1(n3692), .A2(n3694), .ZN(n3693) );
  OAI21_X1 U3784 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n4338), .A(n5023), 
        .ZN(n6634) );
  CLKBUF_X1 U3785 ( .A(n4661), .Z(n4662) );
  INV_X1 U3786 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5129) );
  INV_X1 U3787 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U3788 ( .A1(n4390), .A2(REIP_REG_30__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U3789 ( .A1(n4232), .A2(n4231), .ZN(n5927) );
  OR3_X1 U3790 ( .A1(n5414), .A2(n5367), .A3(n4386), .ZN(n5342) );
  AOI21_X1 U3791 ( .B1(n6262), .B2(n3137), .A(n3135), .ZN(n3134) );
  INV_X1 U3792 ( .A(n5708), .ZN(n3137) );
  OR2_X1 U3793 ( .A1(n3136), .A2(n5341), .ZN(n3135) );
  NAND2_X1 U3794 ( .A1(n5357), .A2(REIP_REG_27__SCAN_IN), .ZN(n3133) );
  NOR2_X1 U3795 ( .A1(n4398), .A2(n5263), .ZN(n4370) );
  AND2_X1 U3796 ( .A1(n5557), .A2(n4372), .ZN(n6305) );
  AND2_X1 U3797 ( .A1(n5628), .A2(n4693), .ZN(n6341) );
  OR2_X1 U3798 ( .A1(n4411), .A2(n5296), .ZN(n4135) );
  INV_X2 U3799 ( .A(n6341), .ZN(n7064) );
  OR2_X1 U3800 ( .A1(n4416), .A2(n4412), .ZN(n5070) );
  OAI21_X1 U3801 ( .B1(n5336), .B2(n5337), .A(n5325), .ZN(n5715) );
  OR2_X1 U3802 ( .A1(n5976), .A2(n5914), .ZN(n5955) );
  NAND2_X1 U3803 ( .A1(n4589), .A2(n4586), .ZN(n6440) );
  NAND2_X1 U3804 ( .A1(n4338), .A2(n6632), .ZN(n6636) );
  AND2_X1 U3805 ( .A1(n6582), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4073)
         );
  XNOR2_X1 U3806 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4097) );
  INV_X1 U3807 ( .A(n4276), .ZN(n4268) );
  NAND2_X1 U3808 ( .A1(n4078), .A2(n4297), .ZN(n4114) );
  AND2_X2 U3809 ( .A1(n3264), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3271)
         );
  NAND2_X1 U3810 ( .A1(n4633), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3627) );
  INV_X1 U3811 ( .A(n3694), .ZN(n3144) );
  AOI22_X1 U3812 ( .A1(n3476), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U3813 ( .A1(n3476), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U3814 ( .A1(n3377), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3477), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U3815 ( .A1(n3226), .A2(n3225), .ZN(n4281) );
  INV_X1 U3816 ( .A(n3719), .ZN(n3226) );
  NAND2_X1 U3817 ( .A1(n3198), .A2(n3729), .ZN(n3720) );
  INV_X1 U3818 ( .A(n3628), .ZN(n4133) );
  INV_X1 U3819 ( .A(n3493), .ZN(n3698) );
  NOR2_X1 U3820 ( .A1(n5326), .A2(n3252), .ZN(n3251) );
  INV_X1 U3821 ( .A(n5337), .ZN(n3252) );
  OR2_X1 U3822 ( .A1(n3348), .A2(n3347), .ZN(n4033) );
  NAND2_X1 U3823 ( .A1(n3241), .A2(n5395), .ZN(n3240) );
  NOR2_X1 U3824 ( .A1(n3244), .A2(n3243), .ZN(n3242) );
  INV_X1 U3825 ( .A(n5436), .ZN(n3243) );
  NAND2_X1 U3826 ( .A1(n3245), .A2(n5453), .ZN(n3244) );
  INV_X1 U3827 ( .A(n3247), .ZN(n3245) );
  INV_X1 U3828 ( .A(n3878), .ZN(n3904) );
  NOR2_X2 U3829 ( .A1(n5324), .A2(n5277), .ZN(n5274) );
  AND2_X1 U3830 ( .A1(n3211), .A2(n5339), .ZN(n3210) );
  AND2_X1 U3831 ( .A1(n5359), .A2(n5353), .ZN(n3211) );
  NOR2_X1 U3832 ( .A1(n4324), .A2(n3188), .ZN(n3187) );
  INV_X1 U3833 ( .A(n3220), .ZN(n3164) );
  INV_X1 U3834 ( .A(n3558), .ZN(n4306) );
  INV_X1 U3835 ( .A(n3223), .ZN(n3151) );
  AOI21_X1 U3836 ( .B1(n5771), .B2(n5734), .A(n3154), .ZN(n3153) );
  INV_X1 U3837 ( .A(n5766), .ZN(n3154) );
  OR2_X1 U3838 ( .A1(n6099), .A2(n3217), .ZN(n3216) );
  INV_X1 U3839 ( .A(n5530), .ZN(n3217) );
  INV_X1 U3840 ( .A(n4152), .ZN(n4210) );
  OR2_X1 U3841 ( .A1(n5225), .A2(n4421), .ZN(n3201) );
  INV_X1 U3842 ( .A(n4287), .ZN(n3157) );
  OAI21_X1 U3843 ( .B1(n4288), .B2(n4305), .A(n4294), .ZN(n4296) );
  AND2_X1 U3844 ( .A1(n4688), .A2(n4684), .ZN(n4297) );
  NAND2_X1 U3845 ( .A1(n3236), .A2(n3235), .ZN(n3619) );
  INV_X1 U3846 ( .A(n3730), .ZN(n3729) );
  INV_X1 U3847 ( .A(n4114), .ZN(n4120) );
  AOI221_X1 U3848 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4119), .C1(
        n4113), .C2(n4119), .A(n4118), .ZN(n4363) );
  INV_X1 U3849 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U3850 ( .A1(n3483), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3458)
         );
  AND4_X2 U3851 ( .A1(n3404), .A2(n3403), .A3(n3401), .A4(n3402), .ZN(n3453)
         );
  OR2_X1 U3852 ( .A1(n3638), .A2(n3637), .ZN(n4269) );
  INV_X1 U3853 ( .A(n3683), .ZN(n3684) );
  NOR2_X1 U3854 ( .A1(n6307), .A2(n3140), .ZN(n3136) );
  AND2_X1 U3855 ( .A1(n4159), .A2(n4158), .ZN(n5234) );
  AND2_X1 U3856 ( .A1(n4184), .A2(n4183), .ZN(n5615) );
  NOR2_X1 U3857 ( .A1(n4497), .A2(READY_N), .ZN(n4800) );
  NAND2_X1 U3858 ( .A1(n4684), .A2(n4800), .ZN(n4802) );
  AND2_X1 U3859 ( .A1(n6632), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4352) );
  INV_X1 U3860 ( .A(n3139), .ZN(n4356) );
  AOI21_X1 U3861 ( .B1(n5314), .B2(n3101), .A(n4068), .ZN(n4337) );
  AND2_X1 U3862 ( .A1(n3421), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4038)
         );
  NOR2_X1 U3863 ( .A1(n4011), .A2(n3142), .ZN(n4022) );
  NAND2_X1 U3864 ( .A1(n4022), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4031)
         );
  OAI21_X1 U3865 ( .B1(n5748), .B2(n4019), .A(n4018), .ZN(n5386) );
  NOR2_X1 U3866 ( .A1(n3986), .A2(n5761), .ZN(n4007) );
  NAND2_X1 U3867 ( .A1(n4007), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4011)
         );
  OR2_X1 U3868 ( .A1(n3952), .A2(n3951), .ZN(n3954) );
  OR2_X1 U3869 ( .A1(n3954), .A2(n6962), .ZN(n3986) );
  NAND2_X1 U3870 ( .A1(n3934), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3952)
         );
  AND2_X1 U3871 ( .A1(n3420), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3934)
         );
  INV_X1 U3872 ( .A(n3919), .ZN(n3420) );
  AND2_X1 U3873 ( .A1(n3921), .A2(n3920), .ZN(n5471) );
  NAND2_X1 U3874 ( .A1(n3141), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3919)
         );
  INV_X1 U3875 ( .A(n3256), .ZN(n3246) );
  NAND2_X1 U3876 ( .A1(n3831), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3896)
         );
  AND2_X1 U3877 ( .A1(n3815), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3831)
         );
  AND2_X1 U3878 ( .A1(n3807), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3815)
         );
  AND2_X1 U3879 ( .A1(n3169), .A2(n3750), .ZN(n3166) );
  NAND2_X1 U3880 ( .A1(n3751), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3765)
         );
  INV_X1 U3881 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6809) );
  OR2_X1 U3882 ( .A1(n5624), .A2(n5541), .ZN(n5675) );
  NOR2_X1 U3883 ( .A1(n3792), .A2(n3418), .ZN(n3751) );
  INV_X1 U3884 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U3885 ( .A1(n5067), .A2(n3750), .ZN(n4428) );
  AND2_X1 U3886 ( .A1(n3722), .A2(n3127), .ZN(n3746) );
  AND2_X1 U3887 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3733), .ZN(n3722)
         );
  NOR2_X1 U3888 ( .A1(n3732), .A2(n4711), .ZN(n3733) );
  NAND2_X1 U3889 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3732) );
  AND2_X1 U3890 ( .A1(n4212), .A2(n4211), .ZN(n5376) );
  INV_X1 U3891 ( .A(n3197), .ZN(n5778) );
  AND2_X1 U3892 ( .A1(n4193), .A2(n4192), .ZN(n5469) );
  NOR2_X2 U3893 ( .A1(n5514), .A2(n5498), .ZN(n5497) );
  OR2_X1 U3894 ( .A1(n4327), .A2(n6059), .ZN(n5811) );
  NAND2_X1 U3895 ( .A1(n3189), .A2(n3159), .ZN(n5814) );
  NOR2_X1 U3896 ( .A1(n3188), .A2(n3160), .ZN(n3159) );
  NOR2_X1 U3897 ( .A1(n3224), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3160)
         );
  AND2_X1 U3898 ( .A1(n4186), .A2(n4185), .ZN(n5512) );
  NAND2_X1 U3899 ( .A1(n5864), .A2(n3193), .ZN(n3165) );
  OR2_X1 U3900 ( .A1(n6440), .A2(n5891), .ZN(n6068) );
  NAND2_X1 U3901 ( .A1(n3232), .A2(n3230), .ZN(n5834) );
  OR2_X1 U3902 ( .A1(n3099), .A2(n6963), .ZN(n5854) );
  NAND2_X1 U3903 ( .A1(n4314), .A2(n3254), .ZN(n3232) );
  INV_X1 U3904 ( .A(n5864), .ZN(n4314) );
  INV_X1 U3905 ( .A(n5543), .ZN(n4174) );
  NAND2_X1 U3906 ( .A1(n3173), .A2(n3220), .ZN(n5864) );
  OR2_X1 U3907 ( .A1(n5222), .A2(n5225), .ZN(n5223) );
  NOR2_X1 U3908 ( .A1(n4142), .A2(n3202), .ZN(n4651) );
  NAND2_X1 U3909 ( .A1(n3204), .A2(n3203), .ZN(n3202) );
  NAND2_X1 U3910 ( .A1(n5439), .A2(EBX_REG_3__SCAN_IN), .ZN(n3203) );
  AND2_X1 U3911 ( .A1(n5903), .A2(n4657), .ZN(n5910) );
  XNOR2_X1 U3912 ( .A(n3598), .B(n3590), .ZN(n4522) );
  INV_X1 U3913 ( .A(n3597), .ZN(n3590) );
  NAND2_X1 U3914 ( .A1(n3730), .A2(n4765), .ZN(n4624) );
  OR2_X1 U3916 ( .A1(n3512), .A2(n3514), .ZN(n4852) );
  INV_X1 U3917 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4733) );
  OR2_X1 U3918 ( .A1(n5577), .A2(n5582), .ZN(n6586) );
  INV_X1 U3919 ( .A(n6117), .ZN(n6540) );
  OR2_X1 U3920 ( .A1(n6628), .A2(n3102), .ZN(n5165) );
  INV_X1 U3921 ( .A(n6617), .ZN(n5211) );
  INV_X1 U3922 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6582) );
  AND2_X1 U3923 ( .A1(n3102), .A2(n5164), .ZN(n6539) );
  OR2_X1 U3924 ( .A1(n4893), .A2(n4662), .ZN(n6628) );
  NAND2_X1 U3925 ( .A1(n4632), .A2(n4631), .ZN(n4702) );
  INV_X1 U3926 ( .A(n5023), .ZN(n6192) );
  OR2_X1 U3927 ( .A1(n4499), .A2(n5114), .ZN(n4496) );
  INV_X1 U3928 ( .A(n3520), .ZN(n6753) );
  INV_X1 U3929 ( .A(n6330), .ZN(n6307) );
  OR2_X1 U3930 ( .A1(n5357), .A2(n4389), .ZN(n5327) );
  INV_X1 U3931 ( .A(n5312), .ZN(n5313) );
  INV_X1 U3932 ( .A(n6320), .ZN(n6285) );
  INV_X1 U3933 ( .A(n5554), .ZN(n6299) );
  AND2_X1 U3934 ( .A1(n5557), .A2(n4395), .ZN(n6319) );
  NAND2_X1 U3935 ( .A1(n4198), .A2(n4197), .ZN(n5423) );
  INV_X1 U3936 ( .A(n4693), .ZN(n4413) );
  AND2_X1 U3937 ( .A1(n5070), .A2(n4620), .ZN(n5662) );
  AND2_X1 U3938 ( .A1(n4416), .A2(n4415), .ZN(n5661) );
  NAND2_X2 U3939 ( .A1(n5070), .A2(n4619), .ZN(n5683) );
  NOR2_X1 U3940 ( .A1(n4628), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6376) );
  AND2_X1 U3941 ( .A1(n4598), .A2(n4597), .ZN(n6381) );
  NAND2_X1 U3942 ( .A1(n6398), .A2(n4596), .ZN(n4598) );
  OR2_X1 U3943 ( .A1(n4595), .A2(n4594), .ZN(n4596) );
  NAND2_X1 U3944 ( .A1(n3139), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3138)
         );
  AND2_X1 U3945 ( .A1(n4059), .A2(n4057), .ZN(n5701) );
  INV_X1 U3946 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5761) );
  INV_X1 U3947 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6962) );
  INV_X1 U3948 ( .A(n3141), .ZN(n3864) );
  AND2_X1 U3949 ( .A1(n5501), .A2(n5500), .ZN(n5819) );
  INV_X1 U3950 ( .A(n3172), .ZN(n3171) );
  NAND2_X1 U3951 ( .A1(n6226), .A2(n4340), .ZN(n5868) );
  INV_X1 U3952 ( .A(n5868), .ZN(n6410) );
  OAI21_X1 U3953 ( .B1(n3115), .B2(n5685), .A(n5684), .ZN(n5689) );
  AOI21_X1 U3954 ( .B1(n3178), .B2(n5696), .A(n5700), .ZN(n5949) );
  NAND2_X1 U3955 ( .A1(n3179), .A2(n3184), .ZN(n5728) );
  OR2_X1 U3956 ( .A1(n3189), .A2(n3186), .ZN(n3179) );
  OAI21_X1 U3957 ( .B1(n5770), .B2(n5771), .A(n5734), .ZN(n5765) );
  AND2_X1 U3958 ( .A1(n4198), .A2(n3207), .ZN(n5410) );
  NAND2_X1 U3959 ( .A1(n5246), .A2(n5247), .ZN(n3222) );
  OR2_X1 U3960 ( .A1(n5903), .A2(n4590), .ZN(n6420) );
  AND2_X1 U3961 ( .A1(n4589), .A2(n4581), .ZN(n6432) );
  INV_X1 U3962 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6225) );
  INV_X1 U3963 ( .A(n4662), .ZN(n5010) );
  INV_X1 U3964 ( .A(n6636), .ZN(n6626) );
  CLKBUF_X1 U3965 ( .A(n4543), .Z(n5577) );
  INV_X1 U3966 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5263) );
  NOR2_X1 U3967 ( .A1(n4876), .A2(n4338), .ZN(n5267) );
  NOR2_X1 U3968 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6123) );
  AND2_X1 U3969 ( .A1(n4520), .A2(n4892), .ZN(n6129) );
  INV_X1 U3970 ( .A(n6137), .ZN(n4956) );
  AND3_X1 U3971 ( .A1(n4893), .A2(n5010), .A3(n5073), .ZN(n6478) );
  NOR2_X1 U3972 ( .A1(n4629), .A2(n5164), .ZN(n6513) );
  INV_X1 U3973 ( .A(n6650), .ZN(n6599) );
  INV_X1 U3974 ( .A(n6657), .ZN(n6603) );
  INV_X1 U3975 ( .A(n6149), .ZN(n6179) );
  NOR2_X1 U3976 ( .A1(n5000), .A2(n6192), .ZN(n6673) );
  INV_X1 U3977 ( .A(n6712), .ZN(n6199) );
  OAI21_X1 U3978 ( .B1(n4674), .B2(n4673), .A(n4672), .ZN(n4706) );
  NOR2_X2 U3979 ( .A1(n4666), .A2(n5164), .ZN(n6703) );
  AOI22_X1 U3980 ( .A1(n4670), .A2(n4673), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6194), .ZN(n4709) );
  INV_X1 U3981 ( .A(n6623), .ZN(n6711) );
  INV_X1 U3982 ( .A(n4897), .ZN(n6723) );
  OR4_X1 U3983 ( .A1(n4884), .A2(n4883), .A3(n4882), .A4(n5290), .ZN(n4886) );
  NAND2_X1 U3984 ( .A1(n4129), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5114) );
  AND2_X1 U3985 ( .A1(n4457), .A2(n6750), .ZN(n6741) );
  NOR2_X1 U3986 ( .A1(n4405), .A2(n4404), .ZN(n4406) );
  OAI211_X1 U3987 ( .C1(n5342), .C2(REIP_REG_27__SCAN_IN), .A(n3134), .B(n3133), .ZN(n5343) );
  AOI21_X1 U3988 ( .B1(n4235), .B2(n4234), .A(n4233), .ZN(n4236) );
  NOR2_X1 U3989 ( .A1(n5628), .A2(n4400), .ZN(n4233) );
  OAI21_X1 U3990 ( .B1(n5634), .B2(n7064), .A(n3146), .ZN(U2831) );
  INV_X1 U3991 ( .A(n3147), .ZN(n3146) );
  OAI22_X1 U3992 ( .A1(n5945), .A2(n7065), .B1(n5598), .B2(n5628), .ZN(n3147)
         );
  OR2_X1 U3993 ( .A1(n5411), .A2(n3240), .ZN(n5385) );
  NOR2_X1 U3994 ( .A1(n3248), .A2(n3247), .ZN(n5454) );
  NOR2_X1 U3995 ( .A1(n3248), .A2(n3246), .ZN(n5472) );
  AND2_X1 U3996 ( .A1(n3169), .A2(n5066), .ZN(n5067) );
  NAND2_X1 U3997 ( .A1(n4333), .A2(n3125), .ZN(n3106) );
  AND2_X1 U3998 ( .A1(n5811), .A2(n4326), .ZN(n3107) );
  AND4_X1 U3999 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3108)
         );
  AND4_X1 U4000 ( .A1(n3122), .A2(n3547), .A3(n3545), .A4(n3546), .ZN(n3109)
         );
  NAND2_X1 U4001 ( .A1(n3171), .A2(n3852), .ZN(n5613) );
  AND2_X1 U4002 ( .A1(n3251), .A2(n4337), .ZN(n3110) );
  AND2_X1 U4003 ( .A1(n3970), .A2(n3242), .ZN(n3111) );
  AND2_X1 U4004 ( .A1(n5066), .A2(n3128), .ZN(n3112) );
  AND2_X1 U4005 ( .A1(n3206), .A2(n3132), .ZN(n3113) );
  AND2_X1 U4006 ( .A1(n3711), .A2(n3710), .ZN(n4612) );
  AND2_X1 U4007 ( .A1(n3528), .A2(n3597), .ZN(n3114) );
  OR2_X1 U4008 ( .A1(n5719), .A2(n3177), .ZN(n3115) );
  INV_X1 U4009 ( .A(n4327), .ZN(n3224) );
  AND2_X1 U4010 ( .A1(n3166), .A2(n3112), .ZN(n5526) );
  NAND2_X1 U4011 ( .A1(n3168), .A2(n3167), .ZN(n3750) );
  NAND2_X1 U4012 ( .A1(n4198), .A2(n3206), .ZN(n5401) );
  NAND2_X1 U4013 ( .A1(n5485), .A2(n3242), .ZN(n5420) );
  NAND2_X1 U4014 ( .A1(n3502), .A2(n4633), .ZN(n3520) );
  BUF_X2 U4015 ( .A(n3529), .Z(n3542) );
  AND2_X1 U4016 ( .A1(n3165), .A2(n3227), .ZN(n3116) );
  OAI21_X1 U4017 ( .B1(n3603), .B2(n4733), .A(n3602), .ZN(n3620) );
  AND4_X1 U4018 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3117)
         );
  INV_X1 U4019 ( .A(n3497), .ZN(n4075) );
  NAND2_X1 U4020 ( .A1(n3232), .A2(n4315), .ZN(n5857) );
  NAND2_X1 U4021 ( .A1(n3222), .A2(n4303), .ZN(n5874) );
  INV_X1 U4022 ( .A(n5821), .ZN(n3188) );
  BUF_X2 U4023 ( .A(n3543), .Z(n3544) );
  AND2_X1 U4024 ( .A1(n3852), .A2(n3839), .ZN(n3118) );
  NAND2_X1 U4025 ( .A1(n3682), .A2(n3681), .ZN(n5066) );
  NAND2_X1 U4026 ( .A1(n4327), .A2(n5732), .ZN(n3119) );
  AND2_X1 U4027 ( .A1(n5375), .A2(n5359), .ZN(n5351) );
  NAND2_X1 U4028 ( .A1(n3224), .A2(n4329), .ZN(n3120) );
  AND2_X1 U4029 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3121)
         );
  NOR2_X1 U4030 ( .A1(n5411), .A2(n3239), .ZN(n5373) );
  NAND2_X1 U4031 ( .A1(n5726), .A2(n4331), .ZN(n5719) );
  INV_X1 U4032 ( .A(n5719), .ZN(n3176) );
  AND4_X1 U4033 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3122)
         );
  AND2_X1 U4034 ( .A1(n3587), .A2(n3588), .ZN(n3123) );
  AND2_X1 U4035 ( .A1(n4313), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3124)
         );
  NAND2_X1 U4036 ( .A1(n5375), .A2(n3210), .ZN(n5321) );
  NAND2_X1 U4037 ( .A1(n5375), .A2(n3208), .ZN(n5324) );
  AND2_X1 U4038 ( .A1(n5375), .A2(n3211), .ZN(n5338) );
  NOR2_X1 U4039 ( .A1(n3248), .A2(n3244), .ZN(n5435) );
  AND2_X1 U4040 ( .A1(n4332), .A2(n3195), .ZN(n3125) );
  NOR2_X1 U4041 ( .A1(n5865), .A2(n4321), .ZN(n3126) );
  AND2_X1 U4042 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3127) );
  INV_X1 U4043 ( .A(n3254), .ZN(n3233) );
  AND4_X1 U4044 ( .A1(n5621), .A2(n5539), .A3(n4427), .A4(n5673), .ZN(n3128)
         );
  OR2_X1 U4045 ( .A1(n6100), .A2(n3214), .ZN(n5511) );
  NOR2_X1 U4046 ( .A1(n6100), .A2(n6099), .ZN(n5529) );
  NOR2_X1 U4047 ( .A1(n4759), .A2(n4758), .ZN(n4760) );
  NOR2_X1 U4048 ( .A1(n5222), .A2(n3201), .ZN(n4422) );
  NAND2_X1 U4049 ( .A1(n3158), .A2(n4287), .ZN(n5228) );
  OAI21_X1 U4050 ( .B1(n4281), .B2(n3904), .A(n3728), .ZN(n4995) );
  AND2_X1 U4051 ( .A1(n4332), .A2(n3196), .ZN(n3129) );
  AND2_X1 U4052 ( .A1(n5497), .A2(n5487), .ZN(n5468) );
  AND2_X1 U4053 ( .A1(n3128), .A2(n5527), .ZN(n3130) );
  OR2_X1 U4054 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4019) );
  NAND2_X1 U4055 ( .A1(n3722), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3131)
         );
  NAND2_X1 U4056 ( .A1(n4207), .A2(n4206), .ZN(n3132) );
  INV_X1 U4057 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3142) );
  INV_X1 U4058 ( .A(EBX_REG_3__SCAN_IN), .ZN(n3205) );
  INV_X1 U4059 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3140) );
  INV_X1 U4060 ( .A(n5918), .ZN(n3178) );
  INV_X1 U4061 ( .A(n5919), .ZN(n3175) );
  NOR2_X2 U4062 ( .A1(n3898), .A2(n3881), .ZN(n3141) );
  NAND3_X1 U4063 ( .A1(n3145), .A2(n3597), .A3(n3528), .ZN(n3143) );
  NAND3_X1 U4064 ( .A1(n3528), .A2(n3597), .A3(n5282), .ZN(n3692) );
  MUX2_X1 U4065 ( .A(n3558), .B(n3559), .S(n4253), .Z(n3695) );
  INV_X1 U4066 ( .A(n4320), .ZN(n3229) );
  AOI21_X1 U4067 ( .B1(n3193), .B2(n3164), .A(n3126), .ZN(n3163) );
  NOR2_X1 U4068 ( .A1(n3148), .A2(n4320), .ZN(n3193) );
  OAI21_X2 U4069 ( .B1(n3194), .B2(n3152), .A(n3149), .ZN(n5764) );
  INV_X1 U4070 ( .A(n5764), .ZN(n5735) );
  NAND2_X2 U4071 ( .A1(n3155), .A2(n3156), .ZN(n5246) );
  NAND3_X1 U4072 ( .A1(n5098), .A2(n5099), .A3(n5229), .ZN(n3155) );
  NAND2_X1 U4073 ( .A1(n5098), .A2(n5099), .ZN(n3158) );
  INV_X1 U4074 ( .A(n3173), .ZN(n3162) );
  NAND3_X2 U4075 ( .A1(n3163), .A2(n3227), .A3(n3161), .ZN(n3189) );
  NAND2_X1 U4076 ( .A1(n3162), .A2(n3193), .ZN(n3161) );
  NAND4_X1 U4077 ( .A1(n3169), .A2(n3130), .A3(n5066), .A4(n3750), .ZN(n3838)
         );
  INV_X1 U4078 ( .A(n3750), .ZN(n5220) );
  INV_X1 U4079 ( .A(n3749), .ZN(n3167) );
  NAND2_X1 U4080 ( .A1(n4298), .A2(n3878), .ZN(n3168) );
  NAND2_X1 U4081 ( .A1(n3189), .A2(n3184), .ZN(n3182) );
  NAND2_X1 U4082 ( .A1(n3189), .A2(n3187), .ZN(n3183) );
  AND2_X2 U4083 ( .A1(n4718), .A2(n4537), .ZN(n3536) );
  AND2_X2 U4084 ( .A1(n4718), .A2(n4538), .ZN(n3462) );
  AND2_X2 U4085 ( .A1(n3270), .A2(n4718), .ZN(n3377) );
  AND2_X2 U4086 ( .A1(n3272), .A2(n4718), .ZN(n3564) );
  NAND2_X1 U4087 ( .A1(n4333), .A2(n3129), .ZN(n5686) );
  NAND2_X1 U4088 ( .A1(n4333), .A2(n4332), .ZN(n5710) );
  INV_X1 U4089 ( .A(n5686), .ZN(n4349) );
  OR2_X2 U4090 ( .A1(n5222), .A2(n3199), .ZN(n5625) );
  NAND2_X1 U4091 ( .A1(n4198), .A2(n3113), .ZN(n5402) );
  AND2_X2 U4092 ( .A1(n3218), .A2(n4538), .ZN(n3372) );
  AND2_X2 U4093 ( .A1(n3270), .A2(n3218), .ZN(n3482) );
  AND2_X4 U4094 ( .A1(n3272), .A2(n3218), .ZN(n3840) );
  AND2_X2 U4095 ( .A1(n3265), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3218)
         );
  OR2_X1 U4096 ( .A1(n4281), .A2(n4305), .ZN(n4284) );
  NAND2_X1 U4097 ( .A1(n3720), .A2(n3721), .ZN(n3225) );
  NAND3_X1 U4098 ( .A1(n3233), .A2(n3229), .A3(n3230), .ZN(n3228) );
  NAND2_X1 U4099 ( .A1(n3589), .A2(n3597), .ZN(n3235) );
  NAND2_X2 U4100 ( .A1(n3527), .A2(n3526), .ZN(n3597) );
  NAND2_X1 U4101 ( .A1(n3236), .A2(n3589), .ZN(n3598) );
  INV_X1 U4102 ( .A(n3619), .ZN(n3621) );
  OR2_X2 U4103 ( .A1(n5411), .A2(n3237), .ZN(n5361) );
  NOR2_X1 U4104 ( .A1(n5411), .A2(n5412), .ZN(n5394) );
  INV_X1 U4105 ( .A(n5412), .ZN(n3241) );
  NAND2_X1 U4106 ( .A1(n5336), .A2(n3110), .ZN(n4069) );
  AND2_X1 U4107 ( .A1(n5336), .A2(n3251), .ZN(n4336) );
  OAI211_X1 U4108 ( .C1(n3493), .C2(n4239), .A(n4128), .B(n4693), .ZN(n3508)
         );
  AND2_X1 U4109 ( .A1(n4558), .A2(n4257), .ZN(n6403) );
  OR2_X1 U4110 ( .A1(n5686), .A2(n4348), .ZN(n5687) );
  INV_X1 U4111 ( .A(n4258), .ZN(n4259) );
  NAND2_X1 U4112 ( .A1(n4243), .A2(n4242), .ZN(n4258) );
  XNOR2_X1 U4113 ( .A(n4335), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5942)
         );
  NAND2_X1 U4114 ( .A1(n3115), .A2(n3106), .ZN(n4335) );
  OR2_X1 U4115 ( .A1(n5312), .A2(n5873), .ZN(n4347) );
  OR2_X2 U4116 ( .A1(n3383), .A2(n3382), .ZN(n3497) );
  INV_X1 U4117 ( .A(n3579), .ZN(n3580) );
  NAND2_X1 U4118 ( .A1(n5291), .A2(n4414), .ZN(n4418) );
  NAND2_X2 U4119 ( .A1(n4136), .A2(n4135), .ZN(n5628) );
  INV_X2 U4120 ( .A(n6398), .ZN(n4837) );
  INV_X2 U4121 ( .A(n4801), .ZN(n6396) );
  AND3_X1 U4122 ( .A1(n4726), .A2(n4221), .A3(n6730), .ZN(n3253) );
  INV_X1 U4123 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4338) );
  OR2_X1 U4124 ( .A1(n3099), .A2(n6438), .ZN(n3254) );
  INV_X1 U4125 ( .A(n5927), .ZN(n4235) );
  AND2_X1 U4126 ( .A1(n4353), .A2(EAX_REG_5__SCAN_IN), .ZN(n3255) );
  AND2_X1 U4127 ( .A1(n3260), .A2(n5516), .ZN(n3256) );
  AND2_X1 U4128 ( .A1(n3099), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3257)
         );
  NAND2_X2 U4129 ( .A1(n5628), .A2(n4413), .ZN(n7065) );
  INV_X1 U4130 ( .A(n7065), .ZN(n4234) );
  INV_X1 U4131 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4447) );
  AND2_X1 U4132 ( .A1(n4447), .A2(STATE_REG_1__SCAN_IN), .ZN(n6751) );
  INV_X1 U4133 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4113) );
  INV_X1 U4134 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U4135 ( .A1(n4239), .A2(n3554), .ZN(n3258) );
  AND2_X1 U4136 ( .A1(n3453), .A2(n4693), .ZN(n3259) );
  NOR2_X1 U4137 ( .A1(n5486), .A2(n5499), .ZN(n3260) );
  AND3_X1 U4138 ( .A1(n3780), .A2(n3779), .A3(n3778), .ZN(n3261) );
  AND3_X1 U4139 ( .A1(n3764), .A2(n3763), .A3(n3762), .ZN(n3262) );
  OR2_X1 U4140 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  INV_X1 U4141 ( .A(n3712), .ZN(n3651) );
  NOR2_X1 U4142 ( .A1(n3613), .A2(n3612), .ZN(n4240) );
  XNOR2_X1 U4143 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4101) );
  OR2_X1 U4144 ( .A1(n4021), .A2(n4020), .ZN(n4026) );
  AND2_X1 U4145 ( .A1(n3389), .A2(n3388), .ZN(n3392) );
  OR2_X1 U4146 ( .A1(n3661), .A2(n3660), .ZN(n4289) );
  INV_X1 U4147 ( .A(n3526), .ZN(n3524) );
  AOI22_X1 U4148 ( .A1(n3476), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3481) );
  OR2_X1 U4149 ( .A1(n3650), .A2(n3649), .ZN(n4273) );
  AND4_X1 U4150 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3442)
         );
  AND4_X1 U4151 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  AND2_X1 U4152 ( .A1(n4199), .A2(n5440), .ZN(n4200) );
  AND2_X1 U4153 ( .A1(n4167), .A2(n4166), .ZN(n4421) );
  NOR2_X1 U4154 ( .A1(n3255), .A2(n3727), .ZN(n3728) );
  INV_X1 U4155 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3951) );
  INV_X1 U4156 ( .A(n5442), .ZN(n4197) );
  NAND2_X1 U4157 ( .A1(n3626), .A2(n3625), .ZN(n5075) );
  NAND2_X1 U4158 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  AND2_X1 U4159 ( .A1(n4662), .A2(n4663), .ZN(n4667) );
  INV_X1 U4160 ( .A(n4702), .ZN(n4692) );
  INV_X1 U4161 ( .A(n4343), .ZN(n5284) );
  INV_X1 U4162 ( .A(n4401), .ZN(n4402) );
  AND2_X1 U4163 ( .A1(n6278), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5557) );
  AND2_X1 U4164 ( .A1(n4651), .A2(n5573), .ZN(n4147) );
  OR2_X1 U4165 ( .A1(n4800), .A2(n4837), .ZN(n4801) );
  INV_X1 U4166 ( .A(n3970), .ZN(n5422) );
  INV_X1 U4167 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4711) );
  AND2_X1 U4168 ( .A1(n5686), .A2(n4348), .ZN(n5684) );
  AND2_X1 U4169 ( .A1(n4220), .A2(n4219), .ZN(n5339) );
  AND2_X1 U4170 ( .A1(n5905), .A2(n5904), .ZN(n6098) );
  OR2_X1 U4171 ( .A1(n5888), .A2(n5256), .ZN(n6425) );
  OR2_X1 U4172 ( .A1(n4343), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6443) );
  NOR2_X1 U4173 ( .A1(n4894), .A2(n6225), .ZN(n6116) );
  OR2_X1 U4174 ( .A1(n4927), .A2(n5163), .ZN(n5197) );
  AND2_X1 U4175 ( .A1(n3623), .A2(n6710), .ZN(n6578) );
  NOR2_X1 U4176 ( .A1(n6117), .A2(n3102), .ZN(n4634) );
  AND3_X1 U4177 ( .A1(n5129), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6546) );
  OR2_X1 U4178 ( .A1(n4624), .A2(n4623), .ZN(n6117) );
  AND2_X1 U4179 ( .A1(n6631), .A2(n6682), .ZN(n6633) );
  INV_X1 U4180 ( .A(n4667), .ZN(n4666) );
  NAND2_X1 U4181 ( .A1(n4667), .A2(n5164), .ZN(n5027) );
  NOR2_X1 U4182 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4630), .ZN(n5023) );
  NAND2_X1 U4183 ( .A1(n4578), .A2(n3554), .ZN(n4874) );
  INV_X1 U4184 ( .A(n4435), .ZN(n5281) );
  NAND2_X1 U4185 ( .A1(n4403), .A2(n4402), .ZN(n4404) );
  AND2_X1 U4186 ( .A1(n6278), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6330) );
  INV_X1 U4187 ( .A(n5628), .ZN(n5607) );
  OR2_X1 U4188 ( .A1(n5662), .A2(n5661), .ZN(n5681) );
  INV_X1 U4189 ( .A(n6343), .ZN(n6353) );
  INV_X1 U4190 ( .A(n6383), .ZN(n6374) );
  INV_X1 U4191 ( .A(n4802), .ZN(n6395) );
  INV_X1 U4192 ( .A(n6418), .ZN(n5870) );
  OR2_X1 U4193 ( .A1(n4876), .A2(n5114), .ZN(n4595) );
  INV_X1 U4194 ( .A(n6226), .ZN(n6414) );
  OR2_X1 U4195 ( .A1(n5955), .A2(n5915), .ZN(n5940) );
  OR2_X1 U4196 ( .A1(n5996), .A2(n5913), .ZN(n5976) );
  AND2_X1 U4197 ( .A1(n4196), .A2(n4195), .ZN(n5442) );
  NAND2_X1 U4198 ( .A1(n5892), .A2(n6068), .ZN(n6105) );
  INV_X1 U4199 ( .A(n6422), .ZN(n6456) );
  INV_X1 U4200 ( .A(n6443), .ZN(n6399) );
  NOR2_X1 U4201 ( .A1(n4880), .A2(n3502), .ZN(n5261) );
  INV_X1 U4202 ( .A(n5163), .ZN(n5164) );
  OAI211_X1 U4203 ( .C1(n6626), .C2(n4933), .A(n4932), .B(n6543), .ZN(n4957)
         );
  OAI21_X1 U4204 ( .B1(n4895), .B2(n6636), .A(n6121), .ZN(n4931) );
  OAI211_X1 U4205 ( .C1(n5126), .C2(n5198), .A(n5125), .B(n6590), .ZN(n5204)
         );
  OAI21_X1 U4206 ( .B1(n5009), .B2(n5008), .A(n5007), .ZN(n6479) );
  OAI21_X1 U4207 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(n6514) );
  INV_X1 U4208 ( .A(n4962), .ZN(n4991) );
  AND2_X1 U4209 ( .A1(n4634), .A2(n5164), .ZN(n6534) );
  INV_X1 U4210 ( .A(n6643), .ZN(n6595) );
  NOR2_X1 U4211 ( .A1(n5165), .A2(n5164), .ZN(n6617) );
  OAI21_X1 U4212 ( .B1(n5172), .B2(n5171), .A(n5170), .ZN(n5214) );
  OAI21_X1 U4213 ( .B1(n6148), .B2(n6630), .A(n6147), .ZN(n6183) );
  OAI21_X1 U4214 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6686) );
  INV_X1 U4215 ( .A(n6683), .ZN(n6700) );
  AND2_X1 U4216 ( .A1(n5001), .A2(n6626), .ZN(n4670) );
  INV_X1 U4217 ( .A(n5027), .ZN(n5062) );
  NOR2_X1 U4218 ( .A1(n4647), .A2(n6192), .ZN(n6712) );
  INV_X1 U4219 ( .A(n6664), .ZN(n6718) );
  AND2_X1 U4220 ( .A1(n5263), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4129) );
  OR2_X1 U4221 ( .A1(n4595), .A2(n4874), .ZN(n4497) );
  INV_X1 U4222 ( .A(n5819), .ZN(n5667) );
  INV_X1 U4223 ( .A(n5842), .ZN(n5672) );
  INV_X1 U4224 ( .A(n5681), .ZN(n5072) );
  INV_X2 U4225 ( .A(n6362), .ZN(n6380) );
  NAND2_X1 U4226 ( .A1(n6381), .A2(n3554), .ZN(n6343) );
  OR2_X1 U4227 ( .A1(n6381), .A2(n6374), .ZN(n6362) );
  INV_X1 U4228 ( .A(n6381), .ZN(n6378) );
  INV_X1 U4229 ( .A(n6376), .ZN(n6383) );
  OR2_X1 U4230 ( .A1(n4595), .A2(n4851), .ZN(n6398) );
  NAND2_X1 U4231 ( .A1(n4437), .A2(n6626), .ZN(n5873) );
  NAND2_X1 U4232 ( .A1(n5868), .A2(n5884), .ZN(n6418) );
  INV_X1 U4233 ( .A(n6432), .ZN(n6455) );
  NAND2_X1 U4234 ( .A1(n4589), .A2(n4577), .ZN(n6422) );
  INV_X1 U4235 ( .A(n6465), .ZN(n4754) );
  INV_X1 U4236 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6466) );
  OR2_X1 U4237 ( .A1(n4927), .A2(n5164), .ZN(n6137) );
  AOI22_X1 U4238 ( .A1(n4931), .A2(n4926), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4933), .ZN(n4960) );
  NAND3_X1 U4239 ( .A1(n4893), .A2(n5010), .A3(n6539), .ZN(n6517) );
  INV_X1 U4240 ( .A(n4961), .ZN(n4994) );
  NAND2_X1 U4241 ( .A1(n6540), .A2(n5073), .ZN(n6576) );
  NAND2_X1 U4242 ( .A1(n6540), .A2(n6539), .ZN(n6621) );
  AOI22_X1 U4243 ( .A1(n5168), .A2(n5171), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6583), .ZN(n5217) );
  AOI21_X1 U4244 ( .B1(n6146), .B2(n6630), .A(n6145), .ZN(n6186) );
  OR2_X1 U4245 ( .A1(n6628), .A2(n6138), .ZN(n6690) );
  OR2_X1 U4246 ( .A1(n6628), .A2(n6187), .ZN(n6708) );
  INV_X1 U4247 ( .A(n6673), .ZN(n6219) );
  INV_X1 U4248 ( .A(n6694), .ZN(n5192) );
  NOR2_X1 U4249 ( .A1(n5026), .A2(n5025), .ZN(n5065) );
  NAND2_X1 U4250 ( .A1(n4766), .A2(n4662), .ZN(n6713) );
  INV_X1 U4251 ( .A(n6741), .ZN(n6737) );
  OAI21_X1 U4252 ( .B1(n5631), .B2(n5554), .A(n4406), .ZN(U2797) );
  INV_X1 U4253 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3263) );
  AND2_X2 U4254 ( .A1(n3263), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3270)
         );
  AND2_X4 U4255 ( .A1(n3270), .A2(n4717), .ZN(n3541) );
  INV_X1 U4256 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4257 ( .A1(n3541), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3269) );
  INV_X1 U4258 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4259 ( .A1(n3840), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3268) );
  NOR2_X4 U4260 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U4261 ( .A1(n3971), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3267) );
  BUF_X2 U4262 ( .A(n3536), .Z(n3997) );
  AOI22_X1 U4263 ( .A1(n3998), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3266) );
  NAND4_X1 U4264 ( .A1(n3269), .A2(n3268), .A3(n3267), .A4(n3266), .ZN(n3278)
         );
  AOI22_X1 U4265 ( .A1(n3353), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3431), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4266 ( .A1(n3956), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3275) );
  AND2_X2 U4267 ( .A1(n3270), .A2(n3271), .ZN(n3476) );
  AOI22_X1 U4268 ( .A1(n3476), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3274) );
  AND2_X4 U4269 ( .A1(n3272), .A2(n3271), .ZN(n3529) );
  AOI22_X1 U4270 ( .A1(n3529), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3273) );
  NAND4_X1 U4271 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3277)
         );
  NOR2_X1 U4272 ( .A1(n3278), .A2(n3277), .ZN(n3361) );
  AOI22_X1 U4273 ( .A1(n3818), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4274 ( .A1(n3905), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3281) );
  INV_X2 U4275 ( .A(n4725), .ZN(n3976) );
  AOI22_X1 U4276 ( .A1(n3353), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4277 ( .A1(n3990), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3279) );
  NAND4_X1 U4278 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3288)
         );
  AOI22_X1 U4279 ( .A1(n3956), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3541), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4280 ( .A1(n3544), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3285) );
  INV_X2 U4281 ( .A(n4720), .ZN(n3992) );
  AOI22_X1 U4282 ( .A1(n3992), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4283 ( .A1(n3431), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4284 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3287)
         );
  NOR2_X1 U4285 ( .A1(n3288), .A2(n3287), .ZN(n4060) );
  AOI22_X1 U4286 ( .A1(n3956), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4287 ( .A1(n3544), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4288 ( .A1(n3353), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4289 ( .A1(n3971), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3289) );
  NAND4_X1 U4290 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3298)
         );
  AOI22_X1 U4291 ( .A1(n3818), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4292 ( .A1(n3905), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3541), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4293 ( .A1(n3431), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4294 ( .A1(n3992), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3293) );
  NAND4_X1 U4295 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3297)
         );
  NOR2_X1 U4296 ( .A1(n3298), .A2(n3297), .ZN(n4043) );
  AOI22_X1 U4297 ( .A1(n3956), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4298 ( .A1(n3977), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4299 ( .A1(n3544), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4300 ( .A1(n3353), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3299) );
  NAND4_X1 U4301 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3308)
         );
  AOI22_X1 U4302 ( .A1(n3818), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4303 ( .A1(n3541), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4304 ( .A1(n3989), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4305 ( .A1(n3992), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3303) );
  NAND4_X1 U4306 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3307)
         );
  NOR2_X1 U4307 ( .A1(n3308), .A2(n3307), .ZN(n4027) );
  AOI22_X1 U4308 ( .A1(n3956), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4309 ( .A1(n3905), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4310 ( .A1(n3992), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4311 ( .A1(n3353), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3309) );
  NAND4_X1 U4312 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3318)
         );
  AOI22_X1 U4313 ( .A1(n3476), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4314 ( .A1(n3530), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4315 ( .A1(n3431), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4316 ( .A1(n3544), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3313) );
  NAND4_X1 U4317 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  NOR2_X1 U4318 ( .A1(n3318), .A2(n3317), .ZN(n4013) );
  AOI22_X1 U4319 ( .A1(n3818), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4320 ( .A1(n3998), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4321 ( .A1(n3353), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4322 ( .A1(n3544), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3319) );
  NAND4_X1 U4323 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3328)
         );
  AOI22_X1 U4324 ( .A1(n3956), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4325 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3530), .B1(n3372), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4326 ( .A1(n3977), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4327 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3992), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4328 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3327)
         );
  NOR2_X1 U4329 ( .A1(n3328), .A2(n3327), .ZN(n4012) );
  OR2_X1 U4330 ( .A1(n4013), .A2(n4012), .ZN(n4021) );
  AOI22_X1 U4331 ( .A1(n3989), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3332) );
  INV_X1 U4332 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U4333 ( .A1(n3818), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4334 ( .A1(n3431), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4335 ( .A1(n3991), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4336 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3338)
         );
  AOI22_X1 U4337 ( .A1(n3905), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4338 ( .A1(n3353), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4339 ( .A1(n3956), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4340 ( .A1(n3971), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4341 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3337)
         );
  NOR2_X1 U4342 ( .A1(n3338), .A2(n3337), .ZN(n4020) );
  NOR2_X1 U4343 ( .A1(n4027), .A2(n4026), .ZN(n4034) );
  AOI22_X1 U4344 ( .A1(n3818), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4345 ( .A1(n3541), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4346 ( .A1(n3989), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3340) );
  INV_X1 U4347 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n7043) );
  AOI22_X1 U4348 ( .A1(n3992), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3339) );
  NAND4_X1 U4349 ( .A1(n3342), .A2(n3341), .A3(n3340), .A4(n3339), .ZN(n3348)
         );
  AOI22_X1 U4350 ( .A1(n3956), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4351 ( .A1(n3431), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4352 ( .A1(n3544), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4353 ( .A1(n3353), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3343) );
  NAND4_X1 U4354 ( .A1(n3346), .A2(n3345), .A3(n3344), .A4(n3343), .ZN(n3347)
         );
  NAND2_X1 U4355 ( .A1(n4034), .A2(n4033), .ZN(n4044) );
  NOR2_X1 U4356 ( .A1(n4043), .A2(n4044), .ZN(n4051) );
  AOI22_X1 U4357 ( .A1(n3818), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4358 ( .A1(n3541), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4359 ( .A1(n3989), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4360 ( .A1(n3992), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3349) );
  NAND4_X1 U4361 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3359)
         );
  AOI22_X1 U4362 ( .A1(n3956), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3357) );
  INV_X1 U4363 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U4364 ( .A1(n3431), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4365 ( .A1(n3544), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4366 ( .A1(n3353), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3354) );
  NAND4_X1 U4367 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3358)
         );
  OR2_X1 U4368 ( .A1(n3359), .A2(n3358), .ZN(n4050) );
  NAND2_X1 U4369 ( .A1(n4051), .A2(n4050), .ZN(n4061) );
  NOR2_X1 U4370 ( .A1(n4060), .A2(n4061), .ZN(n3360) );
  XOR2_X1 U4371 ( .A(n3361), .B(n3360), .Z(n3416) );
  AOI22_X1 U4372 ( .A1(n3541), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4373 ( .A1(n3840), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3564), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4374 ( .A1(n3531), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4375 ( .A1(n3431), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4376 ( .A1(n3543), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4377 ( .A1(n3482), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3366) );
  NAND2_X2 U4378 ( .A1(n3371), .A2(n3370), .ZN(n3493) );
  AOI22_X1 U4379 ( .A1(n3372), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3541), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4380 ( .A1(n3543), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4381 ( .A1(n3840), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3564), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4382 ( .A1(n3431), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3373) );
  NAND4_X1 U4383 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3383)
         );
  AOI22_X1 U4384 ( .A1(n3482), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4385 ( .A1(n3531), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4386 ( .A1(n3377), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3477), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3378) );
  NAND4_X1 U4387 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3382)
         );
  NAND2_X1 U4388 ( .A1(n3698), .A2(n3497), .ZN(n3496) );
  NAND2_X1 U4389 ( .A1(n3372), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4390 ( .A1(n3840), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4391 ( .A1(n3531), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3385)
         );
  NAND2_X1 U4392 ( .A1(n3462), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4393 ( .A1(n3482), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4394 ( .A1(n3477), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4395 ( .A1(n3483), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3391)
         );
  NAND2_X1 U4396 ( .A1(n3377), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4397 ( .A1(n3431), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4398 ( .A1(n3543), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4399 ( .A1(n3565), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3394)
         );
  NAND2_X1 U4400 ( .A1(n3536), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4401 ( .A1(n3476), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3400) );
  NAND2_X1 U4402 ( .A1(n3541), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3399)
         );
  NAND2_X1 U4403 ( .A1(n3529), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3398)
         );
  NAND2_X1 U4404 ( .A1(n3564), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4405 ( .A1(n3482), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3543), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4406 ( .A1(n3372), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4407 ( .A1(n3840), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3564), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4408 ( .A1(n3431), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3477), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4409 ( .A1(n3377), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4410 ( .A1(n3565), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4411 ( .A1(n3541), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4412 ( .A1(n3476), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4413 ( .A1(n4579), .A2(n4693), .ZN(n3514) );
  AOI22_X1 U4414 ( .A1(n4353), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6632), .ZN(n3415) );
  OAI21_X1 U4415 ( .B1(n3416), .B2(n4036), .A(n3415), .ZN(n3417) );
  INV_X1 U4416 ( .A(n3417), .ZN(n3422) );
  INV_X1 U4417 ( .A(n4031), .ZN(n3421) );
  INV_X1 U4418 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4344) );
  XNOR2_X1 U4419 ( .A(n4356), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5690)
         );
  MUX2_X1 U4420 ( .A(n3422), .B(n5690), .S(n3101), .Z(n4070) );
  NAND2_X1 U4421 ( .A1(n3543), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4422 ( .A1(n3476), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4423 ( .A1(n3840), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4424 ( .A1(n3564), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4425 ( .A1(n3372), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4426 ( .A1(n3529), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3429)
         );
  NAND2_X1 U4427 ( .A1(n3531), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3428)
         );
  NAND2_X1 U4428 ( .A1(n3462), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U4429 ( .A1(n3377), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4430 ( .A1(n3431), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3434) );
  NAND2_X1 U4431 ( .A1(n3477), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3433)
         );
  NAND2_X1 U4432 ( .A1(n3483), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3432)
         );
  NAND2_X1 U4433 ( .A1(n3482), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4434 ( .A1(n3541), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3438)
         );
  NAND2_X1 U4435 ( .A1(n3565), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3437)
         );
  NAND2_X1 U4436 ( .A1(n3536), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4437 ( .A1(n3476), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4438 ( .A1(n3541), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4439 ( .A1(n3840), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3564), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4440 ( .A1(n3531), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3443) );
  NAND4_X1 U4441 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n3452)
         );
  AOI22_X1 U4442 ( .A1(n3482), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4443 ( .A1(n3431), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4444 ( .A1(n3543), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4445 ( .A1(n3377), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3477), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4446 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3451)
         );
  NAND2_X1 U4447 ( .A1(n4703), .A2(n4668), .ZN(n4524) );
  NAND2_X1 U4448 ( .A1(n3840), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3457) );
  NAND2_X1 U4449 ( .A1(n3476), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4450 ( .A1(n3372), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4451 ( .A1(n3564), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3454) );
  NAND2_X1 U4452 ( .A1(n3377), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U4453 ( .A1(n3431), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U4454 ( .A1(n3477), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3459)
         );
  NAND2_X1 U4455 ( .A1(n3541), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3466)
         );
  NAND2_X1 U4456 ( .A1(n3529), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3465)
         );
  NAND2_X1 U4457 ( .A1(n3531), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3464)
         );
  NAND2_X1 U4458 ( .A1(n3462), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3463) );
  NAND2_X1 U4459 ( .A1(n3482), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U4460 ( .A1(n3543), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4461 ( .A1(n3565), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3468)
         );
  NAND2_X1 U4462 ( .A1(n3536), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3467) );
  AND4_X2 U4463 ( .A1(n3470), .A2(n3469), .A3(n3468), .A4(n3467), .ZN(n3471)
         );
  AND4_X4 U4464 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n4633)
         );
  AND2_X1 U4465 ( .A1(n3512), .A2(n3554), .ZN(n3475) );
  NAND2_X1 U4466 ( .A1(n3492), .A2(n3475), .ZN(n4506) );
  AOI22_X1 U4467 ( .A1(n3564), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4468 ( .A1(n3541), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4469 ( .A1(n3377), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3477), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4470 ( .A1(n3482), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4471 ( .A1(n3431), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3483), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4472 ( .A1(n3543), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4473 ( .A1(n3529), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3484) );
  NAND2_X2 U4474 ( .A1(n3489), .A2(n3488), .ZN(n4134) );
  NAND2_X1 U4475 ( .A1(n4633), .A2(n4684), .ZN(n5555) );
  NAND2_X1 U4476 ( .A1(n5555), .A2(n4688), .ZN(n3490) );
  NAND2_X1 U4477 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4442) );
  OAI21_X1 U4478 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n4442), .ZN(n4373) );
  NAND2_X1 U4479 ( .A1(n3502), .A2(n4373), .ZN(n3576) );
  NAND2_X1 U4480 ( .A1(n3490), .A2(n3576), .ZN(n3491) );
  NAND3_X1 U4481 ( .A1(n4238), .A2(n4506), .A3(n3491), .ZN(n3505) );
  INV_X1 U4482 ( .A(n3492), .ZN(n3578) );
  OAI21_X1 U4483 ( .B1(n4075), .B2(n3494), .A(n3519), .ZN(n3501) );
  OAI21_X1 U4484 ( .B1(n3494), .B2(n3493), .A(n4693), .ZN(n3495) );
  INV_X1 U4485 ( .A(n3495), .ZN(n3500) );
  NAND2_X1 U4486 ( .A1(n3496), .A2(n4668), .ZN(n3499) );
  NAND3_X1 U4487 ( .A1(n4703), .A2(n3497), .A3(n3493), .ZN(n3498) );
  NAND4_X1 U4488 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3579)
         );
  NAND2_X1 U4489 ( .A1(n3579), .A2(n6753), .ZN(n4532) );
  INV_X1 U4490 ( .A(n4239), .ZN(n3503) );
  NAND2_X1 U4491 ( .A1(n3503), .A2(n5439), .ZN(n3504) );
  OAI211_X1 U4492 ( .C1(n3578), .C2(n4391), .A(n4532), .B(n3504), .ZN(n3518)
         );
  OAI21_X1 U4493 ( .B1(n3505), .B2(n3518), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3586) );
  OR2_X1 U4494 ( .A1(n3586), .A2(n5262), .ZN(n3507) );
  NAND2_X1 U4495 ( .A1(n6123), .A2(n5282), .ZN(n4343) );
  MUX2_X1 U4496 ( .A(n4129), .B(n4343), .S(n6582), .Z(n3506) );
  NAND2_X1 U4497 ( .A1(n3507), .A2(n3506), .ZN(n3527) );
  INV_X1 U4498 ( .A(n3527), .ZN(n3525) );
  INV_X1 U4499 ( .A(n3508), .ZN(n3510) );
  AOI21_X1 U4500 ( .B1(n3512), .B2(n4579), .A(n4130), .ZN(n3509) );
  NAND2_X1 U4501 ( .A1(n3510), .A2(n3509), .ZN(n3511) );
  NAND2_X1 U4502 ( .A1(n3511), .A2(n4684), .ZN(n3517) );
  INV_X1 U4503 ( .A(n3512), .ZN(n3513) );
  NAND2_X1 U4504 ( .A1(n3513), .A2(n5280), .ZN(n4505) );
  INV_X1 U4505 ( .A(n3514), .ZN(n3516) );
  NOR2_X1 U4506 ( .A1(n4680), .A2(n4668), .ZN(n3515) );
  NAND3_X1 U4507 ( .A1(n3516), .A2(n3515), .A3(n4703), .ZN(n4726) );
  AND2_X1 U4508 ( .A1(n6123), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6730) );
  INV_X1 U4509 ( .A(n3518), .ZN(n3522) );
  MUX2_X1 U4510 ( .A(n4239), .B(n3519), .S(n3554), .Z(n3521) );
  NAND2_X1 U4511 ( .A1(n3521), .A2(n4871), .ZN(n4529) );
  NAND3_X1 U4512 ( .A1(n3523), .A2(n3522), .A3(n4529), .ZN(n3526) );
  NAND2_X1 U4513 ( .A1(n3525), .A2(n3524), .ZN(n3528) );
  AOI22_X1 U4514 ( .A1(n3476), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4515 ( .A1(n3530), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4516 ( .A1(n3840), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3564), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3533) );
  INV_X1 U4517 ( .A(n3531), .ZN(n4720) );
  AOI22_X1 U4518 ( .A1(n3992), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4519 ( .A1(n3956), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3565), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4520 ( .A1(n3977), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4521 ( .A1(n3544), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4522 ( .A1(n3353), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3977), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4523 ( .A1(n3956), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4524 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3530), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4525 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3544), .B1(n3565), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4526 ( .A1(n3476), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4527 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3564), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4528 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3992), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4529 ( .A1(n3971), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3549) );
  INV_X1 U4530 ( .A(n3695), .ZN(n3553) );
  INV_X1 U4531 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3557) );
  AOI21_X1 U4532 ( .B1(n4697), .B2(n4308), .A(n5282), .ZN(n3556) );
  NAND2_X1 U4533 ( .A1(n4633), .A2(n4253), .ZN(n3555) );
  INV_X1 U4534 ( .A(n3559), .ZN(n3575) );
  NAND2_X1 U4535 ( .A1(n4078), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3574) );
  INV_X1 U4536 ( .A(n3627), .ZN(n3572) );
  AOI22_X1 U4537 ( .A1(n3353), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3977), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4538 ( .A1(n3956), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4539 ( .A1(n3476), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4540 ( .A1(n3530), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4541 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3571)
         );
  AOI22_X1 U4542 ( .A1(n3840), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4543 ( .A1(n3905), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4544 ( .A1(n3998), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4545 ( .A1(n3971), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3566) );
  NAND4_X1 U4546 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(n3570)
         );
  NAND2_X1 U4547 ( .A1(n3572), .A2(n4245), .ZN(n3573) );
  XNOR2_X1 U4548 ( .A(n6582), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6197)
         );
  INV_X1 U4549 ( .A(n4129), .ZN(n3624) );
  AOI22_X1 U4550 ( .A1(n5284), .A2(n6197), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3624), .ZN(n3588) );
  INV_X1 U4551 ( .A(n3588), .ZN(n3585) );
  INV_X1 U4552 ( .A(n3576), .ZN(n3582) );
  NOR2_X1 U4553 ( .A1(n4524), .A2(n4688), .ZN(n3577) );
  NOR2_X1 U4554 ( .A1(n4688), .A2(n4668), .ZN(n3581) );
  NAND3_X1 U4555 ( .A1(n6753), .A2(n4703), .A3(n3581), .ZN(n4533) );
  NAND2_X1 U4556 ( .A1(n4680), .A2(n4693), .ZN(n4617) );
  OAI211_X1 U4557 ( .C1(n3582), .C2(n4874), .A(n4736), .B(n4580), .ZN(n3583)
         );
  NAND2_X1 U4558 ( .A1(n3583), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3587) );
  INV_X1 U4559 ( .A(n3587), .ZN(n3584) );
  OAI21_X1 U4560 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3585), .A(n3584), 
        .ZN(n3589) );
  INV_X1 U4561 ( .A(n3586), .ZN(n3622) );
  INV_X1 U4562 ( .A(n4245), .ZN(n3591) );
  NOR2_X1 U4563 ( .A1(n3628), .A2(n3591), .ZN(n3592) );
  INV_X1 U4564 ( .A(n3593), .ZN(n3594) );
  NOR2_X1 U4565 ( .A1(n3595), .A2(n3594), .ZN(n3596) );
  AOI21_X2 U4566 ( .B1(n3686), .B2(n3687), .A(n3596), .ZN(n3683) );
  AND2_X1 U4567 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U4568 ( .A1(n3599), .A2(n6143), .ZN(n5004) );
  INV_X1 U4569 ( .A(n3599), .ZN(n3600) );
  NAND2_X1 U4570 ( .A1(n3600), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4571 ( .A1(n5004), .A2(n3601), .ZN(n4902) );
  AOI22_X1 U4572 ( .A1(n5284), .A2(n4902), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3624), .ZN(n3602) );
  XNOR2_X1 U4573 ( .A(n3619), .B(n3620), .ZN(n4543) );
  NAND2_X1 U4574 ( .A1(n4543), .A2(n5282), .ZN(n3618) );
  AOI22_X1 U4575 ( .A1(n3818), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4576 ( .A1(n3530), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4577 ( .A1(n3840), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4578 ( .A1(n3992), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3604) );
  NAND4_X1 U4579 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3613)
         );
  AOI22_X1 U4580 ( .A1(n3956), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4581 ( .A1(n3977), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4582 ( .A1(n3544), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4583 ( .A1(n3353), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4584 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3612)
         );
  INV_X1 U4585 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3614) );
  OAI22_X1 U4586 ( .A1(n4240), .A2(n3627), .B1(n4109), .B2(n3614), .ZN(n3616)
         );
  NOR2_X1 U4587 ( .A1(n3628), .A2(n4240), .ZN(n3615) );
  XNOR2_X1 U4588 ( .A(n3616), .B(n3615), .ZN(n3617) );
  NAND2_X1 U4589 ( .A1(n3622), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4590 ( .A1(n6546), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U4591 ( .A1(n6570), .A2(n5129), .ZN(n3623) );
  NAND3_X1 U4592 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5022) );
  INV_X1 U4593 ( .A(n5022), .ZN(n4772) );
  NAND2_X1 U4594 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4772), .ZN(n6710) );
  AOI22_X1 U4595 ( .A1(n6578), .A2(n5284), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3624), .ZN(n3625) );
  AOI22_X1 U4596 ( .A1(n3818), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4597 ( .A1(n3530), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4598 ( .A1(n3840), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4599 ( .A1(n3992), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4600 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3638)
         );
  AOI22_X1 U4601 ( .A1(n3956), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4602 ( .A1(n3977), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4603 ( .A1(n3544), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4604 ( .A1(n3353), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3633) );
  NAND4_X1 U4605 ( .A1(n3636), .A2(n3635), .A3(n3634), .A4(n3633), .ZN(n3637)
         );
  AOI22_X1 U4606 ( .A1(n4123), .A2(n4269), .B1(n4078), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3639) );
  NAND2_X2 U4607 ( .A1(n3640), .A2(n3639), .ZN(n4770) );
  AOI22_X1 U4608 ( .A1(n3818), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4609 ( .A1(n3530), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4610 ( .A1(n3840), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4611 ( .A1(n3992), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4612 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3650)
         );
  AOI22_X1 U4613 ( .A1(n3956), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4614 ( .A1(n3977), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4615 ( .A1(n3544), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4616 ( .A1(n3353), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3645) );
  NAND4_X1 U4617 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(n3649)
         );
  AOI22_X1 U4618 ( .A1(n4123), .A2(n4273), .B1(n4078), .B2(
        INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4619 ( .A1(n3818), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4620 ( .A1(n3530), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4621 ( .A1(n3840), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4622 ( .A1(n3992), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3652) );
  NAND4_X1 U4623 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3661)
         );
  AOI22_X1 U4624 ( .A1(n3956), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4625 ( .A1(n3977), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4626 ( .A1(n3544), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4627 ( .A1(n3353), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4628 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3660)
         );
  AOI22_X1 U4629 ( .A1(n4123), .A2(n4289), .B1(n4078), .B2(
        INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4630 ( .A1(n3353), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3977), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4631 ( .A1(n3956), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4632 ( .A1(n3818), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4633 ( .A1(n3905), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4634 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4635 ( .A1(n3530), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4636 ( .A1(n3992), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4637 ( .A1(n3998), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4638 ( .A1(n3971), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4639 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NAND2_X1 U4640 ( .A1(n4123), .A2(n4292), .ZN(n3673) );
  NAND2_X1 U4641 ( .A1(n4078), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3672) );
  NAND2_X1 U4642 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  INV_X1 U4643 ( .A(n4288), .ZN(n3675) );
  INV_X2 U4644 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U4645 ( .A1(n3675), .A2(n3878), .ZN(n3682) );
  INV_X1 U4646 ( .A(n3746), .ZN(n3678) );
  INV_X1 U4647 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4648 ( .A1(n3131), .A2(n3676), .ZN(n3677) );
  NAND2_X1 U4649 ( .A1(n3678), .A2(n3677), .ZN(n6302) );
  INV_X1 U4650 ( .A(n6302), .ZN(n3680) );
  AOI22_X1 U4651 ( .A1(n4353), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6632), .ZN(n3679) );
  MUX2_X1 U4652 ( .A(n3680), .B(n3679), .S(n4019), .Z(n3681) );
  NAND2_X1 U4653 ( .A1(n4661), .A2(n3878), .ZN(n3685) );
  INV_X1 U4654 ( .A(n4352), .ZN(n3899) );
  NAND2_X1 U4655 ( .A1(n4625), .A2(n3878), .ZN(n3691) );
  AOI22_X1 U4656 ( .A1(n4353), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6632), .ZN(n3689) );
  INV_X1 U4657 ( .A(n4617), .ZN(n4415) );
  NAND2_X1 U4658 ( .A1(n4415), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3738) );
  INV_X1 U4659 ( .A(n3738), .ZN(n3702) );
  NAND2_X1 U4660 ( .A1(n3702), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3688) );
  AND2_X1 U4661 ( .A1(n3689), .A2(n3688), .ZN(n3690) );
  NAND2_X1 U4662 ( .A1(n3691), .A2(n3690), .ZN(n4608) );
  AND2_X1 U4663 ( .A1(n3698), .A2(n4693), .ZN(n3699) );
  AOI21_X1 U4664 ( .B1(n5163), .B2(n3699), .A(n6632), .ZN(n4607) );
  INV_X1 U4665 ( .A(n3114), .ZN(n6629) );
  AOI22_X1 U4666 ( .A1(n4353), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6632), .ZN(n3701) );
  NAND2_X1 U4667 ( .A1(n3702), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3700) );
  OAI211_X1 U4668 ( .C1(n6629), .C2(n3904), .A(n3701), .B(n3700), .ZN(n4606)
         );
  MUX2_X1 U4669 ( .A(n3101), .B(n4607), .S(n4606), .Z(n4609) );
  NAND2_X1 U4670 ( .A1(n3708), .A2(n3709), .ZN(n3707) );
  NAND2_X1 U4671 ( .A1(n3702), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3706) );
  INV_X1 U4672 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5572) );
  OAI21_X1 U4673 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3732), .ZN(n6408) );
  NAND2_X1 U4674 ( .A1(n3101), .A2(n6408), .ZN(n3703) );
  OAI21_X1 U4675 ( .B1(n5572), .B2(n3899), .A(n3703), .ZN(n3704) );
  AOI21_X1 U4676 ( .B1(n4353), .B2(EAX_REG_2__SCAN_IN), .A(n3704), .ZN(n3705)
         );
  AND2_X1 U4677 ( .A1(n3706), .A2(n3705), .ZN(n4613) );
  NAND2_X1 U4678 ( .A1(n3707), .A2(n4613), .ZN(n3711) );
  INV_X1 U4679 ( .A(n3708), .ZN(n4615) );
  INV_X1 U4680 ( .A(n3709), .ZN(n4614) );
  NAND2_X1 U4681 ( .A1(n4615), .A2(n4614), .ZN(n3710) );
  NAND2_X1 U4682 ( .A1(n4268), .A2(n3878), .ZN(n3718) );
  NAND2_X1 U4683 ( .A1(n6632), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3714)
         );
  NAND2_X1 U4684 ( .A1(n4353), .A2(EAX_REG_4__SCAN_IN), .ZN(n3713) );
  OAI211_X1 U4685 ( .C1(n3738), .C2(n4113), .A(n3714), .B(n3713), .ZN(n3715)
         );
  XNOR2_X1 U4686 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .B(n3733), .ZN(n6325) );
  MUX2_X1 U4687 ( .A(n3715), .B(n6325), .S(n3101), .Z(n3716) );
  INV_X1 U4688 ( .A(n3716), .ZN(n3717) );
  NAND2_X1 U4689 ( .A1(n3718), .A2(n3717), .ZN(n4755) );
  INV_X1 U4690 ( .A(n3722), .ZN(n3724) );
  INV_X1 U4691 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3723) );
  NAND2_X1 U4692 ( .A1(n3724), .A2(n3723), .ZN(n3725) );
  NAND2_X1 U4693 ( .A1(n3131), .A2(n3725), .ZN(n6316) );
  AOI22_X1 U4694 ( .A1(n6316), .A2(n3101), .B1(n4352), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3726) );
  INV_X1 U4695 ( .A(n3726), .ZN(n3727) );
  INV_X1 U4696 ( .A(n4770), .ZN(n4765) );
  NAND2_X2 U4697 ( .A1(n3731), .A2(n4624), .ZN(n4893) );
  INV_X1 U4698 ( .A(n3732), .ZN(n3735) );
  INV_X1 U4699 ( .A(n3733), .ZN(n3734) );
  OAI21_X1 U4700 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3735), .A(n3734), 
        .ZN(n5559) );
  AOI22_X1 U4701 ( .A1(n3101), .A2(n5559), .B1(n4352), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4702 ( .A1(n4353), .A2(EAX_REG_3__SCAN_IN), .ZN(n3736) );
  OAI211_X1 U4703 ( .C1(n3738), .C2(n6128), .A(n3737), .B(n3736), .ZN(n3739)
         );
  INV_X1 U4704 ( .A(n3739), .ZN(n3740) );
  NAND2_X1 U4705 ( .A1(n3741), .A2(n3740), .ZN(n4643) );
  INV_X1 U4706 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4707 ( .A1(n4123), .A2(n4308), .ZN(n3743) );
  OAI21_X1 U4708 ( .B1(n3744), .B2(n4109), .A(n3743), .ZN(n3745) );
  INV_X1 U4709 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3748) );
  OAI21_X1 U4710 ( .B1(n3746), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3792), 
        .ZN(n6291) );
  AOI22_X1 U4711 ( .A1(n6291), .A2(n3101), .B1(n4352), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3747) );
  OAI21_X1 U4712 ( .B1(n4064), .B2(n3748), .A(n3747), .ZN(n3749) );
  XOR2_X1 U4713 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3751), .Z(n6271) );
  AOI22_X1 U4714 ( .A1(n3956), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4715 ( .A1(n3542), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4716 ( .A1(n3905), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4717 ( .A1(n3977), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4718 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3761)
         );
  AOI22_X1 U4719 ( .A1(n3818), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3840), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4720 ( .A1(n3544), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4721 ( .A1(n3530), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4722 ( .A1(n3353), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3756) );
  NAND4_X1 U4723 ( .A1(n3759), .A2(n3758), .A3(n3757), .A4(n3756), .ZN(n3760)
         );
  OAI21_X1 U4724 ( .B1(n3761), .B2(n3760), .A(n3878), .ZN(n3764) );
  NAND2_X1 U4725 ( .A1(n4353), .A2(EAX_REG_9__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4726 ( .A1(n4352), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3762)
         );
  OAI21_X1 U4727 ( .B1(n6271), .B2(n4019), .A(n3262), .ZN(n5621) );
  NAND2_X1 U4728 ( .A1(n3765), .A2(n6809), .ZN(n3767) );
  INV_X1 U4729 ( .A(n3807), .ZN(n3766) );
  NAND2_X1 U4730 ( .A1(n3767), .A2(n3766), .ZN(n5860) );
  NAND2_X1 U4731 ( .A1(n5860), .A2(n3101), .ZN(n3781) );
  AOI22_X1 U4732 ( .A1(n3353), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4733 ( .A1(n3840), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4734 ( .A1(n3956), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4735 ( .A1(n3542), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4736 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3777)
         );
  AOI22_X1 U4737 ( .A1(n3530), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4738 ( .A1(n3818), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4739 ( .A1(n3971), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4740 ( .A1(n3977), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4741 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3776)
         );
  OAI21_X1 U4742 ( .B1(n3777), .B2(n3776), .A(n3878), .ZN(n3780) );
  NAND2_X1 U4743 ( .A1(n4353), .A2(EAX_REG_10__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4744 ( .A1(n4352), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3778)
         );
  NAND2_X1 U4745 ( .A1(n3781), .A2(n3261), .ZN(n5539) );
  INV_X1 U4746 ( .A(EAX_REG_8__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4747 ( .A1(n3818), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4748 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3542), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4749 ( .A1(n3544), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4750 ( .A1(n3353), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4751 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AOI22_X1 U4752 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3989), .B1(n3905), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4753 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3530), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4754 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3956), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4755 ( .A1(n3977), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4756 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  OAI21_X1 U4757 ( .B1(n3791), .B2(n3790), .A(n3878), .ZN(n3795) );
  INV_X1 U4758 ( .A(n3792), .ZN(n3793) );
  XNOR2_X1 U4759 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3793), .ZN(n5877) );
  AOI22_X1 U4760 ( .A1(n3101), .A2(n5877), .B1(n4352), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4761 ( .C1(n4064), .C2(n3796), .A(n3795), .B(n3794), .ZN(n4427)
         );
  AOI22_X1 U4762 ( .A1(n3977), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4763 ( .A1(n3989), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4764 ( .A1(n3956), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4765 ( .A1(n3992), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4766 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3806)
         );
  AOI22_X1 U4767 ( .A1(n3818), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4768 ( .A1(n3530), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4769 ( .A1(n3353), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4770 ( .A1(n3971), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4771 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  NOR2_X1 U4772 ( .A1(n3806), .A2(n3805), .ZN(n3811) );
  XOR2_X1 U4773 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3807), .Z(n6261) );
  INV_X1 U4774 ( .A(n6261), .ZN(n3808) );
  AOI22_X1 U4775 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n4352), .B1(n3101), 
        .B2(n3808), .ZN(n3810) );
  NAND2_X1 U4776 ( .A1(n4353), .A2(EAX_REG_11__SCAN_IN), .ZN(n3809) );
  OAI211_X1 U4777 ( .C1(n3904), .C2(n3811), .A(n3810), .B(n3809), .ZN(n5673)
         );
  INV_X1 U4778 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3814) );
  INV_X1 U4779 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5839) );
  AOI21_X1 U4780 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5839), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3812) );
  INV_X1 U4781 ( .A(n3812), .ZN(n3813) );
  OAI21_X1 U4782 ( .B1(n4064), .B2(n3814), .A(n3813), .ZN(n3817) );
  XNOR2_X1 U4783 ( .A(n3815), .B(n5839), .ZN(n5841) );
  NAND2_X1 U4784 ( .A1(n5841), .A2(n3101), .ZN(n3816) );
  NAND2_X1 U4785 ( .A1(n3817), .A2(n3816), .ZN(n3830) );
  AOI22_X1 U4786 ( .A1(n3956), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3818), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4787 ( .A1(n3544), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4788 ( .A1(n3530), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4789 ( .A1(n3997), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4790 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4791 ( .A1(n3840), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4792 ( .A1(n3542), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4793 ( .A1(n3977), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4794 ( .A1(n3353), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4795 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  OAI21_X1 U4796 ( .B1(n3828), .B2(n3827), .A(n3878), .ZN(n3829) );
  NAND2_X1 U4797 ( .A1(n3830), .A2(n3829), .ZN(n5527) );
  NAND2_X1 U4798 ( .A1(n4353), .A2(EAX_REG_13__SCAN_IN), .ZN(n3836) );
  INV_X1 U4799 ( .A(n3831), .ZN(n3833) );
  INV_X1 U4800 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4801 ( .A1(n3833), .A2(n3832), .ZN(n3834) );
  NAND2_X1 U4802 ( .A1(n3896), .A2(n3834), .ZN(n6255) );
  AOI22_X1 U4803 ( .A1(n6255), .A2(n3101), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .B2(n4352), .ZN(n3835) );
  NAND2_X1 U4804 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  AOI22_X1 U4805 ( .A1(n3977), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4806 ( .A1(n3818), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4807 ( .A1(n3840), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4808 ( .A1(n3353), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4809 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3850)
         );
  AOI22_X1 U4810 ( .A1(n3956), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4811 ( .A1(n3905), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3541), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4812 ( .A1(n3971), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4813 ( .A1(n3992), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4814 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3849)
         );
  OR2_X1 U4815 ( .A1(n3850), .A2(n3849), .ZN(n3851) );
  AND2_X1 U4816 ( .A1(n3878), .A2(n3851), .ZN(n5614) );
  AOI22_X1 U4817 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3956), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4818 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3905), .B1(n3530), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3818), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4820 ( .A1(n3977), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4821 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4822 ( .A1(n3989), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4823 ( .A1(n3544), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3992), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4825 ( .A1(n3353), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4826 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  OR2_X1 U4827 ( .A1(n3862), .A2(n3861), .ZN(n3869) );
  INV_X1 U4828 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3867) );
  NAND2_X1 U4829 ( .A1(n4352), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3866)
         );
  INV_X1 U4830 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3863) );
  XNOR2_X1 U4831 ( .A(n3864), .B(n3863), .ZN(n5807) );
  NAND2_X1 U4832 ( .A1(n5807), .A2(n3101), .ZN(n3865) );
  OAI211_X1 U4833 ( .C1(n4064), .C2(n3867), .A(n3866), .B(n3865), .ZN(n3868)
         );
  AOI21_X1 U4834 ( .B1(n4066), .B2(n3869), .A(n3868), .ZN(n5486) );
  AOI22_X1 U4835 ( .A1(n3353), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3977), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4836 ( .A1(n3905), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4837 ( .A1(n3542), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4838 ( .A1(n3956), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4839 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3880)
         );
  AOI22_X1 U4840 ( .A1(n3818), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4841 ( .A1(n3530), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4842 ( .A1(n3544), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4843 ( .A1(n3971), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4844 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3879)
         );
  OAI21_X1 U4845 ( .B1(n3880), .B2(n3879), .A(n3878), .ZN(n3885) );
  NAND2_X1 U4846 ( .A1(n4353), .A2(EAX_REG_15__SCAN_IN), .ZN(n3884) );
  XNOR2_X1 U4847 ( .A(n3898), .B(n3881), .ZN(n5817) );
  NAND2_X1 U4848 ( .A1(n5817), .A2(n3101), .ZN(n3883) );
  NAND2_X1 U4849 ( .A1(n4352), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3882)
         );
  AOI22_X1 U4850 ( .A1(n3977), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4851 ( .A1(n3818), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4852 ( .A1(n3956), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4853 ( .A1(n3971), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4854 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4855 ( .A1(n3905), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4856 ( .A1(n3989), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4857 ( .A1(n3530), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4858 ( .A1(n3353), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4859 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  NOR2_X1 U4860 ( .A1(n3895), .A2(n3894), .ZN(n3903) );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U4862 ( .A1(n3896), .A2(n6980), .ZN(n3897) );
  NAND2_X1 U4863 ( .A1(n3898), .A2(n3897), .ZN(n5825) );
  NOR2_X1 U4864 ( .A1(n3899), .A2(n6980), .ZN(n3900) );
  AOI21_X1 U4865 ( .B1(n5825), .B2(n3101), .A(n3900), .ZN(n3902) );
  NAND2_X1 U4866 ( .A1(n4353), .A2(EAX_REG_14__SCAN_IN), .ZN(n3901) );
  OAI211_X1 U4867 ( .C1(n3904), .C2(n3903), .A(n3902), .B(n3901), .ZN(n5516)
         );
  AOI22_X1 U4868 ( .A1(n3353), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3977), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4869 ( .A1(n3818), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3905), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4870 ( .A1(n3530), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4871 ( .A1(n3990), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4872 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3915)
         );
  AOI22_X1 U4873 ( .A1(n3956), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4874 ( .A1(n3544), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4875 ( .A1(n3542), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4876 ( .A1(n3971), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4877 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  NOR2_X1 U4878 ( .A1(n3915), .A2(n3914), .ZN(n3918) );
  INV_X1 U4879 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5794) );
  AOI21_X1 U4880 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5794), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3916) );
  AOI21_X1 U4881 ( .B1(n4353), .B2(EAX_REG_17__SCAN_IN), .A(n3916), .ZN(n3917)
         );
  OAI21_X1 U4882 ( .B1(n4036), .B2(n3918), .A(n3917), .ZN(n3921) );
  XNOR2_X1 U4883 ( .A(n3919), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5796)
         );
  NAND2_X1 U4884 ( .A1(n5796), .A2(n3101), .ZN(n3920) );
  AOI22_X1 U4885 ( .A1(n3956), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4886 ( .A1(n3542), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4887 ( .A1(n3977), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4888 ( .A1(n3971), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4889 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3931)
         );
  AOI22_X1 U4890 ( .A1(n3818), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3372), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4891 ( .A1(n3544), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4892 ( .A1(n3530), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4893 ( .A1(n3353), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4894 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NOR2_X1 U4895 ( .A1(n3931), .A2(n3930), .ZN(n3933) );
  AOI22_X1 U4896 ( .A1(n4353), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6632), .ZN(n3932) );
  OAI21_X1 U4897 ( .B1(n4036), .B2(n3933), .A(n3932), .ZN(n3938) );
  INV_X1 U4898 ( .A(n3934), .ZN(n3936) );
  INV_X1 U4899 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4900 ( .A1(n3936), .A2(n3935), .ZN(n3937) );
  NAND2_X1 U4901 ( .A1(n3952), .A2(n3937), .ZN(n5787) );
  MUX2_X1 U4902 ( .A(n3938), .B(n5787), .S(n3101), .Z(n5453) );
  AOI22_X1 U4903 ( .A1(n3977), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4904 ( .A1(n3905), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4905 ( .A1(n3956), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4906 ( .A1(n3353), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4907 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3948)
         );
  AOI22_X1 U4908 ( .A1(n3818), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4909 ( .A1(n3989), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4910 ( .A1(n3992), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4911 ( .A1(n3971), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4912 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947)
         );
  NOR2_X1 U4913 ( .A1(n3948), .A2(n3947), .ZN(n3950) );
  AOI22_X1 U4914 ( .A1(n4353), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6632), .ZN(n3949) );
  OAI21_X1 U4915 ( .B1(n4036), .B2(n3950), .A(n3949), .ZN(n3953) );
  XNOR2_X1 U4916 ( .A(n3952), .B(n3951), .ZN(n5779) );
  MUX2_X1 U4917 ( .A(n3953), .B(n5779), .S(n3101), .Z(n5436) );
  NAND2_X1 U4918 ( .A1(n3954), .A2(n6962), .ZN(n3955) );
  NAND2_X1 U4919 ( .A1(n3986), .A2(n3955), .ZN(n5772) );
  AOI22_X1 U4920 ( .A1(n3977), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4921 ( .A1(n3989), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4922 ( .A1(n3956), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4923 ( .A1(n3353), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4924 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3966)
         );
  AOI22_X1 U4925 ( .A1(n3818), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4926 ( .A1(n3905), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3541), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4927 ( .A1(n3997), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4928 ( .A1(n3992), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3961) );
  NAND4_X1 U4929 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3965)
         );
  NOR2_X1 U4930 ( .A1(n3966), .A2(n3965), .ZN(n3968) );
  AOI22_X1 U4931 ( .A1(n4353), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6632), .ZN(n3967) );
  OAI21_X1 U4932 ( .B1(n4036), .B2(n3968), .A(n3967), .ZN(n3969) );
  MUX2_X1 U4933 ( .A(n5772), .B(n3969), .S(n4019), .Z(n3970) );
  AOI22_X1 U4934 ( .A1(n3905), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3542), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4935 ( .A1(n3956), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4936 ( .A1(n3992), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4937 ( .A1(n3544), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4938 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3983)
         );
  AOI22_X1 U4939 ( .A1(n3818), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4940 ( .A1(n3989), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4941 ( .A1(n3353), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4942 ( .A1(n3977), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3978) );
  NAND4_X1 U4943 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3982)
         );
  OAI21_X1 U4944 ( .B1(n3983), .B2(n3982), .A(n4066), .ZN(n3985) );
  AOI22_X1 U4945 ( .A1(n4353), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6632), .ZN(n3984) );
  AND2_X1 U4946 ( .A1(n3985), .A2(n3984), .ZN(n3988) );
  INV_X1 U4947 ( .A(n3986), .ZN(n3987) );
  XOR2_X1 U4948 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3987), .Z(n5763) );
  MUX2_X1 U4949 ( .A(n3988), .B(n5763), .S(n3101), .Z(n5412) );
  AOI22_X1 U4950 ( .A1(n3818), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4951 ( .A1(n3905), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3530), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4952 ( .A1(n3544), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3990), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4953 ( .A1(n3992), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4954 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4004)
         );
  AOI22_X1 U4955 ( .A1(n3956), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3529), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4956 ( .A1(n3353), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3976), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4957 ( .A1(n3431), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3971), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4958 ( .A1(n3998), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3997), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4959 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  OAI21_X1 U4960 ( .B1(n4004), .B2(n4003), .A(n4066), .ZN(n4006) );
  AOI22_X1 U4961 ( .A1(n4353), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6632), .ZN(n4005) );
  NAND2_X1 U4962 ( .A1(n4006), .A2(n4005), .ZN(n4010) );
  INV_X1 U4963 ( .A(n4007), .ZN(n4008) );
  INV_X1 U4964 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U4965 ( .A1(n4008), .A2(n5398), .ZN(n4009) );
  NAND2_X1 U4966 ( .A1(n4011), .A2(n4009), .ZN(n5756) );
  MUX2_X1 U4967 ( .A(n4010), .B(n5756), .S(n3101), .Z(n5395) );
  XNOR2_X1 U4968 ( .A(n4011), .B(n3142), .ZN(n5748) );
  INV_X1 U4969 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4017) );
  XOR2_X1 U4970 ( .A(n4013), .B(n4012), .Z(n4014) );
  NAND2_X1 U4971 ( .A1(n4066), .A2(n4014), .ZN(n4016) );
  OAI21_X1 U4972 ( .B1(n6225), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6632), 
        .ZN(n4015) );
  OAI211_X1 U4973 ( .C1(n4064), .C2(n4017), .A(n4016), .B(n4015), .ZN(n4018)
         );
  XNOR2_X1 U4974 ( .A(n4021), .B(n4020), .ZN(n4025) );
  OAI21_X1 U4975 ( .B1(n4022), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4031), 
        .ZN(n5740) );
  NAND2_X1 U4976 ( .A1(n5740), .A2(n3101), .ZN(n4024) );
  AOI22_X1 U4977 ( .A1(n4353), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4352), .ZN(n4023) );
  OAI211_X1 U4978 ( .C1(n4025), .C2(n4036), .A(n4024), .B(n4023), .ZN(n5374)
         );
  XOR2_X1 U4979 ( .A(n4027), .B(n4026), .Z(n4030) );
  INV_X1 U4980 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4028) );
  INV_X1 U4981 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5723) );
  OAI22_X1 U4982 ( .A1(n4064), .A2(n4028), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5723), .ZN(n4029) );
  AOI21_X1 U4983 ( .B1(n4030), .B2(n4066), .A(n4029), .ZN(n4032) );
  XNOR2_X1 U4984 ( .A(n4031), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5725)
         );
  MUX2_X1 U4985 ( .A(n4032), .B(n5725), .S(n3101), .Z(n5362) );
  XNOR2_X1 U4986 ( .A(n4034), .B(n4033), .ZN(n4037) );
  AOI22_X1 U4987 ( .A1(n4353), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6632), .ZN(n4035) );
  OAI21_X1 U4988 ( .B1(n4037), .B2(n4036), .A(n4035), .ZN(n4042) );
  INV_X1 U4989 ( .A(n4038), .ZN(n4040) );
  INV_X1 U4990 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4039) );
  NAND2_X1 U4991 ( .A1(n4040), .A2(n4039), .ZN(n4041) );
  NAND2_X1 U4992 ( .A1(n4048), .A2(n4041), .ZN(n5716) );
  MUX2_X1 U4993 ( .A(n4042), .B(n5716), .S(n3101), .Z(n5348) );
  XOR2_X1 U4994 ( .A(n4044), .B(n4043), .Z(n4045) );
  NAND2_X1 U4995 ( .A1(n4045), .A2(n4066), .ZN(n4047) );
  AOI22_X1 U4996 ( .A1(n4353), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6632), .ZN(n4046) );
  NAND2_X1 U4997 ( .A1(n4047), .A2(n4046), .ZN(n4049) );
  XOR2_X1 U4998 ( .A(n4048), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .Z(n5708) );
  XOR2_X1 U4999 ( .A(n4051), .B(n4050), .Z(n4054) );
  INV_X1 U5000 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4052) );
  INV_X1 U5001 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5703) );
  OAI22_X1 U5002 ( .A1(n4064), .A2(n4052), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5703), .ZN(n4053) );
  AOI21_X1 U5003 ( .B1(n4054), .B2(n4066), .A(n4053), .ZN(n4058) );
  INV_X1 U5004 ( .A(n4055), .ZN(n4056) );
  NAND2_X1 U5005 ( .A1(n4056), .A2(n5703), .ZN(n4057) );
  MUX2_X1 U5006 ( .A(n4058), .B(n5701), .S(n3101), .Z(n5326) );
  XNOR2_X1 U5007 ( .A(n4059), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5314)
         );
  XOR2_X1 U5008 ( .A(n4061), .B(n4060), .Z(n4067) );
  INV_X1 U5009 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4063) );
  NOR2_X1 U5010 ( .A1(n6225), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4062)
         );
  OAI22_X1 U5011 ( .A1(n4064), .A2(n4063), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4062), .ZN(n4065) );
  AOI21_X1 U5012 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4068) );
  INV_X1 U5013 ( .A(n5694), .ZN(n5631) );
  XNOR2_X1 U5014 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4076) );
  AOI21_X1 U5015 ( .B1(n4239), .B2(n4076), .A(n4633), .ZN(n4072) );
  NAND2_X1 U5016 ( .A1(n3502), .A2(n4688), .ZN(n4071) );
  NAND2_X1 U5017 ( .A1(n4871), .A2(n4071), .ZN(n4089) );
  OR2_X1 U5018 ( .A1(n4072), .A2(n4089), .ZN(n4081) );
  XNOR2_X1 U5019 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U5020 ( .A1(n4073), .A2(n4074), .ZN(n4088) );
  OAI21_X1 U5021 ( .B1(n4074), .B2(n4073), .A(n4088), .ZN(n4361) );
  AOI21_X1 U5022 ( .B1(n4123), .B2(n4684), .A(n4075), .ZN(n4082) );
  NAND2_X1 U5023 ( .A1(n4082), .A2(n4361), .ZN(n4077) );
  NAND4_X1 U5024 ( .A1(n4077), .A2(n4123), .A3(n4076), .A4(n4081), .ZN(n4079)
         );
  NAND2_X1 U5025 ( .A1(n4079), .A2(n4114), .ZN(n4080) );
  OAI21_X1 U5026 ( .B1(n4081), .B2(n4361), .A(n4080), .ZN(n4086) );
  INV_X1 U5027 ( .A(n4082), .ZN(n4084) );
  INV_X1 U5028 ( .A(n4361), .ZN(n4083) );
  NAND3_X1 U5029 ( .A1(n4084), .A2(STATE2_REG_0__SCAN_IN), .A3(n4083), .ZN(
        n4085) );
  NAND2_X1 U5030 ( .A1(n4086), .A2(n4085), .ZN(n4092) );
  NAND2_X1 U5031 ( .A1(n4858), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U5032 ( .A1(n4088), .A2(n4087), .ZN(n4098) );
  XNOR2_X1 U5033 ( .A(n4098), .B(n4097), .ZN(n4360) );
  INV_X1 U5034 ( .A(n4360), .ZN(n4090) );
  NAND2_X1 U5035 ( .A1(n4123), .A2(n4090), .ZN(n4093) );
  INV_X1 U5036 ( .A(n4089), .ZN(n4094) );
  OAI211_X1 U5037 ( .C1(n4090), .C2(n4109), .A(n4093), .B(n4094), .ZN(n4091)
         );
  NAND2_X1 U5038 ( .A1(n4092), .A2(n4091), .ZN(n4096) );
  NAND2_X1 U5039 ( .A1(n4096), .A2(n4095), .ZN(n4105) );
  NAND2_X1 U5040 ( .A1(n4098), .A2(n4097), .ZN(n4100) );
  NAND2_X1 U5041 ( .A1(n6143), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U5042 ( .A1(n4100), .A2(n4099), .ZN(n4102) );
  NOR2_X1 U5043 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  OR2_X1 U5044 ( .A1(n4108), .A2(n4103), .ZN(n4362) );
  NAND2_X1 U5045 ( .A1(n4109), .A2(n4362), .ZN(n4104) );
  NAND2_X1 U5046 ( .A1(n4105), .A2(n4104), .ZN(n4107) );
  NAND2_X1 U5047 ( .A1(n4120), .A2(n4362), .ZN(n4106) );
  NAND2_X1 U5048 ( .A1(n4107), .A2(n4106), .ZN(n4112) );
  NAND3_X1 U5049 ( .A1(n4113), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(n4119), .ZN(n4364) );
  INV_X1 U5050 ( .A(n4364), .ZN(n4110) );
  NAND2_X1 U5051 ( .A1(n4110), .A2(n4109), .ZN(n4111) );
  NAND2_X1 U5052 ( .A1(n4112), .A2(n4111), .ZN(n4117) );
  OAI22_X1 U5053 ( .A1(n4364), .A2(n4114), .B1(STATE2_REG_0__SCAN_IN), .B2(
        n4113), .ZN(n4115) );
  INV_X1 U5054 ( .A(n4115), .ZN(n4116) );
  NAND2_X1 U5055 ( .A1(n4117), .A2(n4116), .ZN(n4122) );
  NOR2_X1 U5056 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6466), .ZN(n4118)
         );
  NAND2_X1 U5057 ( .A1(n4363), .A2(n4120), .ZN(n4121) );
  NOR2_X1 U5058 ( .A1(n4852), .A2(n5424), .ZN(n4126) );
  NAND2_X1 U5059 ( .A1(n4126), .A2(n4529), .ZN(n4878) );
  NOR2_X1 U5060 ( .A1(n4878), .A2(n5114), .ZN(n4127) );
  NAND2_X1 U5061 ( .A1(n4876), .A2(n4127), .ZN(n4136) );
  INV_X1 U5062 ( .A(n4128), .ZN(n4132) );
  AND4_X1 U5063 ( .A1(n4413), .A2(n4130), .A3(n4703), .A4(n4129), .ZN(n4131)
         );
  NAND3_X1 U5064 ( .A1(n4133), .A2(n4132), .A3(n4131), .ZN(n4411) );
  AND2_X4 U5065 ( .A1(n3554), .A2(n4134), .ZN(n6752) );
  INV_X4 U5066 ( .A(n6752), .ZN(n5296) );
  OR2_X1 U5067 ( .A1(n5272), .A2(EBX_REG_1__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U5068 ( .A1(n4221), .A2(n4591), .ZN(n4137) );
  OAI211_X1 U5069 ( .C1(n5296), .C2(EBX_REG_1__SCAN_IN), .A(n5424), .B(n4137), 
        .ZN(n4138) );
  NAND2_X1 U5070 ( .A1(n4139), .A2(n4138), .ZN(n4141) );
  NAND2_X1 U5071 ( .A1(n4221), .A2(EBX_REG_0__SCAN_IN), .ZN(n4140) );
  OAI21_X1 U5072 ( .B1(n5439), .B2(EBX_REG_0__SCAN_IN), .A(n4140), .ZN(n4605)
         );
  XNOR2_X1 U5073 ( .A(n4141), .B(n4605), .ZN(n4582) );
  NAND2_X1 U5074 ( .A1(n4582), .A2(n6752), .ZN(n4583) );
  NAND2_X1 U5075 ( .A1(n4583), .A2(n4141), .ZN(n4650) );
  INV_X1 U5076 ( .A(n4650), .ZN(n4148) );
  NOR2_X1 U5077 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4142)
         );
  OR2_X1 U5078 ( .A1(n5272), .A2(EBX_REG_2__SCAN_IN), .ZN(n4146) );
  INV_X1 U5079 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U5080 ( .A1(n4221), .A2(n4143), .ZN(n4144) );
  OAI211_X1 U5081 ( .C1(n5296), .C2(EBX_REG_2__SCAN_IN), .A(n5424), .B(n4144), 
        .ZN(n4145) );
  NAND2_X1 U5082 ( .A1(n4146), .A2(n4145), .ZN(n5573) );
  NAND2_X1 U5083 ( .A1(n4148), .A2(n4147), .ZN(n4759) );
  OR2_X1 U5084 ( .A1(n5272), .A2(EBX_REG_4__SCAN_IN), .ZN(n4151) );
  INV_X1 U5085 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4277) );
  NAND2_X1 U5086 ( .A1(n4221), .A2(n4277), .ZN(n4149) );
  OAI211_X1 U5087 ( .C1(n5296), .C2(EBX_REG_4__SCAN_IN), .A(n5424), .B(n4149), 
        .ZN(n4150) );
  AND2_X1 U5088 ( .A1(n4151), .A2(n4150), .ZN(n4758) );
  MUX2_X1 U5089 ( .A(n4152), .B(n5439), .S(EBX_REG_5__SCAN_IN), .Z(n4154) );
  NOR2_X1 U5090 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4153)
         );
  NOR2_X1 U5091 ( .A1(n4154), .A2(n4153), .ZN(n4998) );
  NAND2_X1 U5092 ( .A1(n4760), .A2(n4998), .ZN(n4997) );
  INV_X1 U5093 ( .A(n4997), .ZN(n4161) );
  INV_X1 U5094 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4155) );
  MUX2_X1 U5095 ( .A(n4221), .B(n5272), .S(n4155), .Z(n4159) );
  INV_X1 U5096 ( .A(n4221), .ZN(n4156) );
  NAND2_X1 U5097 ( .A1(n4156), .A2(n5296), .ZN(n4179) );
  NAND2_X1 U5098 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5296), .ZN(n4157)
         );
  AND2_X1 U5099 ( .A1(n4179), .A2(n4157), .ZN(n4158) );
  INV_X1 U5100 ( .A(n5234), .ZN(n4160) );
  NAND2_X1 U5101 ( .A1(n4161), .A2(n4160), .ZN(n5222) );
  INV_X1 U5102 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4163) );
  INV_X1 U5103 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U5104 ( .A1(n6752), .A2(n6281), .ZN(n4162) );
  OAI211_X1 U5105 ( .C1(n5439), .C2(n4163), .A(n4162), .B(n4221), .ZN(n4164)
         );
  OAI21_X1 U5106 ( .B1(n4210), .B2(EBX_REG_7__SCAN_IN), .A(n4164), .ZN(n5225)
         );
  OR2_X1 U5107 ( .A1(n5272), .A2(EBX_REG_8__SCAN_IN), .ZN(n4167) );
  INV_X1 U5108 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4312) );
  NAND2_X1 U5109 ( .A1(n4221), .A2(n4312), .ZN(n4165) );
  OAI211_X1 U5110 ( .C1(n5296), .C2(EBX_REG_8__SCAN_IN), .A(n5424), .B(n4165), 
        .ZN(n4166) );
  MUX2_X1 U5111 ( .A(n4152), .B(n5439), .S(EBX_REG_9__SCAN_IN), .Z(n4169) );
  NOR2_X1 U5112 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4168)
         );
  NOR2_X1 U5113 ( .A1(n4169), .A2(n4168), .ZN(n5626) );
  INV_X1 U5114 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4170) );
  MUX2_X1 U5115 ( .A(n4221), .B(n5272), .S(n4170), .Z(n4173) );
  NAND2_X1 U5116 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5296), .ZN(n4171) );
  AND2_X1 U5117 ( .A1(n4179), .A2(n4171), .ZN(n4172) );
  NAND2_X1 U5118 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4176) );
  OAI211_X1 U5119 ( .C1(n5296), .C2(EBX_REG_11__SCAN_IN), .A(n4221), .B(n4176), 
        .ZN(n4177) );
  OAI21_X1 U5120 ( .B1(n4210), .B2(EBX_REG_11__SCAN_IN), .A(n4177), .ZN(n6099)
         );
  MUX2_X1 U5121 ( .A(n5272), .B(n4221), .S(EBX_REG_12__SCAN_IN), .Z(n4181) );
  NAND2_X1 U5122 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5296), .ZN(n4178) );
  AND2_X1 U5123 ( .A1(n4179), .A2(n4178), .ZN(n4180) );
  NAND2_X1 U5124 ( .A1(n4181), .A2(n4180), .ZN(n5530) );
  INV_X1 U5125 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U5126 ( .A1(n4152), .A2(n6246), .ZN(n4184) );
  NAND2_X1 U5127 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4182) );
  OAI211_X1 U5128 ( .C1(n5296), .C2(EBX_REG_13__SCAN_IN), .A(n4221), .B(n4182), 
        .ZN(n4183) );
  INV_X1 U5129 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6825) );
  MUX2_X1 U5130 ( .A(n4221), .B(n5272), .S(n6825), .Z(n4186) );
  NAND2_X1 U5131 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4185) );
  NAND2_X1 U5132 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4187) );
  OAI211_X1 U5133 ( .C1(n5296), .C2(EBX_REG_15__SCAN_IN), .A(n4221), .B(n4187), 
        .ZN(n4188) );
  OAI21_X1 U5134 ( .B1(n4210), .B2(EBX_REG_15__SCAN_IN), .A(n4188), .ZN(n5498)
         );
  MUX2_X1 U5135 ( .A(n5272), .B(n4221), .S(EBX_REG_16__SCAN_IN), .Z(n4190) );
  NAND2_X1 U5136 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4189) );
  NAND2_X1 U5137 ( .A1(n4190), .A2(n4189), .ZN(n5487) );
  INV_X1 U5138 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U5139 ( .A1(n4152), .A2(n5609), .ZN(n4193) );
  NAND2_X1 U5140 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4191) );
  OAI211_X1 U5141 ( .C1(n5296), .C2(EBX_REG_17__SCAN_IN), .A(n4221), .B(n4191), 
        .ZN(n4192) );
  NAND2_X1 U5142 ( .A1(n5468), .A2(n5469), .ZN(n5438) );
  INV_X2 U5143 ( .A(n5438), .ZN(n4198) );
  OR2_X1 U5144 ( .A1(n5272), .A2(EBX_REG_19__SCAN_IN), .ZN(n4196) );
  INV_X1 U5145 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U5146 ( .A1(n4221), .A2(n5732), .ZN(n4194) );
  OAI211_X1 U5147 ( .C1(n5296), .C2(EBX_REG_19__SCAN_IN), .A(n5424), .B(n4194), 
        .ZN(n4195) );
  INV_X1 U5148 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6908) );
  OR2_X1 U5149 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4199)
         );
  OR2_X1 U5150 ( .A1(n5296), .A2(EBX_REG_18__SCAN_IN), .ZN(n5440) );
  OAI22_X1 U5151 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n5296), .B2(EBX_REG_20__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U5152 ( .A1(n4200), .A2(n5425), .ZN(n4202) );
  NAND2_X1 U5153 ( .A1(n5441), .A2(n5424), .ZN(n4201) );
  OAI211_X1 U5154 ( .C1(n5424), .C2(n6908), .A(n4202), .B(n4201), .ZN(n4203)
         );
  MUX2_X1 U5155 ( .A(n4152), .B(n5439), .S(EBX_REG_21__SCAN_IN), .Z(n4205) );
  NOR2_X1 U5156 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4204)
         );
  NOR2_X1 U5157 ( .A1(n4205), .A2(n4204), .ZN(n5409) );
  INV_X1 U5158 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6938) );
  MUX2_X1 U5159 ( .A(n4221), .B(n5272), .S(n6938), .Z(n4207) );
  NAND2_X1 U5160 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5161 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4208) );
  OAI211_X1 U5162 ( .C1(n5296), .C2(EBX_REG_23__SCAN_IN), .A(n4221), .B(n4208), 
        .ZN(n4209) );
  OAI21_X1 U5163 ( .B1(n4210), .B2(EBX_REG_23__SCAN_IN), .A(n4209), .ZN(n5382)
         );
  OR2_X2 U5164 ( .A1(n5402), .A2(n5382), .ZN(n5384) );
  INV_X1 U5165 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6850) );
  MUX2_X1 U5166 ( .A(n4221), .B(n5272), .S(n6850), .Z(n4212) );
  NAND2_X1 U5167 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4211) );
  NOR2_X4 U5168 ( .A1(n5384), .A2(n5376), .ZN(n5375) );
  MUX2_X1 U5169 ( .A(n4152), .B(n5439), .S(EBX_REG_25__SCAN_IN), .Z(n4214) );
  NOR2_X1 U5170 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4213)
         );
  NOR2_X1 U5171 ( .A1(n4214), .A2(n4213), .ZN(n5359) );
  OR2_X1 U5172 ( .A1(n5272), .A2(EBX_REG_26__SCAN_IN), .ZN(n4217) );
  INV_X1 U5173 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U5174 ( .A1(n4221), .A2(n6851), .ZN(n4215) );
  OAI211_X1 U5175 ( .C1(n5296), .C2(EBX_REG_26__SCAN_IN), .A(n5424), .B(n4215), 
        .ZN(n4216) );
  NAND2_X1 U5176 ( .A1(n4217), .A2(n4216), .ZN(n5353) );
  INV_X1 U5177 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5178 ( .A1(n4152), .A2(n5599), .ZN(n4220) );
  NAND2_X1 U5179 ( .A1(n5424), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4218) );
  OAI211_X1 U5180 ( .C1(n5296), .C2(EBX_REG_27__SCAN_IN), .A(n4221), .B(n4218), 
        .ZN(n4219) );
  OR2_X1 U5181 ( .A1(n5272), .A2(EBX_REG_28__SCAN_IN), .ZN(n4224) );
  INV_X1 U5182 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U5183 ( .A1(n4221), .A2(n5697), .ZN(n4222) );
  OAI211_X1 U5184 ( .C1(n5296), .C2(EBX_REG_28__SCAN_IN), .A(n5424), .B(n4222), 
        .ZN(n4223) );
  AND2_X1 U5185 ( .A1(n4224), .A2(n4223), .ZN(n5322) );
  OAI22_X1 U5186 ( .A1(n5297), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n5296), .B2(EBX_REG_29__SCAN_IN), .ZN(n5277) );
  INV_X1 U5187 ( .A(n5274), .ZN(n4230) );
  NAND2_X1 U5188 ( .A1(n4230), .A2(n5424), .ZN(n5292) );
  OR2_X1 U5189 ( .A1(n5274), .A2(n5324), .ZN(n4227) );
  NAND2_X1 U5190 ( .A1(n5297), .A2(EBX_REG_30__SCAN_IN), .ZN(n4226) );
  NAND2_X1 U5191 ( .A1(n5296), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4225) );
  NAND2_X1 U5192 ( .A1(n4226), .A2(n4225), .ZN(n5293) );
  NAND2_X1 U5193 ( .A1(n5292), .A2(n4228), .ZN(n4232) );
  INV_X1 U5194 ( .A(n5324), .ZN(n5273) );
  INV_X1 U5195 ( .A(n5293), .ZN(n4229) );
  OAI211_X1 U5196 ( .C1(n5273), .C2(n5424), .A(n4230), .B(n4229), .ZN(n4231)
         );
  INV_X1 U5197 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4400) );
  OAI21_X1 U5198 ( .B1(n5631), .B2(n7064), .A(n4236), .ZN(U2829) );
  NAND2_X1 U5199 ( .A1(n4852), .A2(n4633), .ZN(n4237) );
  NAND2_X1 U5200 ( .A1(n4238), .A2(n4237), .ZN(n4507) );
  OR2_X1 U5201 ( .A1(n4507), .A2(n4239), .ZN(n4869) );
  NAND2_X1 U5202 ( .A1(n4661), .A2(n4297), .ZN(n4243) );
  NAND2_X1 U5203 ( .A1(n4245), .A2(n4253), .ZN(n4244) );
  NAND2_X1 U5204 ( .A1(n4244), .A2(n4240), .ZN(n4270) );
  OAI21_X1 U5205 ( .B1(n4240), .B2(n4244), .A(n4270), .ZN(n4241) );
  AND2_X1 U5206 ( .A1(n4633), .A2(n4668), .ZN(n4251) );
  AOI21_X1 U5207 ( .B1(n4241), .B2(n5280), .A(n4251), .ZN(n4242) );
  NAND2_X1 U5208 ( .A1(n4258), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6400)
         );
  NAND2_X1 U5209 ( .A1(n4625), .A2(n4297), .ZN(n4250) );
  OAI21_X1 U5210 ( .B1(n4245), .B2(n4253), .A(n4244), .ZN(n4247) );
  INV_X1 U5211 ( .A(n4524), .ZN(n4246) );
  OAI211_X1 U5212 ( .C1(n4247), .C2(n4391), .A(n4246), .B(n4688), .ZN(n4248)
         );
  INV_X1 U5213 ( .A(n4248), .ZN(n4249) );
  NAND2_X1 U5214 ( .A1(n4250), .A2(n4249), .ZN(n4560) );
  INV_X1 U5215 ( .A(n4297), .ZN(n4305) );
  INV_X1 U5216 ( .A(n4251), .ZN(n4252) );
  OAI21_X1 U5217 ( .B1(n4391), .B2(n4253), .A(n4252), .ZN(n4254) );
  INV_X1 U5218 ( .A(n4254), .ZN(n4255) );
  OAI21_X1 U5219 ( .B1(n5163), .B2(n4305), .A(n4255), .ZN(n5883) );
  NAND2_X1 U5220 ( .A1(n5883), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6457)
         );
  XNOR2_X1 U5221 ( .A(n6457), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4559)
         );
  NAND2_X1 U5222 ( .A1(n4560), .A2(n4559), .ZN(n4558) );
  INV_X1 U5223 ( .A(n6457), .ZN(n4256) );
  NAND2_X1 U5224 ( .A1(n4256), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4257)
         );
  NAND2_X1 U5225 ( .A1(n6400), .A2(n6403), .ZN(n4260) );
  NAND2_X1 U5226 ( .A1(n4259), .A2(n4143), .ZN(n6401) );
  INV_X1 U5227 ( .A(n4269), .ZN(n4261) );
  XNOR2_X1 U5228 ( .A(n4270), .B(n4261), .ZN(n4262) );
  NAND2_X1 U5229 ( .A1(n4262), .A2(n5280), .ZN(n4263) );
  OAI21_X2 U5230 ( .B1(n4893), .B2(n4305), .A(n4263), .ZN(n4265) );
  INV_X1 U5231 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4264) );
  XNOR2_X1 U5232 ( .A(n4265), .B(n4264), .ZN(n4648) );
  NAND2_X1 U5233 ( .A1(n4649), .A2(n4648), .ZN(n4267) );
  NAND2_X1 U5234 ( .A1(n4265), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4266)
         );
  NAND2_X1 U5235 ( .A1(n4267), .A2(n4266), .ZN(n4840) );
  NAND2_X1 U5236 ( .A1(n4270), .A2(n4269), .ZN(n4272) );
  INV_X1 U5237 ( .A(n4272), .ZN(n4274) );
  INV_X1 U5238 ( .A(n4273), .ZN(n4271) );
  OR2_X1 U5239 ( .A1(n4272), .A2(n4271), .ZN(n4291) );
  OAI211_X1 U5240 ( .C1(n4274), .C2(n4273), .A(n5280), .B(n4291), .ZN(n4275)
         );
  XNOR2_X1 U5241 ( .A(n4278), .B(n4277), .ZN(n4841) );
  NAND2_X1 U5242 ( .A1(n4840), .A2(n4841), .ZN(n4280) );
  NAND2_X1 U5243 ( .A1(n4278), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4279)
         );
  NAND2_X1 U5244 ( .A1(n4280), .A2(n4279), .ZN(n5098) );
  XNOR2_X1 U5245 ( .A(n4291), .B(n4289), .ZN(n4282) );
  NAND2_X1 U5246 ( .A1(n4282), .A2(n5280), .ZN(n4283) );
  NAND2_X1 U5247 ( .A1(n4284), .A2(n4283), .ZN(n4286) );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4285) );
  XNOR2_X1 U5249 ( .A(n4286), .B(n4285), .ZN(n5099) );
  NAND2_X1 U5250 ( .A1(n4286), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4287)
         );
  INV_X1 U5251 ( .A(n4289), .ZN(n4290) );
  NOR2_X1 U5252 ( .A1(n4291), .A2(n4290), .ZN(n4293) );
  NAND2_X1 U5253 ( .A1(n4293), .A2(n4292), .ZN(n4310) );
  OAI211_X1 U5254 ( .C1(n4293), .C2(n4292), .A(n4310), .B(n5280), .ZN(n4294)
         );
  INV_X1 U5255 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4295) );
  XNOR2_X1 U5256 ( .A(n4296), .B(n4295), .ZN(n5229) );
  NAND2_X1 U5257 ( .A1(n4298), .A2(n4297), .ZN(n4301) );
  XNOR2_X1 U5258 ( .A(n4310), .B(n4308), .ZN(n4299) );
  NAND2_X1 U5259 ( .A1(n4299), .A2(n5280), .ZN(n4300) );
  NAND2_X1 U5260 ( .A1(n4301), .A2(n4300), .ZN(n4302) );
  XNOR2_X1 U5261 ( .A(n4302), .B(n4163), .ZN(n5247) );
  NAND2_X1 U5262 ( .A1(n4302), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4303)
         );
  NOR2_X1 U5263 ( .A1(n4306), .A2(n4305), .ZN(n4307) );
  NAND2_X1 U5264 ( .A1(n5280), .A2(n4308), .ZN(n4309) );
  OR2_X1 U5265 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  NAND2_X1 U5266 ( .A1(n4327), .A2(n4311), .ZN(n4313) );
  XNOR2_X1 U5267 ( .A(n4313), .B(n4312), .ZN(n5875) );
  INV_X1 U5268 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U5269 ( .A1(n3099), .A2(n6438), .ZN(n4315) );
  INV_X1 U5270 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6963) );
  AND2_X1 U5271 ( .A1(n3099), .A2(n6963), .ZN(n5855) );
  INV_X1 U5272 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7032) );
  NAND2_X1 U5273 ( .A1(n3099), .A2(n7032), .ZN(n5845) );
  INV_X1 U5274 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U5275 ( .A1(n3099), .A2(n5835), .ZN(n4316) );
  NAND2_X1 U5276 ( .A1(n5845), .A2(n4316), .ZN(n4320) );
  NOR2_X1 U5277 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4317) );
  OR2_X1 U5278 ( .A1(n3099), .A2(n4317), .ZN(n4318) );
  AND2_X1 U5279 ( .A1(n5854), .A2(n4318), .ZN(n4319) );
  NOR2_X1 U5280 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4321) );
  INV_X1 U5281 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U5282 ( .A1(n4327), .A2(n6086), .ZN(n5821) );
  AND2_X1 U5283 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4322) );
  NAND4_X1 U5284 ( .A1(n4322), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A4(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n4323) );
  AND2_X1 U5285 ( .A1(n3099), .A2(n4323), .ZN(n4324) );
  INV_X1 U5286 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6059) );
  INV_X1 U5287 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6028) );
  INV_X1 U5288 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6048) );
  INV_X1 U5289 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6037) );
  AND3_X1 U5290 ( .A1(n6028), .A2(n6048), .A3(n6037), .ZN(n4325) );
  OR2_X1 U5291 ( .A1(n3099), .A2(n4325), .ZN(n4326) );
  NOR2_X1 U5292 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5978) );
  NOR2_X1 U5293 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6013) );
  INV_X1 U5294 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4328) );
  INV_X1 U5295 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6004) );
  NAND4_X1 U5296 ( .A1(n5978), .A2(n6013), .A3(n4328), .A4(n6004), .ZN(n4329)
         );
  AND2_X1 U5297 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6012) );
  AND2_X1 U5298 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5897) );
  AND2_X1 U5299 ( .A1(n6012), .A2(n5897), .ZN(n5974) );
  AND2_X1 U5300 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U5301 ( .A1(n5974), .A2(n5911), .ZN(n5916) );
  NAND2_X1 U5302 ( .A1(n4327), .A2(n5916), .ZN(n4330) );
  XNOR2_X1 U5303 ( .A(n5865), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5727)
         );
  INV_X1 U5304 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U5305 ( .A1(n3099), .A2(n6899), .ZN(n4331) );
  NAND2_X1 U5306 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5918) );
  INV_X1 U5307 ( .A(n5726), .ZN(n4333) );
  NOR2_X1 U5308 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4332)
         );
  INV_X1 U5309 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U5310 ( .A1(n5697), .A2(n5711), .ZN(n4334) );
  NAND2_X1 U5311 ( .A1(n5282), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4366) );
  NOR2_X1 U5312 ( .A1(n4366), .A2(n6225), .ZN(n4437) );
  NAND2_X1 U5313 ( .A1(n4343), .A2(n6636), .ZN(n4339) );
  NAND2_X1 U5314 ( .A1(n4339), .A2(n5282), .ZN(n4340) );
  NAND2_X1 U5315 ( .A1(n5282), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5316 ( .A1(n6225), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U5317 ( .A1(n4342), .A2(n4341), .ZN(n5884) );
  NAND2_X1 U5318 ( .A1(n6399), .A2(REIP_REG_29__SCAN_IN), .ZN(n5935) );
  OAI21_X1 U5319 ( .B1(n5868), .B2(n4344), .A(n5935), .ZN(n4345) );
  AOI21_X1 U5320 ( .B1(n5314), .B2(n5870), .A(n4345), .ZN(n4346) );
  OAI211_X1 U5321 ( .C1(n6226), .C2(n5942), .A(n4347), .B(n4346), .ZN(U2957)
         );
  INV_X1 U5322 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5685) );
  INV_X1 U5323 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U5324 ( .A1(n4349), .A2(n4348), .ZN(n4350) );
  AND2_X1 U5325 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U5326 ( .A1(n4350), .A2(n5688), .ZN(n4351) );
  XNOR2_X1 U5327 ( .A(n4351), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5926)
         );
  AOI22_X1 U5328 ( .A1(n4353), .A2(EAX_REG_31__SCAN_IN), .B1(n4352), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4354) );
  INV_X1 U5329 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U5330 ( .A1(n6399), .A2(REIP_REG_31__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U5331 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4357)
         );
  OAI211_X1 U5332 ( .C1(n4398), .C2(n6418), .A(n5921), .B(n4357), .ZN(n4358)
         );
  AOI21_X1 U5333 ( .B1(n5291), .B2(n6404), .A(n4358), .ZN(n4359) );
  OAI21_X1 U5334 ( .B1(n5926), .B2(n6226), .A(n4359), .ZN(U2955) );
  NOR3_X1 U5335 ( .A1(n4362), .A2(n4361), .A3(n4360), .ZN(n4365) );
  AOI21_X1 U5336 ( .B1(n4365), .B2(n4364), .A(n4363), .ZN(n4881) );
  NAND2_X1 U5337 ( .A1(n4881), .A2(n4502), .ZN(n4499) );
  INV_X1 U5338 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5339 ( .A1(n4367), .A2(n3101), .ZN(n6734) );
  NOR2_X1 U5340 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4435) );
  NOR2_X1 U5341 ( .A1(n5281), .A2(n4338), .ZN(n4368) );
  NAND2_X1 U5342 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4368), .ZN(n5108) );
  NAND3_X1 U5343 ( .A1(n6443), .A2(n6734), .A3(n5108), .ZN(n4369) );
  OR2_X4 U5344 ( .A1(n6756), .A2(n4369), .ZN(n6278) );
  NAND2_X2 U5345 ( .A1(n4370), .A2(n6278), .ZN(n5554) );
  NAND2_X1 U5346 ( .A1(n7019), .A2(n6225), .ZN(n4392) );
  NAND2_X1 U5347 ( .A1(n4392), .A2(EBX_REG_31__SCAN_IN), .ZN(n4371) );
  NOR2_X1 U5348 ( .A1(n5296), .A2(n4371), .ZN(n4372) );
  NOR2_X1 U5349 ( .A1(n5927), .A2(n6334), .ZN(n4405) );
  NOR2_X1 U5350 ( .A1(n4633), .A2(n4392), .ZN(n4374) );
  OR2_X1 U5351 ( .A1(n4373), .A2(STATE_REG_0__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U5352 ( .A1(n3502), .A2(n4870), .ZN(n4567) );
  AND2_X1 U5353 ( .A1(n4374), .A2(n4567), .ZN(n4375) );
  AND2_X2 U5354 ( .A1(n5557), .A2(n4375), .ZN(n6320) );
  INV_X1 U5355 ( .A(REIP_REG_13__SCAN_IN), .ZN(n4378) );
  INV_X1 U5356 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4376) );
  INV_X1 U5357 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6323) );
  NAND3_X1 U5358 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U5359 ( .A1(n6323), .A2(n5565), .ZN(n6311) );
  NAND2_X1 U5360 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6311), .ZN(n6284) );
  NAND2_X1 U5361 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n6286) );
  NOR2_X1 U5362 ( .A1(n6284), .A2(n6286), .ZN(n4424) );
  NAND2_X1 U5363 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4424), .ZN(n5542) );
  NOR2_X1 U5364 ( .A1(n4376), .A2(n5542), .ZN(n5545) );
  AND2_X1 U5365 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5545), .ZN(n6257) );
  NAND2_X1 U5366 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6257), .ZN(n5536) );
  INV_X1 U5367 ( .A(n5536), .ZN(n4377) );
  NAND2_X1 U5368 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4377), .ZN(n6244) );
  NOR2_X1 U5369 ( .A1(n4378), .A2(n6244), .ZN(n5519) );
  AND2_X1 U5370 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5519), .ZN(n5505) );
  AND2_X1 U5371 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5505), .ZN(n4379) );
  NAND2_X1 U5372 ( .A1(n6320), .A2(n4379), .ZN(n5494) );
  NAND2_X1 U5373 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .ZN(
        n4383) );
  NOR2_X2 U5374 ( .A1(n5494), .A2(n4383), .ZN(n5459) );
  NAND2_X1 U5375 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5445) );
  NOR2_X1 U5376 ( .A1(n5445), .A2(n6817), .ZN(n4380) );
  NAND2_X1 U5377 ( .A1(n5459), .A2(n4380), .ZN(n5414) );
  NAND3_X1 U5378 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5367) );
  NAND3_X1 U5379 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n4386) );
  INV_X1 U5380 ( .A(n5342), .ZN(n4382) );
  AND2_X1 U5381 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4381) );
  NAND2_X1 U5382 ( .A1(n4382), .A2(n4381), .ZN(n4396) );
  NOR2_X1 U5383 ( .A1(n4396), .A2(REIP_REG_29__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U5384 ( .A1(n6285), .A2(n6278), .ZN(n5594) );
  INV_X1 U5385 ( .A(n5445), .ZN(n5427) );
  AND2_X1 U5386 ( .A1(n6278), .A2(n5505), .ZN(n5502) );
  NAND2_X1 U5387 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5502), .ZN(n5491) );
  NOR2_X1 U5388 ( .A1(n5491), .A2(n4383), .ZN(n5443) );
  AND2_X1 U5389 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5443), .ZN(n5396) );
  INV_X1 U5390 ( .A(n5367), .ZN(n4384) );
  NAND3_X1 U5391 ( .A1(n5427), .A2(n5396), .A3(n4384), .ZN(n4385) );
  NAND2_X1 U5392 ( .A1(n5594), .A2(n4385), .ZN(n5387) );
  NAND2_X1 U5393 ( .A1(n5594), .A2(n4386), .ZN(n4387) );
  NAND2_X1 U5394 ( .A1(n5387), .A2(n4387), .ZN(n5357) );
  NAND2_X1 U5395 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4388) );
  AND2_X1 U5396 ( .A1(n6320), .A2(n4388), .ZN(n4389) );
  NOR2_X1 U5397 ( .A1(n5317), .A2(n5327), .ZN(n5301) );
  INV_X1 U5398 ( .A(n5301), .ZN(n4390) );
  NOR2_X1 U5399 ( .A1(n4870), .A2(n4392), .ZN(n4890) );
  NOR2_X1 U5400 ( .A1(n4391), .A2(n4890), .ZN(n5304) );
  INV_X1 U5401 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5402 ( .A1(n4392), .A2(n5596), .ZN(n4393) );
  NOR2_X1 U5403 ( .A1(n4633), .A2(n4393), .ZN(n4394) );
  OR2_X1 U5404 ( .A1(n5304), .A2(n4394), .ZN(n4395) );
  INV_X1 U5405 ( .A(n4396), .ZN(n5303) );
  INV_X1 U5406 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4489) );
  NOR2_X1 U5407 ( .A1(n4489), .A2(REIP_REG_30__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U5408 ( .A1(n5303), .A2(n4397), .ZN(n5300) );
  AOI22_X1 U5409 ( .A1(n6262), .A2(n5690), .B1(PHYADDRPOINTER_REG_30__SCAN_IN), 
        .B2(n6330), .ZN(n4399) );
  OAI211_X1 U5410 ( .C1(n4400), .C2(n6294), .A(n5300), .B(n4399), .ZN(n4401)
         );
  OR2_X1 U5411 ( .A1(n4507), .A2(n4871), .ZN(n4573) );
  INV_X1 U5412 ( .A(n4736), .ZN(n4518) );
  INV_X1 U5413 ( .A(n5114), .ZN(n6729) );
  INV_X1 U5414 ( .A(n4881), .ZN(n4407) );
  NOR2_X1 U5415 ( .A1(n4407), .A2(READY_N), .ZN(n4562) );
  NAND3_X1 U5416 ( .A1(n4518), .A2(n6729), .A3(n4562), .ZN(n4408) );
  OAI21_X1 U5417 ( .B1(n4595), .B2(n4573), .A(n4408), .ZN(n4409) );
  INV_X1 U5418 ( .A(n4409), .ZN(n4410) );
  NAND2_X1 U5419 ( .A1(n4802), .A2(n4410), .ZN(n4416) );
  NOR2_X1 U5420 ( .A1(n4411), .A2(n4871), .ZN(n4412) );
  AND2_X1 U5421 ( .A1(n5070), .A2(n4413), .ZN(n4414) );
  AOI22_X1 U5422 ( .A1(n5680), .A2(EAX_REG_31__SCAN_IN), .B1(n5661), .B2(
        DATAI_31_), .ZN(n4417) );
  NAND2_X1 U5423 ( .A1(n4418), .A2(n4417), .ZN(U2860) );
  INV_X1 U5424 ( .A(EBX_REG_8__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U5425 ( .A1(n6320), .A2(n5542), .ZN(n4425) );
  NAND2_X1 U5426 ( .A1(n6278), .A2(n4425), .ZN(n6267) );
  AOI22_X1 U5427 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6330), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6267), .ZN(n4420) );
  OR2_X1 U5428 ( .A1(n6636), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6755) );
  INV_X1 U5429 ( .A(n6755), .ZN(n4419) );
  NAND2_X1 U5430 ( .A1(n6278), .A2(n4419), .ZN(n6321) );
  OAI211_X1 U5431 ( .C1(n6294), .C2(n7003), .A(n4420), .B(n6321), .ZN(n4432)
         );
  AND2_X1 U5432 ( .A1(n5223), .A2(n4421), .ZN(n4423) );
  OR2_X1 U5433 ( .A1(n4423), .A2(n4422), .ZN(n6109) );
  INV_X1 U5434 ( .A(n4424), .ZN(n4426) );
  OAI22_X1 U5435 ( .A1(n6334), .A2(n6109), .B1(n4426), .B2(n4425), .ZN(n4431)
         );
  INV_X1 U5436 ( .A(n4427), .ZN(n4429) );
  NOR2_X1 U5437 ( .A1(n4428), .A2(n4429), .ZN(n5622) );
  AOI21_X1 U5438 ( .B1(n4429), .B2(n4428), .A(n5622), .ZN(n5879) );
  INV_X1 U5439 ( .A(n5879), .ZN(n5245) );
  OAI22_X1 U5440 ( .A1(n5245), .A2(n5554), .B1(n5877), .B2(n3104), .ZN(n4430)
         );
  OR3_X1 U5441 ( .A1(n4432), .A2(n4431), .A3(n4430), .ZN(U2819) );
  INV_X1 U5442 ( .A(READY_N), .ZN(n7019) );
  INV_X1 U5443 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4456) );
  INV_X1 U5444 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4448) );
  NOR2_X1 U5445 ( .A1(n4447), .A2(n4448), .ZN(n4443) );
  AND2_X1 U5446 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4449) );
  NAND2_X1 U5447 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4433) );
  OAI21_X1 U5448 ( .B1(n4443), .B2(n4449), .A(n4433), .ZN(n4434) );
  OAI211_X1 U5449 ( .C1(n7019), .C2(n4456), .A(n4434), .B(n4870), .ZN(U3182)
         );
  AOI21_X1 U5450 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n7019), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5451 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4628) );
  INV_X1 U5452 ( .A(n4628), .ZN(n4745) );
  AND2_X1 U5453 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4745), .ZN(n5110) );
  NOR3_X1 U5454 ( .A1(n4436), .A2(n5110), .A3(n4435), .ZN(n4438) );
  OR2_X1 U5455 ( .A1(n4438), .A2(n4437), .ZN(U3150) );
  AOI221_X1 U5456 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7019), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4439) );
  AOI221_X1 U5457 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4439), .C2(HOLD), .A(n4447), .ZN(n4446) );
  AND2_X1 U5458 ( .A1(n4442), .A2(n4447), .ZN(n4441) );
  INV_X1 U5459 ( .A(NA_N), .ZN(n4444) );
  NAND2_X1 U5460 ( .A1(n4444), .A2(STATE_REG_2__SCAN_IN), .ZN(n4440) );
  AND2_X1 U5461 ( .A1(n4441), .A2(n4440), .ZN(n4450) );
  AOI22_X1 U5462 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4454) );
  INV_X1 U5463 ( .A(n4442), .ZN(n4453) );
  AOI21_X1 U5464 ( .B1(n4444), .B2(n4443), .A(n4453), .ZN(n4445) );
  OAI22_X1 U5465 ( .A1(n4446), .A2(n4450), .B1(n4454), .B2(n4445), .ZN(U3183)
         );
  OAI21_X1 U5466 ( .B1(n4449), .B2(n4448), .A(n6750), .ZN(n4452) );
  INV_X1 U5467 ( .A(n4450), .ZN(n4451) );
  OAI211_X1 U5468 ( .C1(n4454), .C2(n4453), .A(n4452), .B(n4451), .ZN(U3181)
         );
  AND2_X1 U5469 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6751), .ZN(n4460) );
  INV_X1 U5470 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5707) );
  INV_X1 U5471 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6905) );
  INV_X1 U5472 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5330) );
  INV_X1 U5473 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U5474 ( .A1(n4455), .A2(n6751), .ZN(n4459) );
  OAI222_X1 U5475 ( .A1(n3100), .A2(n5707), .B1(n6751), .B2(n6905), .C1(n5330), 
        .C2(n4459), .ZN(U3210) );
  INV_X1 U5476 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6902) );
  INV_X1 U5477 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4471) );
  INV_X1 U5478 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U5479 ( .A1(n3100), .A2(n6902), .B1(n4459), .B2(n4471), .C1(n6978), 
        .C2(n6751), .ZN(U3189) );
  INV_X1 U5480 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7045) );
  INV_X1 U5481 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5476) );
  INV_X1 U5482 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6887) );
  OAI222_X1 U5483 ( .A1(n3100), .A2(n7045), .B1(n4459), .B2(n5476), .C1(n6887), 
        .C2(n6751), .ZN(U3199) );
  INV_X1 U5484 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6959) );
  OAI21_X1 U5485 ( .B1(n4456), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4457) );
  INV_X2 U5486 ( .A(n6751), .ZN(n6750) );
  OAI21_X1 U5487 ( .B1(n6751), .B2(n6959), .A(n6737), .ZN(U2789) );
  AOI22_X1 U5488 ( .A1(n4460), .A2(REIP_REG_5__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5489 ( .B1(n6902), .B2(n4459), .A(n4458), .ZN(U3188) );
  INV_X2 U5490 ( .A(n4459), .ZN(n4493) );
  AOI222_X1 U5491 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4493), .B1(n4460), .B2(
        REIP_REG_13__SCAN_IN), .C1(n6750), .C2(ADDRESS_REG_12__SCAN_IN), .ZN(
        n4461) );
  INV_X1 U5492 ( .A(n4461), .ZN(U3196) );
  INV_X1 U5493 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U5494 ( .A1(n4493), .A2(REIP_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6750), .ZN(n4462) );
  OAI21_X1 U5495 ( .B1(n4463), .B2(n3100), .A(n4462), .ZN(U3186) );
  AOI22_X1 U5496 ( .A1(n4493), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6750), .ZN(n4464) );
  OAI21_X1 U5497 ( .B1(n4376), .B2(n3100), .A(n4464), .ZN(U3192) );
  INV_X1 U5498 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4466) );
  AOI22_X1 U5499 ( .A1(n4493), .A2(REIP_REG_25__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n4465) );
  OAI21_X1 U5500 ( .B1(n4466), .B2(n3100), .A(n4465), .ZN(U3207) );
  INV_X1 U5501 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U5502 ( .A1(n4493), .A2(REIP_REG_2__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n4467) );
  OAI21_X1 U5503 ( .B1(n6742), .B2(n3100), .A(n4467), .ZN(U3184) );
  INV_X1 U5504 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6444) );
  AOI22_X1 U5505 ( .A1(n4493), .A2(REIP_REG_3__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U5506 ( .B1(n6444), .B2(n3100), .A(n4468), .ZN(U3185) );
  AOI22_X1 U5507 ( .A1(n4493), .A2(REIP_REG_5__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_3__SCAN_IN), .ZN(n4469) );
  OAI21_X1 U5508 ( .B1(n3100), .B2(n6323), .A(n4469), .ZN(U3187) );
  AOI22_X1 U5509 ( .A1(n4493), .A2(REIP_REG_8__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_6__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5510 ( .B1(n4471), .B2(n3100), .A(n4470), .ZN(U3190) );
  INV_X1 U5511 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U5512 ( .A1(n4493), .A2(REIP_REG_9__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5513 ( .B1(n6890), .B2(n3100), .A(n4472), .ZN(U3191) );
  INV_X1 U5514 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U5515 ( .A1(n4493), .A2(REIP_REG_11__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_9__SCAN_IN), .ZN(n4473) );
  OAI21_X1 U5516 ( .B1(n4474), .B2(n3100), .A(n4473), .ZN(U3193) );
  INV_X1 U5517 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5518 ( .A1(n4493), .A2(REIP_REG_12__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n4475) );
  OAI21_X1 U5519 ( .B1(n4476), .B2(n3100), .A(n4475), .ZN(U3194) );
  INV_X1 U5520 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5838) );
  AOI22_X1 U5521 ( .A1(n4493), .A2(REIP_REG_13__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n4477) );
  OAI21_X1 U5522 ( .B1(n5838), .B2(n3100), .A(n4477), .ZN(U3195) );
  INV_X1 U5523 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5518) );
  AOI22_X1 U5524 ( .A1(n4493), .A2(REIP_REG_15__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_13__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U5525 ( .B1(n5518), .B2(n3100), .A(n4478), .ZN(U3197) );
  INV_X1 U5526 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5504) );
  AOI22_X1 U5527 ( .A1(n4493), .A2(REIP_REG_16__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n4479) );
  OAI21_X1 U5528 ( .B1(n5504), .B2(n3100), .A(n4479), .ZN(U3198) );
  AOI22_X1 U5529 ( .A1(n4493), .A2(REIP_REG_18__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_16__SCAN_IN), .ZN(n4480) );
  OAI21_X1 U5530 ( .B1(n5476), .B2(n3100), .A(n4480), .ZN(U3200) );
  INV_X1 U5531 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5461) );
  AOI22_X1 U5532 ( .A1(n4493), .A2(REIP_REG_19__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5533 ( .B1(n5461), .B2(n3100), .A(n4481), .ZN(U3201) );
  INV_X1 U5534 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6811) );
  AOI22_X1 U5535 ( .A1(n4493), .A2(REIP_REG_20__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n4482) );
  OAI21_X1 U5536 ( .B1(n6811), .B2(n3100), .A(n4482), .ZN(U3202) );
  AOI22_X1 U5537 ( .A1(n4493), .A2(REIP_REG_21__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n4483) );
  OAI21_X1 U5538 ( .B1(n6817), .B2(n3100), .A(n4483), .ZN(U3203) );
  INV_X1 U5539 ( .A(REIP_REG_21__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5540 ( .A1(n4493), .A2(REIP_REG_22__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_20__SCAN_IN), .ZN(n4484) );
  OAI21_X1 U5541 ( .B1(n4485), .B2(n3100), .A(n4484), .ZN(U3204) );
  INV_X1 U5542 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5755) );
  AOI22_X1 U5543 ( .A1(n4493), .A2(REIP_REG_23__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n4486) );
  OAI21_X1 U5544 ( .B1(n5755), .B2(n3100), .A(n4486), .ZN(U3205) );
  INV_X1 U5545 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5388) );
  AOI22_X1 U5546 ( .A1(n4493), .A2(REIP_REG_24__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n4487) );
  OAI21_X1 U5547 ( .B1(n5388), .B2(n3100), .A(n4487), .ZN(U3206) );
  AOI22_X1 U5548 ( .A1(n4493), .A2(REIP_REG_30__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U5549 ( .B1(n4489), .B2(n3100), .A(n4488), .ZN(U3212) );
  INV_X1 U5550 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5368) );
  AOI22_X1 U5551 ( .A1(n4493), .A2(REIP_REG_26__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_24__SCAN_IN), .ZN(n4490) );
  OAI21_X1 U5552 ( .B1(n5368), .B2(n3100), .A(n4490), .ZN(U3208) );
  INV_X1 U5553 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6934) );
  AOI22_X1 U5554 ( .A1(n4493), .A2(REIP_REG_27__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_25__SCAN_IN), .ZN(n4491) );
  OAI21_X1 U5555 ( .B1(n6934), .B2(n3100), .A(n4491), .ZN(U3209) );
  AOI22_X1 U5556 ( .A1(n4493), .A2(REIP_REG_29__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_27__SCAN_IN), .ZN(n4492) );
  OAI21_X1 U5557 ( .B1(n5330), .B2(n3100), .A(n4492), .ZN(U3211) );
  INV_X1 U5558 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5559 ( .A1(n4493), .A2(REIP_REG_31__SCAN_IN), .B1(n6750), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U5560 ( .B1(n4495), .B2(n3100), .A(n4494), .ZN(U3213) );
  INV_X1 U5561 ( .A(n4496), .ZN(n4498) );
  INV_X1 U5562 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6856) );
  OAI211_X1 U5563 ( .C1(n4498), .C2(n6856), .A(n4497), .B(n6755), .ZN(U2788)
         );
  AOI22_X1 U5564 ( .A1(n4876), .A2(n4871), .B1(n4874), .B2(n4499), .ZN(n4873)
         );
  INV_X1 U5565 ( .A(n4873), .ZN(n4500) );
  OAI21_X1 U5566 ( .B1(n4500), .B2(n5114), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4501) );
  OAI21_X1 U5567 ( .B1(n6755), .B2(n5282), .A(n4501), .ZN(U2790) );
  OR2_X1 U5568 ( .A1(n4874), .A2(n3502), .ZN(n4574) );
  NAND2_X1 U5569 ( .A1(n4574), .A2(n4870), .ZN(n4503) );
  OAI211_X1 U5570 ( .C1(n5261), .C2(n4578), .A(n7019), .B(n4503), .ZN(n4504)
         );
  MUX2_X1 U5571 ( .A(n4504), .B(n4878), .S(n4876), .Z(n4514) );
  INV_X1 U5572 ( .A(n4876), .ZN(n4512) );
  INV_X1 U5573 ( .A(n4573), .ZN(n4511) );
  INV_X1 U5574 ( .A(n4562), .ZN(n4509) );
  NAND2_X1 U5575 ( .A1(n4506), .A2(n4505), .ZN(n4523) );
  OR2_X1 U5576 ( .A1(n4507), .A2(n4523), .ZN(n4508) );
  NAND2_X1 U5577 ( .A1(n4508), .A2(n4880), .ZN(n4564) );
  OR2_X1 U5578 ( .A1(n5555), .A2(n3519), .ZN(n4525) );
  OAI211_X1 U5579 ( .C1(n4736), .C2(n4509), .A(n4564), .B(n4525), .ZN(n4510)
         );
  AOI21_X1 U5580 ( .B1(n4512), .B2(n4511), .A(n4510), .ZN(n4513) );
  NAND2_X1 U5581 ( .A1(n4514), .A2(n4513), .ZN(n4860) );
  AND2_X1 U5582 ( .A1(n5110), .A2(FLUSH_REG_SCAN_IN), .ZN(n4515) );
  AOI21_X1 U5583 ( .B1(n4860), .B2(n6729), .A(n4515), .ZN(n4520) );
  AND2_X1 U5584 ( .A1(n5282), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4632) );
  INV_X1 U5585 ( .A(n4632), .ZN(n4892) );
  INV_X1 U5586 ( .A(n6129), .ZN(n4521) );
  INV_X1 U5587 ( .A(n5075), .ZN(n6189) );
  NOR2_X1 U5588 ( .A1(n4516), .A2(n6189), .ZN(n4517) );
  XNOR2_X1 U5589 ( .A(n4517), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4737)
         );
  INV_X1 U5590 ( .A(n4737), .ZN(n6317) );
  NAND3_X1 U5591 ( .A1(n6317), .A2(n4518), .A3(n6123), .ZN(n4519) );
  OAI22_X1 U5592 ( .A1(n4521), .A2(n4113), .B1(n4520), .B2(n4519), .ZN(U3455)
         );
  INV_X1 U5593 ( .A(n5582), .ZN(n5003) );
  INV_X1 U5594 ( .A(n4523), .ZN(n4531) );
  NAND2_X1 U5595 ( .A1(n3508), .A2(n5439), .ZN(n4528) );
  NAND2_X1 U5596 ( .A1(n5297), .A2(n4524), .ZN(n4527) );
  NAND2_X1 U5597 ( .A1(n3519), .A2(n4617), .ZN(n4526) );
  AND4_X1 U5598 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4530)
         );
  AND4_X1 U5599 ( .A1(n4532), .A2(n4531), .A3(n4530), .A4(n4529), .ZN(n4584)
         );
  INV_X1 U5600 ( .A(n4533), .ZN(n4534) );
  NOR2_X1 U5601 ( .A1(n4578), .A2(n4534), .ZN(n4535) );
  AND2_X1 U5602 ( .A1(n4736), .A2(n4535), .ZN(n4536) );
  NAND2_X1 U5603 ( .A1(n4584), .A2(n4536), .ZN(n4854) );
  INV_X1 U5604 ( .A(n4854), .ZN(n4540) );
  NAND2_X1 U5605 ( .A1(n5261), .A2(n3263), .ZN(n4544) );
  INV_X1 U5606 ( .A(n4852), .ZN(n4561) );
  INV_X1 U5607 ( .A(n4537), .ZN(n4719) );
  INV_X1 U5608 ( .A(n4538), .ZN(n4742) );
  NAND3_X1 U5609 ( .A1(n4561), .A2(n4719), .A3(n4742), .ZN(n4539) );
  OAI211_X1 U5610 ( .C1(n5003), .C2(n4540), .A(n4544), .B(n4539), .ZN(n4859)
         );
  INV_X1 U5611 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5922) );
  INV_X1 U5612 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5613 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5922), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4591), .ZN(n4552) );
  INV_X1 U5614 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6464) );
  NOR2_X1 U5615 ( .A1(n5263), .A2(n6464), .ZN(n4550) );
  INV_X1 U5616 ( .A(n5267), .ZN(n6124) );
  NOR2_X1 U5617 ( .A1(n6124), .A2(n4537), .ZN(n4555) );
  AOI222_X1 U5618 ( .A1(n4859), .A2(n6123), .B1(n4552), .B2(n4550), .C1(n4742), 
        .C2(n4555), .ZN(n4542) );
  NAND2_X1 U5619 ( .A1(n6129), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4541) );
  OAI21_X1 U5620 ( .B1(n4542), .B2(n6129), .A(n4541), .ZN(U3460) );
  XNOR2_X1 U5621 ( .A(n4537), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4548)
         );
  NAND2_X1 U5622 ( .A1(n5261), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4545) );
  MUX2_X1 U5623 ( .A(n4545), .B(n4544), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4547) );
  NAND2_X1 U5624 ( .A1(n4573), .A2(n4878), .ZN(n4722) );
  NAND2_X1 U5625 ( .A1(n4722), .A2(n4548), .ZN(n4546) );
  OAI211_X1 U5626 ( .C1(n4726), .C2(n4548), .A(n4547), .B(n4546), .ZN(n4549)
         );
  AOI21_X1 U5627 ( .B1(n5577), .B2(n4854), .A(n4549), .ZN(n4732) );
  INV_X1 U5628 ( .A(n4732), .ZN(n4554) );
  INV_X1 U5629 ( .A(n4550), .ZN(n5265) );
  NAND3_X1 U5630 ( .A1(n5267), .A2(n4537), .A3(n4733), .ZN(n4551) );
  OAI21_X1 U5631 ( .B1(n5265), .B2(n4552), .A(n4551), .ZN(n4553) );
  AOI21_X1 U5632 ( .B1(n6123), .B2(n4554), .A(n4553), .ZN(n4557) );
  OAI21_X1 U5633 ( .B1(n6129), .B2(n4555), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4556) );
  OAI21_X1 U5634 ( .B1(n6129), .B2(n4557), .A(n4556), .ZN(U3459) );
  OAI21_X1 U5635 ( .B1(n4560), .B2(n4559), .A(n4558), .ZN(n6412) );
  NAND3_X1 U5636 ( .A1(n4876), .A2(n4561), .A3(n4684), .ZN(n4565) );
  INV_X1 U5637 ( .A(n4870), .ZN(n4597) );
  OAI211_X1 U5638 ( .C1(n3502), .C2(n4597), .A(n3519), .B(n4562), .ZN(n4563)
         );
  NAND3_X1 U5639 ( .A1(n4565), .A2(n4564), .A3(n4563), .ZN(n4566) );
  NAND2_X1 U5640 ( .A1(n4566), .A2(n6729), .ZN(n4572) );
  NAND3_X1 U5641 ( .A1(n4578), .A2(n4567), .A3(n7019), .ZN(n4568) );
  NAND3_X1 U5642 ( .A1(n4568), .A2(n3554), .A3(n4617), .ZN(n4569) );
  NAND2_X1 U5643 ( .A1(n4569), .A2(n4703), .ZN(n4570) );
  NAND2_X2 U5644 ( .A1(n4572), .A2(n4571), .ZN(n4589) );
  AND2_X1 U5645 ( .A1(n4573), .A2(n4869), .ZN(n4875) );
  OAI211_X1 U5646 ( .C1(n4697), .C2(n4580), .A(n4574), .B(n4736), .ZN(n4575)
         );
  INV_X1 U5647 ( .A(n4575), .ZN(n4576) );
  NAND2_X1 U5648 ( .A1(n4875), .A2(n4576), .ZN(n4577) );
  NAND2_X1 U5649 ( .A1(n4578), .A2(n5280), .ZN(n4851) );
  OAI21_X1 U5650 ( .B1(n4580), .B2(n4579), .A(n4851), .ZN(n4581) );
  OAI21_X1 U5651 ( .B1(n4582), .B2(n6752), .A(n4583), .ZN(n4610) );
  NOR2_X1 U5652 ( .A1(n6443), .A2(n6742), .ZN(n6409) );
  OR2_X1 U5653 ( .A1(n4589), .A2(n6399), .ZN(n6462) );
  NAND2_X1 U5654 ( .A1(n4584), .A2(n4726), .ZN(n4585) );
  NAND2_X1 U5655 ( .A1(n4589), .A2(n4585), .ZN(n6069) );
  INV_X1 U5656 ( .A(n4878), .ZN(n4586) );
  NAND2_X1 U5657 ( .A1(n6069), .A2(n6440), .ZN(n4587) );
  NAND2_X1 U5658 ( .A1(n6464), .A2(n4587), .ZN(n6453) );
  AOI21_X1 U5659 ( .B1(n6462), .B2(n6453), .A(n4591), .ZN(n4588) );
  AOI211_X1 U5660 ( .C1(n6432), .C2(n4610), .A(n6409), .B(n4588), .ZN(n4593)
         );
  NAND2_X1 U5661 ( .A1(n4589), .A2(n5261), .ZN(n6463) );
  INV_X1 U5662 ( .A(n6440), .ZN(n4590) );
  NAND2_X1 U5663 ( .A1(n6463), .A2(n6464), .ZN(n4657) );
  NAND3_X1 U5664 ( .A1(n6420), .A2(n4591), .A3(n4657), .ZN(n4592) );
  OAI211_X1 U5665 ( .C1(n6412), .C2(n6422), .A(n4593), .B(n4592), .ZN(U3017)
         );
  INV_X1 U5666 ( .A(n5261), .ZN(n4594) );
  AOI22_X1 U5667 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6376), .B1(n6380), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4599) );
  OAI21_X1 U5668 ( .B1(n3867), .B2(n6343), .A(n4599), .ZN(U2907) );
  INV_X1 U5669 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5670 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6376), .B1(n6380), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4600) );
  OAI21_X1 U5671 ( .B1(n4601), .B2(n6343), .A(n4600), .ZN(U2903) );
  INV_X1 U5672 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6853) );
  AOI22_X1 U5673 ( .A1(n6376), .A2(UWORD_REG_2__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4602) );
  OAI21_X1 U5674 ( .B1(n6853), .B2(n6343), .A(n4602), .ZN(U2905) );
  AOI22_X1 U5675 ( .A1(n6374), .A2(UWORD_REG_9__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4603) );
  OAI21_X1 U5676 ( .B1(n4028), .B2(n6343), .A(n4603), .ZN(U2898) );
  INV_X1 U5677 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7013) );
  AOI22_X1 U5678 ( .A1(n6376), .A2(UWORD_REG_5__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4604) );
  OAI21_X1 U5679 ( .B1(n7013), .B2(n6343), .A(n4604), .ZN(U2902) );
  OAI21_X1 U5680 ( .B1(n5297), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4605), 
        .ZN(n6454) );
  INV_X1 U5681 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U5682 ( .A(n4607), .B(n4606), .ZN(n5881) );
  OAI222_X1 U5683 ( .A1(n6454), .A2(n7065), .B1(n5628), .B2(n5591), .C1(n7064), 
        .C2(n5881), .ZN(U2859) );
  OAI21_X1 U5684 ( .B1(n4609), .B2(n4608), .A(n4614), .ZN(n6411) );
  AOI22_X1 U5685 ( .A1(n4234), .A2(n4610), .B1(n5607), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4611) );
  OAI21_X1 U5686 ( .B1(n6411), .B2(n7064), .A(n4611), .ZN(U2858) );
  AND3_X1 U5687 ( .A1(n4615), .A2(n4614), .A3(n4613), .ZN(n4616) );
  NOR2_X1 U5688 ( .A1(n4612), .A2(n4616), .ZN(n6405) );
  INV_X1 U5689 ( .A(n6405), .ZN(n4621) );
  AND2_X1 U5690 ( .A1(n4075), .A2(n4693), .ZN(n4620) );
  INV_X1 U5691 ( .A(n4620), .ZN(n4618) );
  AND2_X1 U5692 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  INV_X1 U5693 ( .A(DATAI_2_), .ZN(n4701) );
  INV_X1 U5694 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6946) );
  OAI222_X1 U5695 ( .A1(n4621), .A2(n5683), .B1(n5072), .B2(n4701), .C1(n5070), 
        .C2(n6946), .ZN(U2889) );
  INV_X1 U5696 ( .A(DATAI_1_), .ZN(n7025) );
  INV_X1 U5697 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6379) );
  OAI222_X1 U5698 ( .A1(n6411), .A2(n5683), .B1(n5072), .B2(n7025), .C1(n5070), 
        .C2(n6379), .ZN(U2890) );
  NOR2_X1 U5699 ( .A1(n3683), .A2(n4622), .ZN(n4623) );
  AOI21_X1 U5700 ( .B1(n4634), .B2(STATEBS16_REG_SCAN_IN), .A(n6636), .ZN(
        n4639) );
  NAND2_X1 U5701 ( .A1(n5577), .A2(n5003), .ZN(n6486) );
  NOR2_X1 U5702 ( .A1(n6486), .A2(n5075), .ZN(n6495) );
  NOR2_X1 U5703 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4626) );
  AND2_X1 U5704 ( .A1(n4626), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6488)
         );
  NAND2_X1 U5705 ( .A1(n6488), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4636) );
  INV_X1 U5706 ( .A(n4636), .ZN(n4987) );
  AOI21_X1 U5707 ( .B1(n6495), .B2(n3114), .A(n4987), .ZN(n4638) );
  INV_X1 U5708 ( .A(n4638), .ZN(n4627) );
  AOI22_X1 U5709 ( .A1(n4639), .A2(n4627), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6488), .ZN(n4962) );
  INV_X1 U5710 ( .A(DATAI_0_), .ZN(n4647) );
  INV_X2 U5711 ( .A(n5873), .ZN(n6404) );
  NAND2_X1 U5712 ( .A1(n6404), .A2(DATAI_24_), .ZN(n6624) );
  INV_X1 U5713 ( .A(n6624), .ZN(n6715) );
  INV_X1 U5714 ( .A(n4634), .ZN(n4629) );
  INV_X1 U5715 ( .A(n4630), .ZN(n4631) );
  OR2_X1 U5716 ( .A1(n4633), .A2(n4702), .ZN(n6623) );
  NAND2_X1 U5717 ( .A1(n6404), .A2(DATAI_16_), .ZN(n6642) );
  INV_X1 U5718 ( .A(n6642), .ZN(n6714) );
  NAND2_X1 U5719 ( .A1(n6534), .A2(n6714), .ZN(n4635) );
  OAI21_X1 U5720 ( .B1(n4636), .B2(n6623), .A(n4635), .ZN(n4637) );
  AOI21_X1 U5721 ( .B1(n6715), .B2(n6513), .A(n4637), .ZN(n4642) );
  NAND2_X1 U5722 ( .A1(n4639), .A2(n4638), .ZN(n4640) );
  INV_X1 U5723 ( .A(n6634), .ZN(n6543) );
  OAI211_X1 U5724 ( .C1(n6626), .C2(n6488), .A(n4640), .B(n6543), .ZN(n4961)
         );
  NAND2_X1 U5725 ( .A1(n4961), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4641) );
  OAI211_X1 U5726 ( .C1(n4962), .C2(n6199), .A(n4642), .B(n4641), .ZN(U3060)
         );
  INV_X1 U5727 ( .A(n4643), .ZN(n4646) );
  INV_X1 U5728 ( .A(n4612), .ZN(n4645) );
  NAND2_X1 U5729 ( .A1(n4612), .A2(n4643), .ZN(n4756) );
  INV_X1 U5730 ( .A(n4756), .ZN(n4644) );
  AOI21_X1 U5731 ( .B1(n4646), .B2(n4645), .A(n4644), .ZN(n4714) );
  INV_X1 U5732 ( .A(n4714), .ZN(n5571) );
  INV_X1 U5733 ( .A(DATAI_3_), .ZN(n4665) );
  INV_X1 U5734 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6373) );
  OAI222_X1 U5735 ( .A1(n5571), .A2(n5683), .B1(n5072), .B2(n4665), .C1(n5070), 
        .C2(n6373), .ZN(U2888) );
  INV_X1 U5736 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6974) );
  OAI222_X1 U5737 ( .A1(n5683), .A2(n5881), .B1(n5070), .B2(n6974), .C1(n4647), 
        .C2(n5072), .ZN(U2891) );
  XNOR2_X1 U5738 ( .A(n4649), .B(n4648), .ZN(n4716) );
  INV_X1 U5739 ( .A(n5573), .ZN(n4653) );
  INV_X1 U5740 ( .A(n4651), .ZN(n4652) );
  OAI21_X1 U5741 ( .B1(n4650), .B2(n4653), .A(n4652), .ZN(n4654) );
  NAND2_X1 U5742 ( .A1(n4654), .A2(n4759), .ZN(n5560) );
  AOI21_X1 U5743 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5252) );
  INV_X1 U5744 ( .A(n5252), .ZN(n6442) );
  NAND2_X1 U5745 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4656) );
  OR2_X1 U5746 ( .A1(n6069), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4655)
         );
  NAND2_X1 U5747 ( .A1(n4655), .A2(n6462), .ZN(n5908) );
  AOI21_X1 U5748 ( .B1(n5903), .B2(n4656), .A(n5908), .ZN(n6450) );
  OAI21_X1 U5749 ( .B1(n6440), .B2(n6442), .A(n6450), .ZN(n5100) );
  NAND2_X1 U5750 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5910), .ZN(n6451)
         );
  OAI22_X1 U5751 ( .A1(n5252), .A2(n6440), .B1(n4143), .B2(n6451), .ZN(n5235)
         );
  AOI22_X1 U5752 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n5100), .B1(n5235), 
        .B2(n4264), .ZN(n4658) );
  NAND2_X1 U5753 ( .A1(n6399), .A2(REIP_REG_3__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5754 ( .C1(n6455), .C2(n5560), .A(n4658), .B(n4710), .ZN(n4659)
         );
  INV_X1 U5755 ( .A(n4659), .ZN(n4660) );
  OAI21_X1 U5756 ( .B1(n4716), .B2(n6422), .A(n4660), .ZN(U3015) );
  NOR2_X1 U5757 ( .A1(n3102), .A2(n4765), .ZN(n4663) );
  NAND2_X1 U5758 ( .A1(n4667), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5759 ( .A1(n6141), .A2(n3114), .ZN(n5162) );
  AND3_X1 U5760 ( .A1(n4858), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U5761 ( .A1(n6194), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4704) );
  OAI21_X1 U5762 ( .B1(n5162), .B2(n6486), .A(n4704), .ZN(n4673) );
  NOR2_X2 U5763 ( .A1(n4665), .A2(n6192), .ZN(n6660) );
  INV_X1 U5764 ( .A(n6660), .ZN(n6211) );
  NAND2_X1 U5765 ( .A1(n6404), .A2(DATAI_27_), .ZN(n6658) );
  INV_X1 U5766 ( .A(n6658), .ZN(n6527) );
  NAND2_X1 U5767 ( .A1(n6404), .A2(DATAI_19_), .ZN(n6663) );
  NAND2_X1 U5768 ( .A1(n4668), .A2(n4692), .ZN(n6657) );
  OAI22_X1 U5769 ( .A1(n5027), .A2(n6663), .B1(n6657), .B2(n4704), .ZN(n4669)
         );
  AOI21_X1 U5770 ( .B1(n6527), .B2(n6703), .A(n4669), .ZN(n4676) );
  INV_X1 U5771 ( .A(n4670), .ZN(n4674) );
  INV_X1 U5772 ( .A(n6194), .ZN(n4671) );
  AOI21_X1 U5773 ( .B1(n4671), .B2(n6636), .A(n6634), .ZN(n4672) );
  NAND2_X1 U5774 ( .A1(n4706), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4675)
         );
  OAI211_X1 U5775 ( .C1(n4709), .C2(n6211), .A(n4676), .B(n4675), .ZN(U3127)
         );
  OAI22_X1 U5776 ( .A1(n5027), .A2(n6642), .B1(n6623), .B2(n4704), .ZN(n4677)
         );
  AOI21_X1 U5777 ( .B1(n6715), .B2(n6703), .A(n4677), .ZN(n4679) );
  NAND2_X1 U5778 ( .A1(n4706), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4678)
         );
  OAI211_X1 U5779 ( .C1(n4709), .C2(n6199), .A(n4679), .B(n4678), .ZN(U3124)
         );
  INV_X1 U5780 ( .A(DATAI_6_), .ZN(n5071) );
  NOR2_X2 U5781 ( .A1(n5071), .A2(n6192), .ZN(n6694) );
  NAND2_X1 U5782 ( .A1(n6404), .A2(DATAI_30_), .ZN(n6698) );
  INV_X1 U5783 ( .A(n6698), .ZN(n5089) );
  NAND2_X1 U5784 ( .A1(n6404), .A2(DATAI_22_), .ZN(n6678) );
  NAND2_X1 U5785 ( .A1(n4680), .A2(n4692), .ZN(n6677) );
  OAI22_X1 U5786 ( .A1(n5027), .A2(n6678), .B1(n6677), .B2(n4704), .ZN(n4681)
         );
  AOI21_X1 U5787 ( .B1(n5089), .B2(n6703), .A(n4681), .ZN(n4683) );
  NAND2_X1 U5788 ( .A1(n4706), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4682)
         );
  OAI211_X1 U5789 ( .C1(n4709), .C2(n5192), .A(n4683), .B(n4682), .ZN(U3130)
         );
  NOR2_X2 U5790 ( .A1(n7025), .A2(n6192), .ZN(n6646) );
  INV_X1 U5791 ( .A(n6646), .ZN(n6203) );
  NAND2_X1 U5792 ( .A1(n6404), .A2(DATAI_25_), .ZN(n6644) );
  INV_X1 U5793 ( .A(n6644), .ZN(n6521) );
  NAND2_X1 U5794 ( .A1(n6404), .A2(DATAI_17_), .ZN(n6649) );
  NAND2_X1 U5795 ( .A1(n4684), .A2(n4692), .ZN(n6643) );
  OAI22_X1 U5796 ( .A1(n5027), .A2(n6649), .B1(n6643), .B2(n4704), .ZN(n4685)
         );
  AOI21_X1 U5797 ( .B1(n6521), .B2(n6703), .A(n4685), .ZN(n4687) );
  NAND2_X1 U5798 ( .A1(n4706), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4686)
         );
  OAI211_X1 U5799 ( .C1(n4709), .C2(n6203), .A(n4687), .B(n4686), .ZN(U3125)
         );
  INV_X1 U5800 ( .A(DATAI_5_), .ZN(n5000) );
  NAND2_X1 U5801 ( .A1(n6404), .A2(DATAI_29_), .ZN(n6676) );
  INV_X1 U5802 ( .A(n6676), .ZN(n6535) );
  NAND2_X1 U5803 ( .A1(n6404), .A2(DATAI_21_), .ZN(n6671) );
  NAND2_X1 U5804 ( .A1(n4688), .A2(n4692), .ZN(n6670) );
  OAI22_X1 U5805 ( .A1(n5027), .A2(n6671), .B1(n6670), .B2(n4704), .ZN(n4689)
         );
  AOI21_X1 U5806 ( .B1(n6535), .B2(n6703), .A(n4689), .ZN(n4691) );
  NAND2_X1 U5807 ( .A1(n4706), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4690)
         );
  OAI211_X1 U5808 ( .C1(n4709), .C2(n6219), .A(n4691), .B(n4690), .ZN(U3129)
         );
  INV_X1 U5809 ( .A(DATAI_7_), .ZN(n6906) );
  NOR2_X2 U5810 ( .A1(n6906), .A2(n6192), .ZN(n6701) );
  INV_X1 U5811 ( .A(n6701), .ZN(n5175) );
  NAND2_X1 U5812 ( .A1(n6404), .A2(DATAI_31_), .ZN(n6709) );
  INV_X1 U5813 ( .A(n6709), .ZN(n6477) );
  NAND2_X1 U5814 ( .A1(n6404), .A2(DATAI_23_), .ZN(n6684) );
  NAND2_X1 U5815 ( .A1(n4693), .A2(n4692), .ZN(n6683) );
  OAI22_X1 U5816 ( .A1(n5027), .A2(n6684), .B1(n6683), .B2(n4704), .ZN(n4694)
         );
  AOI21_X1 U5817 ( .B1(n6477), .B2(n6703), .A(n4694), .ZN(n4696) );
  NAND2_X1 U5818 ( .A1(n4706), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4695)
         );
  OAI211_X1 U5819 ( .C1(n4709), .C2(n5175), .A(n4696), .B(n4695), .ZN(U3131)
         );
  INV_X1 U5820 ( .A(DATAI_4_), .ZN(n7028) );
  NOR2_X2 U5821 ( .A1(n7028), .A2(n6192), .ZN(n6720) );
  INV_X1 U5822 ( .A(n6720), .ZN(n6215) );
  NAND2_X1 U5823 ( .A1(n6404), .A2(DATAI_28_), .ZN(n6669) );
  INV_X1 U5824 ( .A(n6669), .ZN(n6724) );
  NAND2_X1 U5825 ( .A1(n6404), .A2(DATAI_20_), .ZN(n6665) );
  OR2_X1 U5826 ( .A1(n4697), .A2(n4702), .ZN(n6664) );
  OAI22_X1 U5827 ( .A1(n5027), .A2(n6665), .B1(n6664), .B2(n4704), .ZN(n4698)
         );
  AOI21_X1 U5828 ( .B1(n6724), .B2(n6703), .A(n4698), .ZN(n4700) );
  NAND2_X1 U5829 ( .A1(n4706), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4699)
         );
  OAI211_X1 U5830 ( .C1(n4709), .C2(n6215), .A(n4700), .B(n4699), .ZN(U3128)
         );
  NOR2_X2 U5831 ( .A1(n4701), .A2(n6192), .ZN(n6653) );
  INV_X1 U5832 ( .A(n6653), .ZN(n6207) );
  NAND2_X1 U5833 ( .A1(n6404), .A2(DATAI_26_), .ZN(n6656) );
  INV_X1 U5834 ( .A(n6656), .ZN(n6524) );
  NAND2_X1 U5835 ( .A1(n6404), .A2(DATAI_18_), .ZN(n6651) );
  OR2_X1 U5836 ( .A1(n4703), .A2(n4702), .ZN(n6650) );
  OAI22_X1 U5837 ( .A1(n5027), .A2(n6651), .B1(n6650), .B2(n4704), .ZN(n4705)
         );
  AOI21_X1 U5838 ( .B1(n6524), .B2(n6703), .A(n4705), .ZN(n4708) );
  NAND2_X1 U5839 ( .A1(n4706), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4707)
         );
  OAI211_X1 U5840 ( .C1(n4709), .C2(n6207), .A(n4708), .B(n4707), .ZN(U3126)
         );
  NOR2_X1 U5841 ( .A1(n6418), .A2(n5559), .ZN(n4713) );
  OAI21_X1 U5842 ( .B1(n5868), .B2(n4711), .A(n4710), .ZN(n4712) );
  AOI211_X1 U5843 ( .C1(n4714), .C2(n6404), .A(n4713), .B(n4712), .ZN(n4715)
         );
  OAI21_X1 U5844 ( .B1(n4716), .B2(n6226), .A(n4715), .ZN(U2983) );
  OAI222_X1 U5845 ( .A1(n5560), .A2(n7065), .B1(n3205), .B2(n5628), .C1(n5571), 
        .C2(n7064), .ZN(U2856) );
  NOR2_X1 U5846 ( .A1(FLUSH_REG_SCAN_IN), .A2(n5263), .ZN(n4739) );
  AOI21_X1 U5847 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4721) );
  NAND3_X1 U5848 ( .A1(n4722), .A2(n4721), .A3(n4720), .ZN(n4730) );
  NAND2_X1 U5849 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4723) );
  INV_X1 U5850 ( .A(n4723), .ZN(n4724) );
  MUX2_X1 U5851 ( .A(n4724), .B(n4723), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4728) );
  OAI21_X1 U5852 ( .B1(n3544), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4725), 
        .ZN(n6125) );
  NOR2_X1 U5853 ( .A1(n4726), .A2(n6125), .ZN(n4727) );
  AOI21_X1 U5854 ( .B1(n5261), .B2(n4728), .A(n4727), .ZN(n4729) );
  NAND2_X1 U5855 ( .A1(n4730), .A2(n4729), .ZN(n4731) );
  AOI21_X1 U5856 ( .B1(n6141), .B2(n4854), .A(n4731), .ZN(n6127) );
  MUX2_X1 U5857 ( .A(n6128), .B(n6127), .S(n4860), .Z(n4868) );
  MUX2_X1 U5858 ( .A(n4733), .B(n4732), .S(n4860), .Z(n4863) );
  NOR3_X1 U5859 ( .A1(n4868), .A2(n4863), .A3(STATE2_REG_1__SCAN_IN), .ZN(
        n4734) );
  AOI21_X1 U5860 ( .B1(n4717), .B2(n4739), .A(n4734), .ZN(n4735) );
  INV_X1 U5861 ( .A(n4735), .ZN(n4885) );
  OAI22_X1 U5862 ( .A1(n4737), .A2(n4736), .B1(n4860), .B2(n4113), .ZN(n4738)
         );
  NAND2_X1 U5863 ( .A1(n4738), .A2(n5263), .ZN(n4741) );
  NAND2_X1 U5864 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4739), .ZN(n4740) );
  NAND2_X1 U5865 ( .A1(n4741), .A2(n4740), .ZN(n4884) );
  AOI21_X1 U5866 ( .B1(n4885), .B2(n4742), .A(n4884), .ZN(n5111) );
  INV_X1 U5867 ( .A(n5111), .ZN(n4743) );
  OAI21_X1 U5868 ( .B1(n4743), .B2(FLUSH_REG_SCAN_IN), .A(n5110), .ZN(n4744)
         );
  NAND2_X1 U5869 ( .A1(n4744), .A2(n6192), .ZN(n6465) );
  NAND2_X1 U5870 ( .A1(n4338), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6115) );
  AOI222_X1 U5871 ( .A1(n4745), .A2(n5111), .B1(n5164), .B2(n6626), .C1(n3114), 
        .C2(n6115), .ZN(n4747) );
  NAND2_X1 U5872 ( .A1(n4754), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4746) );
  OAI21_X1 U5873 ( .B1(n4754), .B2(n4747), .A(n4746), .ZN(U3465) );
  INV_X1 U5874 ( .A(n3102), .ZN(n4894) );
  AOI211_X1 U5875 ( .C1(n4894), .C2(n6225), .A(n6636), .B(n6116), .ZN(n4748)
         );
  AOI21_X1 U5876 ( .B1(n5582), .B2(n6115), .A(n4748), .ZN(n4750) );
  NAND2_X1 U5877 ( .A1(n4754), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5878 ( .B1(n4754), .B2(n4750), .A(n4749), .ZN(U3464) );
  XNOR2_X1 U5879 ( .A(n6116), .B(n5010), .ZN(n4751) );
  AOI22_X1 U5880 ( .A1(n4751), .A2(n6626), .B1(n6115), .B2(n5577), .ZN(n4753)
         );
  NAND2_X1 U5881 ( .A1(n4754), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4752) );
  OAI21_X1 U5882 ( .B1(n4754), .B2(n4753), .A(n4752), .ZN(U3463) );
  INV_X1 U5883 ( .A(n4755), .ZN(n4757) );
  NOR2_X1 U5884 ( .A1(n4756), .A2(n4757), .ZN(n4996) );
  AOI21_X1 U5885 ( .B1(n4757), .B2(n4756), .A(n4996), .ZN(n4844) );
  INV_X1 U5886 ( .A(n4844), .ZN(n6327) );
  AND2_X1 U5887 ( .A1(n4759), .A2(n4758), .ZN(n4761) );
  OR2_X1 U5888 ( .A1(n4761), .A2(n4760), .ZN(n6333) );
  INV_X1 U5889 ( .A(n6333), .ZN(n4762) );
  AOI22_X1 U5890 ( .A1(n4234), .A2(n4762), .B1(n5607), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4763) );
  OAI21_X1 U5891 ( .B1(n6327), .B2(n7064), .A(n4763), .ZN(U2855) );
  INV_X1 U5892 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4764) );
  OAI222_X1 U5893 ( .A1(n6327), .A2(n5683), .B1(n5072), .B2(n7028), .C1(n5070), 
        .C2(n4764), .ZN(U2887) );
  NAND2_X1 U5894 ( .A1(n3102), .A2(n5163), .ZN(n6138) );
  NOR2_X1 U5895 ( .A1(n6138), .A2(n4765), .ZN(n4766) );
  NAND3_X1 U5896 ( .A1(n4662), .A2(n4770), .A3(n3102), .ZN(n4767) );
  OR2_X1 U5897 ( .A1(n6636), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6121) );
  INV_X1 U5898 ( .A(n6121), .ZN(n6489) );
  AOI21_X1 U5899 ( .B1(n4767), .B2(n6404), .A(n6489), .ZN(n4768) );
  NAND2_X1 U5900 ( .A1(n5577), .A2(n5582), .ZN(n5076) );
  OAI21_X1 U5901 ( .B1(n5162), .B2(n5076), .A(n6710), .ZN(n4771) );
  NOR2_X1 U5902 ( .A1(n4768), .A2(n4771), .ZN(n4769) );
  AOI211_X1 U5903 ( .C1(n5022), .C2(n6636), .A(n6634), .B(n4769), .ZN(n6728)
         );
  INV_X1 U5904 ( .A(n6728), .ZN(n4795) );
  NAND2_X1 U5905 ( .A1(n4795), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4778)
         );
  NAND3_X1 U5906 ( .A1(n6539), .A2(n4662), .A3(n4770), .ZN(n4897) );
  INV_X1 U5907 ( .A(n6651), .ZN(n6600) );
  NAND2_X1 U5908 ( .A1(n4771), .A2(n6626), .ZN(n4774) );
  NAND2_X1 U5909 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4772), .ZN(n4773) );
  NAND2_X1 U5910 ( .A1(n4774), .A2(n4773), .ZN(n6721) );
  NAND2_X1 U5911 ( .A1(n6721), .A2(n6653), .ZN(n4775) );
  OAI21_X1 U5912 ( .B1(n6650), .B2(n6710), .A(n4775), .ZN(n4776) );
  AOI21_X1 U5913 ( .B1(n6723), .B2(n6600), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5914 ( .C1(n6713), .C2(n6656), .A(n4778), .B(n4777), .ZN(U3142)
         );
  NAND2_X1 U5915 ( .A1(n4795), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4782)
         );
  INV_X1 U5916 ( .A(n6649), .ZN(n6596) );
  NAND2_X1 U5917 ( .A1(n6721), .A2(n6646), .ZN(n4779) );
  OAI21_X1 U5918 ( .B1(n6643), .B2(n6710), .A(n4779), .ZN(n4780) );
  AOI21_X1 U5919 ( .B1(n6723), .B2(n6596), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5920 ( .C1(n6713), .C2(n6644), .A(n4782), .B(n4781), .ZN(U3141)
         );
  NAND2_X1 U5921 ( .A1(n4795), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4786)
         );
  INV_X1 U5922 ( .A(n6678), .ZN(n6695) );
  NAND2_X1 U5923 ( .A1(n6721), .A2(n6694), .ZN(n4783) );
  OAI21_X1 U5924 ( .B1(n6677), .B2(n6710), .A(n4783), .ZN(n4784) );
  AOI21_X1 U5925 ( .B1(n6723), .B2(n6695), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5926 ( .C1(n6713), .C2(n6698), .A(n4786), .B(n4785), .ZN(U3146)
         );
  NAND2_X1 U5927 ( .A1(n4795), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4790)
         );
  INV_X1 U5928 ( .A(n6684), .ZN(n6704) );
  NAND2_X1 U5929 ( .A1(n6721), .A2(n6701), .ZN(n4787) );
  OAI21_X1 U5930 ( .B1(n6683), .B2(n6710), .A(n4787), .ZN(n4788) );
  AOI21_X1 U5931 ( .B1(n6723), .B2(n6704), .A(n4788), .ZN(n4789) );
  OAI211_X1 U5932 ( .C1(n6713), .C2(n6709), .A(n4790), .B(n4789), .ZN(U3147)
         );
  NAND2_X1 U5933 ( .A1(n4795), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4794)
         );
  INV_X1 U5934 ( .A(n6671), .ZN(n6610) );
  NAND2_X1 U5935 ( .A1(n6721), .A2(n6673), .ZN(n4791) );
  OAI21_X1 U5936 ( .B1(n6670), .B2(n6710), .A(n4791), .ZN(n4792) );
  AOI21_X1 U5937 ( .B1(n6723), .B2(n6610), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5938 ( .C1(n6713), .C2(n6676), .A(n4794), .B(n4793), .ZN(U3145)
         );
  NAND2_X1 U5939 ( .A1(n4795), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4799)
         );
  INV_X1 U5940 ( .A(n6663), .ZN(n6604) );
  NAND2_X1 U5941 ( .A1(n6721), .A2(n6660), .ZN(n4796) );
  OAI21_X1 U5942 ( .B1(n6657), .B2(n6710), .A(n4796), .ZN(n4797) );
  AOI21_X1 U5943 ( .B1(n6723), .B2(n6604), .A(n4797), .ZN(n4798) );
  OAI211_X1 U5944 ( .C1(n6713), .C2(n6658), .A(n4799), .B(n4798), .ZN(U3143)
         );
  AOI22_X1 U5945 ( .A1(n6396), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4837), .ZN(n4803) );
  NAND2_X1 U5946 ( .A1(n6395), .A2(DATAI_7_), .ZN(n4807) );
  NAND2_X1 U5947 ( .A1(n4803), .A2(n4807), .ZN(U2931) );
  AOI22_X1 U5948 ( .A1(n6396), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4837), .ZN(n4804) );
  NAND2_X1 U5949 ( .A1(n6395), .A2(DATAI_6_), .ZN(n4809) );
  NAND2_X1 U5950 ( .A1(n4804), .A2(n4809), .ZN(U2930) );
  AOI22_X1 U5951 ( .A1(n6396), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4837), .ZN(n4805) );
  NAND2_X1 U5952 ( .A1(n6395), .A2(DATAI_5_), .ZN(n4811) );
  NAND2_X1 U5953 ( .A1(n4805), .A2(n4811), .ZN(U2929) );
  AOI22_X1 U5954 ( .A1(n6396), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4837), .ZN(n4806) );
  NAND2_X1 U5955 ( .A1(n6395), .A2(DATAI_8_), .ZN(n4813) );
  NAND2_X1 U5956 ( .A1(n4806), .A2(n4813), .ZN(U2947) );
  AOI22_X1 U5957 ( .A1(n6396), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4837), .ZN(n4808) );
  NAND2_X1 U5958 ( .A1(n4808), .A2(n4807), .ZN(U2946) );
  AOI22_X1 U5959 ( .A1(n6396), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4837), .ZN(n4810) );
  NAND2_X1 U5960 ( .A1(n4810), .A2(n4809), .ZN(U2945) );
  AOI22_X1 U5961 ( .A1(n6396), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4837), .ZN(n4812) );
  NAND2_X1 U5962 ( .A1(n4812), .A2(n4811), .ZN(U2944) );
  AOI22_X1 U5963 ( .A1(n6396), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4837), .ZN(n4814) );
  NAND2_X1 U5964 ( .A1(n4814), .A2(n4813), .ZN(U2932) );
  AOI22_X1 U5965 ( .A1(n6396), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4837), .ZN(n4815) );
  NAND2_X1 U5966 ( .A1(n6395), .A2(DATAI_14_), .ZN(n4838) );
  NAND2_X1 U5967 ( .A1(n4815), .A2(n4838), .ZN(U2953) );
  AOI22_X1 U5968 ( .A1(n6396), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4837), .ZN(n4816) );
  NAND2_X1 U5969 ( .A1(n6395), .A2(DATAI_3_), .ZN(n4826) );
  NAND2_X1 U5970 ( .A1(n4816), .A2(n4826), .ZN(U2942) );
  AOI22_X1 U5971 ( .A1(n6396), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4837), .ZN(n4817) );
  NAND2_X1 U5972 ( .A1(n6395), .A2(DATAI_12_), .ZN(n4821) );
  NAND2_X1 U5973 ( .A1(n4817), .A2(n4821), .ZN(U2951) );
  AOI22_X1 U5974 ( .A1(n6396), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4837), .ZN(n4818) );
  NAND2_X1 U5975 ( .A1(n6395), .A2(DATAI_1_), .ZN(n4823) );
  NAND2_X1 U5976 ( .A1(n4818), .A2(n4823), .ZN(U2940) );
  AOI22_X1 U5977 ( .A1(n6396), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n4837), .ZN(n4819) );
  NAND2_X1 U5978 ( .A1(n6395), .A2(DATAI_10_), .ZN(n4833) );
  NAND2_X1 U5979 ( .A1(n4819), .A2(n4833), .ZN(U2949) );
  AOI22_X1 U5980 ( .A1(n6396), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4837), .ZN(n4820) );
  NAND2_X1 U5981 ( .A1(n6395), .A2(DATAI_2_), .ZN(n4831) );
  NAND2_X1 U5982 ( .A1(n4820), .A2(n4831), .ZN(U2926) );
  AOI22_X1 U5983 ( .A1(n6396), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4837), .ZN(n4822) );
  NAND2_X1 U5984 ( .A1(n4822), .A2(n4821), .ZN(U2936) );
  AOI22_X1 U5985 ( .A1(n6396), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4837), .ZN(n4824) );
  NAND2_X1 U5986 ( .A1(n4824), .A2(n4823), .ZN(U2925) );
  AOI22_X1 U5987 ( .A1(n6396), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4837), .ZN(n4825) );
  NAND2_X1 U5988 ( .A1(n6395), .A2(DATAI_0_), .ZN(n4829) );
  NAND2_X1 U5989 ( .A1(n4825), .A2(n4829), .ZN(U2924) );
  AOI22_X1 U5990 ( .A1(n6396), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4837), .ZN(n4827) );
  NAND2_X1 U5991 ( .A1(n4827), .A2(n4826), .ZN(U2927) );
  AOI22_X1 U5992 ( .A1(n6396), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4837), .ZN(n4828) );
  NAND2_X1 U5993 ( .A1(n6395), .A2(DATAI_4_), .ZN(n4835) );
  NAND2_X1 U5994 ( .A1(n4828), .A2(n4835), .ZN(U2928) );
  AOI22_X1 U5995 ( .A1(n6396), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4837), .ZN(n4830) );
  NAND2_X1 U5996 ( .A1(n4830), .A2(n4829), .ZN(U2939) );
  AOI22_X1 U5997 ( .A1(n6396), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4837), .ZN(n4832) );
  NAND2_X1 U5998 ( .A1(n4832), .A2(n4831), .ZN(U2941) );
  AOI22_X1 U5999 ( .A1(n6396), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n4837), .ZN(n4834) );
  NAND2_X1 U6000 ( .A1(n4834), .A2(n4833), .ZN(U2934) );
  AOI22_X1 U6001 ( .A1(n6396), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4837), .ZN(n4836) );
  NAND2_X1 U6002 ( .A1(n4836), .A2(n4835), .ZN(U2943) );
  AOI22_X1 U6003 ( .A1(n6396), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4837), .ZN(n4839) );
  NAND2_X1 U6004 ( .A1(n4839), .A2(n4838), .ZN(U2938) );
  XNOR2_X1 U6005 ( .A(n4840), .B(n4841), .ZN(n4850) );
  NAND2_X1 U6006 ( .A1(n6399), .A2(REIP_REG_4__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U6007 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4842)
         );
  OAI211_X1 U6008 ( .C1(n6418), .C2(n6325), .A(n4846), .B(n4842), .ZN(n4843)
         );
  AOI21_X1 U6009 ( .B1(n4844), .B2(n6404), .A(n4843), .ZN(n4845) );
  OAI21_X1 U6010 ( .B1(n6226), .B2(n4850), .A(n4845), .ZN(U2982) );
  NAND2_X1 U6011 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5102) );
  OAI211_X1 U6012 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5235), .B(n5102), .ZN(n4847) );
  OAI211_X1 U6013 ( .C1(n6455), .C2(n6333), .A(n4847), .B(n4846), .ZN(n4848)
         );
  AOI21_X1 U6014 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n5100), .A(n4848), 
        .ZN(n4849) );
  OAI21_X1 U6015 ( .B1(n6422), .B2(n4850), .A(n4849), .ZN(U3014) );
  INV_X1 U6016 ( .A(n4851), .ZN(n4889) );
  NOR2_X1 U6017 ( .A1(n4852), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4853)
         );
  AOI21_X1 U6018 ( .B1(n3114), .B2(n4854), .A(n4853), .ZN(n5264) );
  AOI21_X1 U6019 ( .B1(n5261), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6582), 
        .ZN(n4856) );
  NAND2_X1 U6020 ( .A1(n5264), .A2(n4856), .ZN(n4857) );
  NOR2_X1 U6021 ( .A1(n4857), .A2(n4858), .ZN(n4862) );
  AOI22_X1 U6022 ( .A1(n4860), .A2(n4859), .B1(n4858), .B2(n4857), .ZN(n4861)
         );
  AOI211_X1 U6023 ( .C1(n4863), .C2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n4862), .B(n4861), .ZN(n4866) );
  NOR2_X1 U6024 ( .A1(n4863), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4865)
         );
  INV_X1 U6025 ( .A(n4868), .ZN(n4864) );
  OAI22_X1 U6026 ( .A1(n4866), .A2(n4865), .B1(n4864), .B2(n5129), .ZN(n4867)
         );
  OAI21_X1 U6027 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4868), .A(n4867), 
        .ZN(n4887) );
  INV_X1 U6028 ( .A(n4869), .ZN(n4883) );
  INV_X1 U6029 ( .A(MORE_REG_SCAN_IN), .ZN(n7018) );
  INV_X1 U6030 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6227) );
  NAND3_X1 U6031 ( .A1(n4871), .A2(n4870), .A3(n5296), .ZN(n4872) );
  NAND2_X1 U6032 ( .A1(n4872), .A2(n7019), .ZN(n5279) );
  NAND2_X1 U6033 ( .A1(n4873), .A2(n5279), .ZN(n5289) );
  AOI21_X1 U6034 ( .B1(n7018), .B2(n6227), .A(n5289), .ZN(n4882) );
  AND2_X1 U6035 ( .A1(n4875), .A2(n4874), .ZN(n4877) );
  MUX2_X1 U6036 ( .A(n4878), .B(n4877), .S(n4876), .Z(n4879) );
  OAI21_X1 U6037 ( .B1(n4881), .B2(n4880), .A(n4879), .ZN(n5290) );
  AOI211_X1 U6038 ( .C1(n6466), .C2(n4887), .A(n4886), .B(n4885), .ZN(n5115)
         );
  AOI22_X1 U6039 ( .A1(n5115), .A2(n6729), .B1(READY_N), .B2(n6374), .ZN(n4888) );
  AOI21_X1 U6040 ( .B1(n4890), .B2(n4889), .A(n4888), .ZN(n6736) );
  INV_X1 U6041 ( .A(n6736), .ZN(n5106) );
  INV_X1 U6042 ( .A(n5110), .ZN(n4891) );
  OAI211_X1 U6043 ( .C1(n5106), .C2(n4338), .A(n4892), .B(n4891), .ZN(U3453)
         );
  NAND3_X1 U6044 ( .A1(n4893), .A2(n5010), .A3(n4894), .ZN(n4927) );
  INV_X1 U6045 ( .A(n4927), .ZN(n4895) );
  NOR2_X1 U6046 ( .A1(n6141), .A2(n6586), .ZN(n4925) );
  INV_X1 U6047 ( .A(n4925), .ZN(n4896) );
  OAI211_X1 U6048 ( .C1(n6489), .C2(n4897), .A(n4931), .B(n4896), .ZN(n4901)
         );
  NOR3_X1 U6049 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4933) );
  INV_X1 U6050 ( .A(n4933), .ZN(n4898) );
  OR2_X1 U6051 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4898), .ZN(n6132)
         );
  NAND2_X1 U6052 ( .A1(n4902), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6590) );
  INV_X1 U6053 ( .A(n6590), .ZN(n5083) );
  OAI21_X1 U6054 ( .B1(n6578), .B2(n6197), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4899) );
  NAND2_X1 U6055 ( .A1(n4899), .A2(n5023), .ZN(n6491) );
  AOI211_X1 U6056 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6132), .A(n5083), .B(
        n6491), .ZN(n4900) );
  NAND2_X1 U6057 ( .A1(n4901), .A2(n4900), .ZN(n6131) );
  NAND2_X1 U6058 ( .A1(n6131), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4906) );
  NOR2_X1 U6059 ( .A1(n4902), .A2(n6632), .ZN(n6492) );
  INV_X1 U6060 ( .A(n6197), .ZN(n6191) );
  NAND2_X1 U6061 ( .A1(n6492), .A2(n6191), .ZN(n6579) );
  NOR2_X1 U6062 ( .A1(n6579), .A2(n6578), .ZN(n4903) );
  AOI21_X1 U6063 ( .B1(n4925), .B2(n6626), .A(n4903), .ZN(n6133) );
  OAI22_X1 U6064 ( .A1(n6133), .A2(n5192), .B1(n6677), .B2(n6132), .ZN(n4904)
         );
  AOI21_X1 U6065 ( .B1(n6723), .B2(n5089), .A(n4904), .ZN(n4905) );
  OAI211_X1 U6066 ( .C1(n6137), .C2(n6678), .A(n4906), .B(n4905), .ZN(U3026)
         );
  NAND2_X1 U6067 ( .A1(n6131), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4909) );
  OAI22_X1 U6068 ( .A1(n6133), .A2(n6203), .B1(n6643), .B2(n6132), .ZN(n4907)
         );
  AOI21_X1 U6069 ( .B1(n6723), .B2(n6521), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6070 ( .C1(n6137), .C2(n6649), .A(n4909), .B(n4908), .ZN(U3021)
         );
  NAND2_X1 U6071 ( .A1(n6131), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6072 ( .A1(n6133), .A2(n6207), .B1(n6650), .B2(n6132), .ZN(n4910)
         );
  AOI21_X1 U6073 ( .B1(n6723), .B2(n6524), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6074 ( .C1(n6137), .C2(n6651), .A(n4912), .B(n4911), .ZN(U3022)
         );
  NAND2_X1 U6075 ( .A1(n6131), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U6076 ( .A1(n6133), .A2(n6215), .B1(n6664), .B2(n6132), .ZN(n4913)
         );
  AOI21_X1 U6077 ( .B1(n6723), .B2(n6724), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6078 ( .C1(n6137), .C2(n6665), .A(n4915), .B(n4914), .ZN(U3024)
         );
  NAND2_X1 U6079 ( .A1(n6131), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4918) );
  OAI22_X1 U6080 ( .A1(n6133), .A2(n5175), .B1(n6683), .B2(n6132), .ZN(n4916)
         );
  AOI21_X1 U6081 ( .B1(n6723), .B2(n6477), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6082 ( .C1(n6137), .C2(n6684), .A(n4918), .B(n4917), .ZN(U3027)
         );
  NAND2_X1 U6083 ( .A1(n6131), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4921) );
  OAI22_X1 U6084 ( .A1(n6133), .A2(n6211), .B1(n6657), .B2(n6132), .ZN(n4919)
         );
  AOI21_X1 U6085 ( .B1(n6723), .B2(n6527), .A(n4919), .ZN(n4920) );
  OAI211_X1 U6086 ( .C1(n6137), .C2(n6663), .A(n4921), .B(n4920), .ZN(U3023)
         );
  NAND2_X1 U6087 ( .A1(n6131), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4924) );
  OAI22_X1 U6088 ( .A1(n6133), .A2(n6219), .B1(n6670), .B2(n6132), .ZN(n4922)
         );
  AOI21_X1 U6089 ( .B1(n6723), .B2(n6535), .A(n4922), .ZN(n4923) );
  OAI211_X1 U6090 ( .C1(n6137), .C2(n6671), .A(n4924), .B(n4923), .ZN(U3025)
         );
  AND2_X1 U6091 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4933), .ZN(n4928)
         );
  AOI21_X1 U6092 ( .B1(n4925), .B2(n3114), .A(n4928), .ZN(n4930) );
  INV_X1 U6093 ( .A(n4930), .ZN(n4926) );
  INV_X1 U6094 ( .A(n4928), .ZN(n4954) );
  OAI22_X1 U6095 ( .A1(n5197), .A2(n6651), .B1(n6650), .B2(n4954), .ZN(n4929)
         );
  AOI21_X1 U6096 ( .B1(n6524), .B2(n4956), .A(n4929), .ZN(n4935) );
  NAND2_X1 U6097 ( .A1(n4931), .A2(n4930), .ZN(n4932) );
  NAND2_X1 U6098 ( .A1(n4957), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4934) );
  OAI211_X1 U6099 ( .C1(n4960), .C2(n6207), .A(n4935), .B(n4934), .ZN(U3030)
         );
  OAI22_X1 U6100 ( .A1(n5197), .A2(n6642), .B1(n6623), .B2(n4954), .ZN(n4936)
         );
  AOI21_X1 U6101 ( .B1(n6715), .B2(n4956), .A(n4936), .ZN(n4938) );
  NAND2_X1 U6102 ( .A1(n4957), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4937) );
  OAI211_X1 U6103 ( .C1(n4960), .C2(n6199), .A(n4938), .B(n4937), .ZN(U3028)
         );
  OAI22_X1 U6104 ( .A1(n5197), .A2(n6671), .B1(n6670), .B2(n4954), .ZN(n4939)
         );
  AOI21_X1 U6105 ( .B1(n6535), .B2(n4956), .A(n4939), .ZN(n4941) );
  NAND2_X1 U6106 ( .A1(n4957), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4940) );
  OAI211_X1 U6107 ( .C1(n4960), .C2(n6219), .A(n4941), .B(n4940), .ZN(U3033)
         );
  OAI22_X1 U6108 ( .A1(n5197), .A2(n6678), .B1(n6677), .B2(n4954), .ZN(n4942)
         );
  AOI21_X1 U6109 ( .B1(n5089), .B2(n4956), .A(n4942), .ZN(n4944) );
  NAND2_X1 U6110 ( .A1(n4957), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4943) );
  OAI211_X1 U6111 ( .C1(n4960), .C2(n5192), .A(n4944), .B(n4943), .ZN(U3034)
         );
  OAI22_X1 U6112 ( .A1(n5197), .A2(n6663), .B1(n6657), .B2(n4954), .ZN(n4945)
         );
  AOI21_X1 U6113 ( .B1(n6527), .B2(n4956), .A(n4945), .ZN(n4947) );
  NAND2_X1 U6114 ( .A1(n4957), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4946) );
  OAI211_X1 U6115 ( .C1(n4960), .C2(n6211), .A(n4947), .B(n4946), .ZN(U3031)
         );
  OAI22_X1 U6116 ( .A1(n5197), .A2(n6665), .B1(n6664), .B2(n4954), .ZN(n4948)
         );
  AOI21_X1 U6117 ( .B1(n6724), .B2(n4956), .A(n4948), .ZN(n4950) );
  NAND2_X1 U6118 ( .A1(n4957), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4949) );
  OAI211_X1 U6119 ( .C1(n4960), .C2(n6215), .A(n4950), .B(n4949), .ZN(U3032)
         );
  OAI22_X1 U6120 ( .A1(n5197), .A2(n6649), .B1(n6643), .B2(n4954), .ZN(n4951)
         );
  AOI21_X1 U6121 ( .B1(n6521), .B2(n4956), .A(n4951), .ZN(n4953) );
  NAND2_X1 U6122 ( .A1(n4957), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4952) );
  OAI211_X1 U6123 ( .C1(n4960), .C2(n6203), .A(n4953), .B(n4952), .ZN(U3029)
         );
  OAI22_X1 U6124 ( .A1(n5197), .A2(n6684), .B1(n6683), .B2(n4954), .ZN(n4955)
         );
  AOI21_X1 U6125 ( .B1(n6477), .B2(n4956), .A(n4955), .ZN(n4959) );
  NAND2_X1 U6126 ( .A1(n4957), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4958) );
  OAI211_X1 U6127 ( .C1(n4960), .C2(n5175), .A(n4959), .B(n4958), .ZN(U3035)
         );
  INV_X1 U6128 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4966) );
  INV_X1 U6129 ( .A(n6513), .ZN(n4989) );
  INV_X1 U6130 ( .A(n6670), .ZN(n6609) );
  AOI22_X1 U6131 ( .A1(n6534), .A2(n6610), .B1(n6609), .B2(n4987), .ZN(n4963)
         );
  OAI21_X1 U6132 ( .B1(n4989), .B2(n6676), .A(n4963), .ZN(n4964) );
  AOI21_X1 U6133 ( .B1(n6673), .B2(n4991), .A(n4964), .ZN(n4965) );
  OAI21_X1 U6134 ( .B1(n4994), .B2(n4966), .A(n4965), .ZN(U3065) );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4970) );
  INV_X1 U6136 ( .A(n6677), .ZN(n6693) );
  AOI22_X1 U6137 ( .A1(n6534), .A2(n6695), .B1(n6693), .B2(n4987), .ZN(n4967)
         );
  OAI21_X1 U6138 ( .B1(n4989), .B2(n6698), .A(n4967), .ZN(n4968) );
  AOI21_X1 U6139 ( .B1(n6694), .B2(n4991), .A(n4968), .ZN(n4969) );
  OAI21_X1 U6140 ( .B1(n4994), .B2(n4970), .A(n4969), .ZN(U3066) );
  INV_X1 U6141 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U6142 ( .A1(n6534), .A2(n6600), .B1(n6599), .B2(n4987), .ZN(n4971)
         );
  OAI21_X1 U6143 ( .B1(n4989), .B2(n6656), .A(n4971), .ZN(n4972) );
  AOI21_X1 U6144 ( .B1(n6653), .B2(n4991), .A(n4972), .ZN(n4973) );
  OAI21_X1 U6145 ( .B1(n4994), .B2(n4974), .A(n4973), .ZN(U3062) );
  INV_X1 U6146 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4978) );
  AOI22_X1 U6147 ( .A1(n6534), .A2(n6604), .B1(n6603), .B2(n4987), .ZN(n4975)
         );
  OAI21_X1 U6148 ( .B1(n4989), .B2(n6658), .A(n4975), .ZN(n4976) );
  AOI21_X1 U6149 ( .B1(n6660), .B2(n4991), .A(n4976), .ZN(n4977) );
  OAI21_X1 U6150 ( .B1(n4994), .B2(n4978), .A(n4977), .ZN(U3063) );
  INV_X1 U6151 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4982) );
  AOI22_X1 U6152 ( .A1(n6534), .A2(n6596), .B1(n6595), .B2(n4987), .ZN(n4979)
         );
  OAI21_X1 U6153 ( .B1(n4989), .B2(n6644), .A(n4979), .ZN(n4980) );
  AOI21_X1 U6154 ( .B1(n6646), .B2(n4991), .A(n4980), .ZN(n4981) );
  OAI21_X1 U6155 ( .B1(n4994), .B2(n4982), .A(n4981), .ZN(U3061) );
  INV_X1 U6156 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4986) );
  INV_X1 U6157 ( .A(n6665), .ZN(n6722) );
  AOI22_X1 U6158 ( .A1(n6534), .A2(n6722), .B1(n6718), .B2(n4987), .ZN(n4983)
         );
  OAI21_X1 U6159 ( .B1(n4989), .B2(n6669), .A(n4983), .ZN(n4984) );
  AOI21_X1 U6160 ( .B1(n6720), .B2(n4991), .A(n4984), .ZN(n4985) );
  OAI21_X1 U6161 ( .B1(n4994), .B2(n4986), .A(n4985), .ZN(U3064) );
  INV_X1 U6162 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U6163 ( .A1(n6534), .A2(n6704), .B1(n6700), .B2(n4987), .ZN(n4988)
         );
  OAI21_X1 U6164 ( .B1(n4989), .B2(n6709), .A(n4988), .ZN(n4990) );
  AOI21_X1 U6165 ( .B1(n6701), .B2(n4991), .A(n4990), .ZN(n4992) );
  OAI21_X1 U6166 ( .B1(n4994), .B2(n4993), .A(n4992), .ZN(U3067) );
  NAND2_X1 U6167 ( .A1(n4996), .A2(n4995), .ZN(n5068) );
  OAI21_X1 U6168 ( .B1(n4996), .B2(n4995), .A(n5068), .ZN(n5116) );
  INV_X1 U6169 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4999) );
  OAI21_X1 U6170 ( .B1(n4760), .B2(n4998), .A(n4997), .ZN(n6303) );
  OAI222_X1 U6171 ( .A1(n5116), .A2(n7064), .B1(n5628), .B2(n4999), .C1(n6303), 
        .C2(n7065), .ZN(U2854) );
  INV_X1 U6172 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6370) );
  OAI222_X1 U6173 ( .A1(n5116), .A2(n5683), .B1(n5072), .B2(n5000), .C1(n5070), 
        .C2(n6370), .ZN(U2886) );
  NAND2_X1 U6174 ( .A1(n6628), .A2(n5001), .ZN(n6118) );
  NAND2_X1 U6175 ( .A1(n6116), .A2(n5010), .ZN(n5002) );
  OAI21_X1 U6176 ( .B1(n6118), .B2(n5002), .A(n6626), .ZN(n5009) );
  INV_X1 U6177 ( .A(n6141), .ZN(n6587) );
  NOR2_X1 U6178 ( .A1(n5577), .A2(n5003), .ZN(n6142) );
  NAND2_X1 U6179 ( .A1(n6587), .A2(n6142), .ZN(n5127) );
  OR2_X1 U6180 ( .A1(n5127), .A2(n6629), .ZN(n5005) );
  INV_X1 U6181 ( .A(n5004), .ZN(n6622) );
  NAND2_X1 U6182 ( .A1(n6622), .A2(n5129), .ZN(n6467) );
  AND2_X1 U6183 ( .A1(n5005), .A2(n6467), .ZN(n5006) );
  NAND3_X1 U6184 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5129), .A3(n6143), .ZN(n5124) );
  OAI22_X1 U6185 ( .A1(n5009), .A2(n5006), .B1(n5124), .B2(n6632), .ZN(n6480)
         );
  INV_X1 U6186 ( .A(n6480), .ZN(n5020) );
  INV_X1 U6187 ( .A(n5006), .ZN(n5008) );
  AOI21_X1 U6188 ( .B1(n6636), .B2(n5124), .A(n6634), .ZN(n5007) );
  NOR2_X1 U6189 ( .A1(n6517), .A2(n6671), .ZN(n5012) );
  INV_X1 U6190 ( .A(n6138), .ZN(n5073) );
  INV_X1 U6191 ( .A(n6478), .ZN(n5201) );
  OAI22_X1 U6192 ( .A1(n5201), .A2(n6676), .B1(n6670), .B2(n6467), .ZN(n5011)
         );
  AOI211_X1 U6193 ( .C1(n6479), .C2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n5012), 
        .B(n5011), .ZN(n5013) );
  OAI21_X1 U6194 ( .B1(n5020), .B2(n6219), .A(n5013), .ZN(U3049) );
  NOR2_X1 U6195 ( .A1(n6517), .A2(n6642), .ZN(n5015) );
  OAI22_X1 U6196 ( .A1(n5201), .A2(n6624), .B1(n6623), .B2(n6467), .ZN(n5014)
         );
  AOI211_X1 U6197 ( .C1(n6479), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n5015), 
        .B(n5014), .ZN(n5016) );
  OAI21_X1 U6198 ( .B1(n5020), .B2(n6199), .A(n5016), .ZN(U3044) );
  NOR2_X1 U6199 ( .A1(n6517), .A2(n6678), .ZN(n5018) );
  OAI22_X1 U6200 ( .A1(n5201), .A2(n6698), .B1(n6677), .B2(n6467), .ZN(n5017)
         );
  AOI211_X1 U6201 ( .C1(n6479), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n5018), 
        .B(n5017), .ZN(n5019) );
  OAI21_X1 U6202 ( .B1(n5020), .B2(n5192), .A(n5019), .ZN(U3050) );
  INV_X1 U6203 ( .A(n5076), .ZN(n5082) );
  AOI21_X1 U6204 ( .B1(n5027), .B2(n6713), .A(n6225), .ZN(n5021) );
  AOI211_X1 U6205 ( .C1(n5082), .C2(n6141), .A(n6636), .B(n5021), .ZN(n5026)
         );
  NOR2_X1 U6206 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5022), .ZN(n5058)
         );
  OR2_X1 U6207 ( .A1(n6197), .A2(n6632), .ZN(n5024) );
  NAND2_X1 U6208 ( .A1(n5024), .A2(n5023), .ZN(n5078) );
  AOI21_X1 U6209 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5129), .A(n5078), .ZN(
        n6144) );
  INV_X1 U6210 ( .A(n6492), .ZN(n5079) );
  OAI211_X1 U6211 ( .C1(n4338), .C2(n5058), .A(n6144), .B(n5079), .ZN(n5025)
         );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5033) );
  AND2_X1 U6213 ( .A1(n6141), .A2(n6626), .ZN(n6577) );
  NAND2_X1 U6214 ( .A1(n6577), .A2(n5082), .ZN(n5029) );
  NAND3_X1 U6215 ( .A1(n5083), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6197), .ZN(n5028) );
  NAND2_X1 U6216 ( .A1(n5029), .A2(n5028), .ZN(n5059) );
  AOI22_X1 U6217 ( .A1(n5059), .A2(n6653), .B1(n6599), .B2(n5058), .ZN(n5030)
         );
  OAI21_X1 U6218 ( .B1(n6713), .B2(n6651), .A(n5030), .ZN(n5031) );
  AOI21_X1 U6219 ( .B1(n6524), .B2(n5062), .A(n5031), .ZN(n5032) );
  OAI21_X1 U6220 ( .B1(n5065), .B2(n5033), .A(n5032), .ZN(U3134) );
  INV_X1 U6221 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5037) );
  AOI22_X1 U6222 ( .A1(n5059), .A2(n6646), .B1(n6595), .B2(n5058), .ZN(n5034)
         );
  OAI21_X1 U6223 ( .B1(n6713), .B2(n6649), .A(n5034), .ZN(n5035) );
  AOI21_X1 U6224 ( .B1(n6521), .B2(n5062), .A(n5035), .ZN(n5036) );
  OAI21_X1 U6225 ( .B1(n5065), .B2(n5037), .A(n5036), .ZN(U3133) );
  INV_X1 U6226 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5041) );
  AOI22_X1 U6227 ( .A1(n5059), .A2(n6712), .B1(n6711), .B2(n5058), .ZN(n5038)
         );
  OAI21_X1 U6228 ( .B1(n6713), .B2(n6642), .A(n5038), .ZN(n5039) );
  AOI21_X1 U6229 ( .B1(n6715), .B2(n5062), .A(n5039), .ZN(n5040) );
  OAI21_X1 U6230 ( .B1(n5065), .B2(n5041), .A(n5040), .ZN(U3132) );
  INV_X1 U6231 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5045) );
  AOI22_X1 U6232 ( .A1(n5059), .A2(n6673), .B1(n6609), .B2(n5058), .ZN(n5042)
         );
  OAI21_X1 U6233 ( .B1(n6713), .B2(n6671), .A(n5042), .ZN(n5043) );
  AOI21_X1 U6234 ( .B1(n6535), .B2(n5062), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6235 ( .B1(n5065), .B2(n5045), .A(n5044), .ZN(U3137) );
  INV_X1 U6236 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5049) );
  AOI22_X1 U6237 ( .A1(n5059), .A2(n6701), .B1(n6700), .B2(n5058), .ZN(n5046)
         );
  OAI21_X1 U6238 ( .B1(n6713), .B2(n6684), .A(n5046), .ZN(n5047) );
  AOI21_X1 U6239 ( .B1(n6477), .B2(n5062), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6240 ( .B1(n5065), .B2(n5049), .A(n5048), .ZN(U3139) );
  INV_X1 U6241 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6242 ( .A1(n5059), .A2(n6720), .B1(n6718), .B2(n5058), .ZN(n5050)
         );
  OAI21_X1 U6243 ( .B1(n6713), .B2(n6665), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6244 ( .B1(n6724), .B2(n5062), .A(n5051), .ZN(n5052) );
  OAI21_X1 U6245 ( .B1(n5065), .B2(n5053), .A(n5052), .ZN(U3136) );
  INV_X1 U6246 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U6247 ( .A1(n5059), .A2(n6660), .B1(n6603), .B2(n5058), .ZN(n5054)
         );
  OAI21_X1 U6248 ( .B1(n6713), .B2(n6663), .A(n5054), .ZN(n5055) );
  AOI21_X1 U6249 ( .B1(n6527), .B2(n5062), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6250 ( .B1(n5065), .B2(n5057), .A(n5056), .ZN(U3135) );
  INV_X1 U6251 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6252 ( .A1(n5059), .A2(n6694), .B1(n6693), .B2(n5058), .ZN(n5060)
         );
  OAI21_X1 U6253 ( .B1(n6713), .B2(n6678), .A(n5060), .ZN(n5061) );
  AOI21_X1 U6254 ( .B1(n5089), .B2(n5062), .A(n5061), .ZN(n5063) );
  OAI21_X1 U6255 ( .B1(n5065), .B2(n5064), .A(n5063), .ZN(U3138) );
  INV_X1 U6256 ( .A(n5066), .ZN(n5069) );
  AOI21_X1 U6257 ( .B1(n5069), .B2(n5068), .A(n5067), .ZN(n6298) );
  INV_X1 U6258 ( .A(n6298), .ZN(n7063) );
  INV_X1 U6259 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U6260 ( .A1(n7063), .A2(n5683), .B1(n5072), .B2(n5071), .C1(n6836), 
        .C2(n5070), .ZN(U2885) );
  INV_X1 U6261 ( .A(n6576), .ZN(n5074) );
  OAI21_X1 U6262 ( .B1(n6534), .B2(n5074), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5077) );
  OR2_X1 U6263 ( .A1(n5076), .A2(n5075), .ZN(n6542) );
  NAND3_X1 U6264 ( .A1(n5077), .A2(n6626), .A3(n6542), .ZN(n5081) );
  INV_X1 U6265 ( .A(n5078), .ZN(n5125) );
  NAND2_X1 U6266 ( .A1(n6546), .A2(n6582), .ZN(n6518) );
  AOI21_X1 U6267 ( .B1(n6518), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5080) );
  NAND4_X1 U6268 ( .A1(n5081), .A2(n5125), .A3(n5080), .A4(n5079), .ZN(n6536)
         );
  INV_X1 U6269 ( .A(n6536), .ZN(n5097) );
  INV_X1 U6270 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5091) );
  NOR2_X1 U6271 ( .A1(n6141), .A2(n6636), .ZN(n6483) );
  NAND2_X1 U6272 ( .A1(n6483), .A2(n5082), .ZN(n5085) );
  NAND3_X1 U6273 ( .A1(n5083), .A2(n6197), .A3(n5129), .ZN(n5084) );
  NAND2_X1 U6274 ( .A1(n5085), .A2(n5084), .ZN(n6533) );
  NOR2_X1 U6275 ( .A1(n6677), .A2(n6518), .ZN(n5086) );
  AOI21_X1 U6276 ( .B1(n6533), .B2(n6694), .A(n5086), .ZN(n5087) );
  OAI21_X1 U6277 ( .B1(n6576), .B2(n6678), .A(n5087), .ZN(n5088) );
  AOI21_X1 U6278 ( .B1(n5089), .B2(n6534), .A(n5088), .ZN(n5090) );
  OAI21_X1 U6279 ( .B1(n5097), .B2(n5091), .A(n5090), .ZN(U3074) );
  INV_X1 U6280 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5096) );
  NOR2_X1 U6281 ( .A1(n6683), .A2(n6518), .ZN(n5092) );
  AOI21_X1 U6282 ( .B1(n6533), .B2(n6701), .A(n5092), .ZN(n5093) );
  OAI21_X1 U6283 ( .B1(n6576), .B2(n6684), .A(n5093), .ZN(n5094) );
  AOI21_X1 U6284 ( .B1(n6477), .B2(n6534), .A(n5094), .ZN(n5095) );
  OAI21_X1 U6285 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(U3075) );
  XNOR2_X1 U6286 ( .A(n5099), .B(n5098), .ZN(n5121) );
  INV_X1 U6287 ( .A(n6420), .ZN(n6010) );
  NOR2_X1 U6288 ( .A1(n4285), .A2(n5102), .ZN(n5251) );
  INV_X1 U6289 ( .A(n5100), .ZN(n5101) );
  OAI21_X1 U6290 ( .B1(n6010), .B2(n5251), .A(n5101), .ZN(n5239) );
  INV_X1 U6291 ( .A(n5235), .ZN(n5256) );
  OAI21_X1 U6292 ( .B1(n5256), .B2(n5102), .A(n4285), .ZN(n5104) );
  NAND2_X1 U6293 ( .A1(n6399), .A2(REIP_REG_5__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U6294 ( .B1(n6455), .B2(n6303), .A(n5117), .ZN(n5103) );
  AOI21_X1 U6295 ( .B1(n5239), .B2(n5104), .A(n5103), .ZN(n5105) );
  OAI21_X1 U6296 ( .B1(n6422), .B2(n5121), .A(n5105), .ZN(U3013) );
  OAI21_X1 U6297 ( .B1(n5281), .B2(n6124), .A(n5106), .ZN(n5107) );
  AOI21_X1 U6298 ( .B1(n6632), .B2(READY_N), .A(n6736), .ZN(n6731) );
  MUX2_X1 U6299 ( .A(n5107), .B(n6731), .S(STATE2_REG_0__SCAN_IN), .Z(n5113)
         );
  INV_X1 U6300 ( .A(n5108), .ZN(n5109) );
  AOI21_X1 U6301 ( .B1(n5111), .B2(n5110), .A(n5109), .ZN(n5112) );
  OAI211_X1 U6302 ( .C1(n5115), .C2(n5114), .A(n5113), .B(n5112), .ZN(U3148)
         );
  INV_X1 U6303 ( .A(n5116), .ZN(n6310) );
  NOR2_X1 U6304 ( .A1(n6418), .A2(n6316), .ZN(n5119) );
  OAI21_X1 U6305 ( .B1(n5868), .B2(n3723), .A(n5117), .ZN(n5118) );
  AOI211_X1 U6306 ( .C1(n6310), .C2(n6404), .A(n5119), .B(n5118), .ZN(n5120)
         );
  OAI21_X1 U6307 ( .B1(n6226), .B2(n5121), .A(n5120), .ZN(U2981) );
  INV_X1 U6308 ( .A(n5197), .ZN(n5122) );
  OAI21_X1 U6309 ( .B1(n5122), .B2(n6478), .A(n6121), .ZN(n5123) );
  AOI21_X1 U6310 ( .B1(n5123), .B2(n5127), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5126) );
  NOR2_X1 U6311 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5124), .ZN(n5198)
         );
  INV_X1 U6312 ( .A(n5127), .ZN(n5128) );
  NAND2_X1 U6313 ( .A1(n5128), .A2(n6626), .ZN(n5131) );
  NAND3_X1 U6314 ( .A1(n6492), .A2(n6197), .A3(n5129), .ZN(n5130) );
  NAND2_X1 U6315 ( .A1(n5131), .A2(n5130), .ZN(n5199) );
  AOI22_X1 U6316 ( .A1(n5199), .A2(n6701), .B1(n6700), .B2(n5198), .ZN(n5133)
         );
  NAND2_X1 U6317 ( .A1(n6478), .A2(n6704), .ZN(n5132) );
  OAI211_X1 U6318 ( .C1(n5197), .C2(n6709), .A(n5133), .B(n5132), .ZN(n5134)
         );
  AOI21_X1 U6319 ( .B1(n5204), .B2(INSTQUEUE_REG_2__7__SCAN_IN), .A(n5134), 
        .ZN(n5135) );
  INV_X1 U6320 ( .A(n5135), .ZN(U3043) );
  AOI22_X1 U6321 ( .A1(n5199), .A2(n6660), .B1(n6603), .B2(n5198), .ZN(n5137)
         );
  NAND2_X1 U6322 ( .A1(n6478), .A2(n6604), .ZN(n5136) );
  OAI211_X1 U6323 ( .C1(n5197), .C2(n6658), .A(n5137), .B(n5136), .ZN(n5138)
         );
  AOI21_X1 U6324 ( .B1(n5204), .B2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n5138), 
        .ZN(n5139) );
  INV_X1 U6325 ( .A(n5139), .ZN(U3039) );
  AOI22_X1 U6326 ( .A1(n5199), .A2(n6653), .B1(n6599), .B2(n5198), .ZN(n5141)
         );
  NAND2_X1 U6327 ( .A1(n6478), .A2(n6600), .ZN(n5140) );
  OAI211_X1 U6328 ( .C1(n5197), .C2(n6656), .A(n5141), .B(n5140), .ZN(n5142)
         );
  AOI21_X1 U6329 ( .B1(n5204), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n5142), 
        .ZN(n5143) );
  INV_X1 U6330 ( .A(n5143), .ZN(U3038) );
  AOI22_X1 U6331 ( .A1(n5199), .A2(n6694), .B1(n6693), .B2(n5198), .ZN(n5145)
         );
  NAND2_X1 U6332 ( .A1(n6478), .A2(n6695), .ZN(n5144) );
  OAI211_X1 U6333 ( .C1(n5197), .C2(n6698), .A(n5145), .B(n5144), .ZN(n5146)
         );
  AOI21_X1 U6334 ( .B1(n5204), .B2(INSTQUEUE_REG_2__6__SCAN_IN), .A(n5146), 
        .ZN(n5147) );
  INV_X1 U6335 ( .A(n5147), .ZN(U3042) );
  AOI22_X1 U6336 ( .A1(n5199), .A2(n6720), .B1(n6718), .B2(n5198), .ZN(n5149)
         );
  NAND2_X1 U6337 ( .A1(n6478), .A2(n6722), .ZN(n5148) );
  OAI211_X1 U6338 ( .C1(n5197), .C2(n6669), .A(n5149), .B(n5148), .ZN(n5150)
         );
  AOI21_X1 U6339 ( .B1(n5204), .B2(INSTQUEUE_REG_2__4__SCAN_IN), .A(n5150), 
        .ZN(n5151) );
  INV_X1 U6340 ( .A(n5151), .ZN(U3040) );
  AOI22_X1 U6341 ( .A1(n5199), .A2(n6673), .B1(n6609), .B2(n5198), .ZN(n5153)
         );
  NAND2_X1 U6342 ( .A1(n6478), .A2(n6610), .ZN(n5152) );
  OAI211_X1 U6343 ( .C1(n5197), .C2(n6676), .A(n5153), .B(n5152), .ZN(n5154)
         );
  AOI21_X1 U6344 ( .B1(n5204), .B2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n5154), 
        .ZN(n5155) );
  INV_X1 U6345 ( .A(n5155), .ZN(U3041) );
  AOI22_X1 U6346 ( .A1(n5199), .A2(n6646), .B1(n6595), .B2(n5198), .ZN(n5157)
         );
  NAND2_X1 U6347 ( .A1(n6478), .A2(n6596), .ZN(n5156) );
  OAI211_X1 U6348 ( .C1(n5197), .C2(n6644), .A(n5157), .B(n5156), .ZN(n5158)
         );
  AOI21_X1 U6349 ( .B1(n5204), .B2(INSTQUEUE_REG_2__1__SCAN_IN), .A(n5158), 
        .ZN(n5159) );
  INV_X1 U6350 ( .A(n5159), .ZN(U3037) );
  INV_X1 U6351 ( .A(n5165), .ZN(n5160) );
  AOI21_X1 U6352 ( .B1(n5160), .B2(STATEBS16_REG_SCAN_IN), .A(n6636), .ZN(
        n5168) );
  NOR2_X1 U6353 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5161) );
  AND2_X1 U6354 ( .A1(n5161), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6583)
         );
  NAND2_X1 U6355 ( .A1(n6583), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5210) );
  OAI21_X1 U6356 ( .B1(n5162), .B2(n6586), .A(n5210), .ZN(n5171) );
  NOR2_X1 U6357 ( .A1(n5165), .A2(n5163), .ZN(n6149) );
  NOR2_X1 U6358 ( .A1(n6683), .A2(n5210), .ZN(n5167) );
  NOR2_X1 U6359 ( .A1(n5211), .A2(n6709), .ZN(n5166) );
  AOI211_X1 U6360 ( .C1(n6704), .C2(n6149), .A(n5167), .B(n5166), .ZN(n5174)
         );
  INV_X1 U6361 ( .A(n5168), .ZN(n5172) );
  INV_X1 U6362 ( .A(n6583), .ZN(n5169) );
  AOI21_X1 U6363 ( .B1(n5169), .B2(n6636), .A(n6634), .ZN(n5170) );
  NAND2_X1 U6364 ( .A1(n5214), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5173) );
  OAI211_X1 U6365 ( .C1(n5217), .C2(n5175), .A(n5174), .B(n5173), .ZN(U3099)
         );
  NOR2_X1 U6366 ( .A1(n6650), .A2(n5210), .ZN(n5177) );
  NOR2_X1 U6367 ( .A1(n5211), .A2(n6656), .ZN(n5176) );
  AOI211_X1 U6368 ( .C1(n6600), .C2(n6149), .A(n5177), .B(n5176), .ZN(n5179)
         );
  NAND2_X1 U6369 ( .A1(n5214), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5178) );
  OAI211_X1 U6370 ( .C1(n5217), .C2(n6207), .A(n5179), .B(n5178), .ZN(U3094)
         );
  NOR2_X1 U6371 ( .A1(n6657), .A2(n5210), .ZN(n5181) );
  NOR2_X1 U6372 ( .A1(n5211), .A2(n6658), .ZN(n5180) );
  AOI211_X1 U6373 ( .C1(n6604), .C2(n6149), .A(n5181), .B(n5180), .ZN(n5183)
         );
  NAND2_X1 U6374 ( .A1(n5214), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5182) );
  OAI211_X1 U6375 ( .C1(n5217), .C2(n6211), .A(n5183), .B(n5182), .ZN(U3095)
         );
  NOR2_X1 U6376 ( .A1(n6643), .A2(n5210), .ZN(n5185) );
  NOR2_X1 U6377 ( .A1(n5211), .A2(n6644), .ZN(n5184) );
  AOI211_X1 U6378 ( .C1(n6596), .C2(n6149), .A(n5185), .B(n5184), .ZN(n5187)
         );
  NAND2_X1 U6379 ( .A1(n5214), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5186) );
  OAI211_X1 U6380 ( .C1(n5217), .C2(n6203), .A(n5187), .B(n5186), .ZN(U3093)
         );
  NOR2_X1 U6381 ( .A1(n6677), .A2(n5210), .ZN(n5189) );
  NOR2_X1 U6382 ( .A1(n5211), .A2(n6698), .ZN(n5188) );
  AOI211_X1 U6383 ( .C1(n6695), .C2(n6149), .A(n5189), .B(n5188), .ZN(n5191)
         );
  NAND2_X1 U6384 ( .A1(n5214), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5190) );
  OAI211_X1 U6385 ( .C1(n5217), .C2(n5192), .A(n5191), .B(n5190), .ZN(U3098)
         );
  NOR2_X1 U6386 ( .A1(n6670), .A2(n5210), .ZN(n5194) );
  NOR2_X1 U6387 ( .A1(n5211), .A2(n6676), .ZN(n5193) );
  AOI211_X1 U6388 ( .C1(n6610), .C2(n6149), .A(n5194), .B(n5193), .ZN(n5196)
         );
  NAND2_X1 U6389 ( .A1(n5214), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5195) );
  OAI211_X1 U6390 ( .C1(n5217), .C2(n6219), .A(n5196), .B(n5195), .ZN(U3097)
         );
  NOR2_X1 U6391 ( .A1(n5197), .A2(n6624), .ZN(n5203) );
  AOI22_X1 U6392 ( .A1(n5199), .A2(n6712), .B1(n6711), .B2(n5198), .ZN(n5200)
         );
  OAI21_X1 U6393 ( .B1(n5201), .B2(n6642), .A(n5200), .ZN(n5202) );
  AOI211_X1 U6394 ( .C1(n5204), .C2(INSTQUEUE_REG_2__0__SCAN_IN), .A(n5203), 
        .B(n5202), .ZN(n5205) );
  INV_X1 U6395 ( .A(n5205), .ZN(U3036) );
  NOR2_X1 U6396 ( .A1(n6623), .A2(n5210), .ZN(n5207) );
  NOR2_X1 U6397 ( .A1(n5211), .A2(n6624), .ZN(n5206) );
  AOI211_X1 U6398 ( .C1(n6714), .C2(n6149), .A(n5207), .B(n5206), .ZN(n5209)
         );
  NAND2_X1 U6399 ( .A1(n5214), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5208) );
  OAI211_X1 U6400 ( .C1(n5217), .C2(n6199), .A(n5209), .B(n5208), .ZN(U3092)
         );
  NOR2_X1 U6401 ( .A1(n6664), .A2(n5210), .ZN(n5213) );
  NOR2_X1 U6402 ( .A1(n5211), .A2(n6669), .ZN(n5212) );
  AOI211_X1 U6403 ( .C1(n6722), .C2(n6149), .A(n5213), .B(n5212), .ZN(n5216)
         );
  NAND2_X1 U6404 ( .A1(n5214), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5215) );
  OAI211_X1 U6405 ( .C1(n5217), .C2(n6215), .A(n5216), .B(n5215), .ZN(U3096)
         );
  INV_X1 U6406 ( .A(n5067), .ZN(n5219) );
  INV_X1 U6407 ( .A(n4428), .ZN(n5218) );
  AOI21_X1 U6408 ( .B1(n5220), .B2(n5219), .A(n5218), .ZN(n6277) );
  INV_X1 U6409 ( .A(n6277), .ZN(n5227) );
  AOI22_X1 U6410 ( .A1(n5681), .A2(DATAI_7_), .B1(EAX_REG_7__SCAN_IN), .B2(
        n5680), .ZN(n5221) );
  OAI21_X1 U6411 ( .B1(n5227), .B2(n5683), .A(n5221), .ZN(U2884) );
  INV_X1 U6412 ( .A(n5223), .ZN(n5224) );
  AOI21_X1 U6413 ( .B1(n5225), .B2(n5222), .A(n5224), .ZN(n6276) );
  AOI22_X1 U6414 ( .A1(n6276), .A2(n4234), .B1(n5607), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5226) );
  OAI21_X1 U6415 ( .B1(n5227), .B2(n7064), .A(n5226), .ZN(U2852) );
  XNOR2_X1 U6416 ( .A(n5228), .B(n5229), .ZN(n5241) );
  NAND2_X1 U6417 ( .A1(n6399), .A2(REIP_REG_6__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6418 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5230)
         );
  OAI211_X1 U6419 ( .C1(n6418), .C2(n6302), .A(n5236), .B(n5230), .ZN(n5231)
         );
  AOI21_X1 U6420 ( .B1(n6298), .B2(n6404), .A(n5231), .ZN(n5232) );
  OAI21_X1 U6421 ( .B1(n6226), .B2(n5241), .A(n5232), .ZN(U2980) );
  INV_X1 U6422 ( .A(n5222), .ZN(n5233) );
  AOI21_X1 U6423 ( .B1(n5234), .B2(n4997), .A(n5233), .ZN(n6293) );
  INV_X1 U6424 ( .A(n6293), .ZN(n7066) );
  NAND3_X1 U6425 ( .A1(n5251), .A2(n4295), .A3(n5235), .ZN(n5237) );
  OAI211_X1 U6426 ( .C1(n6455), .C2(n7066), .A(n5237), .B(n5236), .ZN(n5238)
         );
  AOI21_X1 U6427 ( .B1(n5239), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5238), 
        .ZN(n5240) );
  OAI21_X1 U6428 ( .B1(n6422), .B2(n5241), .A(n5240), .ZN(U3012) );
  INV_X1 U6429 ( .A(n6109), .ZN(n5242) );
  AOI22_X1 U6430 ( .A1(n5242), .A2(n4234), .B1(n5607), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5243) );
  OAI21_X1 U6431 ( .B1(n5245), .B2(n7064), .A(n5243), .ZN(U2851) );
  AOI22_X1 U6432 ( .A1(n5681), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5680), .ZN(n5244) );
  OAI21_X1 U6433 ( .B1(n5245), .B2(n5683), .A(n5244), .ZN(U2883) );
  XNOR2_X1 U6434 ( .A(n5246), .B(n5247), .ZN(n5260) );
  NOR2_X1 U6435 ( .A1(n6418), .A2(n6291), .ZN(n5249) );
  INV_X1 U6436 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U6437 ( .A1(n6399), .A2(REIP_REG_7__SCAN_IN), .ZN(n5254) );
  OAI21_X1 U6438 ( .B1(n5868), .B2(n6280), .A(n5254), .ZN(n5248) );
  AOI211_X1 U6439 ( .C1(n6277), .C2(n6404), .A(n5249), .B(n5248), .ZN(n5250)
         );
  OAI21_X1 U6440 ( .B1(n6226), .B2(n5260), .A(n5250), .ZN(U2979) );
  NAND2_X1 U6441 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5251), .ZN(n5888)
         );
  NOR2_X1 U6442 ( .A1(n5252), .A2(n5888), .ZN(n5253) );
  OAI21_X1 U6443 ( .B1(n6010), .B2(n5253), .A(n6450), .ZN(n6419) );
  INV_X1 U6444 ( .A(n6276), .ZN(n5255) );
  OAI21_X1 U6445 ( .B1(n5255), .B2(n6455), .A(n5254), .ZN(n5258) );
  NOR2_X1 U6446 ( .A1(n6425), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5257)
         );
  AOI211_X1 U6447 ( .C1(n6419), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5258), 
        .B(n5257), .ZN(n5259) );
  OAI21_X1 U6448 ( .B1(n6422), .B2(n5260), .A(n5259), .ZN(U3011) );
  AOI21_X1 U6449 ( .B1(n5261), .B2(n6123), .A(n6129), .ZN(n5269) );
  OAI21_X1 U6450 ( .B1(n5264), .B2(STATE2_REG_3__SCAN_IN), .A(n5263), .ZN(
        n5266) );
  AOI22_X1 U6451 ( .A1(n5267), .A2(n5262), .B1(n5266), .B2(n5265), .ZN(n5268)
         );
  OAI22_X1 U6452 ( .A1(n5269), .A2(n5262), .B1(n6129), .B2(n5268), .ZN(U3461)
         );
  AOI22_X1 U6453 ( .A1(n5680), .A2(EAX_REG_29__SCAN_IN), .B1(n5661), .B2(
        DATAI_29_), .ZN(n5271) );
  NAND2_X1 U6454 ( .A1(n5662), .A2(DATAI_13_), .ZN(n5270) );
  OAI211_X1 U6455 ( .C1(n5312), .C2(n5683), .A(n5271), .B(n5270), .ZN(U2862)
         );
  INV_X1 U6456 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5316) );
  NOR2_X1 U6457 ( .A1(n5272), .A2(EBX_REG_29__SCAN_IN), .ZN(n5275) );
  AOI22_X1 U6458 ( .A1(n5274), .A2(n5424), .B1(n5275), .B2(n5273), .ZN(n5294)
         );
  INV_X1 U6459 ( .A(n5275), .ZN(n5276) );
  OAI211_X1 U6460 ( .C1(n5439), .C2(n5277), .A(n5324), .B(n5276), .ZN(n5278)
         );
  NAND2_X1 U6461 ( .A1(n5294), .A2(n5278), .ZN(n5937) );
  OAI222_X1 U6462 ( .A1(n5316), .A2(n5628), .B1(n7065), .B2(n5937), .C1(n5312), 
        .C2(n7064), .ZN(U2830) );
  AOI211_X1 U6463 ( .C1(n5280), .C2(n6225), .A(n6632), .B(n5279), .ZN(n5283)
         );
  OAI21_X1 U6464 ( .B1(n5283), .B2(n5282), .A(n5281), .ZN(n5288) );
  INV_X1 U6465 ( .A(n6756), .ZN(n5286) );
  AOI211_X1 U6466 ( .C1(n7019), .C2(n6374), .A(n6626), .B(n5284), .ZN(n5285)
         );
  NAND2_X1 U6467 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  MUX2_X1 U6468 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n5288), .S(n5287), .Z(
        U3472) );
  AND2_X1 U6469 ( .A1(n5289), .A2(n6729), .ZN(n6228) );
  MUX2_X1 U6470 ( .A(MORE_REG_SCAN_IN), .B(n5290), .S(n6228), .Z(U3471) );
  INV_X1 U6471 ( .A(n5291), .ZN(n5311) );
  OAI21_X1 U6472 ( .B1(n5294), .B2(n5293), .A(n5292), .ZN(n5295) );
  INV_X1 U6473 ( .A(n5295), .ZN(n5299) );
  AOI22_X1 U6474 ( .A1(n5297), .A2(EBX_REG_31__SCAN_IN), .B1(n5296), .B2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5298) );
  INV_X1 U6475 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5302) );
  AOI21_X1 U6476 ( .B1(n5301), .B2(n5300), .A(n5302), .ZN(n5309) );
  NAND4_X1 U6477 ( .A1(n5303), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n5302), .ZN(n5306) );
  NAND3_X1 U6478 ( .A1(n5557), .A2(EBX_REG_31__SCAN_IN), .A3(n5304), .ZN(n5305) );
  OAI211_X1 U6479 ( .C1(n5307), .C2(n6307), .A(n5306), .B(n5305), .ZN(n5308)
         );
  OAI21_X1 U6480 ( .B1(n5311), .B2(n5554), .A(n5310), .ZN(U2796) );
  NAND2_X1 U6481 ( .A1(n5313), .A2(n6299), .ZN(n5320) );
  INV_X1 U6482 ( .A(n3103), .ZN(n6262) );
  AOI22_X1 U6483 ( .A1(n6262), .A2(n5314), .B1(PHYADDRPOINTER_REG_29__SCAN_IN), 
        .B2(n6330), .ZN(n5315) );
  OAI21_X1 U6484 ( .B1(n6294), .B2(n5316), .A(n5315), .ZN(n5318) );
  AOI211_X1 U6485 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5327), .A(n5318), .B(n5317), .ZN(n5319) );
  OAI211_X1 U6486 ( .C1(n5937), .C2(n6334), .A(n5320), .B(n5319), .ZN(U2798)
         );
  NAND2_X1 U6487 ( .A1(n5321), .A2(n5322), .ZN(n5323) );
  NAND2_X1 U6488 ( .A1(n5324), .A2(n5323), .ZN(n5945) );
  NAND2_X1 U6489 ( .A1(n5705), .A2(n6299), .ZN(n5335) );
  INV_X1 U6490 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6491 ( .A1(n5327), .A2(REIP_REG_28__SCAN_IN), .ZN(n5329) );
  AOI22_X1 U6492 ( .A1(n6262), .A2(n5701), .B1(PHYADDRPOINTER_REG_28__SCAN_IN), 
        .B2(n6330), .ZN(n5328) );
  OAI211_X1 U6493 ( .C1(n5598), .C2(n6294), .A(n5329), .B(n5328), .ZN(n5333)
         );
  NAND2_X1 U6494 ( .A1(n5330), .A2(REIP_REG_27__SCAN_IN), .ZN(n5331) );
  NOR2_X1 U6495 ( .A1(n5342), .A2(n5331), .ZN(n5332) );
  NOR2_X1 U6496 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  OAI211_X1 U6497 ( .C1(n5945), .C2(n6334), .A(n5335), .B(n5334), .ZN(U2799)
         );
  OR2_X1 U6498 ( .A1(n5338), .A2(n5339), .ZN(n5340) );
  NAND2_X1 U6499 ( .A1(n5321), .A2(n5340), .ZN(n5958) );
  INV_X1 U6500 ( .A(n5958), .ZN(n5344) );
  NOR2_X1 U6501 ( .A1(n6294), .A2(n5599), .ZN(n5341) );
  AOI21_X1 U6502 ( .B1(n5344), .B2(n6305), .A(n5343), .ZN(n5345) );
  OAI21_X1 U6503 ( .B1(n5715), .B2(n5554), .A(n5345), .ZN(U2800) );
  INV_X1 U6504 ( .A(n5336), .ZN(n5347) );
  OR3_X1 U6505 ( .A1(n5414), .A2(n5367), .A3(n4466), .ZN(n5366) );
  OAI21_X1 U6506 ( .B1(n5366), .B2(n5368), .A(n6934), .ZN(n5356) );
  NAND2_X1 U6507 ( .A1(n6319), .A2(EBX_REG_26__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6508 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5349)
         );
  OAI211_X1 U6509 ( .C1(n3104), .C2(n5716), .A(n5350), .B(n5349), .ZN(n5355)
         );
  INV_X1 U6510 ( .A(n5338), .ZN(n5352) );
  OAI21_X1 U6511 ( .B1(n5351), .B2(n5353), .A(n5352), .ZN(n5966) );
  NOR2_X1 U6512 ( .A1(n5966), .A2(n6334), .ZN(n5354) );
  AOI211_X1 U6513 ( .C1(n5357), .C2(n5356), .A(n5355), .B(n5354), .ZN(n5358)
         );
  OAI21_X1 U6514 ( .B1(n5722), .B2(n5554), .A(n5358), .ZN(U2801) );
  NOR2_X1 U6515 ( .A1(n5375), .A2(n5359), .ZN(n5360) );
  OR2_X1 U6516 ( .A1(n5351), .A2(n5360), .ZN(n5973) );
  AOI21_X1 U6517 ( .B1(n5362), .B2(n5361), .A(n5346), .ZN(n5600) );
  NAND2_X1 U6518 ( .A1(n5600), .A2(n6299), .ZN(n5372) );
  AOI22_X1 U6519 ( .A1(n6262), .A2(n5725), .B1(PHYADDRPOINTER_REG_25__SCAN_IN), 
        .B2(n6330), .ZN(n5365) );
  NAND2_X1 U6520 ( .A1(n6319), .A2(EBX_REG_25__SCAN_IN), .ZN(n5364) );
  OAI211_X1 U6521 ( .C1(n5366), .C2(REIP_REG_25__SCAN_IN), .A(n5365), .B(n5364), .ZN(n5370) );
  OR3_X1 U6522 ( .A1(n5414), .A2(REIP_REG_24__SCAN_IN), .A3(n5367), .ZN(n5379)
         );
  AOI21_X1 U6523 ( .B1(n5379), .B2(n5387), .A(n5368), .ZN(n5369) );
  NOR2_X1 U6524 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  OAI211_X1 U6525 ( .C1(n5973), .C2(n6334), .A(n5372), .B(n5371), .ZN(U2802)
         );
  OAI21_X1 U6526 ( .B1(n5373), .B2(n5374), .A(n5361), .ZN(n5738) );
  AOI21_X1 U6527 ( .B1(n5376), .B2(n5384), .A(n5375), .ZN(n5982) );
  INV_X1 U6528 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6785) );
  OAI22_X1 U6529 ( .A1(n5740), .A2(n3104), .B1(n6307), .B2(n6785), .ZN(n5377)
         );
  AOI21_X1 U6530 ( .B1(n6319), .B2(EBX_REG_24__SCAN_IN), .A(n5377), .ZN(n5378)
         );
  OAI211_X1 U6531 ( .C1(n5387), .C2(n4466), .A(n5379), .B(n5378), .ZN(n5380)
         );
  AOI21_X1 U6532 ( .B1(n5982), .B2(n6305), .A(n5380), .ZN(n5381) );
  OAI21_X1 U6533 ( .B1(n5738), .B2(n5554), .A(n5381), .ZN(U2803) );
  NAND2_X1 U6534 ( .A1(n5402), .A2(n5382), .ZN(n5383) );
  NAND2_X1 U6535 ( .A1(n5384), .A2(n5383), .ZN(n5987) );
  AOI21_X1 U6536 ( .B1(n5386), .B2(n5385), .A(n5373), .ZN(n5750) );
  NAND2_X1 U6537 ( .A1(n5750), .A2(n6299), .ZN(n5393) );
  OAI22_X1 U6538 ( .A1(n5748), .A2(n3105), .B1(n6307), .B2(n3142), .ZN(n5391)
         );
  INV_X1 U6539 ( .A(n5414), .ZN(n5407) );
  NAND3_X1 U6540 ( .A1(n5407), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5389) );
  AOI21_X1 U6541 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n5390) );
  AOI211_X1 U6542 ( .C1(EBX_REG_23__SCAN_IN), .C2(n6319), .A(n5391), .B(n5390), 
        .ZN(n5392) );
  OAI211_X1 U6543 ( .C1(n5987), .C2(n6334), .A(n5393), .B(n5392), .ZN(U2804)
         );
  OAI21_X1 U6544 ( .B1(n5394), .B2(n5395), .A(n5385), .ZN(n5760) );
  XOR2_X1 U6545 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .Z(n5406) );
  NAND2_X1 U6546 ( .A1(n5427), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U6547 ( .A1(n5594), .A2(n5397), .ZN(n5431) );
  OAI22_X1 U6548 ( .A1(n5756), .A2(n3105), .B1(n6307), .B2(n5398), .ZN(n5399)
         );
  AOI21_X1 U6549 ( .B1(n6319), .B2(EBX_REG_22__SCAN_IN), .A(n5399), .ZN(n5400)
         );
  OAI21_X1 U6550 ( .B1(n5755), .B2(n5431), .A(n5400), .ZN(n5405) );
  INV_X1 U6551 ( .A(n5401), .ZN(n5403) );
  OAI21_X1 U6552 ( .B1(n5403), .B2(n3132), .A(n5402), .ZN(n5999) );
  NOR2_X1 U6553 ( .A1(n5999), .A2(n6334), .ZN(n5404) );
  AOI211_X1 U6554 ( .C1(n5407), .C2(n5406), .A(n5405), .B(n5404), .ZN(n5408)
         );
  OAI21_X1 U6555 ( .B1(n5760), .B2(n5554), .A(n5408), .ZN(U2805) );
  OAI21_X1 U6556 ( .B1(n5410), .B2(n5409), .A(n5401), .ZN(n6008) );
  AOI21_X1 U6557 ( .B1(n5412), .B2(n5411), .A(n5394), .ZN(n5603) );
  NAND2_X1 U6558 ( .A1(n5603), .A2(n6299), .ZN(n5419) );
  INV_X1 U6559 ( .A(n5431), .ZN(n5417) );
  INV_X1 U6560 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5604) );
  AOI22_X1 U6561 ( .A1(n6262), .A2(n5763), .B1(PHYADDRPOINTER_REG_21__SCAN_IN), 
        .B2(n6330), .ZN(n5413) );
  OAI21_X1 U6562 ( .B1(n6294), .B2(n5604), .A(n5413), .ZN(n5416) );
  NOR2_X1 U6563 ( .A1(n5414), .A2(REIP_REG_21__SCAN_IN), .ZN(n5415) );
  AOI211_X1 U6564 ( .C1(n5417), .C2(REIP_REG_21__SCAN_IN), .A(n5416), .B(n5415), .ZN(n5418) );
  OAI211_X1 U6565 ( .C1(n6008), .C2(n6334), .A(n5419), .B(n5418), .ZN(U2806)
         );
  INV_X1 U6566 ( .A(n5411), .ZN(n5421) );
  AOI21_X1 U6567 ( .B1(n5422), .B2(n5420), .A(n5421), .ZN(n5775) );
  INV_X1 U6568 ( .A(n5775), .ZN(n5652) );
  MUX2_X1 U6569 ( .A(n5441), .B(n5424), .S(n5423), .Z(n5426) );
  XNOR2_X1 U6570 ( .A(n5426), .B(n5425), .ZN(n5605) );
  INV_X1 U6571 ( .A(n5605), .ZN(n6016) );
  AOI21_X1 U6572 ( .B1(n5459), .B2(n5427), .A(REIP_REG_20__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6573 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5428)
         );
  OAI21_X1 U6574 ( .B1(n3104), .B2(n5772), .A(n5428), .ZN(n5429) );
  AOI21_X1 U6575 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6319), .A(n5429), .ZN(n5430)
         );
  OAI21_X1 U6576 ( .B1(n5432), .B2(n5431), .A(n5430), .ZN(n5433) );
  AOI21_X1 U6577 ( .B1(n6016), .B2(n6305), .A(n5433), .ZN(n5434) );
  OAI21_X1 U6578 ( .B1(n5652), .B2(n5554), .A(n5434), .ZN(U2807) );
  OR2_X1 U6579 ( .A1(n5435), .A2(n5436), .ZN(n5437) );
  NAND2_X1 U6580 ( .A1(n5420), .A2(n5437), .ZN(n5783) );
  MUX2_X1 U6581 ( .A(n5441), .B(n5440), .S(n5439), .Z(n5458) );
  NOR2_X1 U6582 ( .A1(n5438), .A2(n5458), .ZN(n5457) );
  XOR2_X1 U6583 ( .A(n5442), .B(n5457), .Z(n6027) );
  INV_X1 U6584 ( .A(n6027), .ZN(n5451) );
  INV_X1 U6585 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6586 ( .A1(n5594), .A2(n5444), .ZN(n5475) );
  OAI211_X1 U6587 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5459), .B(n5445), .ZN(n5449) );
  NAND2_X1 U6588 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5446)
         );
  OAI211_X1 U6589 ( .C1(n3104), .C2(n5779), .A(n5446), .B(n6321), .ZN(n5447)
         );
  AOI21_X1 U6590 ( .B1(n6319), .B2(EBX_REG_19__SCAN_IN), .A(n5447), .ZN(n5448)
         );
  OAI211_X1 U6591 ( .C1(n6811), .C2(n5475), .A(n5449), .B(n5448), .ZN(n5450)
         );
  AOI21_X1 U6592 ( .B1(n5451), .B2(n6305), .A(n5450), .ZN(n5452) );
  OAI21_X1 U6593 ( .B1(n5783), .B2(n5554), .A(n5452), .ZN(U2808) );
  INV_X1 U6594 ( .A(n5453), .ZN(n5456) );
  INV_X1 U6595 ( .A(n5454), .ZN(n5455) );
  AOI21_X1 U6596 ( .B1(n5456), .B2(n5455), .A(n5435), .ZN(n5789) );
  INV_X1 U6597 ( .A(n5789), .ZN(n5657) );
  AOI21_X1 U6598 ( .B1(n5438), .B2(n5458), .A(n5457), .ZN(n6034) );
  INV_X1 U6599 ( .A(n5459), .ZN(n5465) );
  NAND2_X1 U6600 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5460)
         );
  OAI211_X1 U6601 ( .C1(n3105), .C2(n5787), .A(n6321), .B(n5460), .ZN(n5463)
         );
  NOR2_X1 U6602 ( .A1(n5475), .A2(n5461), .ZN(n5462) );
  OAI21_X1 U6603 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5465), .A(n5464), .ZN(n5466) );
  AOI21_X1 U6604 ( .B1(n6034), .B2(n6305), .A(n5466), .ZN(n5467) );
  OAI21_X1 U6605 ( .B1(n5657), .B2(n5554), .A(n5467), .ZN(U2809) );
  OR2_X1 U6606 ( .A1(n5468), .A2(n5469), .ZN(n5470) );
  NAND2_X1 U6607 ( .A1(n5438), .A2(n5470), .ZN(n6039) );
  INV_X1 U6608 ( .A(n5471), .ZN(n5474) );
  INV_X1 U6609 ( .A(n5472), .ZN(n5473) );
  AOI21_X1 U6610 ( .B1(n5474), .B2(n5473), .A(n5454), .ZN(n5797) );
  NAND2_X1 U6611 ( .A1(n5797), .A2(n6299), .ZN(n5484) );
  INV_X1 U6612 ( .A(n5475), .ZN(n5482) );
  OAI21_X1 U6613 ( .B1(n7045), .B2(n5494), .A(n5476), .ZN(n5481) );
  INV_X1 U6614 ( .A(n5796), .ZN(n5478) );
  NAND2_X1 U6615 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5477)
         );
  OAI211_X1 U6616 ( .C1(n3105), .C2(n5478), .A(n6321), .B(n5477), .ZN(n5480)
         );
  NOR2_X1 U6617 ( .A1(n6294), .A2(n5609), .ZN(n5479) );
  AOI211_X1 U6618 ( .C1(n5482), .C2(n5481), .A(n5480), .B(n5479), .ZN(n5483)
         );
  OAI211_X1 U6619 ( .C1(n6039), .C2(n6334), .A(n5484), .B(n5483), .ZN(U2810)
         );
  NAND2_X1 U6620 ( .A1(n5485), .A2(n5516), .ZN(n5515) );
  AOI21_X1 U6621 ( .B1(n5486), .B2(n5501), .A(n5472), .ZN(n5809) );
  INV_X1 U6622 ( .A(n5809), .ZN(n5665) );
  NOR2_X1 U6623 ( .A1(n5497), .A2(n5487), .ZN(n5488) );
  OR2_X1 U6624 ( .A1(n5468), .A2(n5488), .ZN(n5611) );
  INV_X1 U6625 ( .A(n5611), .ZN(n6054) );
  NAND2_X1 U6626 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5489)
         );
  OAI211_X1 U6627 ( .C1(n3105), .C2(n5807), .A(n6321), .B(n5489), .ZN(n5490)
         );
  AOI21_X1 U6628 ( .B1(n6319), .B2(EBX_REG_16__SCAN_IN), .A(n5490), .ZN(n5493)
         );
  NAND3_X1 U6629 ( .A1(n5594), .A2(REIP_REG_16__SCAN_IN), .A3(n5491), .ZN(
        n5492) );
  OAI211_X1 U6630 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5494), .A(n5493), .B(n5492), .ZN(n5495) );
  AOI21_X1 U6631 ( .B1(n6054), .B2(n6305), .A(n5495), .ZN(n5496) );
  OAI21_X1 U6632 ( .B1(n5665), .B2(n5554), .A(n5496), .ZN(U2811) );
  AOI21_X1 U6633 ( .B1(n5498), .B2(n5514), .A(n5497), .ZN(n6062) );
  INV_X1 U6634 ( .A(n6062), .ZN(n5612) );
  NAND2_X1 U6635 ( .A1(n5515), .A2(n5499), .ZN(n5500) );
  NAND2_X1 U6636 ( .A1(n5819), .A2(n6299), .ZN(n5510) );
  INV_X1 U6637 ( .A(n5594), .ZN(n5563) );
  NOR2_X1 U6638 ( .A1(n5563), .A2(n5502), .ZN(n5523) );
  NAND2_X1 U6639 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5503)
         );
  OAI211_X1 U6640 ( .C1(n3104), .C2(n5817), .A(n6321), .B(n5503), .ZN(n5508)
         );
  INV_X1 U6641 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6839) );
  NAND3_X1 U6642 ( .A1(n6320), .A2(n5505), .A3(n5504), .ZN(n5506) );
  OAI21_X1 U6643 ( .B1(n6294), .B2(n6839), .A(n5506), .ZN(n5507) );
  AOI211_X1 U6644 ( .C1(n5523), .C2(REIP_REG_15__SCAN_IN), .A(n5508), .B(n5507), .ZN(n5509) );
  OAI211_X1 U6645 ( .C1(n5612), .C2(n6334), .A(n5510), .B(n5509), .ZN(U2812)
         );
  NAND2_X1 U6646 ( .A1(n5511), .A2(n5512), .ZN(n5513) );
  NAND2_X1 U6647 ( .A1(n5514), .A2(n5513), .ZN(n6067) );
  OAI21_X1 U6648 ( .B1(n5485), .B2(n5516), .A(n5515), .ZN(n5669) );
  INV_X1 U6649 ( .A(n5669), .ZN(n5827) );
  NAND2_X1 U6650 ( .A1(n5827), .A2(n6299), .ZN(n5525) );
  NAND2_X1 U6651 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5517)
         );
  OAI211_X1 U6652 ( .C1(n3105), .C2(n5825), .A(n6321), .B(n5517), .ZN(n5522)
         );
  NAND3_X1 U6653 ( .A1(n6320), .A2(n5519), .A3(n5518), .ZN(n5520) );
  OAI21_X1 U6654 ( .B1(n6294), .B2(n6825), .A(n5520), .ZN(n5521) );
  AOI211_X1 U6655 ( .C1(n5523), .C2(REIP_REG_14__SCAN_IN), .A(n5522), .B(n5521), .ZN(n5524) );
  OAI211_X1 U6656 ( .C1(n6067), .C2(n6334), .A(n5525), .B(n5524), .ZN(U2813)
         );
  XOR2_X1 U6657 ( .A(n5527), .B(n5526), .Z(n5842) );
  AND2_X1 U6658 ( .A1(n6320), .A2(n5536), .ZN(n6256) );
  INV_X1 U6659 ( .A(n6256), .ZN(n5528) );
  NAND2_X1 U6660 ( .A1(n5528), .A2(n6278), .ZN(n6260) );
  INV_X1 U6661 ( .A(n5841), .ZN(n5535) );
  INV_X1 U6662 ( .A(n6321), .ZN(n6283) );
  INV_X1 U6663 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5620) );
  NOR2_X1 U6664 ( .A1(n5620), .A2(n6294), .ZN(n5533) );
  NOR2_X1 U6665 ( .A1(n5529), .A2(n5530), .ZN(n5531) );
  OR2_X1 U6666 ( .A1(n5616), .A2(n5531), .ZN(n6088) );
  OAI22_X1 U6667 ( .A1(n5839), .A2(n6307), .B1(n6334), .B2(n6088), .ZN(n5532)
         );
  NOR3_X1 U6668 ( .A1(n6283), .A2(n5533), .A3(n5532), .ZN(n5534) );
  OAI21_X1 U6669 ( .B1(n5535), .B2(n3105), .A(n5534), .ZN(n5537) );
  NOR3_X1 U6670 ( .A1(n6285), .A2(REIP_REG_12__SCAN_IN), .A3(n5536), .ZN(n6252) );
  AOI211_X1 U6671 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6260), .A(n5537), .B(n6252), .ZN(n5538) );
  OAI21_X1 U6672 ( .B1(n5672), .B2(n5554), .A(n5538), .ZN(U2815) );
  INV_X1 U6673 ( .A(n5539), .ZN(n5541) );
  NAND2_X1 U6674 ( .A1(n5622), .A2(n5621), .ZN(n5624) );
  INV_X1 U6675 ( .A(n5675), .ZN(n5540) );
  AOI21_X1 U6676 ( .B1(n5541), .B2(n5624), .A(n5540), .ZN(n5862) );
  NOR3_X1 U6677 ( .A1(n6285), .A2(REIP_REG_9__SCAN_IN), .A3(n5542), .ZN(n6269)
         );
  OAI21_X1 U6678 ( .B1(n6269), .B2(n6267), .A(REIP_REG_10__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6679 ( .A1(n5625), .A2(n5543), .ZN(n5544) );
  NAND2_X1 U6680 ( .A1(n6100), .A2(n5544), .ZN(n6423) );
  OAI22_X1 U6681 ( .A1(n4170), .A2(n6294), .B1(n6334), .B2(n6423), .ZN(n5548)
         );
  NAND3_X1 U6682 ( .A1(n6320), .A2(n4474), .A3(n5545), .ZN(n5546) );
  OAI211_X1 U6683 ( .C1(n6307), .C2(n6809), .A(n6321), .B(n5546), .ZN(n5547)
         );
  NOR2_X1 U6684 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  OAI211_X1 U6685 ( .C1(n3104), .C2(n5860), .A(n5550), .B(n5549), .ZN(n5551)
         );
  AOI21_X1 U6686 ( .B1(n5862), .B2(n6299), .A(n5551), .ZN(n5552) );
  INV_X1 U6687 ( .A(n5552), .ZN(U2817) );
  NAND2_X1 U6688 ( .A1(n5557), .A2(n6753), .ZN(n5553) );
  NAND2_X1 U6689 ( .A1(n5554), .A2(n5553), .ZN(n6309) );
  INV_X1 U6690 ( .A(n5555), .ZN(n5556) );
  AND2_X1 U6691 ( .A1(n5557), .A2(n5556), .ZN(n6318) );
  NAND2_X1 U6692 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5558)
         );
  OAI21_X1 U6693 ( .B1(n3104), .B2(n5559), .A(n5558), .ZN(n5562) );
  OAI22_X1 U6694 ( .A1(n6334), .A2(n5560), .B1(n6294), .B2(n3205), .ZN(n5561)
         );
  AOI211_X1 U6695 ( .C1(n6318), .C2(n6141), .A(n5562), .B(n5561), .ZN(n5570)
         );
  AOI21_X1 U6696 ( .B1(n6278), .B2(REIP_REG_1__SCAN_IN), .A(n5563), .ZN(n5564)
         );
  NOR2_X1 U6697 ( .A1(n5564), .A2(n6444), .ZN(n5581) );
  INV_X1 U6698 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U6699 ( .A1(n6278), .A2(n5566), .ZN(n5567) );
  NAND2_X1 U6700 ( .A1(n5594), .A2(n5567), .ZN(n6322) );
  INV_X1 U6701 ( .A(n6322), .ZN(n5568) );
  OAI21_X1 U6702 ( .B1(n5581), .B2(REIP_REG_3__SCAN_IN), .A(n5568), .ZN(n5569)
         );
  OAI211_X1 U6703 ( .C1(n5571), .C2(n6326), .A(n5570), .B(n5569), .ZN(U2824)
         );
  AOI21_X1 U6704 ( .B1(n6320), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5580) );
  OAI22_X1 U6705 ( .A1(n6408), .A2(n3104), .B1(n6307), .B2(n5572), .ZN(n5576)
         );
  XNOR2_X1 U6706 ( .A(n4650), .B(n5573), .ZN(n6340) );
  INV_X1 U6707 ( .A(n6340), .ZN(n6445) );
  INV_X1 U6708 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5574) );
  OAI22_X1 U6709 ( .A1(n6445), .A2(n6334), .B1(n6294), .B2(n5574), .ZN(n5575)
         );
  AOI211_X1 U6710 ( .C1(n6318), .C2(n5577), .A(n5576), .B(n5575), .ZN(n5579)
         );
  NAND2_X1 U6711 ( .A1(n6405), .A2(n6309), .ZN(n5578) );
  OAI211_X1 U6712 ( .C1(n5581), .C2(n5580), .A(n5579), .B(n5578), .ZN(U2825)
         );
  AOI22_X1 U6713 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6319), .B1(n6305), .B2(n4582), 
        .ZN(n5588) );
  AOI22_X1 U6714 ( .A1(n5582), .A2(n6318), .B1(n6320), .B2(n6742), .ZN(n5585)
         );
  INV_X1 U6715 ( .A(n6278), .ZN(n5583) );
  AOI22_X1 U6716 ( .A1(n6330), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5583), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5584) );
  OAI211_X1 U6717 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n3105), .A(n5585), 
        .B(n5584), .ZN(n5586) );
  INV_X1 U6718 ( .A(n5586), .ZN(n5587) );
  OAI211_X1 U6719 ( .C1(n6411), .C2(n6326), .A(n5588), .B(n5587), .ZN(U2826)
         );
  INV_X1 U6720 ( .A(n6318), .ZN(n5590) );
  OAI21_X1 U6721 ( .B1(n6262), .B2(n6330), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5589) );
  OAI21_X1 U6722 ( .B1(n5590), .B2(n6629), .A(n5589), .ZN(n5593) );
  OAI22_X1 U6723 ( .A1(n5591), .A2(n6294), .B1(n6334), .B2(n6454), .ZN(n5592)
         );
  AOI211_X1 U6724 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5594), .A(n5593), .B(n5592), 
        .ZN(n5595) );
  OAI21_X1 U6725 ( .B1(n6326), .B2(n5881), .A(n5595), .ZN(U2827) );
  INV_X1 U6726 ( .A(n5924), .ZN(n5597) );
  OAI22_X1 U6727 ( .A1(n5597), .A2(n7065), .B1(n5596), .B2(n5628), .ZN(U2828)
         );
  INV_X1 U6728 ( .A(n5705), .ZN(n5634) );
  OAI222_X1 U6729 ( .A1(n5599), .A2(n5628), .B1(n7065), .B2(n5958), .C1(n5715), 
        .C2(n7064), .ZN(U2832) );
  INV_X1 U6730 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6998) );
  OAI222_X1 U6731 ( .A1(n5966), .A2(n7065), .B1(n6998), .B2(n5628), .C1(n5722), 
        .C2(n7064), .ZN(U2833) );
  INV_X1 U6732 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6884) );
  INV_X1 U6733 ( .A(n5600), .ZN(n5731) );
  OAI222_X1 U6734 ( .A1(n5973), .A2(n7065), .B1(n6884), .B2(n5628), .C1(n5731), 
        .C2(n7064), .ZN(U2834) );
  INV_X1 U6735 ( .A(n5982), .ZN(n5601) );
  OAI222_X1 U6736 ( .A1(n6850), .A2(n5628), .B1(n7065), .B2(n5601), .C1(n5738), 
        .C2(n7064), .ZN(U2835) );
  INV_X1 U6737 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5602) );
  INV_X1 U6738 ( .A(n5750), .ZN(n5645) );
  OAI222_X1 U6739 ( .A1(n5602), .A2(n5628), .B1(n7065), .B2(n5987), .C1(n5645), 
        .C2(n7064), .ZN(U2836) );
  OAI222_X1 U6740 ( .A1(n6938), .A2(n5628), .B1(n7065), .B2(n5999), .C1(n5760), 
        .C2(n7064), .ZN(U2837) );
  INV_X1 U6741 ( .A(n5603), .ZN(n5769) );
  OAI222_X1 U6742 ( .A1(n6008), .A2(n7065), .B1(n5604), .B2(n5628), .C1(n5769), 
        .C2(n7064), .ZN(U2838) );
  OAI222_X1 U6743 ( .A1(n5652), .A2(n7064), .B1(n5628), .B2(n6908), .C1(n5605), 
        .C2(n7065), .ZN(U2839) );
  INV_X1 U6744 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5606) );
  OAI222_X1 U6745 ( .A1(n5783), .A2(n7064), .B1(n7065), .B2(n6027), .C1(n5628), 
        .C2(n5606), .ZN(U2840) );
  AOI22_X1 U6746 ( .A1(n6034), .A2(n4234), .B1(n5607), .B2(EBX_REG_18__SCAN_IN), .ZN(n5608) );
  OAI21_X1 U6747 ( .B1(n5657), .B2(n7064), .A(n5608), .ZN(U2841) );
  INV_X1 U6748 ( .A(n5797), .ZN(n5660) );
  OAI222_X1 U6749 ( .A1(n6039), .A2(n7065), .B1(n5609), .B2(n5628), .C1(n5660), 
        .C2(n7064), .ZN(U2842) );
  INV_X1 U6750 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5610) );
  OAI222_X1 U6751 ( .A1(n5611), .A2(n7065), .B1(n5610), .B2(n5628), .C1(n5665), 
        .C2(n7064), .ZN(U2843) );
  OAI222_X1 U6752 ( .A1(n5612), .A2(n7065), .B1(n6839), .B2(n5628), .C1(n5667), 
        .C2(n7064), .ZN(U2844) );
  OAI222_X1 U6753 ( .A1(n6067), .A2(n7065), .B1(n6825), .B2(n5628), .C1(n5669), 
        .C2(n7064), .ZN(U2845) );
  OAI21_X1 U6754 ( .B1(n3118), .B2(n5614), .A(n5613), .ZN(n6243) );
  OR2_X1 U6755 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  NAND2_X1 U6756 ( .A1(n5511), .A2(n5617), .ZN(n6245) );
  OAI22_X1 U6757 ( .A1(n6245), .A2(n7065), .B1(n6246), .B2(n5628), .ZN(n5618)
         );
  INV_X1 U6758 ( .A(n5618), .ZN(n5619) );
  OAI21_X1 U6759 ( .B1(n6243), .B2(n7064), .A(n5619), .ZN(U2846) );
  OAI222_X1 U6760 ( .A1(n6088), .A2(n7065), .B1(n5628), .B2(n5620), .C1(n7064), 
        .C2(n5672), .ZN(U2847) );
  INV_X1 U6761 ( .A(n5862), .ZN(n5679) );
  OAI222_X1 U6762 ( .A1(n6423), .A2(n7065), .B1(n5628), .B2(n4170), .C1(n7064), 
        .C2(n5679), .ZN(U2849) );
  OR2_X1 U6763 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  NAND2_X1 U6764 ( .A1(n5624), .A2(n5623), .ZN(n6270) );
  INV_X1 U6765 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5627) );
  OAI21_X1 U6766 ( .B1(n4422), .B2(n5626), .A(n5625), .ZN(n6266) );
  OAI222_X1 U6767 ( .A1(n6270), .A2(n7064), .B1(n5628), .B2(n5627), .C1(n7065), 
        .C2(n6266), .ZN(U2850) );
  AOI22_X1 U6768 ( .A1(n5680), .A2(EAX_REG_30__SCAN_IN), .B1(n5661), .B2(
        DATAI_30_), .ZN(n5630) );
  NAND2_X1 U6769 ( .A1(n5662), .A2(DATAI_14_), .ZN(n5629) );
  OAI211_X1 U6770 ( .C1(n5631), .C2(n5683), .A(n5630), .B(n5629), .ZN(U2861)
         );
  AOI22_X1 U6771 ( .A1(n5680), .A2(EAX_REG_28__SCAN_IN), .B1(n5661), .B2(
        DATAI_28_), .ZN(n5633) );
  NAND2_X1 U6772 ( .A1(n5662), .A2(DATAI_12_), .ZN(n5632) );
  OAI211_X1 U6773 ( .C1(n5634), .C2(n5683), .A(n5633), .B(n5632), .ZN(U2863)
         );
  AOI22_X1 U6774 ( .A1(n5680), .A2(EAX_REG_27__SCAN_IN), .B1(n5661), .B2(
        DATAI_27_), .ZN(n5636) );
  NAND2_X1 U6775 ( .A1(n5662), .A2(DATAI_11_), .ZN(n5635) );
  OAI211_X1 U6776 ( .C1(n5715), .C2(n5683), .A(n5636), .B(n5635), .ZN(U2864)
         );
  AOI22_X1 U6777 ( .A1(n5680), .A2(EAX_REG_26__SCAN_IN), .B1(n5661), .B2(
        DATAI_26_), .ZN(n5638) );
  NAND2_X1 U6778 ( .A1(n5662), .A2(DATAI_10_), .ZN(n5637) );
  OAI211_X1 U6779 ( .C1(n5722), .C2(n5683), .A(n5638), .B(n5637), .ZN(U2865)
         );
  AOI22_X1 U6780 ( .A1(n5680), .A2(EAX_REG_25__SCAN_IN), .B1(n5661), .B2(
        DATAI_25_), .ZN(n5640) );
  NAND2_X1 U6781 ( .A1(n5662), .A2(DATAI_9_), .ZN(n5639) );
  OAI211_X1 U6782 ( .C1(n5731), .C2(n5683), .A(n5640), .B(n5639), .ZN(U2866)
         );
  AOI22_X1 U6783 ( .A1(n5680), .A2(EAX_REG_24__SCAN_IN), .B1(n5661), .B2(
        DATAI_24_), .ZN(n5642) );
  NAND2_X1 U6784 ( .A1(n5662), .A2(DATAI_8_), .ZN(n5641) );
  OAI211_X1 U6785 ( .C1(n5738), .C2(n5683), .A(n5642), .B(n5641), .ZN(U2867)
         );
  AOI22_X1 U6786 ( .A1(n5680), .A2(EAX_REG_23__SCAN_IN), .B1(n5661), .B2(
        DATAI_23_), .ZN(n5644) );
  NAND2_X1 U6787 ( .A1(n5662), .A2(DATAI_7_), .ZN(n5643) );
  OAI211_X1 U6788 ( .C1(n5645), .C2(n5683), .A(n5644), .B(n5643), .ZN(U2868)
         );
  AOI22_X1 U6789 ( .A1(n5680), .A2(EAX_REG_22__SCAN_IN), .B1(n5661), .B2(
        DATAI_22_), .ZN(n5647) );
  NAND2_X1 U6790 ( .A1(n5662), .A2(DATAI_6_), .ZN(n5646) );
  OAI211_X1 U6791 ( .C1(n5760), .C2(n5683), .A(n5647), .B(n5646), .ZN(U2869)
         );
  AOI22_X1 U6792 ( .A1(n5680), .A2(EAX_REG_21__SCAN_IN), .B1(n5661), .B2(
        DATAI_21_), .ZN(n5649) );
  NAND2_X1 U6793 ( .A1(n5662), .A2(DATAI_5_), .ZN(n5648) );
  OAI211_X1 U6794 ( .C1(n5769), .C2(n5683), .A(n5649), .B(n5648), .ZN(U2870)
         );
  AOI22_X1 U6795 ( .A1(n5680), .A2(EAX_REG_20__SCAN_IN), .B1(n5661), .B2(
        DATAI_20_), .ZN(n5651) );
  NAND2_X1 U6796 ( .A1(n5662), .A2(DATAI_4_), .ZN(n5650) );
  OAI211_X1 U6797 ( .C1(n5652), .C2(n5683), .A(n5651), .B(n5650), .ZN(U2871)
         );
  AOI22_X1 U6798 ( .A1(n5680), .A2(EAX_REG_19__SCAN_IN), .B1(n5661), .B2(
        DATAI_19_), .ZN(n5654) );
  NAND2_X1 U6799 ( .A1(n5662), .A2(DATAI_3_), .ZN(n5653) );
  OAI211_X1 U6800 ( .C1(n5783), .C2(n5683), .A(n5654), .B(n5653), .ZN(U2872)
         );
  AOI22_X1 U6801 ( .A1(n5680), .A2(EAX_REG_18__SCAN_IN), .B1(n5661), .B2(
        DATAI_18_), .ZN(n5656) );
  NAND2_X1 U6802 ( .A1(n5662), .A2(DATAI_2_), .ZN(n5655) );
  OAI211_X1 U6803 ( .C1(n5657), .C2(n5683), .A(n5656), .B(n5655), .ZN(U2873)
         );
  AOI22_X1 U6804 ( .A1(n5680), .A2(EAX_REG_17__SCAN_IN), .B1(n5661), .B2(
        DATAI_17_), .ZN(n5659) );
  NAND2_X1 U6805 ( .A1(n5662), .A2(DATAI_1_), .ZN(n5658) );
  OAI211_X1 U6806 ( .C1(n5660), .C2(n5683), .A(n5659), .B(n5658), .ZN(U2874)
         );
  AOI22_X1 U6807 ( .A1(n5680), .A2(EAX_REG_16__SCAN_IN), .B1(n5661), .B2(
        DATAI_16_), .ZN(n5664) );
  NAND2_X1 U6808 ( .A1(n5662), .A2(DATAI_0_), .ZN(n5663) );
  OAI211_X1 U6809 ( .C1(n5665), .C2(n5683), .A(n5664), .B(n5663), .ZN(U2875)
         );
  AOI22_X1 U6810 ( .A1(n5681), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5680), .ZN(n5666) );
  OAI21_X1 U6811 ( .B1(n5667), .B2(n5683), .A(n5666), .ZN(U2876) );
  AOI22_X1 U6812 ( .A1(n5681), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5680), .ZN(n5668) );
  OAI21_X1 U6813 ( .B1(n5669), .B2(n5683), .A(n5668), .ZN(U2877) );
  AOI22_X1 U6814 ( .A1(n5681), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5680), .ZN(n5670) );
  OAI21_X1 U6815 ( .B1(n6243), .B2(n5683), .A(n5670), .ZN(U2878) );
  AOI22_X1 U6816 ( .A1(n5681), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5680), .ZN(n5671) );
  OAI21_X1 U6817 ( .B1(n5672), .B2(n5683), .A(n5671), .ZN(U2879) );
  INV_X1 U6818 ( .A(n5673), .ZN(n5674) );
  AOI21_X1 U6819 ( .B1(n5675), .B2(n5674), .A(n5526), .ZN(n6337) );
  INV_X1 U6820 ( .A(n6337), .ZN(n5677) );
  AOI22_X1 U6821 ( .A1(n5681), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5680), .ZN(n5676) );
  OAI21_X1 U6822 ( .B1(n5677), .B2(n5683), .A(n5676), .ZN(U2880) );
  AOI22_X1 U6823 ( .A1(n5681), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5680), .ZN(n5678) );
  OAI21_X1 U6824 ( .B1(n5679), .B2(n5683), .A(n5678), .ZN(U2881) );
  AOI22_X1 U6825 ( .A1(n5681), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5680), .ZN(n5682) );
  OAI21_X1 U6826 ( .B1(n6270), .B2(n5683), .A(n5682), .ZN(U2882) );
  NAND3_X1 U6827 ( .A1(n5689), .A2(n5688), .A3(n5687), .ZN(n5933) );
  INV_X1 U6828 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6829 ( .A1(n5870), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U6830 ( .A1(n6399), .A2(REIP_REG_30__SCAN_IN), .ZN(n5928) );
  OAI211_X1 U6831 ( .C1(n5868), .C2(n5692), .A(n5691), .B(n5928), .ZN(n5693)
         );
  AOI21_X1 U6832 ( .B1(n5694), .B2(n6404), .A(n5693), .ZN(n5695) );
  OAI21_X1 U6833 ( .B1(n6226), .B2(n5933), .A(n5695), .ZN(U2956) );
  NAND2_X1 U6834 ( .A1(n5697), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5699) );
  NAND3_X1 U6835 ( .A1(n5710), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5711), .ZN(n5698) );
  OAI211_X1 U6836 ( .C1(n5696), .C2(n5699), .A(n3106), .B(n5698), .ZN(n5700)
         );
  NAND2_X1 U6837 ( .A1(n5870), .A2(n5701), .ZN(n5702) );
  NAND2_X1 U6838 ( .A1(n6399), .A2(REIP_REG_28__SCAN_IN), .ZN(n5943) );
  OAI211_X1 U6839 ( .C1(n5868), .C2(n5703), .A(n5702), .B(n5943), .ZN(n5704)
         );
  AOI21_X1 U6840 ( .B1(n5705), .B2(n6404), .A(n5704), .ZN(n5706) );
  OAI21_X1 U6841 ( .B1(n5949), .B2(n6226), .A(n5706), .ZN(U2958) );
  NOR2_X1 U6842 ( .A1(n6443), .A2(n5707), .ZN(n5951) );
  NOR2_X1 U6843 ( .A1(n6418), .A2(n5708), .ZN(n5709) );
  AOI211_X1 U6844 ( .C1(n6410), .C2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5951), 
        .B(n5709), .ZN(n5714) );
  NAND2_X1 U6845 ( .A1(n5696), .A2(n5710), .ZN(n5712) );
  XNOR2_X1 U6846 ( .A(n5712), .B(n5711), .ZN(n5950) );
  NAND2_X1 U6847 ( .A1(n5950), .A2(n6414), .ZN(n5713) );
  OAI211_X1 U6848 ( .C1(n5715), .C2(n5873), .A(n5714), .B(n5713), .ZN(U2959)
         );
  NOR2_X1 U6849 ( .A1(n6443), .A2(n6934), .ZN(n5963) );
  NOR2_X1 U6850 ( .A1(n6418), .A2(n5716), .ZN(n5717) );
  AOI211_X1 U6851 ( .C1(n6410), .C2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5963), 
        .B(n5717), .ZN(n5721) );
  XNOR2_X1 U6852 ( .A(n5865), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5718)
         );
  XNOR2_X1 U6853 ( .A(n5719), .B(n5718), .ZN(n5959) );
  NAND2_X1 U6854 ( .A1(n5959), .A2(n6414), .ZN(n5720) );
  OAI211_X1 U6855 ( .C1(n5722), .C2(n5873), .A(n5721), .B(n5720), .ZN(U2960)
         );
  NAND2_X1 U6856 ( .A1(n6399), .A2(REIP_REG_25__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U6857 ( .B1(n5868), .B2(n5723), .A(n5968), .ZN(n5724) );
  AOI21_X1 U6858 ( .B1(n5870), .B2(n5725), .A(n5724), .ZN(n5730) );
  OAI21_X1 U6859 ( .B1(n5728), .B2(n5727), .A(n5726), .ZN(n5967) );
  NAND2_X1 U6860 ( .A1(n5967), .A2(n6414), .ZN(n5729) );
  OAI211_X1 U6861 ( .C1(n5731), .C2(n5873), .A(n5730), .B(n5729), .ZN(U2961)
         );
  INV_X1 U6862 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U6863 ( .A(n5865), .B(n5733), .ZN(n5771) );
  NAND2_X1 U6864 ( .A1(n3099), .A2(n5733), .ZN(n5734) );
  XNOR2_X1 U6865 ( .A(n5865), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5766)
         );
  NOR2_X1 U6866 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5752)
         );
  NAND2_X1 U6867 ( .A1(n5735), .A2(n5752), .ZN(n5744) );
  OAI21_X1 U6868 ( .B1(n3224), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5764), 
        .ZN(n5753) );
  NAND3_X1 U6869 ( .A1(n3099), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5736) );
  XNOR2_X1 U6870 ( .A(n5737), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5984)
         );
  INV_X1 U6871 ( .A(n5738), .ZN(n5742) );
  NOR2_X1 U6872 ( .A1(n6443), .A2(n4466), .ZN(n5981) );
  AOI21_X1 U6873 ( .B1(n6410), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5981), 
        .ZN(n5739) );
  OAI21_X1 U6874 ( .B1(n5740), .B2(n6418), .A(n5739), .ZN(n5741) );
  AOI21_X1 U6875 ( .B1(n5742), .B2(n6404), .A(n5741), .ZN(n5743) );
  OAI21_X1 U6876 ( .B1(n5984), .B2(n6226), .A(n5743), .ZN(U2962) );
  NAND2_X1 U6877 ( .A1(n4327), .A2(n5974), .ZN(n5745) );
  OAI21_X1 U6878 ( .B1(n5778), .B2(n5745), .A(n5744), .ZN(n5746) );
  XNOR2_X1 U6879 ( .A(n5746), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5991)
         );
  NAND2_X1 U6880 ( .A1(n6399), .A2(REIP_REG_23__SCAN_IN), .ZN(n5985) );
  NAND2_X1 U6881 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5747)
         );
  OAI211_X1 U6882 ( .C1(n6418), .C2(n5748), .A(n5985), .B(n5747), .ZN(n5749)
         );
  AOI21_X1 U6883 ( .B1(n5750), .B2(n6404), .A(n5749), .ZN(n5751) );
  OAI21_X1 U6884 ( .B1(n5991), .B2(n6226), .A(n5751), .ZN(U2963) );
  AOI21_X1 U6885 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5865), .A(n5752), 
        .ZN(n5754) );
  XOR2_X1 U6886 ( .A(n5754), .B(n5753), .Z(n5992) );
  NAND2_X1 U6887 ( .A1(n5992), .A2(n6414), .ZN(n5759) );
  NOR2_X1 U6888 ( .A1(n6443), .A2(n5755), .ZN(n5995) );
  NOR2_X1 U6889 ( .A1(n6418), .A2(n5756), .ZN(n5757) );
  AOI211_X1 U6890 ( .C1(n6410), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5995), 
        .B(n5757), .ZN(n5758) );
  OAI211_X1 U6891 ( .C1(n5873), .C2(n5760), .A(n5759), .B(n5758), .ZN(U2964)
         );
  NAND2_X1 U6892 ( .A1(n6399), .A2(REIP_REG_21__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U6893 ( .B1(n5868), .B2(n5761), .A(n6001), .ZN(n5762) );
  AOI21_X1 U6894 ( .B1(n5870), .B2(n5763), .A(n5762), .ZN(n5768) );
  OAI21_X1 U6895 ( .B1(n5766), .B2(n5765), .A(n5764), .ZN(n6000) );
  NAND2_X1 U6896 ( .A1(n6000), .A2(n6414), .ZN(n5767) );
  OAI211_X1 U6897 ( .C1(n5769), .C2(n5873), .A(n5768), .B(n5767), .ZN(U2965)
         );
  XOR2_X1 U6898 ( .A(n5771), .B(n5770), .Z(n6019) );
  NOR2_X1 U6899 ( .A1(n6418), .A2(n5772), .ZN(n5774) );
  NAND2_X1 U6900 ( .A1(n6399), .A2(REIP_REG_20__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U6901 ( .B1(n5868), .B2(n6962), .A(n6011), .ZN(n5773) );
  AOI211_X1 U6902 ( .C1(n5775), .C2(n6404), .A(n5774), .B(n5773), .ZN(n5776)
         );
  OAI21_X1 U6903 ( .B1(n6019), .B2(n6226), .A(n5776), .ZN(U2966) );
  XNOR2_X1 U6904 ( .A(n5865), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5777)
         );
  XNOR2_X1 U6905 ( .A(n5778), .B(n5777), .ZN(n6020) );
  NAND2_X1 U6906 ( .A1(n6020), .A2(n6414), .ZN(n5782) );
  NOR2_X1 U6907 ( .A1(n6443), .A2(n6811), .ZN(n6023) );
  NOR2_X1 U6908 ( .A1(n6418), .A2(n5779), .ZN(n5780) );
  AOI211_X1 U6909 ( .C1(n6410), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6023), 
        .B(n5780), .ZN(n5781) );
  OAI211_X1 U6910 ( .C1(n5783), .C2(n5873), .A(n5782), .B(n5781), .ZN(U2967)
         );
  NOR2_X1 U6911 ( .A1(n3224), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5813)
         );
  NOR3_X1 U6912 ( .A1(n5802), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5865), 
        .ZN(n5791) );
  NAND2_X1 U6913 ( .A1(n4327), .A2(n6048), .ZN(n5800) );
  NAND2_X1 U6914 ( .A1(n5802), .A2(n5800), .ZN(n5805) );
  NOR3_X1 U6915 ( .A1(n5805), .A2(n3224), .A3(n6037), .ZN(n5784) );
  AOI21_X1 U6916 ( .B1(n5791), .B2(n6037), .A(n5784), .ZN(n5785) );
  XNOR2_X1 U6917 ( .A(n5785), .B(n6028), .ZN(n6036) );
  NAND2_X1 U6918 ( .A1(n6399), .A2(REIP_REG_18__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U6919 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5786)
         );
  OAI211_X1 U6920 ( .C1(n6418), .C2(n5787), .A(n6030), .B(n5786), .ZN(n5788)
         );
  AOI21_X1 U6921 ( .B1(n5789), .B2(n6404), .A(n5788), .ZN(n5790) );
  OAI21_X1 U6922 ( .B1(n6036), .B2(n6226), .A(n5790), .ZN(U2968) );
  NOR2_X1 U6923 ( .A1(n3224), .A2(n6048), .ZN(n5792) );
  AOI21_X1 U6924 ( .B1(n5792), .B2(n5802), .A(n5791), .ZN(n5793) );
  XNOR2_X1 U6925 ( .A(n5793), .B(n6037), .ZN(n6045) );
  NOR2_X1 U6926 ( .A1(n6443), .A2(n5476), .ZN(n6041) );
  NOR2_X1 U6927 ( .A1(n5868), .A2(n5794), .ZN(n5795) );
  AOI211_X1 U6928 ( .C1(n5870), .C2(n5796), .A(n6041), .B(n5795), .ZN(n5799)
         );
  NAND2_X1 U6929 ( .A1(n5797), .A2(n6404), .ZN(n5798) );
  OAI211_X1 U6930 ( .C1(n6045), .C2(n6226), .A(n5799), .B(n5798), .ZN(U2969)
         );
  NOR2_X1 U6931 ( .A1(n5865), .A2(n6048), .ZN(n5804) );
  INV_X1 U6932 ( .A(n5800), .ZN(n5801) );
  NOR2_X1 U6933 ( .A1(n5804), .A2(n5801), .ZN(n5803) );
  OAI22_X1 U6934 ( .A1(n5805), .A2(n5804), .B1(n5803), .B2(n5802), .ZN(n6056)
         );
  NAND2_X1 U6935 ( .A1(n6399), .A2(REIP_REG_16__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U6936 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5806)
         );
  OAI211_X1 U6937 ( .C1(n6418), .C2(n5807), .A(n6050), .B(n5806), .ZN(n5808)
         );
  AOI21_X1 U6938 ( .B1(n5809), .B2(n6404), .A(n5808), .ZN(n5810) );
  OAI21_X1 U6939 ( .B1(n6056), .B2(n6226), .A(n5810), .ZN(U2970) );
  INV_X1 U6940 ( .A(n5811), .ZN(n5812) );
  NOR2_X1 U6941 ( .A1(n5813), .A2(n5812), .ZN(n5815) );
  XOR2_X1 U6942 ( .A(n5815), .B(n5814), .Z(n6064) );
  NAND2_X1 U6943 ( .A1(n6399), .A2(REIP_REG_15__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U6944 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5816)
         );
  OAI211_X1 U6945 ( .C1(n6418), .C2(n5817), .A(n6057), .B(n5816), .ZN(n5818)
         );
  AOI21_X1 U6946 ( .B1(n5819), .B2(n6404), .A(n5818), .ZN(n5820) );
  OAI21_X1 U6947 ( .B1(n6064), .B2(n6226), .A(n5820), .ZN(U2971) );
  XNOR2_X1 U6948 ( .A(n5865), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5830)
         );
  NAND2_X1 U6949 ( .A1(n3116), .A2(n5830), .ZN(n5829) );
  NAND2_X1 U6950 ( .A1(n5829), .A2(n5821), .ZN(n5823) );
  XNOR2_X1 U6951 ( .A(n3224), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5822)
         );
  XNOR2_X1 U6952 ( .A(n5823), .B(n5822), .ZN(n6077) );
  NAND2_X1 U6953 ( .A1(n6399), .A2(REIP_REG_14__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U6954 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5824)
         );
  OAI211_X1 U6955 ( .C1(n6418), .C2(n5825), .A(n6066), .B(n5824), .ZN(n5826)
         );
  AOI21_X1 U6956 ( .B1(n5827), .B2(n6404), .A(n5826), .ZN(n5828) );
  OAI21_X1 U6957 ( .B1(n6077), .B2(n6226), .A(n5828), .ZN(U2972) );
  OAI21_X1 U6958 ( .B1(n3116), .B2(n5830), .A(n5829), .ZN(n6079) );
  NAND2_X1 U6959 ( .A1(n6079), .A2(n6414), .ZN(n5833) );
  AND2_X1 U6960 ( .A1(n6399), .A2(REIP_REG_13__SCAN_IN), .ZN(n6082) );
  NOR2_X1 U6961 ( .A1(n6418), .A2(n6255), .ZN(n5831) );
  AOI211_X1 U6962 ( .C1(n6410), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6082), 
        .B(n5831), .ZN(n5832) );
  OAI211_X1 U6963 ( .C1(n5873), .C2(n6243), .A(n5833), .B(n5832), .ZN(U2973)
         );
  NAND2_X1 U6964 ( .A1(n5834), .A2(n5854), .ZN(n5849) );
  NOR2_X1 U6965 ( .A1(n5865), .A2(n7032), .ZN(n5847) );
  AOI21_X1 U6966 ( .B1(n5849), .B2(n5845), .A(n5847), .ZN(n5837) );
  XNOR2_X1 U6967 ( .A(n5865), .B(n5835), .ZN(n5836) );
  XNOR2_X1 U6968 ( .A(n5837), .B(n5836), .ZN(n6097) );
  NOR2_X1 U6969 ( .A1(n6443), .A2(n5838), .ZN(n6091) );
  NOR2_X1 U6970 ( .A1(n5868), .A2(n5839), .ZN(n5840) );
  AOI211_X1 U6971 ( .C1(n5870), .C2(n5841), .A(n6091), .B(n5840), .ZN(n5844)
         );
  NAND2_X1 U6972 ( .A1(n5842), .A2(n6404), .ZN(n5843) );
  OAI211_X1 U6973 ( .C1(n6097), .C2(n6226), .A(n5844), .B(n5843), .ZN(U2974)
         );
  INV_X1 U6974 ( .A(n5845), .ZN(n5846) );
  NOR2_X1 U6975 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U6976 ( .A(n5849), .B(n5848), .ZN(n6107) );
  INV_X1 U6977 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U6978 ( .A1(n5870), .A2(n6261), .ZN(n5850) );
  NAND2_X1 U6979 ( .A1(n6399), .A2(REIP_REG_11__SCAN_IN), .ZN(n6102) );
  OAI211_X1 U6980 ( .C1(n5868), .C2(n5851), .A(n5850), .B(n6102), .ZN(n5852)
         );
  AOI21_X1 U6981 ( .B1(n6337), .B2(n6404), .A(n5852), .ZN(n5853) );
  OAI21_X1 U6982 ( .B1(n6107), .B2(n6226), .A(n5853), .ZN(U2975) );
  INV_X1 U6983 ( .A(n5854), .ZN(n5856) );
  NOR2_X1 U6984 ( .A1(n5856), .A2(n5855), .ZN(n5858) );
  XOR2_X1 U6985 ( .A(n5858), .B(n5857), .Z(n6421) );
  AOI22_X1 U6986 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6399), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5859) );
  OAI21_X1 U6987 ( .B1(n5860), .B2(n6418), .A(n5859), .ZN(n5861) );
  AOI21_X1 U6988 ( .B1(n5862), .B2(n6404), .A(n5861), .ZN(n5863) );
  OAI21_X1 U6989 ( .B1(n6421), .B2(n6226), .A(n5863), .ZN(U2976) );
  XNOR2_X1 U6990 ( .A(n5865), .B(n6438), .ZN(n5866) );
  XNOR2_X1 U6991 ( .A(n5864), .B(n5866), .ZN(n6435) );
  NAND2_X1 U6992 ( .A1(n6435), .A2(n6414), .ZN(n5872) );
  INV_X1 U6993 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6994 ( .A1(n6399), .A2(REIP_REG_9__SCAN_IN), .ZN(n6430) );
  OAI21_X1 U6995 ( .B1(n5868), .B2(n5867), .A(n6430), .ZN(n5869) );
  AOI21_X1 U6996 ( .B1(n5870), .B2(n6271), .A(n5869), .ZN(n5871) );
  OAI211_X1 U6997 ( .C1(n5873), .C2(n6270), .A(n5872), .B(n5871), .ZN(U2977)
         );
  XNOR2_X1 U6998 ( .A(n5874), .B(n5875), .ZN(n6114) );
  NAND2_X1 U6999 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5876)
         );
  NAND2_X1 U7000 ( .A1(n6399), .A2(REIP_REG_8__SCAN_IN), .ZN(n6108) );
  OAI211_X1 U7001 ( .C1(n6418), .C2(n5877), .A(n5876), .B(n6108), .ZN(n5878)
         );
  AOI21_X1 U7002 ( .B1(n5879), .B2(n6404), .A(n5878), .ZN(n5880) );
  OAI21_X1 U7003 ( .B1(n6114), .B2(n6226), .A(n5880), .ZN(U2978) );
  INV_X1 U7004 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7005 ( .A1(n5882), .A2(n6404), .ZN(n5887) );
  OR2_X1 U7006 ( .A1(n5883), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6458)
         );
  NAND3_X1 U7007 ( .A1(n6458), .A2(n6414), .A3(n6457), .ZN(n5886) );
  NAND2_X1 U7008 ( .A1(n6399), .A2(REIP_REG_0__SCAN_IN), .ZN(n6452) );
  OAI21_X1 U7009 ( .B1(n6410), .B2(n5884), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5885) );
  NAND4_X1 U7010 ( .A1(n5887), .A2(n5886), .A3(n6452), .A4(n5885), .ZN(U2986)
         );
  NAND2_X1 U7011 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7012 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6427) );
  NOR3_X1 U7013 ( .A1(n5888), .A2(n6426), .A3(n6427), .ZN(n5890) );
  AND2_X1 U7014 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5889) );
  AND2_X1 U7015 ( .A1(n5890), .A2(n5889), .ZN(n5901) );
  NAND2_X1 U7016 ( .A1(n5910), .A2(n5901), .ZN(n5892) );
  AND2_X1 U7017 ( .A1(n6442), .A2(n5890), .ZN(n5899) );
  INV_X1 U7018 ( .A(n5899), .ZN(n5891) );
  NAND2_X1 U7019 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7020 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5893) );
  NOR2_X1 U7021 ( .A1(n6080), .A2(n5893), .ZN(n6049) );
  AND2_X1 U7022 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7023 ( .A1(n6049), .A2(n5894), .ZN(n6038) );
  NOR2_X1 U7024 ( .A1(n6038), .A2(n6037), .ZN(n5895) );
  NAND2_X1 U7025 ( .A1(n6105), .A2(n5895), .ZN(n6031) );
  INV_X1 U7026 ( .A(n6012), .ZN(n5896) );
  NOR2_X1 U7027 ( .A1(n6021), .A2(n5896), .ZN(n6005) );
  INV_X1 U7028 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U7029 ( .A1(n6005), .A2(n5898), .ZN(n5993) );
  NOR2_X1 U7030 ( .A1(n6440), .A2(n5899), .ZN(n5900) );
  NOR2_X1 U7031 ( .A1(n5908), .A2(n5900), .ZN(n5905) );
  INV_X1 U7032 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7033 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  NAND3_X1 U7034 ( .A1(n6012), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U7035 ( .A1(n6038), .A2(n5906), .ZN(n5907) );
  NAND2_X1 U7036 ( .A1(n6098), .A2(n5907), .ZN(n5909) );
  OR2_X1 U7037 ( .A1(n6420), .A2(n5908), .ZN(n6093) );
  NAND2_X1 U7038 ( .A1(n5909), .A2(n6093), .ZN(n6002) );
  NAND2_X1 U7039 ( .A1(n5993), .A2(n6002), .ZN(n5996) );
  INV_X1 U7040 ( .A(n5910), .ZN(n5912) );
  AOI21_X1 U7041 ( .B1(n5912), .B2(n6440), .A(n5911), .ZN(n5913) );
  NAND2_X1 U7042 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5917) );
  AND2_X1 U7043 ( .A1(n6420), .A2(n5917), .ZN(n5914) );
  AND2_X1 U7044 ( .A1(n6420), .A2(n5918), .ZN(n5915) );
  AOI21_X1 U7045 ( .B1(n3175), .B2(n6420), .A(n5940), .ZN(n5930) );
  NOR2_X1 U7046 ( .A1(n6021), .A2(n5916), .ZN(n5960) );
  INV_X1 U7047 ( .A(n5917), .ZN(n5961) );
  NAND2_X1 U7048 ( .A1(n5960), .A2(n5961), .ZN(n5953) );
  NOR2_X1 U7049 ( .A1(n5953), .A2(n5918), .ZN(n5934) );
  NAND3_X1 U7050 ( .A1(n5934), .A2(n5919), .A3(n5922), .ZN(n5920) );
  OAI211_X1 U7051 ( .C1(n5930), .C2(n5922), .A(n5921), .B(n5920), .ZN(n5923)
         );
  AOI21_X1 U7052 ( .B1(n5924), .B2(n6432), .A(n5923), .ZN(n5925) );
  OAI21_X1 U7053 ( .B1(n5926), .B2(n6422), .A(n5925), .ZN(U2987) );
  AOI21_X1 U7054 ( .B1(n5934), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5929) );
  OAI21_X1 U7055 ( .B1(n5930), .B2(n5929), .A(n5928), .ZN(n5931) );
  AOI21_X1 U7056 ( .B1(n4235), .B2(n6432), .A(n5931), .ZN(n5932) );
  OAI21_X1 U7057 ( .B1(n5933), .B2(n6422), .A(n5932), .ZN(U2988) );
  INV_X1 U7058 ( .A(n5934), .ZN(n5936) );
  OAI21_X1 U7059 ( .B1(n5936), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5935), 
        .ZN(n5939) );
  NOR2_X1 U7060 ( .A1(n5937), .A2(n6455), .ZN(n5938) );
  AOI211_X1 U7061 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5940), .A(n5939), .B(n5938), .ZN(n5941) );
  OAI21_X1 U7062 ( .B1(n5942), .B2(n6422), .A(n5941), .ZN(U2989) );
  XNOR2_X1 U7063 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U7064 ( .B1(n5953), .B2(n5944), .A(n5943), .ZN(n5947) );
  NOR2_X1 U7065 ( .A1(n5945), .A2(n6455), .ZN(n5946) );
  AOI211_X1 U7066 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5955), .A(n5947), .B(n5946), .ZN(n5948) );
  OAI21_X1 U7067 ( .B1(n5949), .B2(n6422), .A(n5948), .ZN(U2990) );
  NAND2_X1 U7068 ( .A1(n5950), .A2(n6456), .ZN(n5957) );
  INV_X1 U7069 ( .A(n5951), .ZN(n5952) );
  OAI21_X1 U7070 ( .B1(n5953), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5952), 
        .ZN(n5954) );
  AOI21_X1 U7071 ( .B1(n5955), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5954), 
        .ZN(n5956) );
  OAI211_X1 U7072 ( .C1(n6455), .C2(n5958), .A(n5957), .B(n5956), .ZN(U2991)
         );
  NAND2_X1 U7073 ( .A1(n5959), .A2(n6456), .ZN(n5965) );
  INV_X1 U7074 ( .A(n5960), .ZN(n5969) );
  AOI211_X1 U7075 ( .C1(n6899), .C2(n6851), .A(n5961), .B(n5969), .ZN(n5962)
         );
  AOI211_X1 U7076 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5976), .A(n5963), .B(n5962), .ZN(n5964) );
  OAI211_X1 U7077 ( .C1(n6455), .C2(n5966), .A(n5965), .B(n5964), .ZN(U2992)
         );
  NAND2_X1 U7078 ( .A1(n5967), .A2(n6456), .ZN(n5972) );
  OAI21_X1 U7079 ( .B1(n5969), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5968), 
        .ZN(n5970) );
  AOI21_X1 U7080 ( .B1(n5976), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5970), 
        .ZN(n5971) );
  OAI211_X1 U7081 ( .C1(n6455), .C2(n5973), .A(n5972), .B(n5971), .ZN(U2993)
         );
  INV_X1 U7082 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5979) );
  INV_X1 U7083 ( .A(n6021), .ZN(n5975) );
  NAND2_X1 U7084 ( .A1(n5975), .A2(n5974), .ZN(n5986) );
  INV_X1 U7085 ( .A(n5976), .ZN(n5977) );
  AOI211_X1 U7086 ( .C1(n5979), .C2(n5986), .A(n5978), .B(n5977), .ZN(n5980)
         );
  AOI211_X1 U7087 ( .C1(n5982), .C2(n6432), .A(n5981), .B(n5980), .ZN(n5983)
         );
  OAI21_X1 U7088 ( .B1(n5984), .B2(n6422), .A(n5983), .ZN(U2994) );
  OAI21_X1 U7089 ( .B1(n5986), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5985), 
        .ZN(n5989) );
  NOR2_X1 U7090 ( .A1(n5987), .A2(n6455), .ZN(n5988) );
  AOI211_X1 U7091 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5996), .A(n5989), .B(n5988), .ZN(n5990) );
  OAI21_X1 U7092 ( .B1(n5991), .B2(n6422), .A(n5990), .ZN(U2995) );
  NAND2_X1 U7093 ( .A1(n5992), .A2(n6456), .ZN(n5998) );
  NOR2_X1 U7094 ( .A1(n5993), .A2(n6004), .ZN(n5994) );
  AOI211_X1 U7095 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5996), .A(n5995), .B(n5994), .ZN(n5997) );
  OAI211_X1 U7096 ( .C1(n6455), .C2(n5999), .A(n5998), .B(n5997), .ZN(U2996)
         );
  NAND2_X1 U7097 ( .A1(n6000), .A2(n6456), .ZN(n6007) );
  OAI21_X1 U7098 ( .B1(n6002), .B2(n6004), .A(n6001), .ZN(n6003) );
  AOI21_X1 U7099 ( .B1(n6005), .B2(n6004), .A(n6003), .ZN(n6006) );
  OAI211_X1 U7100 ( .C1(n6455), .C2(n6008), .A(n6007), .B(n6006), .ZN(U2997)
         );
  INV_X1 U7101 ( .A(n6038), .ZN(n6009) );
  OAI211_X1 U7102 ( .C1(n6010), .C2(n6009), .A(n6098), .B(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7103 ( .A1(n6043), .A2(n6093), .ZN(n6029) );
  OAI21_X1 U7104 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6010), .A(n6029), 
        .ZN(n6024) );
  INV_X1 U7105 ( .A(n6011), .ZN(n6015) );
  NOR3_X1 U7106 ( .A1(n6021), .A2(n6013), .A3(n6012), .ZN(n6014) );
  AOI211_X1 U7107 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6024), .A(n6015), .B(n6014), .ZN(n6018) );
  NAND2_X1 U7108 ( .A1(n6016), .A2(n6432), .ZN(n6017) );
  OAI211_X1 U7109 ( .C1(n6019), .C2(n6422), .A(n6018), .B(n6017), .ZN(U2998)
         );
  NAND2_X1 U7110 ( .A1(n6020), .A2(n6456), .ZN(n6026) );
  NOR2_X1 U7111 ( .A1(n6021), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6022)
         );
  AOI211_X1 U7112 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6024), .A(n6023), .B(n6022), .ZN(n6025) );
  OAI211_X1 U7113 ( .C1(n6027), .C2(n6455), .A(n6026), .B(n6025), .ZN(U2999)
         );
  NOR2_X1 U7114 ( .A1(n6029), .A2(n6028), .ZN(n6033) );
  OAI21_X1 U7115 ( .B1(n6031), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6030), 
        .ZN(n6032) );
  AOI211_X1 U7116 ( .C1(n6034), .C2(n6432), .A(n6033), .B(n6032), .ZN(n6035)
         );
  OAI21_X1 U7117 ( .B1(n6036), .B2(n6422), .A(n6035), .ZN(U3000) );
  INV_X1 U7118 ( .A(n6105), .ZN(n6089) );
  OAI21_X1 U7119 ( .B1(n6089), .B2(n6038), .A(n6037), .ZN(n6042) );
  NOR2_X1 U7120 ( .A1(n6039), .A2(n6455), .ZN(n6040) );
  AOI211_X1 U7121 ( .C1(n6043), .C2(n6042), .A(n6041), .B(n6040), .ZN(n6044)
         );
  OAI21_X1 U7122 ( .B1(n6045), .B2(n6422), .A(n6044), .ZN(U3001) );
  INV_X1 U7123 ( .A(n6049), .ZN(n6046) );
  INV_X1 U7124 ( .A(n6098), .ZN(n6094) );
  AOI21_X1 U7125 ( .B1(n6420), .B2(n6046), .A(n6094), .ZN(n6060) );
  AND2_X1 U7126 ( .A1(n6049), .A2(n6059), .ZN(n6047) );
  NAND2_X1 U7127 ( .A1(n6105), .A2(n6047), .ZN(n6058) );
  AOI21_X1 U7128 ( .B1(n6060), .B2(n6058), .A(n6048), .ZN(n6053) );
  NAND4_X1 U7129 ( .A1(n6105), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6049), .A4(n6048), .ZN(n6051) );
  NAND2_X1 U7130 ( .A1(n6051), .A2(n6050), .ZN(n6052) );
  AOI211_X1 U7131 ( .C1(n6054), .C2(n6432), .A(n6053), .B(n6052), .ZN(n6055)
         );
  OAI21_X1 U7132 ( .B1(n6056), .B2(n6422), .A(n6055), .ZN(U3002) );
  OAI211_X1 U7133 ( .C1(n6060), .C2(n6059), .A(n6058), .B(n6057), .ZN(n6061)
         );
  AOI21_X1 U7134 ( .B1(n6062), .B2(n6432), .A(n6061), .ZN(n6063) );
  OAI21_X1 U7135 ( .B1(n6064), .B2(n6422), .A(n6063), .ZN(U3003) );
  NAND2_X1 U7136 ( .A1(n6420), .A2(n6080), .ZN(n6065) );
  OAI211_X1 U7137 ( .C1(INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n6463), .A(n6098), .B(n6065), .ZN(n6078) );
  OAI21_X1 U7138 ( .B1(n6067), .B2(n6455), .A(n6066), .ZN(n6075) );
  INV_X1 U7139 ( .A(n6068), .ZN(n6071) );
  INV_X1 U7140 ( .A(n6069), .ZN(n6070) );
  OAI21_X1 U7141 ( .B1(n6071), .B2(n6070), .A(n6086), .ZN(n6073) );
  AOI21_X1 U7142 ( .B1(n6105), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6072) );
  AOI211_X1 U7143 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6073), .A(n6080), .B(n6072), .ZN(n6074) );
  AOI211_X1 U7144 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6078), .A(n6075), .B(n6074), .ZN(n6076) );
  OAI21_X1 U7145 ( .B1(n6077), .B2(n6422), .A(n6076), .ZN(U3004) );
  INV_X1 U7146 ( .A(n6078), .ZN(n6087) );
  NAND2_X1 U7147 ( .A1(n6079), .A2(n6456), .ZN(n6085) );
  INV_X1 U7148 ( .A(n6245), .ZN(n6083) );
  NOR3_X1 U7149 ( .A1(n6089), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n6080), 
        .ZN(n6081) );
  AOI211_X1 U7150 ( .C1(n6432), .C2(n6083), .A(n6082), .B(n6081), .ZN(n6084)
         );
  OAI211_X1 U7151 ( .C1(n6087), .C2(n6086), .A(n6085), .B(n6084), .ZN(U3005)
         );
  INV_X1 U7152 ( .A(n6088), .ZN(n6092) );
  NOR3_X1 U7153 ( .A1(n6089), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n7032), 
        .ZN(n6090) );
  AOI211_X1 U7154 ( .C1(n6432), .C2(n6092), .A(n6091), .B(n6090), .ZN(n6096)
         );
  OAI211_X1 U7155 ( .C1(n6094), .C2(n7032), .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n6093), .ZN(n6095) );
  OAI211_X1 U7156 ( .C1(n6097), .C2(n6422), .A(n6096), .B(n6095), .ZN(U3006)
         );
  NOR2_X1 U7157 ( .A1(n6098), .A2(n7032), .ZN(n6104) );
  AND2_X1 U7158 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  OR2_X1 U7159 ( .A1(n6101), .A2(n5529), .ZN(n6335) );
  OAI21_X1 U7160 ( .B1(n6335), .B2(n6455), .A(n6102), .ZN(n6103) );
  AOI211_X1 U7161 ( .C1(n7032), .C2(n6105), .A(n6104), .B(n6103), .ZN(n6106)
         );
  OAI21_X1 U7162 ( .B1(n6107), .B2(n6422), .A(n6106), .ZN(U3007) );
  OAI21_X1 U7163 ( .B1(n6455), .B2(n6109), .A(n6108), .ZN(n6112) );
  OAI21_X1 U7164 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6426), .ZN(n6110) );
  NOR2_X1 U7165 ( .A1(n6425), .A2(n6110), .ZN(n6111) );
  AOI211_X1 U7166 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6419), .A(n6112), 
        .B(n6111), .ZN(n6113) );
  OAI21_X1 U7167 ( .B1(n6422), .B2(n6114), .A(n6113), .ZN(U3010) );
  INV_X1 U7168 ( .A(n6115), .ZN(n6120) );
  INV_X1 U7169 ( .A(n6116), .ZN(n6627) );
  NOR2_X1 U7170 ( .A1(n6627), .A2(n6117), .ZN(n6549) );
  NOR2_X1 U7171 ( .A1(n6549), .A2(n6118), .ZN(n6119) );
  OAI222_X1 U7172 ( .A1(n4893), .A2(n6121), .B1(n6587), .B2(n6120), .C1(n6636), 
        .C2(n6119), .ZN(n6122) );
  MUX2_X1 U7173 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6122), .S(n6465), 
        .Z(U3462) );
  INV_X1 U7174 ( .A(n6123), .ZN(n6126) );
  OAI22_X1 U7175 ( .A1(n6127), .A2(n6126), .B1(n6125), .B2(n6124), .ZN(n6130)
         );
  MUX2_X1 U7176 ( .A(n6130), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6129), 
        .Z(U3456) );
  NAND2_X1 U7177 ( .A1(n6131), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6136) );
  OAI22_X1 U7178 ( .A1(n6133), .A2(n6199), .B1(n6623), .B2(n6132), .ZN(n6134)
         );
  AOI21_X1 U7179 ( .B1(n6723), .B2(n6715), .A(n6134), .ZN(n6135) );
  OAI211_X1 U7180 ( .C1(n6137), .C2(n6642), .A(n6136), .B(n6135), .ZN(U3020)
         );
  INV_X1 U7181 ( .A(n6690), .ZN(n6139) );
  OAI21_X1 U7182 ( .B1(n6149), .B2(n6139), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6140) );
  NAND2_X1 U7183 ( .A1(n6140), .A2(n6626), .ZN(n6148) );
  INV_X1 U7184 ( .A(n6148), .ZN(n6146) );
  NAND2_X1 U7185 ( .A1(n6142), .A2(n6141), .ZN(n6630) );
  NAND3_X1 U7186 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6143), .ZN(n6635) );
  NOR2_X1 U7187 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6635), .ZN(n6150)
         );
  OAI211_X1 U7188 ( .C1(n4338), .C2(n6150), .A(n6144), .B(n6590), .ZN(n6145)
         );
  INV_X1 U7189 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6154) );
  NAND3_X1 U7190 ( .A1(n6492), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6197), .ZN(n6147) );
  NOR2_X1 U7191 ( .A1(n6179), .A2(n6624), .ZN(n6152) );
  INV_X1 U7192 ( .A(n6150), .ZN(n6180) );
  OAI22_X1 U7193 ( .A1(n6690), .A2(n6642), .B1(n6180), .B2(n6623), .ZN(n6151)
         );
  AOI211_X1 U7194 ( .C1(n6183), .C2(n6712), .A(n6152), .B(n6151), .ZN(n6153)
         );
  OAI21_X1 U7195 ( .B1(n6186), .B2(n6154), .A(n6153), .ZN(U3100) );
  INV_X1 U7196 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6158) );
  NOR2_X1 U7197 ( .A1(n6179), .A2(n6644), .ZN(n6156) );
  OAI22_X1 U7198 ( .A1(n6690), .A2(n6649), .B1(n6180), .B2(n6643), .ZN(n6155)
         );
  AOI211_X1 U7199 ( .C1(n6183), .C2(n6646), .A(n6156), .B(n6155), .ZN(n6157)
         );
  OAI21_X1 U7200 ( .B1(n6186), .B2(n6158), .A(n6157), .ZN(U3101) );
  INV_X1 U7201 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6162) );
  NOR2_X1 U7202 ( .A1(n6179), .A2(n6656), .ZN(n6160) );
  OAI22_X1 U7203 ( .A1(n6690), .A2(n6651), .B1(n6180), .B2(n6650), .ZN(n6159)
         );
  AOI211_X1 U7204 ( .C1(n6183), .C2(n6653), .A(n6160), .B(n6159), .ZN(n6161)
         );
  OAI21_X1 U7205 ( .B1(n6186), .B2(n6162), .A(n6161), .ZN(U3102) );
  INV_X1 U7206 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6166) );
  NOR2_X1 U7207 ( .A1(n6179), .A2(n6658), .ZN(n6164) );
  OAI22_X1 U7208 ( .A1(n6690), .A2(n6663), .B1(n6180), .B2(n6657), .ZN(n6163)
         );
  AOI211_X1 U7209 ( .C1(n6183), .C2(n6660), .A(n6164), .B(n6163), .ZN(n6165)
         );
  OAI21_X1 U7210 ( .B1(n6186), .B2(n6166), .A(n6165), .ZN(U3103) );
  INV_X1 U7211 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6170) );
  NOR2_X1 U7212 ( .A1(n6179), .A2(n6669), .ZN(n6168) );
  OAI22_X1 U7213 ( .A1(n6690), .A2(n6665), .B1(n6180), .B2(n6664), .ZN(n6167)
         );
  AOI211_X1 U7214 ( .C1(n6183), .C2(n6720), .A(n6168), .B(n6167), .ZN(n6169)
         );
  OAI21_X1 U7215 ( .B1(n6186), .B2(n6170), .A(n6169), .ZN(U3104) );
  INV_X1 U7216 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6174) );
  NOR2_X1 U7217 ( .A1(n6179), .A2(n6676), .ZN(n6172) );
  OAI22_X1 U7218 ( .A1(n6690), .A2(n6671), .B1(n6180), .B2(n6670), .ZN(n6171)
         );
  AOI211_X1 U7219 ( .C1(n6183), .C2(n6673), .A(n6172), .B(n6171), .ZN(n6173)
         );
  OAI21_X1 U7220 ( .B1(n6186), .B2(n6174), .A(n6173), .ZN(U3105) );
  INV_X1 U7221 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6178) );
  NOR2_X1 U7222 ( .A1(n6179), .A2(n6698), .ZN(n6176) );
  OAI22_X1 U7223 ( .A1(n6690), .A2(n6678), .B1(n6180), .B2(n6677), .ZN(n6175)
         );
  AOI211_X1 U7224 ( .C1(n6183), .C2(n6694), .A(n6176), .B(n6175), .ZN(n6177)
         );
  OAI21_X1 U7225 ( .B1(n6186), .B2(n6178), .A(n6177), .ZN(U3106) );
  INV_X1 U7226 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6185) );
  NOR2_X1 U7227 ( .A1(n6179), .A2(n6709), .ZN(n6182) );
  OAI22_X1 U7228 ( .A1(n6690), .A2(n6684), .B1(n6180), .B2(n6683), .ZN(n6181)
         );
  AOI211_X1 U7229 ( .C1(n6183), .C2(n6701), .A(n6182), .B(n6181), .ZN(n6184)
         );
  OAI21_X1 U7230 ( .B1(n6186), .B2(n6185), .A(n6184), .ZN(U3107) );
  INV_X1 U7231 ( .A(n6539), .ZN(n6187) );
  INV_X1 U7232 ( .A(n6708), .ZN(n6188) );
  NOR3_X1 U7233 ( .A1(n6188), .A2(n6703), .A3(n6636), .ZN(n6190) );
  OAI22_X1 U7234 ( .A1(n6190), .A2(n6489), .B1(n6189), .B2(n6486), .ZN(n6196)
         );
  AOI21_X1 U7235 ( .B1(n6578), .B2(n6191), .A(n6632), .ZN(n6193) );
  NOR2_X1 U7236 ( .A1(n6193), .A2(n6192), .ZN(n6591) );
  NAND2_X1 U7237 ( .A1(n6194), .A2(n6582), .ZN(n6692) );
  AOI21_X1 U7238 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6692), .A(n6492), .ZN(
        n6195) );
  NAND3_X1 U7239 ( .A1(n6196), .A2(n6591), .A3(n6195), .ZN(n6705) );
  NAND2_X1 U7240 ( .A1(n6705), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6202)
         );
  INV_X1 U7241 ( .A(n6486), .ZN(n6198) );
  NOR2_X1 U7242 ( .A1(n6590), .A2(n6197), .ZN(n6484) );
  AOI22_X1 U7243 ( .A1(n6577), .A2(n6198), .B1(n6578), .B2(n6484), .ZN(n6691)
         );
  OAI22_X1 U7244 ( .A1(n6691), .A2(n6199), .B1(n6623), .B2(n6692), .ZN(n6200)
         );
  AOI21_X1 U7245 ( .B1(n6703), .B2(n6714), .A(n6200), .ZN(n6201) );
  OAI211_X1 U7246 ( .C1(n6708), .C2(n6624), .A(n6202), .B(n6201), .ZN(U3116)
         );
  NAND2_X1 U7247 ( .A1(n6705), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6206)
         );
  OAI22_X1 U7248 ( .A1(n6691), .A2(n6203), .B1(n6643), .B2(n6692), .ZN(n6204)
         );
  AOI21_X1 U7249 ( .B1(n6703), .B2(n6596), .A(n6204), .ZN(n6205) );
  OAI211_X1 U7250 ( .C1(n6708), .C2(n6644), .A(n6206), .B(n6205), .ZN(U3117)
         );
  NAND2_X1 U7251 ( .A1(n6705), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6210)
         );
  OAI22_X1 U7252 ( .A1(n6691), .A2(n6207), .B1(n6650), .B2(n6692), .ZN(n6208)
         );
  AOI21_X1 U7253 ( .B1(n6703), .B2(n6600), .A(n6208), .ZN(n6209) );
  OAI211_X1 U7254 ( .C1(n6708), .C2(n6656), .A(n6210), .B(n6209), .ZN(U3118)
         );
  NAND2_X1 U7255 ( .A1(n6705), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6214)
         );
  OAI22_X1 U7256 ( .A1(n6691), .A2(n6211), .B1(n6657), .B2(n6692), .ZN(n6212)
         );
  AOI21_X1 U7257 ( .B1(n6703), .B2(n6604), .A(n6212), .ZN(n6213) );
  OAI211_X1 U7258 ( .C1(n6708), .C2(n6658), .A(n6214), .B(n6213), .ZN(U3119)
         );
  NAND2_X1 U7259 ( .A1(n6705), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6218)
         );
  OAI22_X1 U7260 ( .A1(n6691), .A2(n6215), .B1(n6664), .B2(n6692), .ZN(n6216)
         );
  AOI21_X1 U7261 ( .B1(n6703), .B2(n6722), .A(n6216), .ZN(n6217) );
  OAI211_X1 U7262 ( .C1(n6708), .C2(n6669), .A(n6218), .B(n6217), .ZN(U3120)
         );
  NAND2_X1 U7263 ( .A1(n6705), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6222)
         );
  OAI22_X1 U7264 ( .A1(n6691), .A2(n6219), .B1(n6670), .B2(n6692), .ZN(n6220)
         );
  AOI21_X1 U7265 ( .B1(n6703), .B2(n6610), .A(n6220), .ZN(n6221) );
  OAI211_X1 U7266 ( .C1(n6708), .C2(n6676), .A(n6222), .B(n6221), .ZN(U3121)
         );
  AND2_X1 U7267 ( .A1(n6380), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U7268 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6224) );
  OAI21_X1 U7269 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6224), .A(n6750), .ZN(n6223)
         );
  OAI21_X1 U7270 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6750), .A(n6223), .ZN(
        U2791) );
  OAI21_X1 U7271 ( .B1(BS16_N), .B2(n6224), .A(n6741), .ZN(n6739) );
  OAI21_X1 U7272 ( .B1(n6741), .B2(n6225), .A(n6739), .ZN(U2792) );
  OAI21_X1 U7273 ( .B1(n6228), .B2(n6227), .A(n6226), .ZN(U2793) );
  NOR4_X1 U7274 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6232) );
  NOR4_X1 U7275 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6231) );
  NOR4_X1 U7276 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6230) );
  NOR4_X1 U7277 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6229) );
  NAND4_X1 U7278 ( .A1(n6232), .A2(n6231), .A3(n6230), .A4(n6229), .ZN(n6238)
         );
  NOR4_X1 U7279 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6236) );
  AOI211_X1 U7280 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_15__SCAN_IN), .B(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6235) );
  NOR4_X1 U7281 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n6234) );
  NOR4_X1 U7282 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n6233) );
  NAND4_X1 U7283 ( .A1(n6236), .A2(n6235), .A3(n6234), .A4(n6233), .ZN(n6237)
         );
  NOR2_X1 U7284 ( .A1(n6238), .A2(n6237), .ZN(n6749) );
  INV_X1 U7285 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6240) );
  NOR3_X1 U7286 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6241) );
  OAI21_X1 U7287 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6241), .A(n6749), .ZN(n6239)
         );
  OAI21_X1 U7288 ( .B1(n6749), .B2(n6240), .A(n6239), .ZN(U2794) );
  INV_X1 U7289 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6740) );
  AOI21_X1 U7290 ( .B1(n6742), .B2(n6740), .A(n6241), .ZN(n6242) );
  INV_X1 U7291 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6858) );
  INV_X1 U7292 ( .A(n6749), .ZN(n6744) );
  AOI22_X1 U7293 ( .A1(n6749), .A2(n6242), .B1(n6858), .B2(n6744), .ZN(U2795)
         );
  INV_X1 U7294 ( .A(n6243), .ZN(n6251) );
  NOR3_X1 U7295 ( .A1(n6285), .A2(REIP_REG_13__SCAN_IN), .A3(n6244), .ZN(n6250) );
  OAI22_X1 U7296 ( .A1(n6246), .A2(n6294), .B1(n6334), .B2(n6245), .ZN(n6247)
         );
  AOI211_X1 U7297 ( .C1(n6330), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6247), 
        .B(n6283), .ZN(n6248) );
  INV_X1 U7298 ( .A(n6248), .ZN(n6249) );
  AOI211_X1 U7299 ( .C1(n6251), .C2(n6299), .A(n6250), .B(n6249), .ZN(n6254)
         );
  OAI21_X1 U7300 ( .B1(n6252), .B2(n6260), .A(REIP_REG_13__SCAN_IN), .ZN(n6253) );
  OAI211_X1 U7301 ( .C1(n3105), .C2(n6255), .A(n6254), .B(n6253), .ZN(U2814)
         );
  INV_X1 U7302 ( .A(n6335), .ZN(n6258) );
  AOI22_X1 U7303 ( .A1(n6305), .A2(n6258), .B1(n6257), .B2(n6256), .ZN(n6265)
         );
  INV_X1 U7304 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6339) );
  OAI22_X1 U7305 ( .A1(n6339), .A2(n6294), .B1(n5851), .B2(n6307), .ZN(n6259)
         );
  AOI211_X1 U7306 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6260), .A(n6283), .B(n6259), .ZN(n6264) );
  AOI22_X1 U7307 ( .A1(n6337), .A2(n6299), .B1(n6262), .B2(n6261), .ZN(n6263)
         );
  NAND3_X1 U7308 ( .A1(n6265), .A2(n6264), .A3(n6263), .ZN(U2816) );
  INV_X1 U7309 ( .A(n6266), .ZN(n6433) );
  AOI22_X1 U7310 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6330), .B1(n6305), 
        .B2(n6433), .ZN(n6275) );
  AND2_X1 U7311 ( .A1(n6267), .A2(REIP_REG_9__SCAN_IN), .ZN(n6268) );
  AOI211_X1 U7312 ( .C1(n6319), .C2(EBX_REG_9__SCAN_IN), .A(n6269), .B(n6268), 
        .ZN(n6274) );
  INV_X1 U7313 ( .A(n6270), .ZN(n6272) );
  AOI22_X1 U7314 ( .A1(n6272), .A2(n6299), .B1(n6262), .B2(n6271), .ZN(n6273)
         );
  NAND4_X1 U7315 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6321), .ZN(U2818)
         );
  AOI22_X1 U7316 ( .A1(n6277), .A2(n6299), .B1(n6305), .B2(n6276), .ZN(n6289)
         );
  INV_X1 U7317 ( .A(n6284), .ZN(n6279) );
  OAI21_X1 U7318 ( .B1(n6285), .B2(n6279), .A(n6278), .ZN(n6312) );
  OAI22_X1 U7319 ( .A1(n6281), .A2(n6294), .B1(n6280), .B2(n6307), .ZN(n6282)
         );
  AOI211_X1 U7320 ( .C1(REIP_REG_7__SCAN_IN), .C2(n6312), .A(n6283), .B(n6282), 
        .ZN(n6288) );
  NOR2_X1 U7321 ( .A1(n6285), .A2(n6284), .ZN(n6292) );
  OAI211_X1 U7322 ( .C1(REIP_REG_6__SCAN_IN), .C2(REIP_REG_7__SCAN_IN), .A(
        n6292), .B(n6286), .ZN(n6287) );
  AND3_X1 U7323 ( .A1(n6289), .A2(n6288), .A3(n6287), .ZN(n6290) );
  OAI21_X1 U7324 ( .B1(n6291), .B2(n3104), .A(n6290), .ZN(U2820) );
  AOI22_X1 U7325 ( .A1(n6305), .A2(n6293), .B1(n6292), .B2(n6902), .ZN(n6301)
         );
  OAI21_X1 U7326 ( .B1(n6294), .B2(n4155), .A(n6321), .ZN(n6297) );
  AOI22_X1 U7327 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6330), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6312), .ZN(n6295) );
  INV_X1 U7328 ( .A(n6295), .ZN(n6296) );
  AOI211_X1 U7329 ( .C1(n6299), .C2(n6298), .A(n6297), .B(n6296), .ZN(n6300)
         );
  OAI211_X1 U7330 ( .C1(n6302), .C2(n3105), .A(n6301), .B(n6300), .ZN(U2821)
         );
  INV_X1 U7331 ( .A(n6303), .ZN(n6304) );
  AOI22_X1 U7332 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6319), .B1(n6305), .B2(n6304), 
        .ZN(n6306) );
  OAI211_X1 U7333 ( .C1(n6307), .C2(n3723), .A(n6306), .B(n6321), .ZN(n6308)
         );
  AOI21_X1 U7334 ( .B1(n6310), .B2(n6309), .A(n6308), .ZN(n6315) );
  AND2_X1 U7335 ( .A1(n6320), .A2(n6311), .ZN(n6313) );
  OAI21_X1 U7336 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6313), .A(n6312), .ZN(n6314)
         );
  OAI211_X1 U7337 ( .C1(n3104), .C2(n6316), .A(n6315), .B(n6314), .ZN(U2822)
         );
  AOI22_X1 U7338 ( .A1(n6319), .A2(EBX_REG_4__SCAN_IN), .B1(n6318), .B2(n6317), 
        .ZN(n6332) );
  NAND4_X1 U7339 ( .A1(n6320), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .A4(REIP_REG_2__SCAN_IN), .ZN(n6324) );
  OAI221_X1 U7340 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6324), .C1(n6323), .C2(
        n6322), .A(n6321), .ZN(n6329) );
  OAI22_X1 U7341 ( .A1(n6327), .A2(n6326), .B1(n6325), .B2(n3105), .ZN(n6328)
         );
  OAI211_X1 U7342 ( .C1(n6334), .C2(n6333), .A(n6332), .B(n6331), .ZN(U2823)
         );
  NOR2_X1 U7343 ( .A1(n6335), .A2(n7065), .ZN(n6336) );
  AOI21_X1 U7344 ( .B1(n6337), .B2(n6341), .A(n6336), .ZN(n6338) );
  OAI21_X1 U7345 ( .B1(n6339), .B2(n5628), .A(n6338), .ZN(U2848) );
  AOI22_X1 U7346 ( .A1(n6405), .A2(n6341), .B1(n4234), .B2(n6340), .ZN(n6342)
         );
  OAI21_X1 U7347 ( .B1(n5574), .B2(n5628), .A(n6342), .ZN(U2857) );
  INV_X1 U7348 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n7047) );
  AOI22_X1 U7349 ( .A1(n6380), .A2(DATAO_REG_30__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U7350 ( .B1(n7047), .B2(n6383), .A(n6344), .ZN(U2893) );
  INV_X1 U7351 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U7352 ( .A1(n6380), .A2(DATAO_REG_29__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7353 ( .B1(n6814), .B2(n6383), .A(n6345), .ZN(U2894) );
  INV_X1 U7354 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7355 ( .A1(n6353), .A2(EAX_REG_28__SCAN_IN), .B1(n6374), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U7356 ( .B1(n7040), .B2(n6362), .A(n6346), .ZN(U2895) );
  INV_X1 U7357 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7358 ( .A1(n6380), .A2(DATAO_REG_27__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U7359 ( .B1(n6915), .B2(n6383), .A(n6347), .ZN(U2896) );
  INV_X1 U7360 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7361 ( .A1(n6353), .A2(EAX_REG_26__SCAN_IN), .B1(n6374), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7362 ( .B1(n6808), .B2(n6362), .A(n6348), .ZN(U2897) );
  INV_X1 U7363 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7364 ( .A1(n6353), .A2(EAX_REG_24__SCAN_IN), .B1(n6374), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6349) );
  OAI21_X1 U7365 ( .B1(n7026), .B2(n6362), .A(n6349), .ZN(U2899) );
  INV_X1 U7366 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7367 ( .A1(n6380), .A2(DATAO_REG_23__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U7368 ( .B1(n6950), .B2(n6383), .A(n6350), .ZN(U2900) );
  INV_X1 U7369 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6872) );
  AOI22_X1 U7370 ( .A1(n6380), .A2(DATAO_REG_22__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7371 ( .B1(n6872), .B2(n6383), .A(n6351), .ZN(U2901) );
  INV_X1 U7372 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n7000) );
  AOI22_X1 U7373 ( .A1(n6380), .A2(DATAO_REG_19__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6352) );
  OAI21_X1 U7374 ( .B1(n7000), .B2(n6383), .A(n6352), .ZN(U2904) );
  INV_X1 U7375 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U7376 ( .A1(n6380), .A2(DATAO_REG_17__SCAN_IN), .B1(n6353), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U7377 ( .B1(n6869), .B2(n6383), .A(n6354), .ZN(U2906) );
  AOI222_X1 U7378 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6376), .B1(n6381), .B2(
        EAX_REG_15__SCAN_IN), .C1(DATAO_REG_15__SCAN_IN), .C2(n6380), .ZN(
        n6355) );
  INV_X1 U7379 ( .A(n6355), .ZN(U2908) );
  INV_X1 U7380 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6357) );
  AOI22_X1 U7381 ( .A1(n6376), .A2(LWORD_REG_14__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7382 ( .B1(n6357), .B2(n6378), .A(n6356), .ZN(U2909) );
  INV_X1 U7383 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6359) );
  AOI22_X1 U7384 ( .A1(n6376), .A2(LWORD_REG_13__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7385 ( .B1(n6359), .B2(n6378), .A(n6358), .ZN(U2910) );
  AOI22_X1 U7386 ( .A1(n6374), .A2(LWORD_REG_12__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6360) );
  OAI21_X1 U7387 ( .B1(n3814), .B2(n6378), .A(n6360), .ZN(U2911) );
  INV_X1 U7388 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7389 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6381), .B1(n6376), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6361) );
  OAI21_X1 U7390 ( .B1(n7009), .B2(n6362), .A(n6361), .ZN(U2912) );
  INV_X1 U7391 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6364) );
  AOI22_X1 U7392 ( .A1(n6374), .A2(LWORD_REG_10__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U7393 ( .B1(n6364), .B2(n6378), .A(n6363), .ZN(U2913) );
  INV_X1 U7394 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6903) );
  AOI22_X1 U7395 ( .A1(n6374), .A2(LWORD_REG_9__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6365) );
  OAI21_X1 U7396 ( .B1(n6903), .B2(n6378), .A(n6365), .ZN(U2914) );
  INV_X1 U7397 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n7031) );
  AOI22_X1 U7398 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6381), .B1(n6380), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U7399 ( .B1(n7031), .B2(n6383), .A(n6366), .ZN(U2915) );
  AOI222_X1 U7400 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6374), .B1(n6381), .B2(
        EAX_REG_7__SCAN_IN), .C1(DATAO_REG_7__SCAN_IN), .C2(n6380), .ZN(n6367)
         );
  INV_X1 U7401 ( .A(n6367), .ZN(U2916) );
  AOI22_X1 U7402 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6376), .B1(n6380), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6368) );
  OAI21_X1 U7403 ( .B1(n6836), .B2(n6378), .A(n6368), .ZN(U2917) );
  AOI22_X1 U7404 ( .A1(n6374), .A2(LWORD_REG_5__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6369) );
  OAI21_X1 U7405 ( .B1(n6370), .B2(n6378), .A(n6369), .ZN(U2918) );
  AOI222_X1 U7406 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6374), .B1(n6381), .B2(
        EAX_REG_4__SCAN_IN), .C1(DATAO_REG_4__SCAN_IN), .C2(n6380), .ZN(n6371)
         );
  INV_X1 U7407 ( .A(n6371), .ZN(U2919) );
  AOI22_X1 U7408 ( .A1(n6374), .A2(LWORD_REG_3__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6372) );
  OAI21_X1 U7409 ( .B1(n6373), .B2(n6378), .A(n6372), .ZN(U2920) );
  AOI22_X1 U7410 ( .A1(n6374), .A2(LWORD_REG_2__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6375) );
  OAI21_X1 U7411 ( .B1(n6946), .B2(n6378), .A(n6375), .ZN(U2921) );
  AOI22_X1 U7412 ( .A1(n6376), .A2(LWORD_REG_1__SCAN_IN), .B1(n6380), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6377) );
  OAI21_X1 U7413 ( .B1(n6379), .B2(n6378), .A(n6377), .ZN(U2922) );
  INV_X1 U7414 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n7029) );
  AOI22_X1 U7415 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6381), .B1(n6380), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6382) );
  OAI21_X1 U7416 ( .B1(n7029), .B2(n6383), .A(n6382), .ZN(U2923) );
  AOI22_X1 U7417 ( .A1(EAX_REG_25__SCAN_IN), .A2(n4837), .B1(n6396), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U7418 ( .A1(n6395), .A2(DATAI_9_), .ZN(n6389) );
  NAND2_X1 U7419 ( .A1(n6384), .A2(n6389), .ZN(U2933) );
  NAND2_X1 U7420 ( .A1(n6395), .A2(DATAI_11_), .ZN(n6391) );
  INV_X1 U7421 ( .A(n6391), .ZN(n6385) );
  AOI21_X1 U7422 ( .B1(n4837), .B2(EAX_REG_27__SCAN_IN), .A(n6385), .ZN(n6386)
         );
  OAI21_X1 U7423 ( .B1(n6915), .B2(n4801), .A(n6386), .ZN(U2935) );
  NAND2_X1 U7424 ( .A1(n6395), .A2(DATAI_13_), .ZN(n6393) );
  INV_X1 U7425 ( .A(n6393), .ZN(n6387) );
  AOI21_X1 U7426 ( .B1(n4837), .B2(EAX_REG_29__SCAN_IN), .A(n6387), .ZN(n6388)
         );
  OAI21_X1 U7427 ( .B1(n6814), .B2(n4801), .A(n6388), .ZN(U2937) );
  AOI22_X1 U7428 ( .A1(EAX_REG_9__SCAN_IN), .A2(n4837), .B1(n6396), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7429 ( .A1(n6390), .A2(n6389), .ZN(U2948) );
  AOI22_X1 U7430 ( .A1(EAX_REG_11__SCAN_IN), .A2(n4837), .B1(n6396), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U7431 ( .A1(n6392), .A2(n6391), .ZN(U2950) );
  AOI22_X1 U7432 ( .A1(EAX_REG_13__SCAN_IN), .A2(n4837), .B1(n6396), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7433 ( .A1(n6394), .A2(n6393), .ZN(U2952) );
  INV_X1 U7434 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7435 ( .A1(n6396), .A2(LWORD_REG_15__SCAN_IN), .B1(n6395), .B2(
        DATAI_15_), .ZN(n6397) );
  OAI21_X1 U7436 ( .B1(n6936), .B2(n6398), .A(n6397), .ZN(U2954) );
  AOI22_X1 U7437 ( .A1(n6410), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6399), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U7438 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  XOR2_X1 U7439 ( .A(n6403), .B(n6402), .Z(n6448) );
  AOI22_X1 U7440 ( .A1(n6448), .A2(n6414), .B1(n6405), .B2(n6404), .ZN(n6406)
         );
  OAI211_X1 U7441 ( .C1(n6418), .C2(n6408), .A(n6407), .B(n6406), .ZN(U2984)
         );
  AOI21_X1 U7442 ( .B1(n6410), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6409), 
        .ZN(n6417) );
  INV_X1 U7443 ( .A(n6411), .ZN(n6415) );
  INV_X1 U7444 ( .A(n6412), .ZN(n6413) );
  AOI22_X1 U7445 ( .A1(n6415), .A2(n6404), .B1(n6414), .B2(n6413), .ZN(n6416)
         );
  OAI211_X1 U7446 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6418), .A(n6417), 
        .B(n6416), .ZN(U2985) );
  AOI21_X1 U7447 ( .B1(n6420), .B2(n6426), .A(n6419), .ZN(n6439) );
  OAI222_X1 U7448 ( .A1(n6423), .A2(n6455), .B1(n6443), .B2(n4474), .C1(n6422), 
        .C2(n6421), .ZN(n6424) );
  INV_X1 U7449 ( .A(n6424), .ZN(n6429) );
  NOR2_X1 U7450 ( .A1(n6426), .A2(n6425), .ZN(n6434) );
  OAI211_X1 U7451 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6434), .B(n6427), .ZN(n6428) );
  OAI211_X1 U7452 ( .C1(n6439), .C2(n6963), .A(n6429), .B(n6428), .ZN(U3008)
         );
  INV_X1 U7453 ( .A(n6430), .ZN(n6431) );
  AOI21_X1 U7454 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(n6437) );
  AOI22_X1 U7455 ( .A1(n6435), .A2(n6456), .B1(n6434), .B2(n6438), .ZN(n6436)
         );
  OAI211_X1 U7456 ( .C1(n6439), .C2(n6438), .A(n6437), .B(n6436), .ZN(U3009)
         );
  NAND3_X1 U7457 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6441) );
  AOI21_X1 U7458 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(n6447) );
  OAI22_X1 U7459 ( .A1(n6455), .A2(n6445), .B1(n6444), .B2(n6443), .ZN(n6446)
         );
  AOI211_X1 U7460 ( .C1(n6448), .C2(n6456), .A(n6447), .B(n6446), .ZN(n6449)
         );
  OAI221_X1 U7461 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6451), .C1(n4143), .C2(n6450), .A(n6449), .ZN(U3016) );
  OAI211_X1 U7462 ( .C1(n6455), .C2(n6454), .A(n6453), .B(n6452), .ZN(n6460)
         );
  AND3_X1 U7463 ( .A1(n6458), .A2(n6457), .A3(n6456), .ZN(n6459) );
  NOR2_X1 U7464 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  OAI221_X1 U7465 ( .B1(n6464), .B2(n6463), .C1(n6464), .C2(n6462), .A(n6461), 
        .ZN(U3018) );
  NOR2_X1 U7466 ( .A1(n6466), .A2(n6465), .ZN(U3019) );
  INV_X1 U7467 ( .A(n6467), .ZN(n6476) );
  AOI22_X1 U7468 ( .A1(n6478), .A2(n6521), .B1(n6595), .B2(n6476), .ZN(n6469)
         );
  AOI22_X1 U7469 ( .A1(n6646), .A2(n6480), .B1(n6479), .B2(
        INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6468) );
  OAI211_X1 U7470 ( .C1(n6649), .C2(n6517), .A(n6469), .B(n6468), .ZN(U3045)
         );
  AOI22_X1 U7471 ( .A1(n6478), .A2(n6524), .B1(n6599), .B2(n6476), .ZN(n6471)
         );
  AOI22_X1 U7472 ( .A1(n6653), .A2(n6480), .B1(n6479), .B2(
        INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6470) );
  OAI211_X1 U7473 ( .C1(n6651), .C2(n6517), .A(n6471), .B(n6470), .ZN(U3046)
         );
  AOI22_X1 U7474 ( .A1(n6478), .A2(n6527), .B1(n6603), .B2(n6476), .ZN(n6473)
         );
  AOI22_X1 U7475 ( .A1(n6660), .A2(n6480), .B1(n6479), .B2(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6472) );
  OAI211_X1 U7476 ( .C1(n6663), .C2(n6517), .A(n6473), .B(n6472), .ZN(U3047)
         );
  AOI22_X1 U7477 ( .A1(n6478), .A2(n6724), .B1(n6718), .B2(n6476), .ZN(n6475)
         );
  AOI22_X1 U7478 ( .A1(n6720), .A2(n6480), .B1(n6479), .B2(
        INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6474) );
  OAI211_X1 U7479 ( .C1(n6665), .C2(n6517), .A(n6475), .B(n6474), .ZN(U3048)
         );
  AOI22_X1 U7480 ( .A1(n6478), .A2(n6477), .B1(n6700), .B2(n6476), .ZN(n6482)
         );
  AOI22_X1 U7481 ( .A1(n6701), .A2(n6480), .B1(n6479), .B2(
        INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6481) );
  OAI211_X1 U7482 ( .C1(n6684), .C2(n6517), .A(n6482), .B(n6481), .ZN(U3051)
         );
  INV_X1 U7483 ( .A(n6483), .ZN(n6487) );
  INV_X1 U7484 ( .A(n6484), .ZN(n6485) );
  OAI22_X1 U7485 ( .A1(n6487), .A2(n6486), .B1(n6578), .B2(n6485), .ZN(n6512)
         );
  NAND2_X1 U7486 ( .A1(n6488), .A2(n6582), .ZN(n6493) );
  INV_X1 U7487 ( .A(n6493), .ZN(n6511) );
  AOI22_X1 U7488 ( .A1(n6512), .A2(n6712), .B1(n6711), .B2(n6511), .ZN(n6498)
         );
  NOR2_X1 U7489 ( .A1(n6513), .A2(n6636), .ZN(n6490) );
  AOI21_X1 U7490 ( .B1(n6490), .B2(n6517), .A(n6489), .ZN(n6496) );
  AOI211_X1 U7491 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6493), .A(n6492), .B(
        n6491), .ZN(n6494) );
  AOI22_X1 U7492 ( .A1(n6514), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6714), 
        .B2(n6513), .ZN(n6497) );
  OAI211_X1 U7493 ( .C1(n6624), .C2(n6517), .A(n6498), .B(n6497), .ZN(U3052)
         );
  AOI22_X1 U7494 ( .A1(n6512), .A2(n6646), .B1(n6595), .B2(n6511), .ZN(n6500)
         );
  AOI22_X1 U7495 ( .A1(n6514), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6596), 
        .B2(n6513), .ZN(n6499) );
  OAI211_X1 U7496 ( .C1(n6644), .C2(n6517), .A(n6500), .B(n6499), .ZN(U3053)
         );
  AOI22_X1 U7497 ( .A1(n6512), .A2(n6653), .B1(n6599), .B2(n6511), .ZN(n6502)
         );
  AOI22_X1 U7498 ( .A1(n6514), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6600), 
        .B2(n6513), .ZN(n6501) );
  OAI211_X1 U7499 ( .C1(n6656), .C2(n6517), .A(n6502), .B(n6501), .ZN(U3054)
         );
  AOI22_X1 U7500 ( .A1(n6512), .A2(n6660), .B1(n6603), .B2(n6511), .ZN(n6504)
         );
  AOI22_X1 U7501 ( .A1(n6514), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6604), 
        .B2(n6513), .ZN(n6503) );
  OAI211_X1 U7502 ( .C1(n6658), .C2(n6517), .A(n6504), .B(n6503), .ZN(U3055)
         );
  AOI22_X1 U7503 ( .A1(n6512), .A2(n6720), .B1(n6718), .B2(n6511), .ZN(n6506)
         );
  AOI22_X1 U7504 ( .A1(n6514), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6722), 
        .B2(n6513), .ZN(n6505) );
  OAI211_X1 U7505 ( .C1(n6669), .C2(n6517), .A(n6506), .B(n6505), .ZN(U3056)
         );
  AOI22_X1 U7506 ( .A1(n6512), .A2(n6673), .B1(n6609), .B2(n6511), .ZN(n6508)
         );
  AOI22_X1 U7507 ( .A1(n6514), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6610), 
        .B2(n6513), .ZN(n6507) );
  OAI211_X1 U7508 ( .C1(n6676), .C2(n6517), .A(n6508), .B(n6507), .ZN(U3057)
         );
  AOI22_X1 U7509 ( .A1(n6512), .A2(n6694), .B1(n6693), .B2(n6511), .ZN(n6510)
         );
  AOI22_X1 U7510 ( .A1(n6514), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6695), 
        .B2(n6513), .ZN(n6509) );
  OAI211_X1 U7511 ( .C1(n6698), .C2(n6517), .A(n6510), .B(n6509), .ZN(U3058)
         );
  AOI22_X1 U7512 ( .A1(n6512), .A2(n6701), .B1(n6700), .B2(n6511), .ZN(n6516)
         );
  AOI22_X1 U7513 ( .A1(n6514), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6704), 
        .B2(n6513), .ZN(n6515) );
  OAI211_X1 U7514 ( .C1(n6709), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3059)
         );
  INV_X1 U7515 ( .A(n6518), .ZN(n6532) );
  AOI22_X1 U7516 ( .A1(n6533), .A2(n6712), .B1(n6711), .B2(n6532), .ZN(n6520)
         );
  AOI22_X1 U7517 ( .A1(n6536), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6715), 
        .B2(n6534), .ZN(n6519) );
  OAI211_X1 U7518 ( .C1(n6642), .C2(n6576), .A(n6520), .B(n6519), .ZN(U3068)
         );
  AOI22_X1 U7519 ( .A1(n6533), .A2(n6646), .B1(n6595), .B2(n6532), .ZN(n6523)
         );
  AOI22_X1 U7520 ( .A1(n6536), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6521), 
        .B2(n6534), .ZN(n6522) );
  OAI211_X1 U7521 ( .C1(n6649), .C2(n6576), .A(n6523), .B(n6522), .ZN(U3069)
         );
  AOI22_X1 U7522 ( .A1(n6533), .A2(n6653), .B1(n6599), .B2(n6532), .ZN(n6526)
         );
  AOI22_X1 U7523 ( .A1(n6536), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6524), 
        .B2(n6534), .ZN(n6525) );
  OAI211_X1 U7524 ( .C1(n6651), .C2(n6576), .A(n6526), .B(n6525), .ZN(U3070)
         );
  AOI22_X1 U7525 ( .A1(n6533), .A2(n6660), .B1(n6603), .B2(n6532), .ZN(n6529)
         );
  AOI22_X1 U7526 ( .A1(n6536), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6527), 
        .B2(n6534), .ZN(n6528) );
  OAI211_X1 U7527 ( .C1(n6663), .C2(n6576), .A(n6529), .B(n6528), .ZN(U3071)
         );
  AOI22_X1 U7528 ( .A1(n6533), .A2(n6720), .B1(n6718), .B2(n6532), .ZN(n6531)
         );
  AOI22_X1 U7529 ( .A1(n6536), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6724), 
        .B2(n6534), .ZN(n6530) );
  OAI211_X1 U7530 ( .C1(n6665), .C2(n6576), .A(n6531), .B(n6530), .ZN(U3072)
         );
  AOI22_X1 U7531 ( .A1(n6533), .A2(n6673), .B1(n6609), .B2(n6532), .ZN(n6538)
         );
  AOI22_X1 U7532 ( .A1(n6536), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6535), 
        .B2(n6534), .ZN(n6537) );
  OAI211_X1 U7533 ( .C1(n6671), .C2(n6576), .A(n6538), .B(n6537), .ZN(U3073)
         );
  OAI22_X1 U7534 ( .A1(n6576), .A2(n6624), .B1(n6570), .B2(n6623), .ZN(n6541)
         );
  INV_X1 U7535 ( .A(n6541), .ZN(n6551) );
  OAI21_X1 U7536 ( .B1(n6542), .B2(n6629), .A(n6570), .ZN(n6545) );
  OR3_X1 U7537 ( .A1(n6549), .A2(n6636), .A3(n6545), .ZN(n6544) );
  OAI211_X1 U7538 ( .C1(n6546), .C2(n6626), .A(n6544), .B(n6543), .ZN(n6573)
         );
  NAND2_X1 U7539 ( .A1(n6545), .A2(n6626), .ZN(n6548) );
  INV_X1 U7540 ( .A(n6546), .ZN(n6547) );
  OAI22_X1 U7541 ( .A1(n6549), .A2(n6548), .B1(n6547), .B2(n6632), .ZN(n6572)
         );
  AOI22_X1 U7542 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6573), .B1(n6712), 
        .B2(n6572), .ZN(n6550) );
  OAI211_X1 U7543 ( .C1(n6642), .C2(n6621), .A(n6551), .B(n6550), .ZN(U3076)
         );
  OAI22_X1 U7544 ( .A1(n6576), .A2(n6644), .B1(n6570), .B2(n6643), .ZN(n6552)
         );
  INV_X1 U7545 ( .A(n6552), .ZN(n6554) );
  AOI22_X1 U7546 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6573), .B1(n6646), 
        .B2(n6572), .ZN(n6553) );
  OAI211_X1 U7547 ( .C1(n6649), .C2(n6621), .A(n6554), .B(n6553), .ZN(U3077)
         );
  OAI22_X1 U7548 ( .A1(n6621), .A2(n6651), .B1(n6570), .B2(n6650), .ZN(n6555)
         );
  INV_X1 U7549 ( .A(n6555), .ZN(n6557) );
  AOI22_X1 U7550 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6573), .B1(n6653), 
        .B2(n6572), .ZN(n6556) );
  OAI211_X1 U7551 ( .C1(n6656), .C2(n6576), .A(n6557), .B(n6556), .ZN(U3078)
         );
  OAI22_X1 U7552 ( .A1(n6576), .A2(n6658), .B1(n6570), .B2(n6657), .ZN(n6558)
         );
  INV_X1 U7553 ( .A(n6558), .ZN(n6560) );
  AOI22_X1 U7554 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6573), .B1(n6660), 
        .B2(n6572), .ZN(n6559) );
  OAI211_X1 U7555 ( .C1(n6663), .C2(n6621), .A(n6560), .B(n6559), .ZN(U3079)
         );
  OAI22_X1 U7556 ( .A1(n6576), .A2(n6669), .B1(n6570), .B2(n6664), .ZN(n6561)
         );
  INV_X1 U7557 ( .A(n6561), .ZN(n6563) );
  AOI22_X1 U7558 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6573), .B1(n6720), 
        .B2(n6572), .ZN(n6562) );
  OAI211_X1 U7559 ( .C1(n6665), .C2(n6621), .A(n6563), .B(n6562), .ZN(U3080)
         );
  OAI22_X1 U7560 ( .A1(n6576), .A2(n6676), .B1(n6570), .B2(n6670), .ZN(n6564)
         );
  INV_X1 U7561 ( .A(n6564), .ZN(n6566) );
  AOI22_X1 U7562 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6573), .B1(n6673), 
        .B2(n6572), .ZN(n6565) );
  OAI211_X1 U7563 ( .C1(n6671), .C2(n6621), .A(n6566), .B(n6565), .ZN(U3081)
         );
  OAI22_X1 U7564 ( .A1(n6621), .A2(n6678), .B1(n6570), .B2(n6677), .ZN(n6567)
         );
  INV_X1 U7565 ( .A(n6567), .ZN(n6569) );
  AOI22_X1 U7566 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6573), .B1(n6694), 
        .B2(n6572), .ZN(n6568) );
  OAI211_X1 U7567 ( .C1(n6698), .C2(n6576), .A(n6569), .B(n6568), .ZN(U3082)
         );
  OAI22_X1 U7568 ( .A1(n6621), .A2(n6684), .B1(n6570), .B2(n6683), .ZN(n6571)
         );
  INV_X1 U7569 ( .A(n6571), .ZN(n6575) );
  AOI22_X1 U7570 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6573), .B1(n6701), 
        .B2(n6572), .ZN(n6574) );
  OAI211_X1 U7571 ( .C1(n6709), .C2(n6576), .A(n6575), .B(n6574), .ZN(U3083)
         );
  INV_X1 U7572 ( .A(n6577), .ZN(n6581) );
  INV_X1 U7573 ( .A(n6578), .ZN(n6580) );
  OAI22_X1 U7574 ( .A1(n6581), .A2(n6586), .B1(n6580), .B2(n6579), .ZN(n6616)
         );
  NAND2_X1 U7575 ( .A1(n6583), .A2(n6582), .ZN(n6588) );
  INV_X1 U7576 ( .A(n6588), .ZN(n6615) );
  AOI22_X1 U7577 ( .A1(n6616), .A2(n6712), .B1(n6711), .B2(n6615), .ZN(n6594)
         );
  INV_X1 U7578 ( .A(n6621), .ZN(n6584) );
  OAI21_X1 U7579 ( .B1(n6617), .B2(n6584), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6585) );
  OAI211_X1 U7580 ( .C1(n6587), .C2(n6586), .A(n6585), .B(n6626), .ZN(n6592)
         );
  NAND2_X1 U7581 ( .A1(n6588), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6589) );
  NAND4_X1 U7582 ( .A1(n6592), .A2(n6591), .A3(n6590), .A4(n6589), .ZN(n6618)
         );
  AOI22_X1 U7583 ( .A1(n6618), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6714), 
        .B2(n6617), .ZN(n6593) );
  OAI211_X1 U7584 ( .C1(n6624), .C2(n6621), .A(n6594), .B(n6593), .ZN(U3084)
         );
  AOI22_X1 U7585 ( .A1(n6616), .A2(n6646), .B1(n6595), .B2(n6615), .ZN(n6598)
         );
  AOI22_X1 U7586 ( .A1(n6618), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6596), 
        .B2(n6617), .ZN(n6597) );
  OAI211_X1 U7587 ( .C1(n6644), .C2(n6621), .A(n6598), .B(n6597), .ZN(U3085)
         );
  AOI22_X1 U7588 ( .A1(n6616), .A2(n6653), .B1(n6599), .B2(n6615), .ZN(n6602)
         );
  AOI22_X1 U7589 ( .A1(n6618), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6600), 
        .B2(n6617), .ZN(n6601) );
  OAI211_X1 U7590 ( .C1(n6656), .C2(n6621), .A(n6602), .B(n6601), .ZN(U3086)
         );
  AOI22_X1 U7591 ( .A1(n6616), .A2(n6660), .B1(n6603), .B2(n6615), .ZN(n6606)
         );
  AOI22_X1 U7592 ( .A1(n6618), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6604), 
        .B2(n6617), .ZN(n6605) );
  OAI211_X1 U7593 ( .C1(n6658), .C2(n6621), .A(n6606), .B(n6605), .ZN(U3087)
         );
  AOI22_X1 U7594 ( .A1(n6616), .A2(n6720), .B1(n6718), .B2(n6615), .ZN(n6608)
         );
  AOI22_X1 U7595 ( .A1(n6618), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6722), 
        .B2(n6617), .ZN(n6607) );
  OAI211_X1 U7596 ( .C1(n6669), .C2(n6621), .A(n6608), .B(n6607), .ZN(U3088)
         );
  AOI22_X1 U7597 ( .A1(n6616), .A2(n6673), .B1(n6609), .B2(n6615), .ZN(n6612)
         );
  AOI22_X1 U7598 ( .A1(n6618), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6610), 
        .B2(n6617), .ZN(n6611) );
  OAI211_X1 U7599 ( .C1(n6676), .C2(n6621), .A(n6612), .B(n6611), .ZN(U3089)
         );
  AOI22_X1 U7600 ( .A1(n6616), .A2(n6694), .B1(n6693), .B2(n6615), .ZN(n6614)
         );
  AOI22_X1 U7601 ( .A1(n6618), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6695), 
        .B2(n6617), .ZN(n6613) );
  OAI211_X1 U7602 ( .C1(n6698), .C2(n6621), .A(n6614), .B(n6613), .ZN(U3090)
         );
  AOI22_X1 U7603 ( .A1(n6616), .A2(n6701), .B1(n6700), .B2(n6615), .ZN(n6620)
         );
  AOI22_X1 U7604 ( .A1(n6618), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6704), 
        .B2(n6617), .ZN(n6619) );
  OAI211_X1 U7605 ( .C1(n6709), .C2(n6621), .A(n6620), .B(n6619), .ZN(U3091)
         );
  NAND2_X1 U7606 ( .A1(n6622), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6682) );
  OAI22_X1 U7607 ( .A1(n6690), .A2(n6624), .B1(n6623), .B2(n6682), .ZN(n6625)
         );
  INV_X1 U7608 ( .A(n6625), .ZN(n6641) );
  OAI21_X1 U7609 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(n6639) );
  OR2_X1 U7610 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  OAI22_X1 U7611 ( .A1(n6639), .A2(n6633), .B1(n6635), .B2(n6632), .ZN(n6687)
         );
  INV_X1 U7612 ( .A(n6633), .ZN(n6638) );
  AOI21_X1 U7613 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6637) );
  AOI22_X1 U7614 ( .A1(n6712), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6640) );
  OAI211_X1 U7615 ( .C1(n6642), .C2(n6708), .A(n6641), .B(n6640), .ZN(U3108)
         );
  OAI22_X1 U7616 ( .A1(n6690), .A2(n6644), .B1(n6643), .B2(n6682), .ZN(n6645)
         );
  INV_X1 U7617 ( .A(n6645), .ZN(n6648) );
  AOI22_X1 U7618 ( .A1(n6646), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6647) );
  OAI211_X1 U7619 ( .C1(n6649), .C2(n6708), .A(n6648), .B(n6647), .ZN(U3109)
         );
  OAI22_X1 U7620 ( .A1(n6708), .A2(n6651), .B1(n6650), .B2(n6682), .ZN(n6652)
         );
  INV_X1 U7621 ( .A(n6652), .ZN(n6655) );
  AOI22_X1 U7622 ( .A1(n6653), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6654) );
  OAI211_X1 U7623 ( .C1(n6656), .C2(n6690), .A(n6655), .B(n6654), .ZN(U3110)
         );
  OAI22_X1 U7624 ( .A1(n6690), .A2(n6658), .B1(n6657), .B2(n6682), .ZN(n6659)
         );
  INV_X1 U7625 ( .A(n6659), .ZN(n6662) );
  AOI22_X1 U7626 ( .A1(n6660), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6661) );
  OAI211_X1 U7627 ( .C1(n6663), .C2(n6708), .A(n6662), .B(n6661), .ZN(U3111)
         );
  OAI22_X1 U7628 ( .A1(n6708), .A2(n6665), .B1(n6664), .B2(n6682), .ZN(n6666)
         );
  INV_X1 U7629 ( .A(n6666), .ZN(n6668) );
  AOI22_X1 U7630 ( .A1(n6720), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6667) );
  OAI211_X1 U7631 ( .C1(n6669), .C2(n6690), .A(n6668), .B(n6667), .ZN(U3112)
         );
  OAI22_X1 U7632 ( .A1(n6708), .A2(n6671), .B1(n6670), .B2(n6682), .ZN(n6672)
         );
  INV_X1 U7633 ( .A(n6672), .ZN(n6675) );
  AOI22_X1 U7634 ( .A1(n6673), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6674) );
  OAI211_X1 U7635 ( .C1(n6676), .C2(n6690), .A(n6675), .B(n6674), .ZN(U3113)
         );
  OAI22_X1 U7636 ( .A1(n6708), .A2(n6678), .B1(n6677), .B2(n6682), .ZN(n6679)
         );
  INV_X1 U7637 ( .A(n6679), .ZN(n6681) );
  AOI22_X1 U7638 ( .A1(n6694), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6680) );
  OAI211_X1 U7639 ( .C1(n6698), .C2(n6690), .A(n6681), .B(n6680), .ZN(U3114)
         );
  OAI22_X1 U7640 ( .A1(n6708), .A2(n6684), .B1(n6683), .B2(n6682), .ZN(n6685)
         );
  INV_X1 U7641 ( .A(n6685), .ZN(n6689) );
  AOI22_X1 U7642 ( .A1(n6701), .A2(n6687), .B1(n6686), .B2(
        INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6688) );
  OAI211_X1 U7643 ( .C1(n6709), .C2(n6690), .A(n6689), .B(n6688), .ZN(U3115)
         );
  INV_X1 U7644 ( .A(n6691), .ZN(n6702) );
  INV_X1 U7645 ( .A(n6692), .ZN(n6699) );
  AOI22_X1 U7646 ( .A1(n6702), .A2(n6694), .B1(n6693), .B2(n6699), .ZN(n6697)
         );
  AOI22_X1 U7647 ( .A1(n6705), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6695), 
        .B2(n6703), .ZN(n6696) );
  OAI211_X1 U7648 ( .C1(n6698), .C2(n6708), .A(n6697), .B(n6696), .ZN(U3122)
         );
  AOI22_X1 U7649 ( .A1(n6702), .A2(n6701), .B1(n6700), .B2(n6699), .ZN(n6707)
         );
  AOI22_X1 U7650 ( .A1(n6705), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6704), 
        .B2(n6703), .ZN(n6706) );
  OAI211_X1 U7651 ( .C1(n6709), .C2(n6708), .A(n6707), .B(n6706), .ZN(U3123)
         );
  INV_X1 U7652 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6871) );
  INV_X1 U7653 ( .A(n6710), .ZN(n6719) );
  AOI22_X1 U7654 ( .A1(n6721), .A2(n6712), .B1(n6719), .B2(n6711), .ZN(n6717)
         );
  INV_X1 U7655 ( .A(n6713), .ZN(n6725) );
  AOI22_X1 U7656 ( .A1(n6725), .A2(n6715), .B1(n6723), .B2(n6714), .ZN(n6716)
         );
  OAI211_X1 U7657 ( .C1(n6728), .C2(n6871), .A(n6717), .B(n6716), .ZN(U3140)
         );
  INV_X1 U7658 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U7659 ( .A1(n6721), .A2(n6720), .B1(n6719), .B2(n6718), .ZN(n6727)
         );
  AOI22_X1 U7660 ( .A1(n6725), .A2(n6724), .B1(n6723), .B2(n6722), .ZN(n6726)
         );
  OAI211_X1 U7661 ( .C1(n6728), .C2(n6965), .A(n6727), .B(n6726), .ZN(U3144)
         );
  AOI21_X1 U7662 ( .B1(n6730), .B2(n7019), .A(n6729), .ZN(n6735) );
  INV_X1 U7663 ( .A(n6731), .ZN(n6732) );
  OAI211_X1 U7664 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(n6732), .B(STATE2_REG_1__SCAN_IN), .ZN(n6733) );
  OAI211_X1 U7665 ( .C1(n6736), .C2(n6735), .A(n6734), .B(n6733), .ZN(U3149)
         );
  AND2_X1 U7666 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6737), .ZN(U3151) );
  AND2_X1 U7667 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6737), .ZN(U3152) );
  AND2_X1 U7668 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6737), .ZN(U3153) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6737), .ZN(U3154) );
  AND2_X1 U7670 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6737), .ZN(U3155) );
  AND2_X1 U7671 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6737), .ZN(U3156) );
  AND2_X1 U7672 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6737), .ZN(U3157) );
  INV_X1 U7673 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U7674 ( .A1(n6741), .A2(n6994), .ZN(U3158) );
  AND2_X1 U7675 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6737), .ZN(U3159) );
  INV_X1 U7676 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6920) );
  NOR2_X1 U7677 ( .A1(n6741), .A2(n6920), .ZN(U3160) );
  AND2_X1 U7678 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6737), .ZN(U3161) );
  AND2_X1 U7679 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6737), .ZN(U3162) );
  AND2_X1 U7680 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6737), .ZN(U3163) );
  AND2_X1 U7681 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6737), .ZN(U3164) );
  INV_X1 U7682 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6854) );
  NOR2_X1 U7683 ( .A1(n6741), .A2(n6854), .ZN(U3165) );
  INV_X1 U7684 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6885) );
  NOR2_X1 U7685 ( .A1(n6741), .A2(n6885), .ZN(U3166) );
  INV_X1 U7686 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7004) );
  NOR2_X1 U7687 ( .A1(n6741), .A2(n7004), .ZN(U3167) );
  AND2_X1 U7688 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6737), .ZN(U3168) );
  AND2_X1 U7689 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6737), .ZN(U3169) );
  INV_X1 U7690 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6868) );
  NOR2_X1 U7691 ( .A1(n6741), .A2(n6868), .ZN(U3170) );
  AND2_X1 U7692 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6737), .ZN(U3171) );
  AND2_X1 U7693 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6737), .ZN(U3172) );
  AND2_X1 U7694 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6737), .ZN(U3173) );
  AND2_X1 U7695 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6737), .ZN(U3174) );
  AND2_X1 U7696 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6737), .ZN(U3175) );
  AND2_X1 U7697 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6737), .ZN(U3176) );
  AND2_X1 U7698 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6737), .ZN(U3177) );
  AND2_X1 U7699 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6737), .ZN(U3178) );
  AND2_X1 U7700 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6737), .ZN(U3179) );
  AND2_X1 U7701 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6737), .ZN(U3180) );
  INV_X1 U7702 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U7703 ( .A1(n6751), .A2(n6858), .B1(n6888), .B2(n6750), .ZN(U3445)
         );
  MUX2_X1 U7704 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6750), .Z(U3446) );
  MUX2_X1 U7705 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6750), .Z(U3447) );
  INV_X1 U7706 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6748) );
  INV_X1 U7707 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7708 ( .A1(n6751), .A2(n6748), .B1(n6815), .B2(n6750), .ZN(U3448)
         );
  OAI21_X1 U7709 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6741), .A(n6739), .ZN(
        n6738) );
  INV_X1 U7710 ( .A(n6738), .ZN(U3451) );
  OAI21_X1 U7711 ( .B1(n6741), .B2(n6740), .A(n6739), .ZN(U3452) );
  AOI21_X1 U7712 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7713 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6743), .B2(n6742), .ZN(n6746) );
  INV_X1 U7714 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6745) );
  AOI22_X1 U7715 ( .A1(n6749), .A2(n6746), .B1(n6745), .B2(n6744), .ZN(U3468)
         );
  OAI21_X1 U7716 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6749), .ZN(n6747) );
  OAI21_X1 U7717 ( .B1(n6749), .B2(n6748), .A(n6747), .ZN(U3469) );
  INV_X1 U7718 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6953) );
  MUX2_X1 U7719 ( .A(n6953), .B(W_R_N_REG_SCAN_IN), .S(n6750), .Z(U3470) );
  INV_X1 U7720 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7721 ( .A1(n6751), .A2(n6856), .B1(n6968), .B2(n6750), .ZN(U3473)
         );
  OAI21_X1 U7722 ( .B1(n6753), .B2(n6752), .A(n6756), .ZN(n6754) );
  OAI211_X1 U7723 ( .C1(n6756), .C2(n6953), .A(n6755), .B(n6754), .ZN(U3474)
         );
  NOR4_X1 U7724 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(EAX_REG_21__SCAN_IN), 
        .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(
        n6757) );
  NAND4_X1 U7725 ( .A1(EBX_REG_10__SCAN_IN), .A2(DATAO_REG_4__SCAN_IN), .A3(
        n6757), .A4(n7019), .ZN(n6765) );
  INV_X1 U7726 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n7048) );
  NAND4_X1 U7727 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(DATAO_REG_28__SCAN_IN), .A3(UWORD_REG_14__SCAN_IN), .A4(n7048), .ZN(n6764) );
  NAND4_X1 U7728 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(UWORD_REG_3__SCAN_IN), 
        .A3(n4295), .A4(n7043), .ZN(n6763) );
  NOR4_X1 U7729 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(DATAI_29_), .A3(n7003), 
        .A4(n6994), .ZN(n6761) );
  NOR4_X1 U7730 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(MORE_REG_SCAN_IN), 
        .A3(DATAO_REG_7__SCAN_IN), .A4(n6998), .ZN(n6760) );
  NOR4_X1 U7731 ( .A1(LWORD_REG_0__SCAN_IN), .A2(DATAO_REG_24__SCAN_IN), .A3(
        n7025), .A4(n7028), .ZN(n6759) );
  NOR4_X1 U7732 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        REIP_REG_16__SCAN_IN), .A3(n3867), .A4(n7031), .ZN(n6758) );
  NAND4_X1 U7733 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6762)
         );
  NOR4_X1 U7734 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6806)
         );
  INV_X1 U7735 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6875) );
  NAND4_X1 U7736 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(
        INSTQUEUE_REG_15__0__SCAN_IN), .A3(UWORD_REG_6__SCAN_IN), .A4(n6875), 
        .ZN(n6804) );
  NAND4_X1 U7737 ( .A1(EBX_REG_21__SCAN_IN), .A2(BYTEENABLE_REG_3__SCAN_IN), 
        .A3(UWORD_REG_1__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6803)
         );
  NAND4_X1 U7738 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTQUEUE_REG_12__3__SCAN_IN), .A3(n6903), .A4(n6902), .ZN(n6766) );
  NOR3_X1 U7739 ( .A1(DATAI_7_), .A2(ADDRESS_REG_26__SCAN_IN), .A3(n6766), 
        .ZN(n6774) );
  INV_X1 U7740 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6878) );
  NAND4_X1 U7741 ( .A1(EBX_REG_25__SCAN_IN), .A2(UWORD_REG_0__SCAN_IN), .A3(
        n6878), .A4(n6885), .ZN(n6772) );
  NAND4_X1 U7742 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        REIP_REG_8__SCAN_IN), .A3(BE_N_REG_3__SCAN_IN), .A4(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6771) );
  INV_X1 U7743 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6769) );
  INV_X1 U7744 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6921) );
  NAND4_X1 U7745 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(
        INSTQUEUE_REG_2__4__SCAN_IN), .A3(ADDRESS_REG_3__SCAN_IN), .A4(n6908), 
        .ZN(n6767) );
  NOR2_X1 U7746 ( .A1(DATAI_31_), .A2(n6767), .ZN(n6768) );
  NAND4_X1 U7747 ( .A1(n6769), .A2(n6921), .A3(UWORD_REG_11__SCAN_IN), .A4(
        n6768), .ZN(n6770) );
  NOR3_X1 U7748 ( .A1(n6772), .A2(n6771), .A3(n6770), .ZN(n6773) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6893) );
  NAND4_X1 U7750 ( .A1(BS16_N), .A2(n6774), .A3(n6773), .A4(n6893), .ZN(n6802)
         );
  INV_X1 U7751 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6817) );
  NOR4_X1 U7752 ( .A1(STATE_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A3(EBX_REG_6__SCAN_IN), .A4(n6817), 
        .ZN(n6775) );
  INV_X1 U7753 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6824) );
  NAND3_X1 U7754 ( .A1(DATAI_10_), .A2(n6775), .A3(n6824), .ZN(n6784) );
  NAND4_X1 U7755 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), 
        .A3(BE_N_REG_0__SCAN_IN), .A4(UWORD_REG_13__SCAN_IN), .ZN(n6776) );
  NOR3_X1 U7756 ( .A1(DATAO_REG_26__SCAN_IN), .A2(n6809), .A3(n6776), .ZN(
        n6782) );
  INV_X1 U7757 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6842) );
  NAND4_X1 U7758 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        INSTQUEUE_REG_13__6__SCAN_IN), .A3(n6842), .A4(n6839), .ZN(n6780) );
  INV_X1 U7759 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6835) );
  NAND4_X1 U7760 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n6835), .A3(n6825), 
        .A4(n6836), .ZN(n6779) );
  NAND4_X1 U7761 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(MEMORYFETCH_REG_SCAN_IN), .A3(n4312), .A4(n6853), .ZN(n6778) );
  NAND4_X1 U7762 ( .A1(EBX_REG_24__SCAN_IN), .A2(DATAI_28_), .A3(n6851), .A4(
        n4285), .ZN(n6777) );
  NOR4_X1 U7763 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6781)
         );
  NAND4_X1 U7764 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(
        INSTQUEUE_REG_7__5__SCAN_IN), .A3(n6782), .A4(n6781), .ZN(n6783) );
  NOR4_X1 U7765 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6785), .A3(n6784), 
        .A4(n6783), .ZN(n6800) );
  INV_X1 U7766 ( .A(DATAI_8_), .ZN(n6947) );
  NOR4_X1 U7767 ( .A1(EAX_REG_2__SCAN_IN), .A2(DATAI_12_), .A3(n6947), .A4(
        n6953), .ZN(n6799) );
  INV_X1 U7768 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6975) );
  INV_X1 U7769 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6977) );
  NOR4_X1 U7770 ( .A1(EAX_REG_0__SCAN_IN), .A2(ADDRESS_REG_5__SCAN_IN), .A3(
        n6975), .A4(n6977), .ZN(n6789) );
  NOR4_X1 U7771 ( .A1(STATE2_REG_2__SCAN_IN), .A2(EAX_REG_15__SCAN_IN), .A3(
        UWORD_REG_4__SCAN_IN), .A4(n4039), .ZN(n6788) );
  NOR4_X1 U7772 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A3(ADS_N_REG_SCAN_IN), .A4(
        M_IO_N_REG_SCAN_IN), .ZN(n6787) );
  NOR4_X1 U7773 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(PHYADDRPOINTER_REG_20__SCAN_IN), 
        .A4(n6980), .ZN(n6786) );
  NAND4_X1 U7774 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6797)
         );
  INV_X1 U7775 ( .A(DATAI_14_), .ZN(n6791) );
  INV_X1 U7776 ( .A(DATAI_18_), .ZN(n6790) );
  NAND4_X1 U7777 ( .A1(n6791), .A2(n6790), .A3(n6938), .A4(
        REIP_REG_26__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U7778 ( .A1(n4701), .A2(DATAO_REG_15__SCAN_IN), .ZN(n6795) );
  INV_X1 U7779 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6793) );
  NOR3_X1 U7780 ( .A1(n4143), .A2(n6950), .A3(n6178), .ZN(n6792) );
  NAND4_X1 U7781 ( .A1(n6793), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .A3(
        INSTQUEUE_REG_9__7__SCAN_IN), .A4(n6792), .ZN(n6794) );
  NOR4_X1 U7782 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6798)
         );
  NAND3_X1 U7783 ( .A1(n6800), .A2(n6799), .A3(n6798), .ZN(n6801) );
  NOR4_X1 U7784 ( .A1(n6804), .A2(n6803), .A3(n6802), .A4(n6801), .ZN(n6805)
         );
  AOI21_X1 U7785 ( .B1(n6806), .B2(n6805), .A(DATAO_REG_11__SCAN_IN), .ZN(
        n7062) );
  AOI22_X1 U7786 ( .A1(n6809), .A2(keyinput23), .B1(keyinput4), .B2(n6808), 
        .ZN(n6807) );
  OAI221_X1 U7787 ( .B1(n6809), .B2(keyinput23), .C1(n6808), .C2(keyinput4), 
        .A(n6807), .ZN(n6821) );
  INV_X1 U7788 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6812) );
  AOI22_X1 U7789 ( .A1(n6812), .A2(keyinput53), .B1(keyinput20), .B2(n6811), 
        .ZN(n6810) );
  OAI221_X1 U7790 ( .B1(n6812), .B2(keyinput53), .C1(n6811), .C2(keyinput20), 
        .A(n6810), .ZN(n6820) );
  AOI22_X1 U7791 ( .A1(n6815), .A2(keyinput10), .B1(keyinput30), .B2(n6814), 
        .ZN(n6813) );
  OAI221_X1 U7792 ( .B1(n6815), .B2(keyinput10), .C1(n6814), .C2(keyinput30), 
        .A(n6813), .ZN(n6819) );
  AOI22_X1 U7793 ( .A1(n6817), .A2(keyinput26), .B1(n4155), .B2(keyinput79), 
        .ZN(n6816) );
  OAI221_X1 U7794 ( .B1(n6817), .B2(keyinput26), .C1(n4155), .C2(keyinput79), 
        .A(n6816), .ZN(n6818) );
  NOR4_X1 U7795 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6866)
         );
  INV_X1 U7796 ( .A(DATAI_10_), .ZN(n6823) );
  AOI22_X1 U7797 ( .A1(n6824), .A2(keyinput105), .B1(keyinput33), .B2(n6823), 
        .ZN(n6822) );
  OAI221_X1 U7798 ( .B1(n6824), .B2(keyinput105), .C1(n6823), .C2(keyinput33), 
        .A(n6822), .ZN(n6833) );
  XNOR2_X1 U7799 ( .A(n6825), .B(keyinput83), .ZN(n6832) );
  XOR2_X1 U7800 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .B(keyinput1), .Z(n6831) );
  XNOR2_X1 U7801 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .B(keyinput28), .ZN(
        n6829) );
  XNOR2_X1 U7802 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput52), .ZN(
        n6828) );
  XNOR2_X1 U7803 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(keyinput92), .ZN(
        n6827) );
  XNOR2_X1 U7804 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput21), .ZN(n6826) );
  NAND4_X1 U7805 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6830)
         );
  NOR4_X1 U7806 ( .A1(n6833), .A2(n6832), .A3(n6831), .A4(n6830), .ZN(n6865)
         );
  AOI22_X1 U7807 ( .A1(n6836), .A2(keyinput120), .B1(n6835), .B2(keyinput74), 
        .ZN(n6834) );
  OAI221_X1 U7808 ( .B1(n6836), .B2(keyinput120), .C1(n6835), .C2(keyinput74), 
        .A(n6834), .ZN(n6848) );
  INV_X1 U7809 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7810 ( .A1(n6839), .A2(keyinput51), .B1(n6838), .B2(keyinput103), 
        .ZN(n6837) );
  OAI221_X1 U7811 ( .B1(n6839), .B2(keyinput51), .C1(n6838), .C2(keyinput103), 
        .A(n6837), .ZN(n6847) );
  INV_X1 U7812 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6841) );
  AOI22_X1 U7813 ( .A1(n6842), .A2(keyinput34), .B1(keyinput27), .B2(n6841), 
        .ZN(n6840) );
  OAI221_X1 U7814 ( .B1(n6842), .B2(keyinput34), .C1(n6841), .C2(keyinput27), 
        .A(n6840), .ZN(n6846) );
  INV_X1 U7815 ( .A(DATAI_28_), .ZN(n6844) );
  AOI22_X1 U7816 ( .A1(n6844), .A2(keyinput72), .B1(n4285), .B2(keyinput55), 
        .ZN(n6843) );
  OAI221_X1 U7817 ( .B1(n6844), .B2(keyinput72), .C1(n4285), .C2(keyinput55), 
        .A(n6843), .ZN(n6845) );
  NOR4_X1 U7818 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6864)
         );
  AOI22_X1 U7819 ( .A1(n6851), .A2(keyinput41), .B1(keyinput119), .B2(n6850), 
        .ZN(n6849) );
  OAI221_X1 U7820 ( .B1(n6851), .B2(keyinput41), .C1(n6850), .C2(keyinput119), 
        .A(n6849), .ZN(n6862) );
  AOI22_X1 U7821 ( .A1(n6854), .A2(keyinput88), .B1(n6853), .B2(keyinput65), 
        .ZN(n6852) );
  OAI221_X1 U7822 ( .B1(n6854), .B2(keyinput88), .C1(n6853), .C2(keyinput65), 
        .A(n6852), .ZN(n6861) );
  AOI22_X1 U7823 ( .A1(n4312), .A2(keyinput112), .B1(keyinput93), .B2(n6856), 
        .ZN(n6855) );
  OAI221_X1 U7824 ( .B1(n4312), .B2(keyinput112), .C1(n6856), .C2(keyinput93), 
        .A(n6855), .ZN(n6860) );
  AOI22_X1 U7825 ( .A1(n5604), .A2(keyinput16), .B1(keyinput96), .B2(n6858), 
        .ZN(n6857) );
  OAI221_X1 U7826 ( .B1(n5604), .B2(keyinput16), .C1(n6858), .C2(keyinput96), 
        .A(n6857), .ZN(n6859) );
  NOR4_X1 U7827 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6863)
         );
  NAND4_X1 U7828 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n7060)
         );
  AOI22_X1 U7829 ( .A1(n6869), .A2(keyinput43), .B1(keyinput11), .B2(n6868), 
        .ZN(n6867) );
  OAI221_X1 U7830 ( .B1(n6869), .B2(keyinput43), .C1(n6868), .C2(keyinput11), 
        .A(n6867), .ZN(n6882) );
  AOI22_X1 U7831 ( .A1(n6872), .A2(keyinput80), .B1(n6871), .B2(keyinput39), 
        .ZN(n6870) );
  OAI221_X1 U7832 ( .B1(n6872), .B2(keyinput80), .C1(n6871), .C2(keyinput39), 
        .A(n6870), .ZN(n6881) );
  INV_X1 U7833 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6874) );
  AOI22_X1 U7834 ( .A1(n6875), .A2(keyinput100), .B1(keyinput18), .B2(n6874), 
        .ZN(n6873) );
  OAI221_X1 U7835 ( .B1(n6875), .B2(keyinput100), .C1(n6874), .C2(keyinput18), 
        .A(n6873), .ZN(n6880) );
  INV_X1 U7836 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6877) );
  AOI22_X1 U7837 ( .A1(n6878), .A2(keyinput14), .B1(keyinput31), .B2(n6877), 
        .ZN(n6876) );
  OAI221_X1 U7838 ( .B1(n6878), .B2(keyinput14), .C1(n6877), .C2(keyinput31), 
        .A(n6876), .ZN(n6879) );
  NOR4_X1 U7839 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n6931)
         );
  AOI22_X1 U7840 ( .A1(n6885), .A2(keyinput73), .B1(n6884), .B2(keyinput82), 
        .ZN(n6883) );
  OAI221_X1 U7841 ( .B1(n6885), .B2(keyinput73), .C1(n6884), .C2(keyinput82), 
        .A(n6883), .ZN(n6897) );
  AOI22_X1 U7842 ( .A1(n6888), .A2(keyinput35), .B1(keyinput2), .B2(n6887), 
        .ZN(n6886) );
  OAI221_X1 U7843 ( .B1(n6888), .B2(keyinput35), .C1(n6887), .C2(keyinput2), 
        .A(n6886), .ZN(n6896) );
  AOI22_X1 U7844 ( .A1(n6890), .A2(keyinput17), .B1(n4113), .B2(keyinput24), 
        .ZN(n6889) );
  OAI221_X1 U7845 ( .B1(n6890), .B2(keyinput17), .C1(n4113), .C2(keyinput24), 
        .A(n6889), .ZN(n6895) );
  INV_X1 U7846 ( .A(BS16_N), .ZN(n6892) );
  AOI22_X1 U7847 ( .A1(n6893), .A2(keyinput127), .B1(keyinput60), .B2(n6892), 
        .ZN(n6891) );
  OAI221_X1 U7848 ( .B1(n6893), .B2(keyinput127), .C1(n6892), .C2(keyinput60), 
        .A(n6891), .ZN(n6894) );
  NOR4_X1 U7849 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6930)
         );
  INV_X1 U7850 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U7851 ( .A1(n6900), .A2(keyinput116), .B1(keyinput5), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7852 ( .B1(n6900), .B2(keyinput116), .C1(n6899), .C2(keyinput5), 
        .A(n6898), .ZN(n6913) );
  AOI22_X1 U7853 ( .A1(n6903), .A2(keyinput61), .B1(keyinput121), .B2(n6902), 
        .ZN(n6901) );
  OAI221_X1 U7854 ( .B1(n6903), .B2(keyinput61), .C1(n6902), .C2(keyinput121), 
        .A(n6901), .ZN(n6912) );
  AOI22_X1 U7855 ( .A1(n6906), .A2(keyinput110), .B1(keyinput13), .B2(n6905), 
        .ZN(n6904) );
  OAI221_X1 U7856 ( .B1(n6906), .B2(keyinput110), .C1(n6905), .C2(keyinput13), 
        .A(n6904), .ZN(n6911) );
  INV_X1 U7857 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7858 ( .A1(n6909), .A2(keyinput68), .B1(keyinput95), .B2(n6908), 
        .ZN(n6907) );
  OAI221_X1 U7859 ( .B1(n6909), .B2(keyinput68), .C1(n6908), .C2(keyinput95), 
        .A(n6907), .ZN(n6910) );
  NOR4_X1 U7860 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n6929)
         );
  AOI22_X1 U7861 ( .A1(n6915), .A2(keyinput59), .B1(n4170), .B2(keyinput81), 
        .ZN(n6914) );
  OAI221_X1 U7862 ( .B1(n6915), .B2(keyinput59), .C1(n4170), .C2(keyinput81), 
        .A(n6914), .ZN(n6927) );
  INV_X1 U7863 ( .A(DATAI_31_), .ZN(n6917) );
  AOI22_X1 U7864 ( .A1(n4966), .A2(keyinput66), .B1(keyinput32), .B2(n6917), 
        .ZN(n6916) );
  OAI221_X1 U7865 ( .B1(n4966), .B2(keyinput66), .C1(n6917), .C2(keyinput32), 
        .A(n6916), .ZN(n6926) );
  INV_X1 U7866 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U7867 ( .A1(n6920), .A2(keyinput25), .B1(keyinput77), .B2(n6919), 
        .ZN(n6918) );
  OAI221_X1 U7868 ( .B1(n6920), .B2(keyinput25), .C1(n6919), .C2(keyinput77), 
        .A(n6918), .ZN(n6925) );
  XOR2_X1 U7869 ( .A(n6921), .B(keyinput85), .Z(n6923) );
  XNOR2_X1 U7870 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .B(keyinput64), .ZN(n6922)
         );
  NAND2_X1 U7871 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  NOR4_X1 U7872 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(n6928)
         );
  NAND4_X1 U7873 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n7059)
         );
  INV_X1 U7874 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n6933) );
  AOI22_X1 U7875 ( .A1(n6934), .A2(keyinput123), .B1(keyinput91), .B2(n6933), 
        .ZN(n6932) );
  OAI221_X1 U7876 ( .B1(n6934), .B2(keyinput123), .C1(n6933), .C2(keyinput91), 
        .A(n6932), .ZN(n6944) );
  AOI22_X1 U7877 ( .A1(n6936), .A2(keyinput6), .B1(n4039), .B2(keyinput125), 
        .ZN(n6935) );
  OAI221_X1 U7878 ( .B1(n6936), .B2(keyinput6), .C1(n4039), .C2(keyinput125), 
        .A(n6935), .ZN(n6943) );
  AOI22_X1 U7879 ( .A1(n4143), .A2(keyinput71), .B1(n6938), .B2(keyinput9), 
        .ZN(n6937) );
  OAI221_X1 U7880 ( .B1(n4143), .B2(keyinput71), .C1(n6938), .C2(keyinput9), 
        .A(n6937), .ZN(n6942) );
  XOR2_X1 U7881 ( .A(n6790), .B(keyinput63), .Z(n6940) );
  XNOR2_X1 U7882 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput62), .ZN(n6939)
         );
  NAND2_X1 U7883 ( .A1(n6940), .A2(n6939), .ZN(n6941) );
  NOR4_X1 U7884 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6992)
         );
  AOI22_X1 U7885 ( .A1(n6947), .A2(keyinput84), .B1(n6946), .B2(keyinput76), 
        .ZN(n6945) );
  OAI221_X1 U7886 ( .B1(n6947), .B2(keyinput84), .C1(n6946), .C2(keyinput76), 
        .A(n6945), .ZN(n6957) );
  AOI22_X1 U7887 ( .A1(n6178), .A2(keyinput98), .B1(keyinput94), .B2(n6791), 
        .ZN(n6948) );
  OAI221_X1 U7888 ( .B1(n6178), .B2(keyinput98), .C1(n6791), .C2(keyinput94), 
        .A(n6948), .ZN(n6956) );
  AOI22_X1 U7889 ( .A1(n6950), .A2(keyinput42), .B1(n6793), .B2(keyinput15), 
        .ZN(n6949) );
  OAI221_X1 U7890 ( .B1(n6950), .B2(keyinput42), .C1(n6793), .C2(keyinput15), 
        .A(n6949), .ZN(n6955) );
  INV_X1 U7891 ( .A(DATAI_12_), .ZN(n6952) );
  AOI22_X1 U7892 ( .A1(n6953), .A2(keyinput108), .B1(n6952), .B2(keyinput78), 
        .ZN(n6951) );
  OAI221_X1 U7893 ( .B1(n6953), .B2(keyinput108), .C1(n6952), .C2(keyinput78), 
        .A(n6951), .ZN(n6954) );
  NOR4_X1 U7894 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6991)
         );
  AOI22_X1 U7895 ( .A1(n6960), .A2(keyinput107), .B1(keyinput22), .B2(n6959), 
        .ZN(n6958) );
  OAI221_X1 U7896 ( .B1(n6960), .B2(keyinput107), .C1(n6959), .C2(keyinput22), 
        .A(n6958), .ZN(n6972) );
  AOI22_X1 U7897 ( .A1(n6963), .A2(keyinput111), .B1(keyinput37), .B2(n6962), 
        .ZN(n6961) );
  OAI221_X1 U7898 ( .B1(n6963), .B2(keyinput111), .C1(n6962), .C2(keyinput37), 
        .A(n6961), .ZN(n6971) );
  INV_X1 U7899 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6966) );
  AOI22_X1 U7900 ( .A1(n6966), .A2(keyinput86), .B1(n6965), .B2(keyinput40), 
        .ZN(n6964) );
  OAI221_X1 U7901 ( .B1(n6966), .B2(keyinput86), .C1(n6965), .C2(keyinput40), 
        .A(n6964), .ZN(n6970) );
  AOI22_X1 U7902 ( .A1(n4348), .A2(keyinput7), .B1(keyinput69), .B2(n6968), 
        .ZN(n6967) );
  OAI221_X1 U7903 ( .B1(n4348), .B2(keyinput7), .C1(n6968), .C2(keyinput69), 
        .A(n6967), .ZN(n6969) );
  NOR4_X1 U7904 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n6990)
         );
  AOI22_X1 U7905 ( .A1(n6975), .A2(keyinput101), .B1(keyinput124), .B2(n6974), 
        .ZN(n6973) );
  OAI221_X1 U7906 ( .B1(n6975), .B2(keyinput101), .C1(n6974), .C2(keyinput124), 
        .A(n6973), .ZN(n6988) );
  AOI22_X1 U7907 ( .A1(n6978), .A2(keyinput47), .B1(n6977), .B2(keyinput45), 
        .ZN(n6976) );
  OAI221_X1 U7908 ( .B1(n6978), .B2(keyinput47), .C1(n6977), .C2(keyinput45), 
        .A(n6976), .ZN(n6987) );
  INV_X1 U7909 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6981) );
  AOI22_X1 U7910 ( .A1(n6981), .A2(keyinput58), .B1(keyinput122), .B2(n6980), 
        .ZN(n6979) );
  OAI221_X1 U7911 ( .B1(n6981), .B2(keyinput58), .C1(n6980), .C2(keyinput122), 
        .A(n6979), .ZN(n6986) );
  INV_X1 U7912 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6982) );
  XOR2_X1 U7913 ( .A(n6982), .B(keyinput44), .Z(n6984) );
  XNOR2_X1 U7914 ( .A(STATE2_REG_2__SCAN_IN), .B(keyinput89), .ZN(n6983) );
  NAND2_X1 U7915 ( .A1(n6984), .A2(n6983), .ZN(n6985) );
  NOR4_X1 U7916 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n6989)
         );
  NAND4_X1 U7917 ( .A1(n6992), .A2(n6991), .A3(n6990), .A4(n6989), .ZN(n7058)
         );
  INV_X1 U7918 ( .A(DATAI_29_), .ZN(n6995) );
  AOI22_X1 U7919 ( .A1(n6995), .A2(keyinput49), .B1(keyinput70), .B2(n6994), 
        .ZN(n6993) );
  OAI221_X1 U7920 ( .B1(n6995), .B2(keyinput49), .C1(n6994), .C2(keyinput70), 
        .A(n6993), .ZN(n7008) );
  INV_X1 U7921 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U7922 ( .A1(n6998), .A2(keyinput106), .B1(n6997), .B2(keyinput46), 
        .ZN(n6996) );
  OAI221_X1 U7923 ( .B1(n6998), .B2(keyinput106), .C1(n6997), .C2(keyinput46), 
        .A(n6996), .ZN(n7007) );
  INV_X1 U7924 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n7001) );
  AOI22_X1 U7925 ( .A1(n7001), .A2(keyinput48), .B1(keyinput0), .B2(n7000), 
        .ZN(n6999) );
  OAI221_X1 U7926 ( .B1(n7001), .B2(keyinput48), .C1(n7000), .C2(keyinput0), 
        .A(n6999), .ZN(n7006) );
  AOI22_X1 U7927 ( .A1(n7004), .A2(keyinput102), .B1(n7003), .B2(keyinput109), 
        .ZN(n7002) );
  OAI221_X1 U7928 ( .B1(n7004), .B2(keyinput102), .C1(n7003), .C2(keyinput109), 
        .A(n7002), .ZN(n7005) );
  NOR4_X1 U7929 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), .ZN(n7056)
         );
  INV_X1 U7930 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7931 ( .A1(keyinput117), .A2(n7011), .B1(keyinput99), .B2(n7009), 
        .ZN(n7010) );
  OAI21_X1 U7932 ( .B1(n7011), .B2(keyinput117), .A(n7010), .ZN(n7023) );
  AOI22_X1 U7933 ( .A1(n7013), .A2(keyinput50), .B1(n4986), .B2(keyinput54), 
        .ZN(n7012) );
  OAI221_X1 U7934 ( .B1(n7013), .B2(keyinput50), .C1(n4986), .C2(keyinput54), 
        .A(n7012), .ZN(n7022) );
  INV_X1 U7935 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n7015) );
  AOI22_X1 U7936 ( .A1(n7016), .A2(keyinput57), .B1(keyinput56), .B2(n7015), 
        .ZN(n7014) );
  OAI221_X1 U7937 ( .B1(n7016), .B2(keyinput57), .C1(n7015), .C2(keyinput56), 
        .A(n7014), .ZN(n7021) );
  AOI22_X1 U7938 ( .A1(n7019), .A2(keyinput97), .B1(keyinput115), .B2(n7018), 
        .ZN(n7017) );
  OAI221_X1 U7939 ( .B1(n7019), .B2(keyinput97), .C1(n7018), .C2(keyinput115), 
        .A(n7017), .ZN(n7020) );
  NOR4_X1 U7940 ( .A1(n7023), .A2(n7022), .A3(n7021), .A4(n7020), .ZN(n7055)
         );
  AOI22_X1 U7941 ( .A1(n7026), .A2(keyinput104), .B1(n7025), .B2(keyinput67), 
        .ZN(n7024) );
  OAI221_X1 U7942 ( .B1(n7026), .B2(keyinput104), .C1(n7025), .C2(keyinput67), 
        .A(n7024), .ZN(n7038) );
  AOI22_X1 U7943 ( .A1(n7029), .A2(keyinput38), .B1(n7028), .B2(keyinput113), 
        .ZN(n7027) );
  OAI221_X1 U7944 ( .B1(n7029), .B2(keyinput38), .C1(n7028), .C2(keyinput113), 
        .A(n7027), .ZN(n7037) );
  AOI22_X1 U7945 ( .A1(n7032), .A2(keyinput12), .B1(keyinput126), .B2(n7031), 
        .ZN(n7030) );
  OAI221_X1 U7946 ( .B1(n7032), .B2(keyinput12), .C1(n7031), .C2(keyinput126), 
        .A(n7030), .ZN(n7036) );
  XNOR2_X1 U7947 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .B(keyinput8), .ZN(n7034)
         );
  XNOR2_X1 U7948 ( .A(keyinput29), .B(DATAI_2_), .ZN(n7033) );
  NAND2_X1 U7949 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  NOR4_X1 U7950 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .ZN(n7054)
         );
  INV_X1 U7951 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n7041) );
  AOI22_X1 U7952 ( .A1(n7041), .A2(keyinput3), .B1(keyinput19), .B2(n7040), 
        .ZN(n7039) );
  OAI221_X1 U7953 ( .B1(n7041), .B2(keyinput3), .C1(n7040), .C2(keyinput19), 
        .A(n7039), .ZN(n7052) );
  AOI22_X1 U7954 ( .A1(n7043), .A2(keyinput114), .B1(keyinput118), .B2(n4295), 
        .ZN(n7042) );
  OAI221_X1 U7955 ( .B1(n7043), .B2(keyinput114), .C1(n4295), .C2(keyinput118), 
        .A(n7042), .ZN(n7051) );
  AOI22_X1 U7956 ( .A1(n3867), .A2(keyinput90), .B1(keyinput36), .B2(n7045), 
        .ZN(n7044) );
  OAI221_X1 U7957 ( .B1(n3867), .B2(keyinput90), .C1(n7045), .C2(keyinput36), 
        .A(n7044), .ZN(n7050) );
  AOI22_X1 U7958 ( .A1(n7048), .A2(keyinput75), .B1(keyinput87), .B2(n7047), 
        .ZN(n7046) );
  OAI221_X1 U7959 ( .B1(n7048), .B2(keyinput75), .C1(n7047), .C2(keyinput87), 
        .A(n7046), .ZN(n7049) );
  NOR4_X1 U7960 ( .A1(n7052), .A2(n7051), .A3(n7050), .A4(n7049), .ZN(n7053)
         );
  NAND4_X1 U7961 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), .ZN(n7057)
         );
  NOR4_X1 U7962 ( .A1(n7060), .A2(n7059), .A3(n7058), .A4(n7057), .ZN(n7061)
         );
  OAI21_X1 U7963 ( .B1(keyinput99), .B2(n7062), .A(n7061), .ZN(n7068) );
  OAI222_X1 U7964 ( .A1(n7066), .A2(n7065), .B1(n5628), .B2(n4155), .C1(n7064), 
        .C2(n7063), .ZN(n7067) );
  XNOR2_X1 U7965 ( .A(n7068), .B(n7067), .ZN(U2853) );
  CLKBUF_X2 U3552 ( .A(n3377), .Z(n3353) );
  CLKBUF_X1 U3562 ( .A(n3496), .Z(n3512) );
  CLKBUF_X1 U3570 ( .A(n3494), .Z(n4579) );
  CLKBUF_X1 U3571 ( .A(n4134), .Z(n4684) );
  CLKBUF_X1 U3581 ( .A(n5363), .Z(n3103) );
  CLKBUF_X2 U3636 ( .A(n3520), .Z(n4871) );
  CLKBUF_X1 U3691 ( .A(n4625), .Z(n3102) );
endmodule

